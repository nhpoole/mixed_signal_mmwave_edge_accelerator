* NGSPICE file created from analog_top_level_flat.ext - technology: sky130A

.subckt analog_top_level_flat vintp vintm vfiltp vfiltm vlowA vrefA q7A q6A q5A q4A
+ q3A q2A q1A q0A adc_clk sample vlowB vrefB q7B q6B q5B q4B q3B q2B q1B q0B adc_compA
+ adc_compB vcp vcp_sampled vpeak_sampled vpeak vse vcomp vhpf VDD VSS vincm vocm
+ vocm_filt gain_ctrl_0 gain_ctrl_1 vbiasp vbiasn peak_detector_rst vampm vampp adc_vcaparrayB
+ adc_vcaparrayA rst_n
X0 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1 dac_8bit_1/latched_comparator_folded_0/vtailp dac_8bit_1/latched_comparator_folded_0/vtailp dac_8bit_1/latched_comparator_folded_0/vtailp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4 vlowA VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5 input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vbias3 a_163060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6 VDD a_338356_n185269# a_338285_n185243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X7 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X9 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X10 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X11 a_242085_n122799# a_241919_n122799# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X13 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X14 biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail2 vocm_filt biquad_gm_c_filter_0/gm_c_stage_0/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X16 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X17 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X18 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X19 a_275374_n146348# sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X20 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X21 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X22 comparator_0/vo1 comparator_0/vo1 comparator_0/vo1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X23 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X24 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X25 input_amplifier_0/diff_fold_casc_ota_1/M2d input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X26 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X27 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X28 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X29 dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X30 peak_detector_0/verr VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X31 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X32 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X33 VDD vbiasp dac_8bit_0/ibiasn VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X34 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1.2e+07u w=2e+06u
X35 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X36 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 a_356329_n164260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X37 a_228020_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_227562_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X38 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X39 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X40 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X41 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X42 peak_detector_0/verr peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X43 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X44 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X45 VSS a_245481_n123343# a_245649_n123369# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X46 a_242526_n123369# a_242358_n123343# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X47 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 vocm input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X48 input_amplifier_0/vip2 input_amplifier_0/rst input_amplifier_0/vom1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X49 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X50 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X51 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X52 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X53 VSS input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X54 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X55 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X56 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X57 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X58 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X59 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X60 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X61 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X62 input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X63 vintm VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X64 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X65 vpeak VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X66 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X67 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X68 VSS a_242526_n121193# a_242484_n120789# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X69 input_amplifier_0/diff_fold_casc_ota_0/vcascnm input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X70 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X71 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X72 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X73 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X74 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X75 a_338149_n185569# adc_clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X76 adc_vcaparrayA dac_8bit_0/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X77 dac_8bit_1/c0m dac_8bit_1/amux_2to1_8/SELB vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X78 peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X79 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X80 VDD vbiasp low_freq_pll_0/ibiasn VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X81 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X82 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X83 VSS dac_8bit_0/ibiasn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X84 vfiltp vintp biquad_gm_c_filter_0/gm_c_stage_3/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X85 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X86 vpeak_sampled sample sample_and_hold_1/vholdm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X87 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X88 a_222498_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_222040_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X89 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X90 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/vcom_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X91 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X92 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X93 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X94 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X95 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X96 a_241786_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_241328_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X97 VSS low_freq_pll_0/freq_div_0/vin a_241919_n120623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X98 VDD VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X99 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 a_356329_n113250# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X100 input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vfoldm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X101 dac_8bit_0/latched_comparator_folded_0/vtailp vlowA dac_8bit_0/latched_comparator_folded_0/vlatchm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X102 a_338505_n185243# a_338285_n185243# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X103 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X104 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 a_189446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X105 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X106 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X107 vse VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X108 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X109 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X110 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 vse VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X111 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X112 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X113 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X114 vrefB dac_8bit_1/amux_2to1_10/SELB dac_8bit_1/amux_2to1_7/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X115 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X116 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X117 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X118 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X119 vcp_sampled VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X120 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X121 VDD a_245224_n123369# a_245151_n123343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X122 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X123 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X124 input_amplifier_0/txgate_0/txb gain_ctrl_0 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X125 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X126 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X127 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X128 dac_8bit_1/latched_comparator_folded_0/vlatchp dac_8bit_1/vcom_buf dac_8bit_1/latched_comparator_folded_0/vtailp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X129 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X130 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X131 peak_detector_0/verr peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X132 input_amplifier_0/diff_fold_casc_ota_1/vcascnm input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X133 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X134 dac_8bit_0/amux_2to1_10/SELB q1A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X135 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X136 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X137 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/vip2 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X138 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X139 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X140 vampm VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X141 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 vocm input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X142 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X143 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X144 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 a_189446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X145 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X146 VSS VSS vampm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X147 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X148 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X149 vrefB dac_8bit_1/amux_2to1_13/SELB dac_8bit_1/amux_2to1_4/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X150 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X151 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X152 vrefA VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X153 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X154 VDD a_242526_n120511# a_242453_n120257# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X155 a_239048_n115125# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X156 adc_vcaparrayB dac_8bit_1/c3m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X157 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X158 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X159 vlowB VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X160 vpeak sample sample_and_hold_1/vhold VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X161 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X162 VDD a_242951_n121443# a_243382_n121389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X163 a_245056_n123343# a_244617_n123337# a_244971_n123343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X164 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X165 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X166 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X167 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X168 biquad_gm_c_filter_0/gm_c_stage_0/vbiasp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X169 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X170 a_241481_n130007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_241023_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X171 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X172 VDD VDD low_freq_pll_0/pfd_cp_lpf_0/vpbias VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X173 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X174 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X175 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X176 dac_8bit_0/amux_2to1_13/SELB q3A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X177 biquad_gm_c_filter_0/ibiasn1 biquad_gm_c_filter_0/ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X178 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X179 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X180 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X181 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X182 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X183 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X184 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 vpeak_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X185 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X186 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/csinvn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X187 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X188 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X189 vrefB dac_8bit_1/amux_2to1_16/SELB dac_8bit_1/amux_2to1_1/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X190 vrefA VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X191 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X192 a_241785_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_241327_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X193 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X194 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q a_242951_n123369# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X195 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X196 input_amplifier_0/diff_fold_casc_ota_0/vcascnm input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/vom1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X197 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X198 vlowB VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X199 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X200 VDD input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X201 input_amplifier_0/diff_fold_casc_ota_0/vcascnm input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/vom1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X202 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X203 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X204 a_275374_n180872# sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X205 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X206 VDD biquad_gm_c_filter_0/gm_c_stage_0/vcmcn1 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X207 a_243770_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_243312_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X208 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X209 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X210 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X211 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X212 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X213 vampm vampm vampm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X214 a_338356_n185510# a_338149_n185569# a_338532_n185787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X215 a_245481_n122433# a_244783_n122799# a_245224_n122687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X216 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X217 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X218 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X219 a_163060_n102324# input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X220 dac_8bit_0/amux_2to1_16/SELB q6A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X221 diff_to_se_converter_0/vim vfiltm sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X222 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X223 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X224 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X225 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X226 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X227 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X228 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X229 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X230 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X231 VDD VDD dac_8bit_1/latched_comparator_folded_0/vlatchp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X232 dac_8bit_0/amux_2to1_0/SELB sample VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X233 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X234 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X235 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 a_162668_n147576# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X236 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 a_275374_n146348# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X237 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X238 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X239 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X240 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X241 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X242 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X243 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 a_162668_n147576# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X244 VSS diff_to_se_converter_0/ibiasn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X245 biquad_gm_c_filter_0/gm_c_stage_1/vbiasp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X246 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X247 vcp_sampled sample dac_8bit_0/c0m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X248 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X249 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X250 VDD vbiasp input_amplifier_0/ibiasn2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X251 VSS VSS diff_to_se_converter_0/vim VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X252 VSS input_amplifier_0/ibiasn2 input_amplifier_0/ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X253 input_amplifier_0/diff_fold_casc_ota_0/vcascnp input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X254 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X255 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X256 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X257 a_245182_n121877# a_244783_n122249# a_245056_n122255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X258 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X259 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X260 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X261 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X262 input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X263 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X264 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X265 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X266 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X267 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X268 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X269 a_222396_n131500# low_freq_pll_0/cs_ring_osc_0/vosc a_221938_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X270 input_amplifier_0/ibiasn1 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X271 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X272 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X273 a_246786_n134960# vcp a_246328_n134960# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X274 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X275 VDD input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X276 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X277 a_242562_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_242104_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X278 input_amplifier_0/vim2 input_amplifier_0/rst input_amplifier_0/vop1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X279 dac_8bit_0/latched_comparator_folded_0/vlatchp VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X280 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X281 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X282 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X283 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X284 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X285 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X286 VDD biquad_gm_c_filter_0/gm_c_stage_1/vcmcn1 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X287 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X288 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X289 VSS VSS biquad_gm_c_filter_0/gm_c_stage_0/vtail_diff VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X290 VDD a_245649_n121193# a_246080_n121167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X291 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X292 dac_8bit_0/amux_2to1_9/Y dac_8bit_0/amux_2to1_9/SELB vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X293 VSS input_amplifier_0/ibiasn1 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X294 dac_8bit_1/c2m sample dac_8bit_1/amux_2to1_5/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X295 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X296 dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X297 a_228313_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_227855_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X298 dac_8bit_0/c2m dac_8bit_0/amux_2to1_5/SELB vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X299 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X300 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X301 a_239708_n115125# a_238627_n115125# a_239361_n114883# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X302 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X303 input_amplifier_0/venp1 input_amplifier_0/txgate_1/txb input_amplifier_0/vim2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X304 input_amplifier_0/vom1 input_amplifier_0/vip1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X305 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X306 a_356329_n113250# dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X307 a_242085_n122249# a_241919_n122249# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X308 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X309 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_244617_n122249# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X310 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X311 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X312 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X313 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X314 VSS input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X315 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X316 VDD input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X317 a_244971_n123343# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X318 comparator_0/ibiasn vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X319 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X320 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X321 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X322 input_amplifier_0/venm1 input_amplifier_0/txgate_0/txb input_amplifier_0/vip2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X323 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X324 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X325 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X326 diff_to_se_converter_0/vim diff_to_se_converter_0/txgate_1/txb vfiltm VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X327 a_236582_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X328 input_amplifier_0/diff_fold_casc_ota_0/vcascnm input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/vom1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X329 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X330 dac_8bit_1/c5m sample dac_8bit_1/amux_2to1_2/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X331 dac_8bit_0/c5m dac_8bit_0/amux_2to1_2/SELB vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X332 vlowA dac_8bit_0/adc_run adc_vcaparrayA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X333 input_amplifier_0/vim1 vincm sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X334 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X335 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X336 input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X337 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X338 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X339 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 a_230446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X340 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X341 dac_8bit_0/amux_2to1_6/SELB sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X342 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X343 input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/diff_fold_casc_ota_0/M2d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X344 VDD vbiasp vcp_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X345 vlowB q2B dac_8bit_1/amux_2to1_5/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X346 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X347 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X348 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X349 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/csinvn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X350 VDD vbiasp biquad_gm_c_filter_0/ibiasn3 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X351 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X352 biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail1 vfiltp biquad_gm_c_filter_0/gm_c_stage_3/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X353 vrefB VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X354 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X355 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X356 peak_detector_0/verr peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X357 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X358 a_275374_n146348# sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X359 a_243478_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X360 a_189446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X361 VSS a_336608_n185269# a_336537_n185243# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X362 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X363 VSS peak_detector_0/ibiasn1 peak_detector_0/ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X364 a_227412_n119618# vcp low_freq_pll_0/cs_ring_osc_0/vpbias VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X365 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X366 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X367 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X368 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X369 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X370 input_amplifier_0/vim1 vincm sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X371 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.4e+07u
X372 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 vpeak VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X373 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X374 biquad_gm_c_filter_0/gm_c_stage_1/vtail_diff biquad_gm_c_filter_0/ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X375 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X376 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X377 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X378 dac_8bit_0/amux_2to1_3/SELB sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X379 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/vip2 input_amplifier_0/diff_fold_casc_ota_1/vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X380 dac_8bit_1/amux_2to1_11/SELB VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X381 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X382 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X383 VDD dac_8bit_0/latched_comparator_folded_0/vcompp dac_8bit_0/latched_comparator_folded_0/vcomppb VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X384 vlowB q5B dac_8bit_1/amux_2to1_2/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X385 input_amplifier_0/vim1 input_amplifier_0/rst vincm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X386 adc_vcaparrayA dac_8bit_0/c2m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X387 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X388 VDD input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X389 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X390 a_223872_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_223414_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X391 VDD VDD vcp_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X392 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_5/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X393 vampm vampm vampm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X394 VDD a_245649_n122281# a_245565_n122255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X395 vrefB VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X396 dac_8bit_0/vcom_buf dac_8bit_0/vcom_buf dac_8bit_0/vcom_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X397 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X398 VSS low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_242702_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X399 VDD peak_detector_0/verr peak_detector_0/verr VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X400 dac_8bit_0/latched_comparator_folded_0/vlatchp adc_clk dac_8bit_0/latched_comparator_folded_0/vlatchm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X401 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 a_189446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X402 vampm input_amplifier_0/vip2 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X403 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X404 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X405 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X406 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_1/A a_243382_n121167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X407 a_222854_n132168# vcp a_222396_n132168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X408 VDD dac_8bit_0/comp_outm adc_compA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X409 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X410 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X411 biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail2 vocm_filt biquad_gm_c_filter_0/gm_c_stage_1/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X412 VSS VSS low_freq_pll_0/pfd_cp_lpf_0/vpbias VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X413 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X414 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X415 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X416 peak_detector_0/verr peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X417 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X418 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X419 VDD a_245224_n122687# a_245151_n122433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X420 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X421 a_242867_n123343# a_242085_n123337# a_242783_n123343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X422 dac_8bit_1/amux_2to1_14/SELB q4B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X423 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 vcp_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X424 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X425 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q a_244617_n121161# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X426 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X427 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X428 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X429 VDD input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X430 VDD pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A a_338703_n185409# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X431 peak_detector_0/vpeak VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X432 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X433 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X434 a_237396_n132168# vcp a_236938_n132168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X435 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X436 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/vcom_buf VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X437 vrefB VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X438 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X439 dac_8bit_0/amux_2to1_9/SELB q0A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X440 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X441 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X442 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X443 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/diff_fold_casc_ota_0/vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X444 a_356329_n113250# dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X445 dac_8bit_1/vcom_buf VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X446 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X447 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X448 comparator_0/vmirror comparator_0/vcompm VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X449 VDD input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/M1d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X450 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X451 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X452 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X453 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X454 vampp input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X455 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X456 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 a_356329_n113250# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X457 a_229244_n119618# vcp a_228786_n119618# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X458 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 a_189446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X459 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X460 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X461 vse diff_to_se_converter_0/vim sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X462 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X463 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X464 a_242783_n120257# a_242085_n120623# a_242526_n120511# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X465 biquad_gm_c_filter_0/ibiasn1 biquad_gm_c_filter_0/ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X466 vcp_sampled dac_8bit_0/amux_2to1_0/SELB dac_8bit_0/c7m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X467 VDD biquad_gm_c_filter_0/gm_c_stage_2/vcmcn biquad_gm_c_filter_0/gm_c_stage_2/vcmc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X468 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X469 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X470 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X471 VDD input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vfoldm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X472 adc_vcaparrayB dac_8bit_1/c2m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X473 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X474 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_6/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X475 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X476 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 vse VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X477 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X478 a_242453_n121167# a_241919_n121161# a_242358_n121167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X479 biquad_gm_c_filter_0/gm_c_stage_1/vtail_diff vintp vintp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X480 a_338285_n185409# a_338149_n185569# a_337864_n185555# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X481 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X482 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X483 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X484 vpeak_sampled sample sample_and_hold_1/vholdm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X485 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X486 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X487 VSS VSS dac_8bit_0/amux_2to1_6/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X488 comparator_0/vtail comparator_0/ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X489 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X490 VSS peak_detector_0/verr sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X491 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X492 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X493 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X494 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X495 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X496 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X497 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X498 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X499 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn vse peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X500 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/vim2 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X501 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X502 VDD adc_clk dac_8bit_0/latched_comparator_folded_0/vcompm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X503 a_236938_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin a_236480_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X504 dac_8bit_1/c7m dac_8bit_1/amux_2to1_0/SELB vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X505 dac_8bit_0/c7m sample dac_8bit_0/amux_2to1_0/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X506 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X507 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X508 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X509 dac_8bit_1/c1m dac_8bit_1/amux_2to1_7/SELB vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X510 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X511 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_4/A a_243382_n122477# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X512 a_242085_n122799# a_241919_n122799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X513 VDD input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X514 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X515 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X516 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X517 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X518 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X519 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn vintm biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X520 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X521 input_amplifier_0/diff_fold_casc_ota_0/M6d input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X522 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 vpeak_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X523 a_338356_n185269# a_338149_n185269# a_338532_n184877# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X524 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X525 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X526 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X527 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 a_189446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X528 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X529 VSS VSS dac_8bit_0/amux_2to1_3/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X530 dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X531 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X532 VSS vpeak sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X533 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X534 dac_8bit_0/amux_2to1_6/B VSS vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X535 a_239251_n114759# low_freq_pll_0/pfd_cp_lpf_0/vRSTN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X536 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X537 a_245481_n121167# a_244617_n121161# a_245224_n121193# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X538 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X539 VDD dac_8bit_1/ibiasp dac_8bit_1/ibiasp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X540 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn1 vocm_filt biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X541 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X542 VDD adc_clk dac_8bit_0/latched_comparator_folded_0/vcompp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X543 vincm input_amplifier_0/txgate_4/txb input_amplifier_0/vim1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X544 a_245607_n120789# a_244617_n121161# a_245481_n121167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X545 a_189446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X546 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X547 dac_8bit_1/c3m dac_8bit_1/amux_2to1_4/SELB vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X548 a_242855_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_242397_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X549 VDD biquad_gm_c_filter_0/gm_c_stage_3/vcmcn biquad_gm_c_filter_0/gm_c_stage_3/vcmc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X550 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X551 VDD input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X552 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X553 a_239143_n115125# a_238793_n115125# a_239048_n115125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X554 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X555 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X556 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X557 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X558 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 vse VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X559 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X560 dac_8bit_1/amux_2to1_8/SELB sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X561 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X562 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X563 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X564 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X565 a_230446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X566 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X567 a_221938_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin a_221480_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X568 input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vfoldp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X569 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs low_freq_pll_0/cs_ring_osc_0/vosc a_223770_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X570 dac_8bit_0/ibiasp VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=2e+06u
X571 VSS VSS dac_8bit_0/amux_2to1_0/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X572 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_9/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X573 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X574 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X575 VSS biquad_gm_c_filter_0/ibiasn1 biquad_gm_c_filter_0/ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X576 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X577 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X578 dac_8bit_0/amux_2to1_3/B q4A vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X579 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X580 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X581 low_freq_pll_0/pfd_cp_lpf_0/vpbias low_freq_pll_0/pfd_cp_lpf_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X582 VSS VSS low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/csinvn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X583 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X584 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X585 a_217060_n102324# input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X586 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X587 a_275374_n180872# sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X588 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X589 vfiltp diff_to_se_converter_0/txgate_0/txb diff_to_se_converter_0/vip VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X590 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 a_189446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X591 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X592 input_amplifier_0/diff_fold_casc_ota_1/M3d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X593 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X594 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X595 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X596 adc_vcaparrayB dac_8bit_1/adc_run vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X597 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X598 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X599 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X600 dac_8bit_1/c6m dac_8bit_1/amux_2to1_1/SELB vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X601 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X602 VSS VSS sample_and_hold_0/vhold VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X603 vpeak_sampled vpeak_sampled vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X604 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X605 vrefA q0A dac_8bit_0/amux_2to1_9/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X606 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/csinvn vcp a_247702_n134960# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X607 input_amplifier_0/diff_fold_casc_ota_1/M6d input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X608 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X609 vlowB VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X610 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X611 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X612 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X613 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X614 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X615 a_227854_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_227396_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X616 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X617 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X618 comparator_0/vtail comparator_0/ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X619 input_amplifier_0/rst rst_n VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X620 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X621 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X622 VSS diff_to_se_converter_0/ibiasn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X623 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 a_162668_n147576# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X624 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X625 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X626 low_freq_pll_0/freq_div_0/vin low_freq_pll_0/cs_ring_osc_0/vosc2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X627 low_freq_pll_0/pfd_cp_lpf_0/vswitchl VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X628 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X629 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X630 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X631 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_4/A a_243382_n122477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X632 a_275374_n146348# sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X633 a_244971_n122799# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X634 VDD input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X635 VSS biquad_gm_c_filter_0/ibiasn4 biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X636 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X637 diff_to_se_converter_0/vip VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X638 a_238414_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_237956_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X639 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X640 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X641 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X642 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp vse peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X643 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X644 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X645 adc_vcaparrayA dac_8bit_0/c2m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X646 input_amplifier_0/diff_fold_casc_ota_1/vcascnp input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X647 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X648 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 a_162668_n147576# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X649 vlowB VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X650 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X651 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X652 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X653 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 a_217060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X654 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X655 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X656 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X657 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X658 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X659 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X660 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X661 peak_detector_0/verr peak_detector_0/verr peak_detector_0/verr VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X662 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X663 input_amplifier_0/diff_fold_casc_ota_0/M6d input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X664 a_241646_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_242104_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X665 dac_8bit_0/amux_2to1_9/Y dac_8bit_0/amux_2to1_8/SELB dac_8bit_0/c0m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X666 a_245056_n122433# a_244617_n122799# a_244971_n122799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X667 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X668 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X669 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X670 VDD pulse_generator_0/sky130_fd_sc_hd__inv_1_1/A peak_detector_rst VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X671 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X672 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X673 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X674 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X675 VDD a_242783_n121167# a_242951_n121193# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X676 input_amplifier_0/diff_fold_casc_ota_0/M13d input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/M6d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X677 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X678 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X679 input_amplifier_0/diff_fold_casc_ota_0/vcascnm input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X680 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X681 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X682 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X683 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X684 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X685 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X686 adc_vcaparrayB dac_8bit_1/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X687 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X688 input_amplifier_0/vip2 input_amplifier_0/vom1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X689 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X690 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_9/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X691 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X692 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X693 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X694 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X695 a_275374_n146348# sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X696 a_227396_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_226938_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X697 a_242419_n114983# vcomp VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X698 a_223872_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_224330_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X699 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X700 vcp_sampled sample dac_8bit_0/c1m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X701 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X702 input_amplifier_0/diff_fold_casc_ota_0/vcascnp input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X703 VSS VSS dac_8bit_1/amux_2to1_9/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X704 dac_8bit_1/latched_comparator_folded_0/vcompm_buf dac_8bit_1/latched_comparator_folded_0/vcompmb VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X705 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X706 peak_detector_0/verr peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X707 dac_8bit_0/amux_2to1_5/B dac_8bit_0/amux_2to1_5/SELB dac_8bit_0/c2m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X708 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X709 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X710 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X711 VDD a_245649_n121443# a_245565_n121345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X712 VSS input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X713 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X714 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X715 a_239330_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X716 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X717 a_337497_n185813# a_337592_n185460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X718 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X719 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X720 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X721 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X722 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/M2d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X723 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X724 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X725 a_242720_n114759# a_242506_n114759# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X726 dac_8bit_0/amux_2to1_7/B dac_8bit_0/amux_2to1_10/SELB vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X727 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 a_275374_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X728 vcp_sampled sample dac_8bit_0/c3m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X729 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X730 VDD dac_8bit_0/ibiasp dac_8bit_0/ibiasp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X731 dac_8bit_0/latched_comparator_folded_0/vtailp dac_8bit_0/vcom_buf dac_8bit_0/latched_comparator_folded_0/vlatchp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X732 VSS vcp a_238770_n132168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X733 input_amplifier_0/diff_fold_casc_ota_1/M6d input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X734 a_275374_n146348# sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X735 VSS VSS dac_8bit_1/amux_2to1_5/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X736 a_242867_n122433# a_242085_n122799# a_242783_n122433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X737 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X738 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X739 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X740 VSS a_241634_n115151# low_freq_pll_0/pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/Q_N VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X741 dac_8bit_1/amux_2to1_9/Y q0B vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X742 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X743 VSS peak_detector_0/ibiasn1 peak_detector_0/ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X744 VDD pulse_generator_0/sky130_fd_sc_hd__inv_1_0/Y a_338703_n185243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X745 input_amplifier_0/diff_fold_casc_ota_1/M13d input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/M6d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X746 biquad_gm_c_filter_0/gm_c_stage_0/vcmc VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X747 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X748 input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X749 VSS VSS input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X750 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X751 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X752 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X753 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X754 a_245151_n123343# a_244617_n123337# a_245056_n123343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X755 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 vcp_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X756 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X757 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X758 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X759 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X760 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_3/A a_243382_n121389# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X761 VDD VDD low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X762 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X763 VSS VSS dac_8bit_1/ibiasp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=2e+06u
X764 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X765 dac_8bit_0/latched_comparator_folded_0/vlatchp dac_8bit_0/latched_comparator_folded_0/vlatchm VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X766 vintm vfiltp biquad_gm_c_filter_0/gm_c_stage_2/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X767 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X768 a_226188_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_225730_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X769 VSS vpeak_sampled vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X770 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X771 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X772 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X773 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X774 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X775 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X776 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X777 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X778 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X779 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X780 input_amplifier_0/diff_fold_casc_ota_1/vcascnp input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X781 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X782 VSS a_336401_n185269# a_336408_n184969# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X783 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X784 dac_8bit_0/amux_2to1_4/B dac_8bit_0/amux_2to1_13/SELB vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X785 vcp_sampled sample dac_8bit_0/c6m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X786 dac_8bit_1/latched_comparator_folded_0/vtailp dac_8bit_1/vcom_buf dac_8bit_1/latched_comparator_folded_0/vlatchp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X787 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X788 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X789 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X790 a_242453_n120257# a_241919_n120623# a_242358_n120257# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X791 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X792 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X793 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X794 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X795 dac_8bit_0/amux_2to1_5/SELB sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X796 a_338285_n185243# a_338149_n185269# a_337864_n185269# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X797 vampp VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X798 VDD VDD vincm VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X799 VSS VSS vampp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X800 input_amplifier_0/diff_fold_casc_ota_1/vcascnp input_amplifier_0/diff_fold_casc_ota_1/vbias3 vampp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X801 VDD VDD input_amplifier_0/diff_fold_casc_ota_1/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X802 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X803 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X804 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/M2d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X805 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X806 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X807 a_224954_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X808 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X809 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X810 a_244783_n123337# a_244617_n123337# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X811 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X812 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X813 dac_8bit_1/vcom_buf dac_8bit_1/vcom_buf dac_8bit_1/vcom_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X814 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X815 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X816 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 vse VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X817 dac_8bit_0/amux_2to1_1/B dac_8bit_0/amux_2to1_16/SELB vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X818 VDD VDD peak_detector_0/vpeak VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X819 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X820 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X821 VSS dac_8bit_1/latched_comparator_folded_0/vcomppb dac_8bit_1/latched_comparator_folded_0/vcompp_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X822 a_236022_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/csinvn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X823 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X824 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X825 a_238312_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin a_237854_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X826 input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X827 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X828 input_amplifier_0/venp2 input_amplifier_0/vim2 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X829 sample_and_hold_1/vhold sample vpeak VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X830 dac_8bit_0/amux_2to1_2/SELB sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X831 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X832 dac_8bit_1/amux_2to1_12/SELB q2B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X833 a_335749_n185269# a_335844_n185269# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X834 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X835 VSS VSS vlowA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X836 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X837 a_236175_n122049# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X838 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp vse peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X839 low_freq_pll_0/pfd_cp_lpf_0/vQB a_239883_n115151# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X840 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X841 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X842 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X843 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X844 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X845 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X846 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 vocm input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X847 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X848 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X849 a_230446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X850 a_221023_n130007# low_freq_pll_0/cs_ring_osc_0/vosc low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X851 a_338532_n185787# a_338285_n185409# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X852 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X853 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X854 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X855 input_amplifier_0/diff_fold_casc_ota_0/vcascnp input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X856 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X857 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X858 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/vim1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X859 a_275374_n180872# sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X860 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X861 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X862 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X863 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X864 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q a_244617_n122799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X865 dac_8bit_1/amux_2to1_15/SELB q5B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X866 VSS VSS vlowA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X867 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X868 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X869 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn biquad_gm_c_filter_0/gm_c_stage_0/vcmcn VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X870 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X871 VDD VDD biquad_gm_c_filter_0/gm_c_stage_2/vcmcn VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X872 VDD a_242783_n122433# a_242951_n122531# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X873 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X874 a_243138_n114759# a_242419_n114983# a_242575_n114888# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X875 dac_8bit_0/amux_2to1_10/SELB q1A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X876 a_223312_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin a_222854_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X877 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X878 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X879 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X880 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X881 VDD vbiasp dac_8bit_0/ibiasn VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X882 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X883 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X884 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X885 dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X886 biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail2 vocm_filt biquad_gm_c_filter_0/gm_c_stage_3/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X887 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X888 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X889 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X890 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X891 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X892 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X893 biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail2 biquad_gm_c_filter_0/ibiasn3 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X894 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X895 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X896 VSS VSS biquad_gm_c_filter_0/ibiasn4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X897 VSS peak_detector_0/vpeak sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X898 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X899 a_224953_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X900 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X901 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X902 peak_detector_0/verr VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X903 VSS VSS vlowA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X904 a_242358_n120257# a_241919_n120623# a_242273_n120623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X905 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X906 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X907 comparator_0/vo1 comparator_0/vo1 comparator_0/vo1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X908 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X909 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X910 input_amplifier_0/diff_fold_casc_ota_1/M1d input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X911 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X912 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X913 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/diff_fold_casc_ota_1/vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X914 a_242273_n120623# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X915 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X916 a_162668_n147576# diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X917 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X918 dac_8bit_0/amux_2to1_13/SELB q3A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X919 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X920 a_338149_n185569# adc_clk VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X921 a_275374_n146348# sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X922 input_amplifier_0/diff_fold_casc_ota_1/vcascnp input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X923 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X924 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X925 VSS input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X926 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X927 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/M1d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X928 a_356329_n113250# dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X929 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X930 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X931 a_337864_n185269# a_338149_n185269# a_338084_n185243# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X932 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X933 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X934 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X935 vpeak_sampled sample dac_8bit_1/cdumm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X936 input_amplifier_0/diff_fold_casc_ota_0/vcascnp input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/vop1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X937 input_amplifier_0/vom1 input_amplifier_0/vip1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X938 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X939 a_226939_n130007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_226481_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X940 input_amplifier_0/venm1 input_amplifier_0/txgate_0/txb input_amplifier_0/vip2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X941 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X942 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X943 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X944 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X945 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X946 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_1/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X947 adc_vcaparrayA dac_8bit_0/c1m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X948 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X949 vpeak VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X950 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X951 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X952 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn biquad_gm_c_filter_0/gm_c_stage_1/vcmcn VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X953 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X954 VDD VDD biquad_gm_c_filter_0/gm_c_stage_3/vcmcn VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X955 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X956 dac_8bit_1/latched_comparator_folded_0/vcompp dac_8bit_1/latched_comparator_folded_0/vcompm VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X957 VSS VSS diff_to_se_converter_0/vip VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X958 dac_8bit_0/amux_2to1_16/SELB q6A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X959 VSS VSS dac_8bit_0/amux_2to1_2/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X960 input_amplifier_0/diff_fold_casc_ota_1/vfoldm VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X961 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X962 dac_8bit_0/amux_2to1_5/B q2A vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X963 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/vim2 input_amplifier_0/diff_fold_casc_ota_1/vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X964 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X965 a_238770_n150168# vcp a_238312_n150168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X966 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X967 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X968 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X969 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X970 biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail1 vocm_filt biquad_gm_c_filter_0/gm_c_stage_3/vcmcn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X971 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X972 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X973 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X974 dac_8bit_1/amux_2to1_6/B dac_8bit_1/amux_2to1_11/SELB vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X975 vpeak_sampled sample dac_8bit_1/c4m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X976 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X977 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_228770_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X978 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X979 vse diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X980 a_222040_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_222498_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X981 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X982 a_229954_n134960# vcp VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X983 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X984 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_245649_n122281# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X985 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X986 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/verr VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X987 a_225730_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X988 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X989 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X990 dac_8bit_1/amux_2to1_7/SELB sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X991 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X992 input_amplifier_0/vip2 input_amplifier_0/rst input_amplifier_0/vom1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X993 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X994 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X995 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X996 input_amplifier_0/venp2 input_amplifier_0/vim2 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X997 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X998 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X999 vlowA dac_8bit_0/amux_2to1_9/SELB dac_8bit_0/amux_2to1_9/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1000 dac_8bit_0/latched_comparator_folded_0/vlatchp dac_8bit_0/vcom_buf dac_8bit_0/latched_comparator_folded_0/vtailp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1001 VDD a_242783_n121345# a_242951_n121443# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1002 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1003 VDD vbiasp comparator_0/ibiasn VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X1004 dac_8bit_0/amux_2to1_2/B q5A vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1005 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1006 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1007 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1008 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1009 comparator_0/vcompp comparator_0/vcompm VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1010 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1011 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1012 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 a_163060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1013 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1014 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1015 a_238464_n119618# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout a_238006_n119618# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1016 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1017 dac_8bit_1/amux_2to1_3/B dac_8bit_1/amux_2to1_14/SELB vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1018 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X1019 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1020 a_237498_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_237956_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1021 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1022 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X1023 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1024 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1025 VSS a_245649_n121443# a_245607_n121711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1026 vrefA q1A dac_8bit_0/amux_2to1_7/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1027 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1028 dac_8bit_1/amux_2to1_4/SELB sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1029 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1030 biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail2 vintm biquad_gm_c_filter_0/gm_c_stage_1/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1031 VSS VSS vlowB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1032 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1033 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X1034 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 a_230446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1035 VSS biquad_gm_c_filter_0/ibiasn2 biquad_gm_c_filter_0/ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1036 vcp_sampled sample sample_and_hold_0/vholdm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1037 vlowA dac_8bit_0/amux_2to1_12/SELB dac_8bit_0/amux_2to1_5/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1038 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1039 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1040 vcp_sampled VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1041 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1042 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1043 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1044 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1045 a_245151_n122433# a_244617_n122799# a_245056_n122433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1046 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1047 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1048 input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vbias3 a_217060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1049 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X1050 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X1051 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1052 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1053 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1054 VSS input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1055 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 a_275374_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1056 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1057 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1058 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1059 vrefA q3A dac_8bit_0/amux_2to1_4/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1060 VDD vbiasp dac_8bit_1/ibiasn VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X1061 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1062 dac_8bit_1/amux_2to1_1/SELB sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1063 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1064 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1065 VSS VSS vlowB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1066 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1067 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1068 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1069 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1070 input_amplifier_0/vom1 input_amplifier_0/txgate_7/txb input_amplifier_0/vip2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1071 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1072 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn vintm biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1073 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1074 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1075 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1076 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1077 VSS VSS biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1078 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1079 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X1080 biquad_gm_c_filter_0/gm_c_stage_1/vtail_diff vintm vintm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1081 input_amplifier_0/vom1 VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X1082 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1083 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1084 dac_8bit_0/amux_2to1_7/B dac_8bit_0/amux_2to1_7/SELB dac_8bit_0/c1m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1085 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1086 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/vbias2 vampm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1087 input_amplifier_0/diff_fold_casc_ota_1/vcascnp input_amplifier_0/diff_fold_casc_ota_1/vbias3 vampp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1088 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X1089 dac_8bit_0/cdumm sample vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1090 biquad_gm_c_filter_0/ibiasn3 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X1091 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1092 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1093 dac_8bit_1/latched_comparator_folded_0/vlatchp adc_clk dac_8bit_1/latched_comparator_folded_0/vlatchm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X1094 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1095 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X1096 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1097 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1098 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1099 input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1100 vrefA q6A dac_8bit_0/amux_2to1_1/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1101 VSS biquad_gm_c_filter_0/gm_c_stage_0/vcmc biquad_gm_c_filter_0/gm_c_stage_0/vtail_diff VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1102 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/verr VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1103 vcp_sampled vcp_sampled vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1104 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1105 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1106 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1107 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1108 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1109 a_238007_n122049# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout a_237549_n122049# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1110 input_amplifier_0/venp1 input_amplifier_0/vop1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X1111 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1112 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1113 input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1114 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1115 dac_8bit_1/amux_2to1_11/SELB VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1116 VSS VSS dac_8bit_1/amux_2to1_7/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1117 VDD VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1118 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1119 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X1120 dac_8bit_0/amux_2to1_4/B dac_8bit_0/amux_2to1_4/SELB dac_8bit_0/c3m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1121 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1122 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X1123 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1124 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1125 dac_8bit_0/c4m sample vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1126 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X1127 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1128 sample_and_hold_1/vholdm sample vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1129 VDD a_239883_n115151# a_240447_n115125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1130 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1131 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1132 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1133 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1134 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1135 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1136 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1137 a_338532_n184877# a_338285_n185243# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1138 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn vse peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1139 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1140 adc_vcaparrayA dac_8bit_0/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1141 VDD VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1142 input_amplifier_0/diff_fold_casc_ota_0/M1d input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1143 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1144 VSS VSS vintp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1145 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1146 a_217060_n102324# input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1147 a_275374_n180872# sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1148 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/M6d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1149 dac_8bit_1/vcom_buf dac_8bit_1/vcom_buf dac_8bit_1/vcom_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1150 dac_8bit_1/amux_2to1_0/B VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1151 vcp_sampled VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1152 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1153 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_244617_n122249# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1154 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1155 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1156 a_337497_n185813# a_337592_n185460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1157 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1158 dac_8bit_1/amux_2to1_14/SELB q4B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1159 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1160 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1161 a_241480_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_241022_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1162 VSS VSS dac_8bit_1/amux_2to1_4/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1163 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1164 dac_8bit_0/amux_2to1_0/B dac_8bit_0/amux_2to1_17/SELB vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1165 a_243770_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_243312_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1166 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1167 dac_8bit_1/amux_2to1_7/B q1B vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1168 dac_8bit_0/amux_2to1_1/B dac_8bit_0/amux_2to1_1/SELB dac_8bit_0/c6m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1169 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 vocm input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X1170 biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail1 vintm biquad_gm_c_filter_0/gm_c_stage_0/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1171 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1172 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1173 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1174 input_amplifier_0/txgate_5/txb input_amplifier_0/rst VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1175 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1176 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1177 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1178 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1179 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1180 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 vocm input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X1181 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1182 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1183 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1184 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1185 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1186 adc_vcaparrayB VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1187 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1188 vampm input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1189 VDD low_freq_pll_0/pfd_cp_lpf_0/vpbias low_freq_pll_0/pfd_cp_lpf_0/vpbias VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1190 VDD vbiasp input_amplifier_0/ibiasn1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X1191 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1192 a_245224_n122281# a_245056_n122255# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1193 VSS VSS dac_8bit_1/amux_2to1_1/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1194 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1195 a_356329_n164260# dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1196 low_freq_pll_0/pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/Q_N a_240447_n115125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1197 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X1198 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1199 dac_8bit_1/amux_2to1_4/B q3B vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1200 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1201 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1202 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1203 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1204 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/verr VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1205 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1206 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1207 input_amplifier_0/diff_fold_casc_ota_1/vcascnp input_amplifier_0/diff_fold_casc_ota_1/vbias3 vampp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1208 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1209 a_275374_n180872# sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1210 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1211 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1212 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1213 dac_8bit_0/comp_outm adc_compA VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1214 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1215 input_amplifier_0/diff_fold_casc_ota_1/M1d input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1216 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1217 a_163060_n102324# input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1218 VDD a_242951_n123369# a_243382_n123343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1219 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1220 VSS a_242783_n123343# a_242951_n123369# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1221 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1222 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1223 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X1224 vcp_sampled vcp_sampled VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1225 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1226 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/vip2 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X1227 VDD VDD dac_8bit_1/latched_comparator_folded_0/vlatchp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1228 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1229 dac_8bit_0/latched_comparator_folded_0/vcompmb dac_8bit_0/latched_comparator_folded_0/vcompm VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1230 dac_8bit_1/amux_2to1_1/B q6B vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1231 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1232 a_226023_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1233 a_237956_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_238414_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1234 a_228313_n130007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_227855_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1235 input_amplifier_0/vop1 VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X1236 VSS VSS input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1237 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1238 a_356329_n113250# dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1239 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1240 pulse_generator_0/sky130_fd_sc_hd__inv_1_1/A pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1241 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1242 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1243 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1244 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1245 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1246 a_245056_n122255# a_244783_n122249# a_244971_n122255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1247 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1248 biquad_gm_c_filter_0/ibiasn4 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1249 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1250 a_245182_n121711# a_244783_n121711# a_245056_n121345# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1251 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1252 input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc vocm input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X1253 VDD VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1254 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1255 vrefB VSS dac_8bit_1/amux_2to1_6/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1256 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1257 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1258 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1259 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1260 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1261 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1262 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1263 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1264 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1265 input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1266 vcp sample sample_and_hold_0/vhold VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1267 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1268 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1269 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1270 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vfoldm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1271 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1272 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1273 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1274 a_231786_n134960# vcp a_231328_n134960# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1275 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1276 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1277 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1278 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1279 VSS VSS vlowA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1280 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1281 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1282 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1283 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1284 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.4e+07u
X1285 dac_8bit_1/c0m sample vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1286 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/vop1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1287 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1288 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X1289 low_freq_pll_0/pfd_cp_lpf_0/vswitchh low_freq_pll_0/pfd_cp_lpf_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1290 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn2 vocm_filt biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1291 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1292 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1293 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1294 dac_8bit_0/c0m dac_8bit_0/amux_2to1_8/SELB dac_8bit_0/amux_2to1_9/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1295 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/vim1 input_amplifier_0/diff_fold_casc_ota_0/vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X1296 input_amplifier_0/vip2 input_amplifier_0/vom1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X1297 VSS input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1298 vrefB q4B dac_8bit_1/amux_2to1_3/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1299 diff_to_se_converter_0/vim diff_to_se_converter_0/rst vfiltm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1300 a_275374_n146348# sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1301 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1302 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1303 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1304 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1305 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1306 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1307 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1308 VSS a_245649_n121193# a_245607_n120789# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1309 vincm VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1310 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1311 input_amplifier_0/ibiasn2 input_amplifier_0/ibiasn2 input_amplifier_0/ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1312 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1313 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X1314 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1315 dac_8bit_1/amux_2to1_6/B dac_8bit_1/amux_2to1_6/SELB dac_8bit_1/cdumm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1316 VDD vbiasp dac_8bit_1/ibiasn VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X1317 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1318 biquad_gm_c_filter_0/gm_c_stage_3/vtail_diff VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1319 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1320 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1321 VDD input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/M2d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1322 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1323 dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1324 a_221582_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1325 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1326 biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail2 vintm biquad_gm_c_filter_0/gm_c_stage_2/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1327 dac_8bit_1/latched_comparator_folded_0/vcompm dac_8bit_1/latched_comparator_folded_0/vcompp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1328 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1329 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1330 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1331 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1332 dac_8bit_1/amux_2to1_0/B sample dac_8bit_1/c7m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1333 a_240870_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_240412_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1334 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1335 input_amplifier_0/diff_fold_casc_ota_1/M2d input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1336 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1337 VSS biquad_gm_c_filter_0/ibiasn4 biquad_gm_c_filter_0/ibiasn4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1338 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1339 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 a_217060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1340 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q a_244617_n122799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1341 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1342 VSS peak_detector_0/verr sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X1343 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/csinvn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1344 vpeak_sampled sample dac_8bit_1/c2m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1345 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1346 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1347 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1348 VSS VSS low_freq_pll_0/pfd_cp_lpf_0/vpdiode VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1349 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X1350 dac_8bit_1/amux_2to1_3/B dac_8bit_1/amux_2to1_3/SELB dac_8bit_1/c4m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1351 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/vcom_buf VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1352 VSS a_337497_n185269# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_0/Q_N VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1353 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1354 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1355 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1356 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1357 input_amplifier_0/diff_fold_casc_ota_0/M1d input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1358 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1359 VSS input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1360 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1361 VDD vbiasp peak_detector_0/ibiasn1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X1362 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1363 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1364 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1365 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1366 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1367 VDD dac_8bit_1/latched_comparator_folded_0/vcompm dac_8bit_1/latched_comparator_folded_0/vcompp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1368 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1369 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1370 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1371 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1372 dac_8bit_1/amux_2to1_5/B dac_8bit_1/amux_2to1_12/SELB vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1373 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X1374 a_217060_n102324# input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1375 VSS vpeak sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X1376 vpeak_sampled sample dac_8bit_1/c5m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1377 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1378 low_freq_pll_0/cs_ring_osc_0/vpbias VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1379 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1380 dac_8bit_1/amux_2to1_0/B dac_8bit_1/amux_2to1_0/SELB dac_8bit_1/c7m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1381 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1382 dac_8bit_1/latched_comparator_folded_0/vlatchm dac_8bit_1/latched_comparator_folded_0/vlatchp VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1383 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1384 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X1385 low_freq_pll_0/pfd_cp_lpf_0/vQB a_239883_n115151# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1386 input_amplifier_0/diff_fold_casc_ota_1/vcascnp input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1387 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X1388 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1389 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vfoldp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1390 VSS VSS sample_and_hold_1/vholdm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1391 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1392 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X1393 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1394 vlowA dac_8bit_0/amux_2to1_10/SELB dac_8bit_0/amux_2to1_7/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1395 vampp VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X1396 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1397 dac_8bit_0/amux_2to1_6/B VSS vrefA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1398 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1399 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1400 input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vfoldp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1401 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1402 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1403 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1404 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1405 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1406 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1407 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1408 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 vpeak_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1409 input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X1410 dac_8bit_1/amux_2to1_2/B dac_8bit_1/amux_2to1_15/SELB vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1411 diff_to_se_converter_0/vip vocm_filt sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X1412 VSS input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1413 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1414 a_222396_n132168# vcp a_221938_n132168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1415 adc_compA dac_8bit_0/latched_comparator_folded_0/vcompm_buf VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1416 sample_and_hold_1/vholdm vpeak_sampled sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X1417 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1418 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1419 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1420 dac_8bit_0/latched_comparator_folded_0/vlatchm adc_clk dac_8bit_0/latched_comparator_folded_0/vcompm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1421 a_246786_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin a_246328_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1422 VSS low_freq_pll_0/ibiasn low_freq_pll_0/ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1423 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1424 input_amplifier_0/diff_fold_casc_ota_0/vcascnm input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1425 VSS VSS vlowB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1426 peak_detector_0/verr peak_detector_0/verr VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1427 a_242783_n123343# a_241919_n123337# a_242526_n123369# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1428 VDD input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X1429 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1430 biquad_gm_c_filter_0/ibiasn3 biquad_gm_c_filter_0/ibiasn3 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1431 VSS peak_detector_0/ibiasn2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1432 vlowA dac_8bit_0/amux_2to1_13/SELB dac_8bit_0/amux_2to1_4/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1433 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1434 input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1435 VSS vbiasn dac_8bit_1/ibiasp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=2e+06u
X1436 dac_8bit_0/latched_comparator_folded_0/vcompp dac_8bit_0/latched_comparator_folded_0/vcompm VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1437 VDD low_freq_pll_0/pfd_cp_lpf_0/vpbias low_freq_pll_0/pfd_cp_lpf_0/vswitchh VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1438 a_230446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1439 dac_8bit_0/amux_2to1_3/B q4A vrefA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1440 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1441 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1442 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/verr VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1443 a_242909_n122965# a_241919_n123337# a_242783_n123343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1444 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1445 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1446 biquad_gm_c_filter_0/gm_c_stage_0/vcmc VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1447 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1448 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1449 VSS input_amplifier_0/ibiasn1 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1450 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1451 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X1452 input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vbias3 a_217060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1453 dac_8bit_0/ibiasn dac_8bit_0/ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1454 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1455 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1456 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1457 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1458 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1459 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1460 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1461 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1462 VSS VSS biquad_gm_c_filter_0/gm_c_stage_1/vbiasp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1463 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1464 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1465 a_242855_n130007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_242397_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1466 VSS VSS vlowB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1467 VDD comparator_0/vcompp comparator_0/vo1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1468 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1469 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1470 vlowA dac_8bit_0/amux_2to1_16/SELB dac_8bit_0/amux_2to1_1/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1471 a_242273_n123343# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1472 VDD VDD peak_detector_0/verr VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1473 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1474 a_337864_n185555# a_338156_n185665# a_338107_n185787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1475 a_221938_n131500# low_freq_pll_0/cs_ring_osc_0/vosc a_221480_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1476 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X1477 VSS input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1478 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 a_356329_n113250# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1479 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1480 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1481 VDD low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_242701_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1482 dac_8bit_0/c7m sample dac_8bit_0/amux_2to1_0/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1483 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1484 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1485 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1486 vampp VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X1487 dac_8bit_0/c2m sample vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1488 VDD VDD vpeak_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1489 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X1490 vlowA sample adc_vcaparrayA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1491 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1492 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1493 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1494 vintp vintp biquad_gm_c_filter_0/gm_c_stage_1/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1495 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1496 adc_vcaparrayB dac_8bit_1/c3m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1497 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X1498 VDD input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X1499 VDD low_freq_pll_0/cs_ring_osc_0/vpbias a_236582_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1500 VSS VSS vlowB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1501 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1502 a_245870_n134960# vcp a_245412_n134960# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1503 VSS a_242951_n121443# a_243382_n121389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1504 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1505 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1506 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1507 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1508 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1509 diff_to_se_converter_0/vip vocm_filt sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X1510 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1511 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1512 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1513 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1514 dac_8bit_1/amux_2to1_12/SELB q2B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1515 biquad_gm_c_filter_0/gm_c_stage_1/vcmc VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1516 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X1517 input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vbias3 a_163060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1518 vampp vampp vampp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1519 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1520 a_246785_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin a_246327_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1521 vfiltp diff_to_se_converter_0/rst diff_to_se_converter_0/vip VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1522 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1523 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1524 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1525 VDD input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X1526 input_amplifier_0/diff_fold_casc_ota_0/vcascnp input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/vop1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1527 dac_8bit_0/c5m sample vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1528 a_245056_n121345# a_244783_n121711# a_244971_n121711# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1529 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1530 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X1531 biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail1 vocm_filt biquad_gm_c_filter_0/gm_c_stage_0/vcmcn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1532 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1533 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1534 peak_detector_0/ibiasn1 peak_detector_0/ibiasn1 peak_detector_0/ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1535 input_amplifier_0/vip1 input_amplifier_0/rst vincm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1536 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1537 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1538 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1539 vlowA q7A dac_8bit_0/amux_2to1_0/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1540 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1541 VDD input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X1542 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 a_356329_n113250# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1543 a_242397_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_241939_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1544 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X1545 VSS VSS low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/csinvn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1546 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1547 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X1548 biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail1 vintp biquad_gm_c_filter_0/gm_c_stage_1/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1549 VDD VDD dac_8bit_0/amux_2to1_9/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1550 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1551 vpeak_sampled VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1552 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1553 vampm VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X1554 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X1555 dac_8bit_1/amux_2to1_15/SELB q5B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1556 a_189446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1557 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1558 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1559 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1560 VSS a_245649_n123369# a_246080_n123343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1561 VSS input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1562 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1563 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/csinvn vcp a_232702_n134960# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1564 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/csinvp low_freq_pll_0/cs_ring_osc_0/vpbias a_243478_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1565 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1566 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1567 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1568 dac_8bit_1/amux_2to1_0/B q7B vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1569 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 a_189446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1570 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1571 VDD vbiasp vpeak_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X1572 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X1573 dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1574 input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vbias3 a_217060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1575 comparator_0/vcompm comparator_0/vcompp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1576 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1577 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1578 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1579 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1580 vse diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1581 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 a_162668_n147576# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1582 input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1583 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1584 VDD VDD dac_8bit_0/amux_2to1_5/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1585 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1586 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1587 input_amplifier_0/venp2 input_amplifier_0/vim2 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X1588 a_223414_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_222956_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1589 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1590 a_227396_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_226938_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1591 dac_8bit_1/amux_2to1_9/Y q0B vrefB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1592 VDD input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X1593 a_335844_n185269# a_336116_n185269# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1594 VSS VSS biquad_gm_c_filter_0/gm_c_stage_2/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1595 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1596 comparator_0/vtail comparator_0/vtail comparator_0/vtail VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1597 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1598 a_275374_n146348# sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1599 sample_and_hold_0/vhold sample vcp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1600 a_242702_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_242244_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1601 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1602 dac_8bit_0/amux_2to1_9/Y dac_8bit_0/amux_2to1_9/SELB vlowA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1603 VSS low_freq_pll_0/cs_ring_osc_0/vosc2 low_freq_pll_0/freq_div_0/vin VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1604 dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1605 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1606 sample_and_hold_0/vhold VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X1607 VDD input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X1608 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1609 adc_vcaparrayB dac_8bit_1/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1610 VDD VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1611 vse VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X1612 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1613 a_244783_n123337# a_244617_n123337# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1614 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/vcom_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1615 a_237956_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_237498_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1616 VDD a_242951_n121193# a_242867_n121167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1617 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1618 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1619 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X1620 VDD vbiasp diff_to_se_converter_0/ibiasn VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X1621 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1622 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1623 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1624 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X1625 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1626 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1627 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1628 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X1629 a_226646_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_227104_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1630 vcp_sampled VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X1631 biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail1 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1632 vlowB dac_8bit_1/amux_2to1_11/SELB dac_8bit_1/amux_2to1_6/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1633 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1634 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1635 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1636 a_236938_n132168# vcp a_236480_n132168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1637 VDD input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X1638 biquad_gm_c_filter_0/gm_c_stage_0/vbiasp biquad_gm_c_filter_0/ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1639 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1640 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1641 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1642 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1643 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn2 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1644 VSS vse sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X1645 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X1646 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1647 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1648 VSS VSS sample_and_hold_0/vhold VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1649 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1650 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1651 vampm VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X1652 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1653 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1654 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1655 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_10/A a_246080_n123343# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1656 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1657 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1658 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1659 a_239239_n115125# a_238793_n115125# a_239143_n115125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1660 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X1661 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1662 VDD VDD low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1663 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1664 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1665 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1666 vrefB q2B dac_8bit_1/amux_2to1_5/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1667 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1668 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X1669 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 a_356329_n164260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1670 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X1671 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1672 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 vse VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1673 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1674 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1675 vlowB dac_8bit_1/amux_2to1_14/SELB dac_8bit_1/amux_2to1_3/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1676 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1677 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1678 vpeak_sampled VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X1679 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1680 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1681 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1682 a_224330_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1683 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1684 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1685 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1686 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1687 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/vim2 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X1688 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 a_217060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1689 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1690 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1691 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1692 dac_8bit_1/c1m sample vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1693 VDD low_freq_pll_0/cs_ring_osc_0/vpbias a_225580_n122869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1694 VDD VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1695 a_356329_n164260# dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1696 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1697 VSS vcp a_223770_n132168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1698 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1699 VSS input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1700 low_freq_pll_0/pfd_cp_lpf_0/vswitchl low_freq_pll_0/pfd_cp_lpf_0/vQB vcp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1701 dac_8bit_0/c1m dac_8bit_0/amux_2to1_7/SELB dac_8bit_0/amux_2to1_7/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1702 VSS VSS sample_and_hold_1/vhold VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1703 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1704 vrefB q5B dac_8bit_1/amux_2to1_2/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1705 VSS a_242951_n123369# a_242909_n122965# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1706 dac_8bit_0/amux_2to1_6/B VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1707 VSS VSS low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/csinvn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1708 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1709 a_242701_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_242243_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1710 VSS VSS biquad_gm_c_filter_0/gm_c_stage_2/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1711 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1712 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1713 vlowB dac_8bit_1/amux_2to1_17/SELB dac_8bit_1/amux_2to1_0/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1714 VDD input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X1715 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1716 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1717 VDD VDD low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1718 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X1719 VSS low_freq_pll_0/pfd_cp_lpf_0/vRSTN a_242137_n115125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1720 biquad_gm_c_filter_0/ibiasn4 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X1721 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X1722 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1723 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1724 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 vse VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1725 a_236022_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/csinvn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1726 a_242783_n122433# a_241919_n122799# a_242526_n122687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1727 VSS biquad_gm_c_filter_0/ibiasn2 biquad_gm_c_filter_0/ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1728 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/csinvn low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin a_247702_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1729 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1730 a_245224_n122687# a_245056_n122433# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1731 VDD vbiasp biquad_gm_c_filter_0/ibiasn3 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X1732 dac_8bit_1/c3m sample vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1733 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1734 input_amplifier_0/diff_fold_casc_ota_0/vcascnp input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1735 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X1736 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1737 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1738 input_amplifier_0/vop1 VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X1739 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1740 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1741 dac_8bit_1/ibiasp vbiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=2e+06u
X1742 dac_8bit_0/c3m dac_8bit_0/amux_2to1_4/SELB dac_8bit_0/amux_2to1_4/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1743 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/M2d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1744 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1745 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1746 peak_detector_0/verr peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1747 VSS a_242526_n122687# a_242484_n122799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1748 input_amplifier_0/diff_fold_casc_ota_1/M1d input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1749 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1750 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1751 dac_8bit_0/amux_2to1_3/B VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1752 input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vbias3 a_217060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1753 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1754 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X1755 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1756 a_162668_n147576# diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1757 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/M1d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1758 VSS input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1759 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X1760 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1761 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X1762 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1763 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1764 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1765 dac_8bit_1/amux_2to1_2/B dac_8bit_1/amux_2to1_2/SELB dac_8bit_1/c5m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1766 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1767 biquad_gm_c_filter_0/gm_c_stage_2/vtail_diff vfiltm vintp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1768 a_242273_n122799# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1769 dac_8bit_1/c6m sample vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1770 a_337864_n185269# a_338156_n184969# a_338107_n184877# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1771 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1772 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1773 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1774 vlowA VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1775 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1776 dac_8bit_1/latched_comparator_folded_0/vlatchp dac_8bit_1/vcom_buf dac_8bit_1/latched_comparator_folded_0/vtailp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1777 dac_8bit_0/c6m dac_8bit_0/amux_2to1_1/SELB dac_8bit_0/amux_2to1_1/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1778 a_221022_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/csinvn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1779 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1780 a_335844_n185269# a_336116_n185269# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1781 a_223312_n131500# low_freq_pll_0/cs_ring_osc_0/vosc a_222854_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1782 VSS peak_detector_0/ibiasn2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1783 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1784 input_amplifier_0/diff_fold_casc_ota_1/vcascnm input_amplifier_0/diff_fold_casc_ota_1/vbias3 vampm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1785 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X1786 a_247702_n134960# vcp a_247244_n134960# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1787 VSS biquad_gm_c_filter_0/ibiasn3 biquad_gm_c_filter_0/ibiasn3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1788 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1789 a_356329_n113250# dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1790 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1791 input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1792 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1793 VSS a_242951_n121193# a_243382_n121167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1794 dac_8bit_1/latched_comparator_folded_0/vtailp vlowB dac_8bit_1/latched_comparator_folded_0/vlatchm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1795 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1796 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1797 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 a_356329_n113250# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1798 VDD VDD low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1799 a_275374_n180872# sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1800 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X1801 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1802 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X1803 adc_vcaparrayB dac_8bit_1/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1804 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1805 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1806 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1807 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1808 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1809 input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vbias3 a_163060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1810 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1811 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1812 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1813 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1814 dac_8bit_0/amux_2to1_5/B q2A vrefA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1815 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1816 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1817 diff_to_se_converter_0/txgate_1/txb diff_to_se_converter_0/rst VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1818 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1819 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1820 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X1821 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_243771_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1822 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1823 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1824 vpeak VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1825 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1826 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1827 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 input_amplifier_0/ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1828 vse diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1829 VSS a_338356_n185510# a_338285_n185409# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1830 input_amplifier_0/vop1 VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X1831 a_239817_n115125# a_238627_n115125# a_239708_n115125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1832 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1833 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1834 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X1835 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1836 VSS a_338149_n185269# a_338156_n184969# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1837 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1838 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1839 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1840 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1841 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.4e+07u
X1842 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/verr VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1843 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1844 input_amplifier_0/diff_fold_casc_ota_1/vcascnm input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1845 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1846 input_amplifier_0/diff_fold_casc_ota_0/vcascnp input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1847 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1848 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1849 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1850 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1851 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1852 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1853 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1854 dac_8bit_0/amux_2to1_2/B q5A vrefA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1855 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1856 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1857 dac_8bit_1/latched_comparator_folded_0/vlatchm adc_clk dac_8bit_1/latched_comparator_folded_0/vlatchp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X1858 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1859 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1860 a_236480_n150168# vcp a_236022_n150168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1861 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1862 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vfoldp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1863 VDD a_241731_n115151# low_freq_pll_0/pfd_cp_lpf_0/vQA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1864 a_242562_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_243020_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1865 VDD VDD input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1866 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1867 a_226938_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_226480_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1868 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1869 input_amplifier_0/vom1 input_amplifier_0/rst input_amplifier_0/vip2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1870 a_189446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1871 peak_detector_0/verr VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X1872 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_228770_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1873 input_amplifier_0/diff_fold_casc_ota_0/vcascnm input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1874 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X1875 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1876 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1877 VSS VSS adc_vcaparrayA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1878 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1879 VDD vbiasp input_amplifier_0/ibiasn2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X1880 VSS biquad_gm_c_filter_0/gm_c_stage_2/vcmc biquad_gm_c_filter_0/gm_c_stage_2/vcmc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1881 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X1882 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1883 VSS low_freq_pll_0/freq_div_0/vout a_238627_n115125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1884 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1885 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1886 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1887 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1888 vse diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1889 input_amplifier_0/vom1 VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X1890 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1891 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1892 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1893 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1894 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1895 VDD VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1896 a_242575_n114888# a_242419_n114983# a_242720_n114759# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1897 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/csinvp low_freq_pll_0/cs_ring_osc_0/vpbias a_239330_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1898 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1899 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1900 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1901 dac_8bit_1/amux_2to1_9/Y VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1902 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1903 VDD VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1904 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1905 comparator_0/vo1 comparator_0/vcompp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1906 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1907 VDD a_242951_n120355# a_242867_n120257# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1908 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1909 a_242909_n122799# a_241919_n122799# a_242783_n122433# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1910 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1911 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1912 VDD VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1913 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1914 input_amplifier_0/diff_fold_casc_ota_1/vcascnp input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1915 vpeak VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X1916 input_amplifier_0/vim2 input_amplifier_0/vop1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X1917 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/vcom_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1918 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1919 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1920 a_239330_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_238872_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1921 a_223770_n150168# vcp a_223312_n150168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1922 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1923 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.4e+07u
X1924 input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1925 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1926 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X1927 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1928 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1929 diff_to_se_converter_0/txgate_1/txb diff_to_se_converter_0/rst VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1930 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1931 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1932 vpeak vpeak vpeak VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1933 VSS input_amplifier_0/ibiasn1 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1934 a_242526_n122281# a_242358_n122255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1935 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1936 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/diff_fold_casc_ota_0/vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X1937 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1938 a_242085_n123337# a_241919_n123337# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1939 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1940 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1941 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X1942 dac_8bit_1/cdumm dac_8bit_1/amux_2to1_6/SELB dac_8bit_1/amux_2to1_6/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1943 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1944 a_238312_n132168# vcp a_237854_n132168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1945 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X1946 dac_8bit_1/vcom_buf VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X1947 a_242526_n121599# a_242358_n121345# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1948 a_241731_n115151# a_242102_n114873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1949 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1950 a_242783_n122255# a_242085_n122249# a_242526_n122281# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1951 biquad_gm_c_filter_0/ibiasn4 biquad_gm_c_filter_0/ibiasn4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1952 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1953 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1954 VDD dac_8bit_1/latched_comparator_folded_0/vcompp dac_8bit_1/latched_comparator_folded_0/vcompm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1955 diff_to_se_converter_0/vip diff_to_se_converter_0/rst vfiltp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1956 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1957 VSS vcp a_230160_n119618# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1958 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1959 a_238771_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_238313_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1960 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1961 a_222498_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_222956_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1962 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1963 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1964 VDD a_245481_n122255# a_245649_n122281# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1965 vrefB dac_8bit_1/amux_2to1_17/SELB dac_8bit_1/amux_2to1_0/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1966 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1967 a_242526_n120511# a_242358_n120257# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1968 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1969 VDD VDD dac_8bit_0/amux_2to1_7/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1970 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1971 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1972 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn1 vocm_filt biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1973 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1974 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1975 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1976 dac_8bit_1/c4m dac_8bit_1/amux_2to1_3/SELB dac_8bit_1/amux_2to1_3/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1977 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X1978 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1979 input_amplifier_0/vop1 input_amplifier_0/vim1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X1980 a_245565_n122255# a_244783_n122249# a_245481_n122255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1981 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1982 VDD VDD dac_8bit_0/vcom_buf VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1983 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1984 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1985 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1986 input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1987 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1988 input_amplifier_0/vom1 VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X1989 dac_8bit_0/amux_2to1_17/SELB q7A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1990 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1991 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/vcom_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1992 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1993 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1994 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1995 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X1996 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1997 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1998 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/vim2 input_amplifier_0/diff_fold_casc_ota_1/vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X1999 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2000 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2001 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2002 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vfoldm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2003 peak_detector_0/verr peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2004 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2005 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2006 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2007 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2008 a_241634_n115151# a_241731_n115151# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2009 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2010 VDD VDD dac_8bit_0/amux_2to1_4/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2011 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2012 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2013 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2014 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2015 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2016 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2017 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2018 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X2019 low_freq_pll_0/pfd_cp_lpf_0/vswitchh low_freq_pll_0/pfd_cp_lpf_0/vQAb vcp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2020 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2021 dac_8bit_1/amux_2to1_7/B q1B vrefB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2022 peak_detector_0/vpeak VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2023 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2024 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2025 input_amplifier_0/vip2 input_amplifier_0/txgate_7/txb input_amplifier_0/vom1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2026 vampm vampm vampm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2027 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/vim1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X2028 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2029 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2030 dac_8bit_0/amux_2to1_7/B dac_8bit_0/amux_2to1_10/SELB vlowA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2031 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2032 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2033 a_336608_n185510# a_336408_n185665# a_336757_n185421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2034 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2035 vlowA VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2036 VSS a_242526_n122281# a_242484_n121877# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2037 sample_and_hold_0/vholdm VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2038 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X2039 comparator_0/vtail vfiltm comparator_0/vcompp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2040 vampm gain_ctrl_1 input_amplifier_0/venm2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2041 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2042 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2043 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2044 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2045 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2046 VDD VDD dac_8bit_0/amux_2to1_1/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2047 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2048 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2049 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2050 dac_8bit_1/amux_2to1_4/B q3B vrefB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2051 a_162668_n147576# diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2052 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X2053 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2054 a_241480_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_241022_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2055 input_amplifier_0/diff_fold_casc_ota_1/M2d input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2056 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X2057 low_freq_pll_0/pfd_cp_lpf_0/vswitchh low_freq_pll_0/pfd_cp_lpf_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2058 a_226328_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_225870_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2059 vpeak_sampled sample sample_and_hold_1/vholdm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2060 dac_8bit_0/amux_2to1_4/B dac_8bit_0/amux_2to1_13/SELB vlowA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2061 vampm VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X2062 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2063 vlowA VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2064 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2065 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X2066 VDD VDD vintp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2067 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2068 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2069 vintp biquad_gm_c_filter_0/gm_c_stage_2/vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2070 VSS vcp_sampled sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X2071 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2072 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2073 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2074 input_amplifier_0/diff_fold_casc_ota_0/vcascnm input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/vom1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2075 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2076 comparator_0/vmirror comparator_0/vmirror comparator_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2077 a_230446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2078 vintm VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2079 vampp input_amplifier_0/vim2 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X2080 VSS peak_detector_0/ibiasn2 peak_detector_0/ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2081 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2082 low_freq_pll_0/cs_ring_osc_0/vpbias low_freq_pll_0/cs_ring_osc_0/vpbias a_228328_n122869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X2083 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2084 vlowB dac_8bit_1/amux_2to1_15/SELB dac_8bit_1/amux_2to1_2/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2085 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2086 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2087 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X2088 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2089 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2090 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2091 dac_8bit_1/amux_2to1_1/B q6B vrefB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2092 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2093 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2094 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2095 vse vse vse VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2096 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2097 a_229954_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2098 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2099 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2100 dac_8bit_0/amux_2to1_1/B dac_8bit_0/amux_2to1_16/SELB vlowA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2101 vampp input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vfoldp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2102 comparator_0/ibiasn comparator_0/ibiasn comparator_0/ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2103 adc_vcaparrayB dac_8bit_1/c3m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2104 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2105 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q a_242951_n122281# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2106 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2107 input_amplifier_0/diff_fold_casc_ota_0/M1d input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2108 a_356329_n113250# dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2109 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X2110 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/vop1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2111 input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2112 VSS vpeak_sampled sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X2113 VDD VDD vampm VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2114 dac_8bit_0/amux_2to1_5/B VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2115 a_189446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2116 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2117 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2118 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2119 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2120 VSS VSS low_freq_pll_0/pfd_cp_lpf_0/vswitchl VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2121 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2122 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2123 vpeak_sampled VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2124 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2125 vse diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2126 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2127 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2128 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2129 dac_8bit_0/c0m dac_8bit_0/amux_2to1_8/SELB vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2130 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2131 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2132 a_226023_n130007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X2133 biquad_gm_c_filter_0/ibiasn3 biquad_gm_c_filter_0/ibiasn3 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2134 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2135 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2136 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 vpeak VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2137 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2138 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X2139 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X2140 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X2141 VDD VDD vintm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2142 vfiltp biquad_gm_c_filter_0/gm_c_stage_3/vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2143 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2144 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2145 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 vpeak VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2146 a_338703_n185409# a_338149_n185569# a_338356_n185510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2147 diff_to_se_converter_0/vip vfiltp sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X2148 dac_8bit_0/amux_2to1_2/B VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2149 a_226327_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_225869_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X2150 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2151 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2152 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2153 a_189446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2154 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2155 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2156 a_242085_n120623# a_241919_n120623# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2157 dac_8bit_0/amux_2to1_6/B sample dac_8bit_0/cdumm VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2158 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2159 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2160 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2161 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2162 input_amplifier_0/venm2 gain_ctrl_1 vampm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2163 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2164 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_6/A a_246080_n121167# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2165 a_228312_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_227854_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2166 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2167 input_amplifier_0/diff_fold_casc_ota_0/vcascnm input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2168 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2169 a_222956_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_223414_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X2170 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2171 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2172 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2173 input_amplifier_0/diff_fold_casc_ota_1/M1d input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2174 a_217060_n102324# input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2175 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2176 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2177 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X2178 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2179 input_amplifier_0/diff_fold_casc_ota_0/M1d input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2180 a_229953_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X2181 a_244971_n121711# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2182 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2183 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2184 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2185 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2186 vrefB VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2187 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2188 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2189 VDD VDD dac_8bit_1/amux_2to1_6/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2190 VDD VDD vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2191 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2192 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2193 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2194 vse diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2195 VDD comparator_0/vcompm comparator_0/vcompm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2196 dac_8bit_0/amux_2to1_3/B sample dac_8bit_0/c4m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2197 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2198 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2199 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2200 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2201 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2202 VSS dac_8bit_1/latched_comparator_folded_0/vcompp_buf a_383508_n152139# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2203 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2204 dac_8bit_0/latched_comparator_folded_0/vlatchm VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X2205 a_238414_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_238872_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X2206 adc_vcaparrayB dac_8bit_1/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2207 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2208 vampp VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X2209 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2210 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 a_275374_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2211 VDD VDD diff_to_se_converter_0/vim VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2212 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2213 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2214 vlowB VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2215 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2216 VSS low_freq_pll_0/ibiasn low_freq_pll_0/ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2217 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2218 input_amplifier_0/diff_fold_casc_ota_1/vfoldp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2219 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2220 a_189446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2221 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2222 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2223 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2224 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2225 VDD VDD input_amplifier_0/diff_fold_casc_ota_1/vfoldp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2226 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn1 vocm_filt biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2227 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2228 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 a_163060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2229 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2230 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2231 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2232 VSS vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2233 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2234 VDD VDD dac_8bit_1/amux_2to1_3/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2235 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2236 a_227104_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_226646_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X2237 VDD VDD vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2238 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2239 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2240 dac_8bit_0/amux_2to1_0/B sample dac_8bit_0/c7m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2241 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2242 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2243 VDD VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2244 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2245 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2246 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X2247 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2248 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2249 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X2250 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2251 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2252 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2253 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2254 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2255 dac_8bit_1/amux_2to1_6/B dac_8bit_1/amux_2to1_11/SELB vlowB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2256 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2257 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2258 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2259 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2260 a_162668_n147576# diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2261 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2262 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2263 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2264 diff_to_se_converter_0/vip vfiltp sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X2265 VSS VSS low_freq_pll_0/cs_ring_osc_0/vosc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2266 a_245565_n121345# a_244783_n121711# a_245481_n121345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2267 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2268 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2269 sample_and_hold_0/vhold VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2270 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2271 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2272 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2273 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2274 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2275 low_freq_pll_0/pfd_cp_lpf_0/vswitchh low_freq_pll_0/pfd_cp_lpf_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2276 VDD VDD dac_8bit_1/amux_2to1_0/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2277 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2278 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2279 VDD VDD vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2280 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2281 VSS VSS biquad_gm_c_filter_0/ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2282 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2283 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2284 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2285 low_freq_pll_0/cs_ring_osc_0/vosc low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout a_238922_n119618# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2286 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn vintp biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2287 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2288 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2289 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2290 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2291 VDD VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2292 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2293 dac_8bit_1/amux_2to1_3/B dac_8bit_1/amux_2to1_14/SELB vlowB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2294 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X2295 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X2296 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2297 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2298 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 input_amplifier_0/ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2299 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2300 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/vcom_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2301 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2302 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2303 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2304 input_amplifier_0/diff_fold_casc_ota_1/M1d input_amplifier_0/diff_fold_casc_ota_1/M1d input_amplifier_0/diff_fold_casc_ota_1/M1d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2305 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 a_356329_n113250# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2306 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2307 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2308 dac_8bit_1/amux_2to1_7/B VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2309 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2310 VSS peak_detector_0/verr sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X2311 VSS input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2312 low_freq_pll_0/pfd_cp_lpf_0/vpbias low_freq_pll_0/pfd_cp_lpf_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2313 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X2314 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2315 VDD a_242526_n122281# a_242453_n122255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2316 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2317 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2318 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2319 input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc vocm input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X2320 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2321 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2322 VSS dac_8bit_0/latched_comparator_folded_0/vlatchm dac_8bit_0/latched_comparator_folded_0/vlatchp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2323 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/vim1 input_amplifier_0/diff_fold_casc_ota_0/vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X2324 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2325 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2326 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2327 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2328 biquad_gm_c_filter_0/ibiasn2 biquad_gm_c_filter_0/ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2329 input_amplifier_0/vim2 input_amplifier_0/vop1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X2330 dac_8bit_1/c7m dac_8bit_1/amux_2to1_0/SELB vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2331 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2332 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2333 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2334 a_230446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2335 input_amplifier_0/diff_fold_casc_ota_1/vcascnm input_amplifier_0/diff_fold_casc_ota_1/vbias3 vampm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2336 dac_8bit_0/vcom_buf dac_8bit_0/vcom_buf dac_8bit_0/vcom_buf VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2337 vintp vampp biquad_gm_c_filter_0/gm_c_stage_0/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2338 biquad_gm_c_filter_0/gm_c_stage_2/vtail_diff vfiltp vintm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2339 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X2340 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2341 dac_8bit_1/c2m dac_8bit_1/amux_2to1_5/SELB dac_8bit_1/amux_2to1_5/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2342 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2343 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2344 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2345 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2346 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X2347 a_336116_n185269# a_336401_n185269# a_336336_n185243# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2348 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2349 dac_8bit_1/amux_2to1_4/B VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2350 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2351 diff_to_se_converter_0/ibiasn vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X2352 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2353 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2354 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2355 VSS vpeak sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X2356 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/diff_fold_casc_ota_1/vbias2 vampp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2357 dac_8bit_1/latched_comparator_folded_0/vlatchm VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2358 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 a_275374_n146348# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2359 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2360 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2361 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2362 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2363 a_242358_n122255# a_241919_n122249# a_242273_n122255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2364 low_freq_pll_0/freq_div_0/vout a_245649_n121193# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2365 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2366 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X2367 vpeak sample sample_and_hold_1/vhold VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2368 dac_8bit_1/amux_2to1_9/Y sample dac_8bit_1/c0m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2369 vcp_sampled dac_8bit_0/amux_2to1_8/SELB dac_8bit_0/c0m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2370 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2371 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2372 VSS peak_detector_0/vpeak sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X2373 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2374 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2375 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 a_189446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2376 dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2377 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X2378 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X2379 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2380 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2381 biquad_gm_c_filter_0/ibiasn2 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X2382 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X2383 peak_detector_0/ibiasn1 peak_detector_0/ibiasn1 peak_detector_0/ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2384 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2385 a_227412_n122869# low_freq_pll_0/cs_ring_osc_0/vpbias a_227870_n122869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X2386 VSS dac_8bit_1/vcom_buf sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X2387 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2388 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2389 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2390 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2391 dac_8bit_1/c5m dac_8bit_1/amux_2to1_2/SELB dac_8bit_1/amux_2to1_2/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2392 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2393 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2394 dac_8bit_1/amux_2to1_1/B VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2395 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2396 a_231786_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin a_231328_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2397 input_amplifier_0/vop1 input_amplifier_0/vim1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X2398 a_240869_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_240411_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X2399 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2400 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X2401 input_amplifier_0/vom1 VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X2402 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2403 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2404 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2405 VDD VDD vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2406 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2407 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2408 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2409 a_163060_n102324# input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2410 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2411 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc vampp input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X2412 dac_8bit_1/amux_2to1_5/B sample dac_8bit_1/c2m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2413 dac_8bit_1/latched_comparator_folded_0/vlatchm adc_clk dac_8bit_1/latched_comparator_folded_0/vlatchp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X2414 sample_and_hold_1/vholdm sample vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2415 vcp_sampled dac_8bit_0/amux_2to1_5/SELB dac_8bit_0/c2m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2416 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2417 dac_8bit_0/vcom_buf VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X2418 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2419 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_242951_n120355# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2420 input_amplifier_0/vim1 input_amplifier_0/txgate_4/txb vincm VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2421 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2422 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2423 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2424 adc_vcaparrayB dac_8bit_1/cdumm sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2425 a_242854_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_242396_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2426 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2427 a_189446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2428 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2429 a_162668_n147576# diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2430 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2431 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vfoldp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2432 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X2433 VDD a_336608_n185269# a_336537_n185243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X2434 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/vip2 input_amplifier_0/diff_fold_casc_ota_1/vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X2435 VDD VDD dac_8bit_0/latched_comparator_folded_0/vlatchm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2436 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2437 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2438 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2439 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2440 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2441 dac_8bit_1/latched_comparator_folded_0/vcompm_buf dac_8bit_1/latched_comparator_folded_0/vcompmb VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2442 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X2443 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2444 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2445 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2446 VDD VDD low_freq_pll_0/pfd_cp_lpf_0/vswitchh VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2447 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2448 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2449 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2450 VDD VDD vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2451 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2452 VSS a_337497_n185813# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/D VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2453 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2454 comparator_0/vcompm comparator_0/vcompm VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2455 vlowA VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2456 VSS VSS sample_and_hold_1/vholdm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2457 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2458 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2459 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2460 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2461 input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X2462 dac_8bit_0/vcom_buf dac_8bit_0/vcom_buf dac_8bit_0/vcom_buf VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2463 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2464 input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2465 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2466 VSS a_241731_n115151# low_freq_pll_0/pfd_cp_lpf_0/vQA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2467 a_242397_n130007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_241939_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X2468 VDD VDD vintm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2469 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2470 a_242484_n120789# a_242085_n121161# a_242358_n121167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2471 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2472 VSS input_amplifier_0/diff_fold_casc_ota_1/M13d input_amplifier_0/diff_fold_casc_ota_1/M13d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2473 vcp_sampled VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X2474 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2475 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2476 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2477 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2478 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2479 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X2480 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn vse peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2481 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2482 VDD a_241634_n115151# low_freq_pll_0/pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2483 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2484 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2485 vse diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2486 a_230870_n134960# vcp a_230412_n134960# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2487 a_241646_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_241188_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X2488 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2489 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X2490 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2491 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2492 a_275374_n146348# sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2493 vlowA VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2494 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2495 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2496 a_244971_n121167# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2497 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2498 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2499 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2500 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2501 a_231785_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin a_231327_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X2502 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2503 input_amplifier_0/vop1 VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X2504 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2505 a_236582_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_237040_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X2506 a_336401_n185569# adc_clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2507 adc_vcaparrayB sample vlowB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2508 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2509 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2510 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2511 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X2512 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2513 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2514 adc_vcaparrayA sample vlowA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2515 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2516 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2517 vcp_sampled sample dac_8bit_0/c7m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2518 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2519 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2520 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2521 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2522 dac_8bit_0/latched_comparator_folded_0/vlatchm VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2523 a_240412_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_239954_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2524 input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X2525 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 a_275374_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2526 a_356329_n164260# dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2527 vampp input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2528 a_336757_n185243# a_336537_n185243# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2529 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2530 input_amplifier_0/vim2 input_amplifier_0/vop1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X2531 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2532 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2533 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2534 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2535 VDD VDD vintp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2536 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_5/A a_243382_n123343# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2537 dac_8bit_0/amux_2to1_6/SELB sample VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2538 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2539 a_163060_n102324# input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2540 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2541 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2542 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X2543 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2544 diff_to_se_converter_0/vip diff_to_se_converter_0/rst vfiltp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2545 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2546 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2547 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2548 VSS dac_8bit_1/latched_comparator_folded_0/vlatchp dac_8bit_1/latched_comparator_folded_0/vlatchm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X2549 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2550 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2551 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q a_241919_n121711# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2552 VSS biquad_gm_c_filter_0/ibiasn1 biquad_gm_c_filter_0/ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2553 vincm input_amplifier_0/txgate_4/txb input_amplifier_0/vim1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2554 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X2555 VDD dac_8bit_1/latched_comparator_folded_0/vcomppb dac_8bit_1/latched_comparator_folded_0/vcompp_buf VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2556 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2557 dac_8bit_0/c1m dac_8bit_0/amux_2to1_7/SELB vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2558 dac_8bit_0/amux_2to1_0/B dac_8bit_0/amux_2to1_17/SELB vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2559 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q a_241919_n121711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2560 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X2561 adc_vcaparrayA dac_8bit_0/c2m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2562 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2563 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2564 input_amplifier_0/vop1 VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X2565 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X2566 VSS vcp_sampled vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2567 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 a_230446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2568 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2569 input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X2570 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2571 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/vom1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2572 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2573 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2574 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2575 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X2576 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2577 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2578 dac_8bit_0/amux_2to1_3/SELB sample VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2579 a_338285_n185409# a_338156_n185665# a_337864_n185555# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2580 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2581 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2582 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 a_217060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2583 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2584 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2585 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X2586 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 a_275374_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2587 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2588 input_amplifier_0/vim2 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2589 a_189446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2590 input_amplifier_0/diff_fold_casc_ota_1/M1d input_amplifier_0/diff_fold_casc_ota_1/M1d input_amplifier_0/diff_fold_casc_ota_1/M1d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2591 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2592 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2593 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2594 vincm input_amplifier_0/rst input_amplifier_0/vip1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2595 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2596 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2597 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2598 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_10/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2599 dac_8bit_0/c3m dac_8bit_0/amux_2to1_4/SELB vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2600 a_222956_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_222498_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X2601 VDD comparator_0/vcompp comparator_0/vcompp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2602 VSS a_335844_n185269# pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2603 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2604 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/M1d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2605 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2606 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2607 diff_to_se_converter_0/vip vfiltp sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X2608 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2609 dac_8bit_1/latched_comparator_folded_0/vlatchp adc_clk dac_8bit_1/latched_comparator_folded_0/vlatchm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X2610 a_242244_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_241786_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2611 low_freq_pll_0/freq_div_0/vin low_freq_pll_0/cs_ring_osc_0/vosc2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2612 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2613 dac_8bit_0/latched_comparator_folded_0/vlatchp dac_8bit_0/vcom_buf dac_8bit_0/latched_comparator_folded_0/vtailp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2614 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2615 VSS VSS low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2616 a_221938_n132168# vcp a_221480_n132168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2617 biquad_gm_c_filter_0/ibiasn2 biquad_gm_c_filter_0/ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2618 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2619 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2620 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2621 VDD a_242526_n121599# a_242453_n121345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2622 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2623 VDD VDD vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2624 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn vintp biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2625 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X2626 a_240411_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_239953_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X2627 a_337497_n185269# a_337592_n185269# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2628 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2629 input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X2630 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 a_275374_n146348# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2631 VDD a_242951_n122531# a_243382_n122477# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2632 dac_8bit_0/amux_2to1_2/B sample dac_8bit_0/c5m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2633 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2634 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2635 dac_8bit_0/c6m dac_8bit_0/amux_2to1_1/SELB vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2636 input_amplifier_0/diff_fold_casc_ota_1/vcascnm input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2637 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2638 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2639 VDD VDD low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X2640 a_162668_n147576# diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2641 input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X2642 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2643 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2644 VSS input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2645 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X2646 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2647 a_245870_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin a_245412_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2648 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2649 adc_vcaparrayB dac_8bit_1/c2m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2650 vlowB VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2651 dac_8bit_0/latched_comparator_folded_0/vtailp dac_8bit_0/latched_comparator_folded_0/vtailp dac_8bit_0/latched_comparator_folded_0/vtailp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2652 dac_8bit_0/ibiasn vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X2653 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2654 VDD a_242419_n114983# a_242380_n114857# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2655 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2656 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2657 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2658 vampp gain_ctrl_1 input_amplifier_0/venp2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2659 a_228328_n119618# vcp a_227870_n119618# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2660 a_338356_n185269# a_338156_n184969# a_338505_n185243# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2661 VDD VDD vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2662 VDD VDD dac_8bit_1/amux_2to1_2/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2663 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X2664 sample_and_hold_0/vhold sample vcp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2665 VDD VDD vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2666 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2667 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2668 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2669 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2670 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2671 vse vse vse VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2672 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2673 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2674 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2675 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X2676 adc_vcaparrayA dac_8bit_0/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2677 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2678 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2679 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2680 a_337592_n185269# a_337864_n185269# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2681 VSS VSS low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/csinvn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2682 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X2683 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2684 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2685 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn2 vocm_filt biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2686 dac_8bit_1/amux_2to1_5/B dac_8bit_1/amux_2to1_12/SELB vlowB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2687 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2688 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2689 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2690 dac_8bit_1/vcom_buf dac_8bit_1/vcom_buf dac_8bit_1/vcom_buf VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2691 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2692 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2693 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2694 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 a_275374_n146348# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2695 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2696 vlowB VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2697 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2698 a_225580_n122869# low_freq_pll_0/cs_ring_osc_0/vpbias a_226038_n122869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X2699 input_amplifier_0/diff_fold_casc_ota_0/vcascnm input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/vom1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2700 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2701 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X2702 a_217060_n102324# input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2703 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2704 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2705 a_221022_n131500# low_freq_pll_0/cs_ring_osc_0/vosc low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/csinvn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2706 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2707 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2708 dac_8bit_0/amux_2to1_17/SELB q7A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2709 a_335844_n185460# a_336116_n185555# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2710 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2711 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2712 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2713 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/csinvn low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin a_232702_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2714 a_242243_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_241785_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X2715 a_245412_n134960# vcp a_244954_n134960# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2716 input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2717 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2718 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2719 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2720 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2721 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2722 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X2723 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2724 vcp VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2725 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2726 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2727 dac_8bit_1/amux_2to1_2/B dac_8bit_1/amux_2to1_15/SELB vlowB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2728 sample_and_hold_1/vhold sample vpeak VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2729 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2730 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2731 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2732 a_245182_n122965# a_244783_n123337# a_245056_n123343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2733 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2734 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X2735 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.4e+07u
X2736 vlowB VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2737 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2738 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 a_356329_n164260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2739 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2740 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vfoldp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2741 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2742 VDD VDD vampp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2743 vintm vampm biquad_gm_c_filter_0/gm_c_stage_0/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2744 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2745 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/vim2 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X2746 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2747 dac_8bit_1/amux_2to1_8/SELB sample VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2748 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2749 a_241939_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_241481_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X2750 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2751 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_243771_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X2752 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2753 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2754 vampp vampp vampp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2755 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2756 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2757 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2758 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2759 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2760 VDD a_245649_n122281# a_246080_n122255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2761 vpeak_sampled vpeak_sampled VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2762 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2763 vintm vintm biquad_gm_c_filter_0/gm_c_stage_1/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2764 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2765 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X2766 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2767 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2768 VSS VSS sample_and_hold_1/vhold VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2769 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2770 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 vcp_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2771 vcp_sampled dac_8bit_0/amux_2to1_6/SELB dac_8bit_0/cdumm VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2772 a_242085_n123337# a_241919_n123337# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2773 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2774 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q a_244617_n123337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2775 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2776 input_amplifier_0/vim2 input_amplifier_0/vop1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X2777 a_232702_n134960# vcp a_232244_n134960# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2778 a_163060_n102324# input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2779 input_amplifier_0/diff_fold_casc_ota_0/M6d input_amplifier_0/diff_fold_casc_ota_0/M6d input_amplifier_0/diff_fold_casc_ota_0/M6d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2780 VDD VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2781 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2782 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2783 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X2784 VSS biquad_gm_c_filter_0/ibiasn3 biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2785 dac_8bit_0/amux_2to1_9/Y VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2786 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2787 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X2788 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2789 dac_8bit_0/latched_comparator_folded_0/vlatchm adc_clk dac_8bit_0/latched_comparator_folded_0/vlatchp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X2790 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2791 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2792 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2793 input_amplifier_0/diff_fold_casc_ota_0/M13d input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/M6d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2794 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2795 VDD a_335844_n185269# pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2796 VDD VDD low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X2797 vincm VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2798 dac_8bit_1/vcom_buf VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X2799 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2800 dac_8bit_0/latched_comparator_folded_0/vtailp dac_8bit_0/vcom_buf dac_8bit_0/latched_comparator_folded_0/vlatchp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2801 a_247244_n134960# vcp a_246786_n134960# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2802 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X2803 dac_8bit_0/ibiasp dac_8bit_0/ibiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2804 a_243020_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_242562_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X2805 dac_8bit_1/amux_2to1_7/B sample dac_8bit_1/c1m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2806 vcp_sampled dac_8bit_0/amux_2to1_7/SELB dac_8bit_0/c1m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2807 input_amplifier_0/venp2 gain_ctrl_1 vampp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2808 dac_8bit_1/cdumm dac_8bit_1/amux_2to1_6/SELB vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2809 a_226938_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_226480_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2810 dac_8bit_1/latched_comparator_folded_0/vtailp vlowB dac_8bit_1/latched_comparator_folded_0/vlatchm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2811 dac_8bit_0/cdumm sample dac_8bit_0/amux_2to1_6/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2812 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2813 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2814 vcp_sampled dac_8bit_0/amux_2to1_3/SELB dac_8bit_0/c4m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2815 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/csinvp low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin a_247701_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X2816 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2817 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2818 dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2819 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2820 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2821 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2822 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2823 dac_8bit_1/amux_2to1_0/SELB sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2824 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2825 VDD VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2826 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2827 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2828 input_amplifier_0/venp1 input_amplifier_0/vop1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X2829 a_237498_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_237040_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X2830 dac_8bit_1/latched_comparator_folded_0/vlatchm vlowB dac_8bit_1/latched_comparator_folded_0/vtailp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2831 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2832 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X2833 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2834 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2835 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2836 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2837 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2838 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2839 VDD VDD vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2840 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2841 VDD VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2842 dac_8bit_1/amux_2to1_4/B sample dac_8bit_1/c3m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2843 vcp_sampled dac_8bit_0/amux_2to1_4/SELB dac_8bit_0/c3m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2844 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2845 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2846 input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vbias3 a_217060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2847 vampm VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X2848 dac_8bit_1/ibiasn dac_8bit_1/ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2849 dac_8bit_1/c4m dac_8bit_1/amux_2to1_3/SELB vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2850 dac_8bit_0/c4m sample dac_8bit_0/amux_2to1_3/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2851 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2852 input_amplifier_0/diff_fold_casc_ota_1/M6d input_amplifier_0/diff_fold_casc_ota_1/M6d input_amplifier_0/diff_fold_casc_ota_1/M6d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2853 a_237040_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_236582_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X2854 a_221480_n150168# vcp a_221022_n150168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2855 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2856 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/vcom_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2857 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X2858 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2859 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2860 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X2861 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2862 VDD VDD vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2863 vrefA q7A dac_8bit_0/amux_2to1_0/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2864 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2865 vampp input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2866 input_amplifier_0/diff_fold_casc_ota_1/M13d input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/M6d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2867 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2868 input_amplifier_0/diff_fold_casc_ota_0/M6d input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2869 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2870 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_241919_n121161# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2871 VSS sample dac_8bit_0/adc_run VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2872 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2873 VDD a_245649_n123369# a_245565_n123343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2874 a_338505_n185421# a_338285_n185409# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2875 a_236022_n132168# vcp low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/csinvn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2876 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X2877 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2878 a_337592_n185269# a_337864_n185269# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2879 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vfoldm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2880 biquad_gm_c_filter_0/gm_c_stage_3/vbiasp biquad_gm_c_filter_0/ibiasn3 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2881 VDD VDD vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2882 dac_8bit_1/amux_2to1_1/B sample dac_8bit_1/c6m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2883 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2884 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 a_356329_n164260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2885 vcp_sampled dac_8bit_0/amux_2to1_1/SELB dac_8bit_0/c6m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2886 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2887 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_2/A a_243382_n122255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2888 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X2889 adc_vcaparrayA dac_8bit_0/c1m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2890 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2891 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2892 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2893 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2894 a_236481_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_236023_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X2895 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/csinvp low_freq_pll_0/cs_ring_osc_0/vpbias a_224330_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X2896 a_356329_n113250# dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2897 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X2898 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2899 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2900 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2901 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2902 a_238771_n130007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin a_238313_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X2903 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2904 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2905 biquad_gm_c_filter_0/gm_c_stage_1/vcmc VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2906 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2907 VDD VDD vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2908 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2909 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2910 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2911 peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2912 a_338084_n185243# a_337592_n185269# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2913 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2914 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2915 VDD VDD diff_to_se_converter_0/vip VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2916 a_336537_n185409# a_336401_n185569# a_336116_n185555# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2917 a_224330_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_223872_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X2918 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2919 VDD VDD vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2920 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2921 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2922 biquad_gm_c_filter_0/gm_c_stage_0/vtail_diff biquad_gm_c_filter_0/ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2923 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2924 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 a_162668_n147576# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2925 VDD biquad_gm_c_filter_0/gm_c_stage_2/vbiasp biquad_gm_c_filter_0/gm_c_stage_2/vbiasp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2926 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2927 VDD VDD input_amplifier_0/diff_fold_casc_ota_0/M6d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2928 adc_vcaparrayB dac_8bit_1/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2929 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2930 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2931 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2932 vpeak_sampled vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X2933 a_223312_n132168# vcp a_222854_n132168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2934 a_242783_n121345# a_242085_n121711# a_242526_n121599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2935 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2936 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2937 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2938 VDD VDD vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2939 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2940 a_247702_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin a_247244_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2941 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_8/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2942 vampm VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X2943 a_242453_n122255# a_241919_n122249# a_242358_n122255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2944 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2945 VDD comparator_0/vcompm comparator_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2946 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2947 VSS low_freq_pll_0/pfd_cp_lpf_0/vQA low_freq_pll_0/pfd_cp_lpf_0/vQAb VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2948 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2949 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2950 input_amplifier_0/vip2 input_amplifier_0/txgate_7/txb input_amplifier_0/vom1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2951 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2952 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2953 a_223771_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin a_223313_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X2954 VSS vbiasn dac_8bit_0/ibiasp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=2e+06u
X2955 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2956 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2957 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2958 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2959 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X2960 adc_vcaparrayB dac_8bit_1/c0m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2961 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2962 vampp vampp vampp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2963 dac_8bit_0/amux_2to1_5/SELB sample VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2964 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2965 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X2966 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X2967 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2968 VSS a_245649_n122531# a_245607_n122799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2969 vcp_sampled vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X2970 VDD sample dac_8bit_0/adc_run VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2971 vpeak_sampled dac_8bit_1/amux_2to1_8/SELB dac_8bit_1/c0m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2972 dac_8bit_0/amux_2to1_9/Y sample dac_8bit_0/c0m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2973 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 a_217060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2974 sample_and_hold_1/vholdm vpeak_sampled sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X2975 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2976 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2977 input_amplifier_0/vim2 gain_ctrl_0 input_amplifier_0/venp1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2978 dac_8bit_1/latched_comparator_folded_0/vcompm VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2979 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2980 a_245481_n122255# a_244617_n122249# a_245224_n122281# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2981 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X2982 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2983 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2984 dac_8bit_1/amux_2to1_0/B q7B vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2985 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2986 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2987 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2988 vintp vfiltm biquad_gm_c_filter_0/gm_c_stage_2/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2989 VDD biquad_gm_c_filter_0/gm_c_stage_3/vbiasp biquad_gm_c_filter_0/gm_c_stage_3/vbiasp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2990 a_245607_n121877# a_244617_n122249# a_245481_n122255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2991 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2992 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X2993 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2994 low_freq_pll_0/pfd_cp_lpf_0/vpbias low_freq_pll_0/pfd_cp_lpf_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2995 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2996 dac_8bit_0/amux_2to1_2/SELB sample VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2997 dac_8bit_1/c0m sample dac_8bit_1/amux_2to1_9/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2998 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2999 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3000 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3001 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3002 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc vampp input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X3003 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3004 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X3005 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3006 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3007 a_163060_n102324# input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3008 a_226496_n122869# low_freq_pll_0/cs_ring_osc_0/vpbias a_226038_n122869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X3009 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 a_275374_n146348# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3010 diff_to_se_converter_0/vip vfiltp sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X3011 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3012 vlowA q0A dac_8bit_0/amux_2to1_9/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3013 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3014 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3015 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3016 dac_8bit_0/latched_comparator_folded_0/vtailp dac_8bit_0/vcom_buf dac_8bit_0/latched_comparator_folded_0/vlatchp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3017 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3018 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X3019 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3020 a_230446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3021 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3022 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3023 a_247701_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin a_247243_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X3024 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3025 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3026 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3027 dac_8bit_1/latched_comparator_folded_0/vtailp dac_8bit_1/ibiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3028 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3029 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X3030 vpeak_sampled dac_8bit_1/amux_2to1_6/SELB dac_8bit_1/cdumm VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3031 biquad_gm_c_filter_0/ibiasn4 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X3032 vcp VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3033 VDD VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3034 VDD VDD low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X3035 VSS VSS biquad_gm_c_filter_0/ibiasn3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3036 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vfoldm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3037 comparator_0/vcompp comparator_0/vcompp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3038 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3039 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3040 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3041 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3042 a_217060_n102324# input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3043 VDD VDD vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3044 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3045 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3046 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3047 a_243313_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_242855_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X3048 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3049 VDD VDD vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3050 a_275374_n180872# sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3051 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 a_356329_n164260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3052 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3053 vlowA q2A dac_8bit_0/amux_2to1_5/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3054 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3055 dac_8bit_1/latched_comparator_folded_0/vlatchm vlowB dac_8bit_1/latched_comparator_folded_0/vtailp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3056 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3057 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3058 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3059 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3060 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3061 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X3062 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3063 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3064 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3065 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3066 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc vampm input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X3067 vpeak_sampled dac_8bit_1/amux_2to1_3/SELB dac_8bit_1/c4m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3068 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3069 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3070 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3071 VSS biquad_gm_c_filter_0/gm_c_stage_0/vcmc biquad_gm_c_filter_0/gm_c_stage_0/vcmc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3072 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3073 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/vim1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X3074 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3075 VDD VDD vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3076 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3077 input_amplifier_0/diff_fold_casc_ota_1/vcascnm input_amplifier_0/diff_fold_casc_ota_1/vbias3 vampm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3078 sample_and_hold_1/vholdm VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3079 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3080 VDD VDD vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3081 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3082 input_amplifier_0/vop1 input_amplifier_0/vop1 input_amplifier_0/vop1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3083 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3084 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3085 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3086 VSS comparator_0/ibiasn comparator_0/ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3087 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X3088 vintp biquad_gm_c_filter_0/gm_c_stage_0/vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3089 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3090 a_239251_n114759# a_238627_n115125# a_239143_n115125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3091 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3092 a_226022_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3093 peak_detector_0/verr peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3094 a_228312_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_227854_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3095 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3096 VDD a_337497_n185269# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_0/Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3097 adc_vcaparrayA VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3098 adc_vcaparrayA dac_8bit_0/c3m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3099 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X3100 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3101 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3102 vpeak_sampled dac_8bit_1/amux_2to1_0/SELB dac_8bit_1/c7m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3103 VDD VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3104 VDD a_242783_n122255# a_242951_n122281# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3105 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3106 peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3107 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3108 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3109 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3110 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 vpeak VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3111 VDD VDD vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3112 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3113 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3114 peak_detector_0/ibiasn2 peak_detector_0/ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3115 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3116 a_238872_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_238414_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X3117 a_335749_n185813# a_335844_n185460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3118 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3119 VDD VDD biquad_gm_c_filter_0/gm_c_stage_0/vcmcn2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3120 vse diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3121 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3122 low_freq_pll_0/ibiasn vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X3123 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X3124 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3125 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3126 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3127 VSS dac_8bit_0/ibiasn dac_8bit_0/ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3128 vlowB sample adc_vcaparrayB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3129 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3130 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3131 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3132 input_amplifier_0/diff_fold_casc_ota_0/vcascnm input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3133 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3134 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3135 a_237854_n150168# vcp a_237396_n150168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3136 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3137 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3138 adc_vcaparrayB dac_8bit_1/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3139 VDD a_245649_n122531# a_245565_n122433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3140 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3141 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn vfiltm biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3142 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3143 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3144 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3145 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3146 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3147 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 a_163060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3148 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 a_189446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3149 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3150 dac_8bit_1/amux_2to1_7/SELB sample VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3151 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3152 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3153 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn1 vocm_filt biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3154 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/M1d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3155 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3156 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X3157 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3158 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 a_162668_n147576# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3159 vintm biquad_gm_c_filter_0/gm_c_stage_1/vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3160 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3161 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/vip2 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X3162 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3163 input_amplifier_0/vom1 VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X3164 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3165 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3166 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3167 dac_8bit_1/latched_comparator_folded_0/vcompm dac_8bit_1/latched_comparator_folded_0/vcompp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3168 vcp_sampled dac_8bit_0/amux_2to1_5/SELB dac_8bit_0/c2m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3169 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3170 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3171 a_223414_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_223872_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X3172 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3173 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3174 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3175 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3176 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3177 vampp input_amplifier_0/vim2 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X3178 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3179 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 a_356329_n164260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3180 dac_8bit_0/amux_2to1_7/B VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3181 a_336537_n185243# a_336401_n185269# a_336116_n185269# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3182 a_237548_n119618# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout a_237090_n119618# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3183 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3184 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3185 a_242419_n114983# vcomp VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3186 dac_8bit_1/amux_2to1_4/SELB sample VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3187 peak_detector_0/verr peak_detector_0/verr peak_detector_0/verr VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3188 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3189 a_245182_n122799# a_244783_n122799# a_245056_n122433# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3190 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3191 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3192 vampp input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3193 VSS a_242951_n120355# a_242909_n120623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3194 input_amplifier_0/vip2 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3195 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/vcom_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3196 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3197 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3198 vfiltm vintm biquad_gm_c_filter_0/gm_c_stage_3/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3199 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X3200 vpeak_sampled vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X3201 VDD VDD biquad_gm_c_filter_0/gm_c_stage_1/vcmcn2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3202 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp vse peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3203 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3204 dac_8bit_0/amux_2to1_9/Y q0A vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3205 input_amplifier_0/diff_fold_casc_ota_1/vcascnm input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3206 adc_vcaparrayB dac_8bit_1/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3207 vpeak_sampled vpeak_sampled vpeak_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3208 a_237090_n119618# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout a_236632_n119618# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3209 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3210 dac_8bit_1/c2m dac_8bit_1/amux_2to1_5/SELB vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3211 dac_8bit_0/c2m sample dac_8bit_0/amux_2to1_5/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3212 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X3213 VSS VSS biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3214 vcp_sampled dac_8bit_0/amux_2to1_2/SELB dac_8bit_0/c5m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3215 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3216 VSS low_freq_pll_0/ibiasn low_freq_pll_0/ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3217 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3218 a_242453_n121345# a_241919_n121711# a_242358_n121345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3219 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3220 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3221 peak_detector_0/ibiasn2 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X3222 biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail1 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3223 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3224 dac_8bit_0/amux_2to1_4/B VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3225 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3226 comparator_0/vcompm comparator_0/vcompp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3227 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3228 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3229 dac_8bit_1/amux_2to1_1/SELB sample VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3230 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3231 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3232 input_amplifier_0/venm2 input_amplifier_0/vip2 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X3233 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3234 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X3235 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/vcom_buf VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3236 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3237 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3238 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3239 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3240 VDD VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3241 vrefA dac_8bit_0/amux_2to1_11/SELB dac_8bit_0/amux_2to1_6/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3242 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3243 diff_to_se_converter_0/vim diff_to_se_converter_0/txgate_1/txb vfiltm VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3244 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3245 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3246 dac_8bit_1/c5m dac_8bit_1/amux_2to1_2/SELB vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3247 a_242102_n114873# a_242419_n114983# a_242377_n115125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3248 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3249 dac_8bit_0/c5m sample dac_8bit_0/amux_2to1_2/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3250 VSS a_245649_n122281# a_245607_n121877# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3251 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3252 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3253 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3254 biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail1 vintp biquad_gm_c_filter_0/gm_c_stage_2/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3255 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3256 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3257 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3258 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3259 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3260 comparator_0/vcompp vfiltm comparator_0/vtail VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3261 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3262 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3263 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/diff_fold_casc_ota_0/vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X3264 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/vcom_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3265 input_amplifier_0/vom1 VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X3266 dac_8bit_0/amux_2to1_1/B VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3267 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3268 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3269 input_amplifier_0/venm2 input_amplifier_0/vip2 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X3270 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3271 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3272 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3273 a_245481_n121345# a_244617_n121711# a_245224_n121599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3274 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/M6d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3275 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3276 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3277 a_163060_n102324# input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3278 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3279 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3280 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3281 VDD VDD vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3282 vrefA dac_8bit_0/amux_2to1_14/SELB dac_8bit_0/amux_2to1_3/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3283 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3284 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3285 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3286 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3287 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3288 input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/diff_fold_casc_ota_0/M2d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3289 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3290 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3291 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3292 vcp sample sample_and_hold_0/vhold VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3293 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3294 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 a_275374_n146348# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3295 VSS VSS vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3296 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3297 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3298 VDD VDD vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3299 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3300 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3301 a_227870_n122869# low_freq_pll_0/cs_ring_osc_0/vpbias a_227412_n122869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X3302 input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vbias3 a_217060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3303 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3304 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3305 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3306 input_amplifier_0/diff_fold_casc_ota_1/M3d VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3307 biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail2 vocm_filt biquad_gm_c_filter_0/gm_c_stage_0/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3308 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3309 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3310 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3311 VDD VDD vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3312 a_336401_n185569# adc_clk VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3313 vrefA dac_8bit_0/amux_2to1_17/SELB dac_8bit_0/amux_2to1_0/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3314 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3315 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3316 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3317 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/vcom_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3318 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X3319 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3320 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3321 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X3322 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3323 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3324 input_amplifier_0/txgate_5/txb input_amplifier_0/rst VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3325 biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail2 vintm biquad_gm_c_filter_0/gm_c_stage_1/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3326 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3327 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3328 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3329 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3330 a_242854_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_242396_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3331 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X3332 a_242358_n121345# a_241919_n121711# a_242273_n121711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3333 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3334 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3335 a_217060_n102324# input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3336 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3337 peak_detector_0/ibiasn1 peak_detector_0/ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3338 a_242273_n121711# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3339 VSS input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3340 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3341 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3342 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3343 VDD VDD vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3344 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3345 peak_detector_0/vpeak VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X3346 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3347 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/M2d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3348 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3349 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X3350 VSS a_245481_n121167# a_245649_n121193# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3351 a_242526_n121193# a_242358_n121167# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3352 biquad_gm_c_filter_0/gm_c_stage_0/vtail_diff vampm vintm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3353 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3354 input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/diff_fold_casc_ota_0/M2d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3355 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_2/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3356 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3357 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.4e+07u
X3358 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3359 input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vbias3 a_163060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3360 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3361 vpeak_sampled dac_8bit_1/amux_2to1_7/SELB dac_8bit_1/c1m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3362 dac_8bit_0/amux_2to1_7/B sample dac_8bit_0/c1m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3363 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3364 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3365 sample_and_hold_1/vhold VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3366 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3367 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3368 VSS dac_8bit_1/latched_comparator_folded_0/vcompp dac_8bit_1/latched_comparator_folded_0/vcomppb VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3369 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3370 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3371 low_freq_pll_0/freq_div_0/vin low_freq_pll_0/cs_ring_osc_0/vosc2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3372 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3373 vampm input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vfoldm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3374 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3375 adc_vcaparrayA dac_8bit_0/c2m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3376 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3377 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3378 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3379 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/vom1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3380 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1.2e+07u w=2e+06u
X3381 VSS a_242783_n120257# a_242951_n120355# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3382 dac_8bit_1/c1m sample dac_8bit_1/amux_2to1_7/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3383 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3384 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3385 a_189446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3386 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3387 adc_compB dac_8bit_1/comp_outm a_383050_n152139# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3388 a_242396_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_241938_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3389 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q a_245649_n123369# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3390 input_amplifier_0/vop1 VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3391 vpeak_sampled dac_8bit_1/amux_2to1_4/SELB dac_8bit_1/c3m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3392 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3393 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3394 a_238872_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_239330_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X3395 biquad_gm_c_filter_0/ibiasn3 biquad_gm_c_filter_0/ibiasn3 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3396 dac_8bit_0/amux_2to1_4/B sample dac_8bit_0/c3m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3397 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3398 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3399 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3400 vampp vampp vampp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3401 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn1 vocm_filt biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3402 input_amplifier_0/diff_fold_casc_ota_1/vcascnm input_amplifier_0/diff_fold_casc_ota_1/vbias3 vampm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3403 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3404 dac_8bit_1/amux_2to1_6/B VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3405 vcp_sampled VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3406 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3407 a_242358_n121167# a_242085_n121161# a_242273_n121167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3408 peak_detector_0/verr peak_detector_0/verr peak_detector_0/verr VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3409 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 vpeak VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3410 vlowA q1A dac_8bit_0/amux_2to1_7/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3411 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3412 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3413 dac_8bit_1/latched_comparator_folded_0/vtailp vlowB dac_8bit_1/latched_comparator_folded_0/vlatchm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3414 a_242484_n120623# a_242085_n120623# a_242358_n120257# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3415 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3416 dac_8bit_0/amux_2to1_6/B dac_8bit_0/amux_2to1_11/SELB vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3417 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3418 input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vbias3 a_217060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3419 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3420 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3421 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3422 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X3423 vrefB dac_8bit_1/amux_2to1_9/SELB dac_8bit_1/amux_2to1_9/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3424 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3425 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3426 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3427 input_amplifier_0/diff_fold_casc_ota_1/M2d input_amplifier_0/diff_fold_casc_ota_1/M2d input_amplifier_0/diff_fold_casc_ota_1/M2d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3428 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 a_230446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3429 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3430 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3431 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3432 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X3433 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3434 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3435 dac_8bit_1/c3m sample dac_8bit_1/amux_2to1_4/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3436 vse diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3437 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3438 dac_8bit_0/latched_comparator_folded_0/vcompm dac_8bit_0/latched_comparator_folded_0/vcompp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3439 vlowA dac_8bit_0/adc_run adc_vcaparrayA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3440 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3441 vpeak_sampled dac_8bit_1/amux_2to1_1/SELB dac_8bit_1/c6m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3442 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3443 VSS dac_8bit_0/ibiasn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3444 dac_8bit_0/amux_2to1_1/B sample dac_8bit_0/c6m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3445 input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3446 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 a_162668_n147576# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3447 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3448 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3449 VSS a_242951_n122531# a_243382_n122477# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3450 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3451 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X3452 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 a_275374_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3453 VDD VDD vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3454 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3455 dac_8bit_1/amux_2to1_3/B VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3456 vcp_sampled VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3457 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3458 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3459 a_338149_n185269# adc_clk VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3460 vlowA q3A dac_8bit_0/amux_2to1_4/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3461 sample_and_hold_1/vholdm sample vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3462 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3463 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3464 dac_8bit_0/amux_2to1_3/B dac_8bit_0/amux_2to1_14/SELB vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3465 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3466 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/vip2 input_amplifier_0/diff_fold_casc_ota_1/vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X3467 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3468 vintm biquad_gm_c_filter_0/gm_c_stage_0/vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3469 adc_vcaparrayA dac_8bit_0/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3470 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3471 a_245224_n121193# a_245056_n121167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X3472 VSS biquad_gm_c_filter_0/ibiasn3 biquad_gm_c_filter_0/ibiasn3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3473 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3474 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3475 vrefB dac_8bit_1/amux_2to1_12/SELB dac_8bit_1/amux_2to1_5/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3476 a_241188_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_240730_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X3477 vfiltp diff_to_se_converter_0/txgate_0/txb diff_to_se_converter_0/vip VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3478 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/vip2 input_amplifier_0/diff_fold_casc_ota_1/vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X3479 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 vocm input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X3480 VSS input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3481 vpeak_sampled dac_8bit_1/amux_2to1_2/SELB dac_8bit_1/c5m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3482 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3483 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3484 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3485 VDD VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3486 a_356329_n113250# dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3487 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3488 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3489 VSS VSS dac_8bit_1/latched_comparator_folded_0/vlatchp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3490 dac_8bit_1/c6m sample dac_8bit_1/amux_2to1_1/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3491 a_238922_n119618# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout a_238464_n119618# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3492 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/verr VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3493 sample_and_hold_1/vholdm vpeak_sampled sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X3494 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3495 a_245481_n121167# a_244783_n121161# a_245224_n121193# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3496 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3497 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3498 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3499 vampp input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3500 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3501 VSS a_336401_n185569# a_336408_n185665# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3502 vampp VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X3503 VDD VDD vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3504 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X3505 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3506 input_amplifier_0/venm1 input_amplifier_0/vom1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X3507 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3508 vlowA q6A dac_8bit_0/amux_2to1_1/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3509 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3510 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X3511 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X3512 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3513 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3514 vpeak_sampled VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X3515 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3516 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3517 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q a_242951_n121193# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3518 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X3519 input_amplifier_0/ibiasn2 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X3520 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3521 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3522 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X3523 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3524 dac_8bit_1/latched_comparator_folded_0/vcompp adc_clk dac_8bit_1/latched_comparator_folded_0/vlatchp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3525 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_7/A a_246080_n121389# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3526 dac_8bit_1/c7m sample vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3527 VDD VDD input_amplifier_0/diff_fold_casc_ota_1/vfoldm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3528 VSS VSS low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3529 VSS biquad_gm_c_filter_0/ibiasn1 biquad_gm_c_filter_0/ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3530 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X3531 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3532 input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3533 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3534 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3535 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3536 dac_8bit_0/c7m dac_8bit_0/amux_2to1_0/SELB dac_8bit_0/amux_2to1_0/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3537 input_amplifier_0/venm1 input_amplifier_0/vom1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X3538 VDD VDD vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3539 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3540 comparator_0/vo1 comparator_0/vo1 comparator_0/vo1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3541 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3542 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3543 a_356329_n113250# dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3544 a_335749_n185813# a_335844_n185460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3545 vintp biquad_gm_c_filter_0/gm_c_stage_1/vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3546 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3547 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3548 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3549 VDD VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3550 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3551 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 a_189446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3552 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3553 dac_8bit_1/latched_comparator_folded_0/vcompp dac_8bit_1/latched_comparator_folded_0/vcompm VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3554 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3555 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3556 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3557 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3558 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3559 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3560 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3561 input_amplifier_0/diff_fold_casc_ota_1/vcascnp input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3562 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X3563 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 a_356329_n113250# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3564 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3565 a_189446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3566 VSS dac_8bit_1/ibiasn dac_8bit_1/ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3567 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3568 a_240062_n115125# low_freq_pll_0/pfd_cp_lpf_0/vRSTN VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3569 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3570 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3571 a_227870_n122869# low_freq_pll_0/cs_ring_osc_0/vpbias a_228328_n122869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X3572 input_amplifier_0/vip2 gain_ctrl_0 input_amplifier_0/venm1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3573 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3574 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3575 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3576 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q a_244617_n123337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3577 vfiltp vintp biquad_gm_c_filter_0/gm_c_stage_3/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3578 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3579 VSS VSS low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3580 input_amplifier_0/vip2 input_amplifier_0/vom1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X3581 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3582 a_162668_n147576# diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3583 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3584 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X3585 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3586 vrefA dac_8bit_0/amux_2to1_9/SELB dac_8bit_0/amux_2to1_9/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3587 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3588 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3589 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3590 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3591 VDD dac_8bit_1/latched_comparator_folded_0/vcompp dac_8bit_1/latched_comparator_folded_0/vcompm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3592 a_217060_n102324# input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3593 VSS VSS biquad_gm_c_filter_0/gm_c_stage_1/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3594 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3595 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3596 comparator_0/vcompp comparator_0/vcompm VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3597 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3598 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 a_275374_n146348# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3599 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3600 dac_8bit_1/amux_2to1_6/B sample dac_8bit_1/cdumm VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3601 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3602 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 a_189446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3603 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3604 biquad_gm_c_filter_0/ibiasn2 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3605 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3606 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3607 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3608 a_230870_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin a_230412_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3609 input_amplifier_0/diff_fold_casc_ota_0/M13d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3610 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3611 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3612 sample_and_hold_0/vholdm vcp_sampled sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X3613 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3614 a_242575_n114888# a_242380_n114857# a_242885_n115125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3615 biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail2 biquad_gm_c_filter_0/ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3616 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3617 dac_8bit_0/amux_2to1_7/B q1A vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3618 vcp_sampled vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X3619 vpeak_sampled VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3620 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3621 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3622 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3623 dac_8bit_1/amux_2to1_9/Y dac_8bit_1/amux_2to1_9/SELB vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3624 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3625 a_242273_n121167# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3626 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3627 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3628 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X3629 comparator_0/vcompm vfiltp comparator_0/vtail VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3630 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3631 VSS input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3632 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3633 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 a_356329_n164260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3634 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3635 input_amplifier_0/vom1 input_amplifier_0/vom1 input_amplifier_0/vom1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3636 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3637 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3638 dac_8bit_1/amux_2to1_3/B sample dac_8bit_1/c4m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3639 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3640 a_241939_n130007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_241481_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X3641 peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3642 dac_8bit_0/amux_2to1_4/B q3A vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3643 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3644 VDD comparator_0/vcompm comparator_0/vcompp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3645 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3646 vlowB VSS dac_8bit_1/amux_2to1_6/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3647 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3648 input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X3649 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3650 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3651 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3652 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3653 VSS a_337592_n185269# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/D VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3654 vcp sample sample_and_hold_0/vhold VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3655 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3656 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3657 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3658 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3659 a_230412_n134960# vcp a_229954_n134960# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3660 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3661 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 vse VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3662 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3663 VSS input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3664 a_245056_n123343# a_244783_n123337# a_244971_n123343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3665 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3666 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3667 input_amplifier_0/diff_fold_casc_ota_1/M13d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3668 vincm input_amplifier_0/txgate_5/txb input_amplifier_0/vip1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3669 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3670 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3671 peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3672 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_243770_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3673 VSS a_335844_n185460# pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3674 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3675 VDD vbiasp input_amplifier_0/ibiasn1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X3676 a_237040_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_237498_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X3677 vrefA dac_8bit_0/amux_2to1_15/SELB dac_8bit_0/amux_2to1_2/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3678 input_amplifier_0/txgate_4/txb input_amplifier_0/rst VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3679 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X3680 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 vcp_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3681 a_244954_n134960# vcp VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3682 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3683 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3684 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3685 dac_8bit_0/amux_2to1_1/B q6A vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3686 a_240730_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X3687 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3688 vlowB q4B dac_8bit_1/amux_2to1_3/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3689 adc_vcaparrayA dac_8bit_0/c3m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3690 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3691 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3692 VDD low_freq_pll_0/cs_ring_osc_0/vpbias a_221582_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X3693 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3694 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3695 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3696 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3697 a_245869_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin a_245411_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X3698 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q a_245649_n121443# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3699 VSS VSS biquad_gm_c_filter_0/gm_c_stage_1/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3700 a_242358_n120257# a_242085_n120623# a_242273_n120623# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3701 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3702 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 input_amplifier_0/ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3703 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3704 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3705 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3706 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3707 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 a_230446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3708 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3709 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3710 VDD VDD vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3711 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn2 vocm_filt biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3712 a_189446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3713 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3714 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3715 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3716 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3717 input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X3718 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3719 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3720 vlowB q7B dac_8bit_1/amux_2to1_0/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3721 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3722 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3723 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3724 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3725 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 vpeak VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3726 adc_vcaparrayB dac_8bit_1/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3727 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3728 input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3729 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3730 VSS a_242951_n122281# a_243382_n122255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3731 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3732 input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc vocm input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X3733 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/vip2 input_amplifier_0/diff_fold_casc_ota_1/vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X3734 biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail2 vocm_filt biquad_gm_c_filter_0/gm_c_stage_2/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3735 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 a_162668_n147576# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3736 a_232244_n134960# vcp a_231786_n134960# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3737 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3738 VSS a_335749_n185269# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/Q_N VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3739 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3740 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3741 biquad_gm_c_filter_0/gm_c_stage_1/vtail_diff vintp vintp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3742 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X3743 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X3744 sample_and_hold_1/vhold sample vpeak VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3745 low_freq_pll_0/pfd_cp_lpf_0/vpbias low_freq_pll_0/pfd_cp_lpf_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3746 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/csinvp low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin a_232701_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X3747 dac_8bit_0/cdumm sample dac_8bit_0/amux_2to1_6/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3748 a_337592_n185460# a_337864_n185555# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3749 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3750 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3751 input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X3752 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3753 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3754 VSS low_freq_pll_0/cs_ring_osc_0/vosc2 low_freq_pll_0/freq_div_0/vin VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3755 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3756 VSS a_245224_n121599# a_245182_n121711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3757 VSS vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3758 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3759 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3760 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 a_230446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3761 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3762 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3763 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/vim2 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X3764 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3765 a_222498_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_222040_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X3766 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3767 a_163060_n102324# input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3768 a_236481_n130007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin a_236023_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X3769 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X3770 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3771 VSS comparator_0/ibiasn comparator_0/vtail VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3772 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3773 input_amplifier_0/vim1 vincm sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X3774 input_amplifier_0/vop1 input_amplifier_0/txgate_6/txb input_amplifier_0/vim2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3775 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3776 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3777 a_356329_n113250# dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3778 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X3779 a_222040_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_221582_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X3780 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X3781 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3782 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3783 dac_8bit_0/c4m sample dac_8bit_0/amux_2to1_3/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3784 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3785 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3786 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3787 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3788 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3789 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3790 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3791 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X3792 vampp input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3793 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X3794 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3795 VSS vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3796 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3797 input_amplifier_0/vom1 input_amplifier_0/vom1 input_amplifier_0/vom1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3798 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3799 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3800 VDD VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3801 biquad_gm_c_filter_0/gm_c_stage_2/vtail_diff VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3802 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3803 vlowA VSS dac_8bit_0/amux_2to1_6/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3804 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3805 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3806 a_238770_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_238312_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3807 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3808 a_221022_n132168# vcp low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/csinvn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3809 VSS input_amplifier_0/ibiasn1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3810 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X3811 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3812 input_amplifier_0/vom1 input_amplifier_0/txgate_7/txb input_amplifier_0/vip2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3813 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3814 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3815 VDD VDD adc_vcaparrayA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3816 input_amplifier_0/vop1 VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X3817 vrefA VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3818 a_245412_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin a_244954_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3819 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3820 biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail1 vocm_filt biquad_gm_c_filter_0/gm_c_stage_2/vcmcn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3821 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3822 dac_8bit_1/amux_2to1_5/B VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3823 vcp_sampled VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3824 vse diff_to_se_converter_0/vim sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X3825 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3826 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3827 VDD VDD a_243138_n114759# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3828 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3829 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3830 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3831 dac_8bit_0/amux_2to1_5/B dac_8bit_0/amux_2to1_12/SELB vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3832 input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X3833 a_217060_n102324# input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3834 VDD VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3835 a_221481_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin a_221023_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X3836 dac_8bit_1/amux_2to1_0/B q7B vrefB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3837 a_223771_n130007# low_freq_pll_0/cs_ring_osc_0/vosc a_223313_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X3838 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3839 VDD a_337592_n185269# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/D VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3840 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3841 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3842 vrefB dac_8bit_1/amux_2to1_10/SELB dac_8bit_1/amux_2to1_7/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3843 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3844 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3845 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3846 dac_8bit_1/amux_2to1_6/B VSS vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3847 dac_8bit_0/amux_2to1_0/B dac_8bit_0/amux_2to1_17/SELB vlowA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3848 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3849 input_amplifier_0/venm1 input_amplifier_0/vom1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X3850 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3851 vlowA q4A dac_8bit_0/amux_2to1_3/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3852 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3853 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3854 VSS low_freq_pll_0/ibiasn low_freq_pll_0/ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3855 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3856 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3857 VDD a_245224_n121193# a_245151_n121167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3858 dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3859 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/M1d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3860 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X3861 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3862 VDD low_freq_pll_0/pfd_cp_lpf_0/vpbias low_freq_pll_0/pfd_cp_lpf_0/vpbias VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3863 dac_8bit_1/amux_2to1_2/B VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3864 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3865 input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3866 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3867 sample_and_hold_0/vholdm sample vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3868 vcp_sampled VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3869 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3870 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3871 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3872 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3873 a_226038_n122869# low_freq_pll_0/cs_ring_osc_0/vpbias a_226496_n122869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X3874 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 a_189446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3875 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3876 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3877 dac_8bit_0/amux_2to1_2/B dac_8bit_0/amux_2to1_15/SELB vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3878 input_amplifier_0/vom1 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3879 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3880 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vfoldm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3881 a_336116_n185555# a_336408_n185665# a_336359_n185787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3882 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3883 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3884 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3885 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3886 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 vse VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3887 a_242526_n122687# a_242358_n122433# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3888 vrefB dac_8bit_1/amux_2to1_13/SELB dac_8bit_1/amux_2to1_4/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3889 a_232702_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin a_232244_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3890 biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail2 vintp biquad_gm_c_filter_0/gm_c_stage_0/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3891 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3892 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3893 dac_8bit_1/amux_2to1_3/B q4B vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3894 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3895 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3896 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3897 a_335844_n185460# a_336116_n185555# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3898 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3899 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3900 comparator_0/vmirror comparator_0/vmirror VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3901 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3902 diff_to_se_converter_0/vip diff_to_se_converter_0/txgate_0/txb vfiltp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3903 dac_8bit_1/ibiasn vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X3904 a_245056_n121167# a_244617_n121161# a_244971_n121167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3905 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3906 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3907 a_247244_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin a_246786_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3908 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 a_189446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3909 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3910 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3911 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3912 a_163060_n102324# input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3913 VSS low_freq_pll_0/ibiasn low_freq_pll_0/pfd_cp_lpf_0/vswitchl VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3914 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3915 dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3916 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3917 dac_8bit_0/ibiasp vbiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=2e+06u
X3918 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3919 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3920 biquad_gm_c_filter_0/ibiasn4 biquad_gm_c_filter_0/ibiasn4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3921 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3922 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3923 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3924 vrefB dac_8bit_1/amux_2to1_16/SELB dac_8bit_1/amux_2to1_1/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3925 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3926 a_162668_n147576# diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3927 dac_8bit_1/latched_comparator_folded_0/vlatchp VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X3928 a_245411_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin a_244953_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X3929 a_230446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3930 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3931 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn vintp biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3932 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3933 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3934 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3935 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3936 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 a_356329_n113250# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3937 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3938 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X3939 VSS a_239883_n115151# a_240447_n115125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3940 VDD VDD low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X3941 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3942 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3943 biquad_gm_c_filter_0/gm_c_stage_0/vtail_diff vampp vintp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3944 VSS comparator_0/vmirror comparator_0/vo1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3945 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/verr VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3946 VSS input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3947 VSS vpeak_sampled sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X3948 a_245607_n121711# a_244617_n121711# a_245481_n121345# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3949 a_241023_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X3950 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 a_275374_n146348# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3951 a_243313_n130007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_242855_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X3952 vcp_sampled VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X3953 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3954 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3955 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3956 VDD dac_8bit_1/latched_comparator_folded_0/vcompp_buf dac_8bit_1/comp_outm VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3957 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3958 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 a_356329_n164260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3959 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3960 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3961 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3962 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3963 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3964 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q a_241919_n122249# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3965 dac_8bit_1/c0m sample dac_8bit_1/amux_2to1_9/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3966 VSS VSS biquad_gm_c_filter_0/gm_c_stage_0/vbiasp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3967 dac_8bit_0/c0m dac_8bit_0/amux_2to1_8/SELB vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3968 a_245056_n122433# a_244783_n122799# a_244971_n122799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3969 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3970 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3971 VDD VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3972 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3973 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3974 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3975 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3976 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/vim2 input_amplifier_0/diff_fold_casc_ota_1/vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X3977 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3978 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3979 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3980 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3981 input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vbias3 a_163060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3982 vampm input_amplifier_0/txgate_2/txb input_amplifier_0/venm2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3983 a_232701_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin a_232243_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X3984 input_amplifier_0/diff_fold_casc_ota_0/M3d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3985 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3986 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3987 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3988 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3989 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3990 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3991 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3992 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X3993 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3994 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3995 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X3996 vpeak_sampled VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X3997 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3998 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3999 vampm input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4000 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4001 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4002 adc_vcaparrayA dac_8bit_0/c2m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4003 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4004 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4005 VDD vbiasp biquad_gm_c_filter_0/ibiasn2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X4006 input_amplifier_0/vip2 input_amplifier_0/vom1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X4007 VSS sample pulse_generator_0/sky130_fd_sc_hd__inv_1_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4008 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4009 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4010 a_226022_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4011 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4012 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4013 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4014 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4015 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4016 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4017 vrefA dac_8bit_0/amux_2to1_10/SELB dac_8bit_0/amux_2to1_7/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4018 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4019 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4020 a_247243_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin a_246785_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X4021 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 vcp_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4022 input_amplifier_0/ibiasn2 input_amplifier_0/ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4023 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4024 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4025 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4026 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4027 input_amplifier_0/venm2 input_amplifier_0/vip2 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X4028 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1.2e+07u w=2e+06u
X4029 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4030 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4031 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4032 input_amplifier_0/vop1 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4033 VSS input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4034 vlowB q0B dac_8bit_1/amux_2to1_9/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4035 a_338107_n185787# a_337592_n185460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4036 VSS dac_8bit_0/vcom_buf sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X4037 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4038 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X4039 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X4040 dac_8bit_1/amux_2to1_5/B sample dac_8bit_1/c2m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4041 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4042 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4043 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4044 dac_8bit_0/latched_comparator_folded_0/vlatchp dac_8bit_0/vcom_buf dac_8bit_0/latched_comparator_folded_0/vtailp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4045 VSS biquad_gm_c_filter_0/gm_c_stage_3/vcmc biquad_gm_c_filter_0/gm_c_stage_3/vcmc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4046 a_236582_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X4047 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4048 low_freq_pll_0/pfd_cp_lpf_0/vswitchh low_freq_pll_0/pfd_cp_lpf_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4049 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X4050 vpeak_sampled VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4051 input_amplifier_0/vim2 VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4052 input_amplifier_0/vom1 VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X4053 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4054 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4055 input_amplifier_0/diff_fold_casc_ota_0/vcascnp input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4056 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4057 dac_8bit_1/amux_2to1_7/B dac_8bit_1/amux_2to1_10/SELB vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4058 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4059 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4060 VDD comparator_0/vcompp comparator_0/vcompm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4061 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4062 vampm gain_ctrl_1 input_amplifier_0/venm2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4063 vrefA dac_8bit_0/amux_2to1_13/SELB dac_8bit_0/amux_2to1_4/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4064 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/csinvn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4065 a_245224_n123369# a_245056_n123343# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4066 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 input_amplifier_0/ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4067 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4068 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4069 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4070 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4071 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 a_162668_n147576# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4072 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4073 a_244971_n121167# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4074 vlowA VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4075 VDD a_242951_n122281# a_242867_n122255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4076 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4077 input_amplifier_0/diff_fold_casc_ota_0/M6d input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4078 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4079 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4080 dac_8bit_1/amux_2to1_2/B sample dac_8bit_1/c5m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4081 VDD a_239361_n114883# a_239251_n114759# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4082 VDD dac_8bit_0/ibiasp dac_8bit_0/latched_comparator_folded_0/vtailp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4083 VSS a_245224_n121193# a_245182_n120789# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4084 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4085 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 a_162668_n147576# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4086 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4087 vpeak_sampled VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4088 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 a_275374_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4089 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4090 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4091 a_242336_n114759# a_241731_n115151# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4092 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4093 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4094 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4095 dac_8bit_1/amux_2to1_4/B dac_8bit_1/amux_2to1_13/SELB vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4096 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4097 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 a_230446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4098 vrefA dac_8bit_0/amux_2to1_16/SELB dac_8bit_0/amux_2to1_1/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4099 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4100 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4101 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4102 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4103 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4104 a_223872_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_223414_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X4105 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4106 input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc vocm input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X4107 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X4108 VSS VSS vpeak VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4109 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_241919_n121161# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4110 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4111 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4112 input_amplifier_0/diff_fold_casc_ota_1/M6d input_amplifier_0/diff_fold_casc_ota_1/M6d input_amplifier_0/diff_fold_casc_ota_1/M6d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4113 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X4114 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4115 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4116 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4117 vlowA VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4118 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4119 VDD VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4120 VSS vpeak_sampled vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4121 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 a_162668_n147576# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4122 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4123 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4124 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4125 VSS pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/D a_336955_n185243# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4126 a_222854_n150168# vcp a_222396_n150168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4127 input_amplifier_0/diff_fold_casc_ota_1/M2d input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/M3d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4128 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4129 vpeak_sampled VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4130 vlowB q5B dac_8bit_1/amux_2to1_2/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4131 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4132 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4133 biquad_gm_c_filter_0/gm_c_stage_3/vtail_diff biquad_gm_c_filter_0/ibiasn3 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4134 dac_8bit_1/amux_2to1_1/B dac_8bit_1/amux_2to1_16/SELB vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4135 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4136 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4137 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/M2d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4138 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/vim1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X4139 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4140 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4141 VDD VDD dac_8bit_0/latched_comparator_folded_0/vlatchp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X4142 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X4143 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp vse peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4144 input_amplifier_0/venm2 input_amplifier_0/txgate_2/txb vampm VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4145 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4146 a_237396_n150168# vcp a_236938_n150168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4147 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4148 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4149 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4150 input_amplifier_0/diff_fold_casc_ota_1/M6d input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4151 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 a_230446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4152 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4153 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn2 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn2 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4154 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4155 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4156 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4157 a_237855_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_237397_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X4158 a_244971_n122799# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4159 VDD low_freq_pll_0/pfd_cp_lpf_0/vpbias low_freq_pll_0/pfd_cp_lpf_0/vswitchh VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4160 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X4161 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4162 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4163 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4164 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4165 dac_8bit_1/amux_2to1_0/B VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4166 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4167 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4168 biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail2 vocm_filt biquad_gm_c_filter_0/gm_c_stage_3/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4169 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4170 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4171 a_242867_n121167# a_242085_n121161# a_242783_n121167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4172 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 a_275374_n146348# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4173 VDD a_245649_n121443# a_246080_n121389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4174 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4175 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X4176 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4177 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4178 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4179 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4180 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4181 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4182 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4183 a_336116_n185269# a_336408_n184969# a_336359_n184877# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4184 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4185 a_383508_n152139# adc_compB dac_8bit_1/comp_outm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4186 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4187 input_amplifier_0/diff_fold_casc_ota_1/M2d input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/M3d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4188 adc_vcaparrayA dac_8bit_0/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4189 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4190 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4191 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4192 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4193 VDD dac_8bit_1/latched_comparator_folded_0/vcompm dac_8bit_1/latched_comparator_folded_0/vcompp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4194 dac_8bit_0/c2m sample dac_8bit_0/amux_2to1_5/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4195 dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4196 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4197 input_amplifier_0/diff_fold_casc_ota_0/vcascnp input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/vop1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4198 a_162668_n147576# diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4199 VDD VDD input_amplifier_0/diff_fold_casc_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4200 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4201 adc_vcaparrayA dac_8bit_0/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4202 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/M2d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4203 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 input_amplifier_0/ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4204 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4205 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4206 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4207 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4208 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4209 dac_8bit_1/latched_comparator_folded_0/vcompmb dac_8bit_1/latched_comparator_folded_0/vcompm VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4210 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4211 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4212 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4213 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4214 biquad_gm_c_filter_0/gm_c_stage_3/vtail_diff vintp vfiltp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4215 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4216 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4217 a_225580_n122869# low_freq_pll_0/cs_ring_osc_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X4218 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/vip2 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X4219 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn2 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn2 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4220 diff_to_se_converter_0/ibiasn vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X4221 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4222 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4223 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4224 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4225 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4226 input_amplifier_0/diff_fold_casc_ota_0/M1d input_amplifier_0/diff_fold_casc_ota_0/M1d input_amplifier_0/diff_fold_casc_ota_0/M1d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4227 VDD VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4228 a_275374_n180872# sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4229 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4230 dac_8bit_0/c5m sample dac_8bit_0/amux_2to1_2/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4231 VSS VSS vincm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4232 VSS vse sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X4233 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4234 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4235 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4236 vampm vampm vampm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4237 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4238 VSS biquad_gm_c_filter_0/ibiasn1 biquad_gm_c_filter_0/ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4239 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X4240 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4241 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4242 a_242137_n115125# a_242102_n114873# a_241731_n115151# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4243 VSS a_336608_n185510# a_336537_n185409# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4244 biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail1 vocm_filt biquad_gm_c_filter_0/gm_c_stage_3/vcmcn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4245 vlowA q2A dac_8bit_0/amux_2to1_5/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4246 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4247 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4248 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4249 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 vcp_sampled VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4250 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4251 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4252 a_228771_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_228313_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X4253 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4254 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4255 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4256 a_242085_n120623# a_241919_n120623# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4257 vrefB dac_8bit_1/amux_2to1_11/SELB dac_8bit_1/amux_2to1_6/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4258 vrefA VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4259 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4260 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4261 VDD low_freq_pll_0/pfd_cp_lpf_0/vRSTN a_242720_n114759# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4262 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4263 vlowB VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4264 a_163060_n102324# input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4265 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4266 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X4267 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4268 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4269 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4270 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4271 dac_8bit_1/vcom_buf VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X4272 VSS diff_to_se_converter_0/ibiasn diff_to_se_converter_0/ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4273 comparator_0/vtail vfiltp comparator_0/vcompm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4274 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4275 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4276 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4277 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4278 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4279 dac_8bit_1/amux_2to1_5/B q2B vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4280 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4281 dac_8bit_0/amux_2to1_11/SELB VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4282 vlowA q5A dac_8bit_0/amux_2to1_2/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4283 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4284 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4285 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4286 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4287 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4288 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/vip2 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X4289 vrefB dac_8bit_1/amux_2to1_14/SELB dac_8bit_1/amux_2to1_3/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4290 vrefA VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4291 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4292 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4293 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4294 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4295 sample_and_hold_0/vhold VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X4296 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4297 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4298 input_amplifier_0/diff_fold_casc_ota_1/M1d input_amplifier_0/diff_fold_casc_ota_1/M1d input_amplifier_0/diff_fold_casc_ota_1/M1d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4299 VSS biquad_gm_c_filter_0/ibiasn4 biquad_gm_c_filter_0/ibiasn4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4300 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4301 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4302 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4303 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4304 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4305 sample_and_hold_0/vhold sample vcp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4306 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4307 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4308 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4309 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4310 input_amplifier_0/diff_fold_casc_ota_0/M1d input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4311 a_238414_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_237956_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X4312 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4313 VDD a_336401_n185569# a_336408_n185665# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4314 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4315 dac_8bit_1/amux_2to1_2/B q5B vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4316 VSS input_amplifier_0/ibiasn1 input_amplifier_0/ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4317 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4318 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp vse peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4319 dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4320 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4321 a_338107_n184877# a_337592_n185269# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4322 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4323 dac_8bit_0/amux_2to1_14/SELB q4A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4324 VDD VDD input_amplifier_0/diff_fold_casc_ota_1/M3d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4325 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4326 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4327 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4328 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/vim1 input_amplifier_0/diff_fold_casc_ota_0/vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X4329 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4330 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4331 VSS VSS dac_8bit_1/latched_comparator_folded_0/vlatchm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X4332 biquad_gm_c_filter_0/ibiasn2 biquad_gm_c_filter_0/ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4333 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4334 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4335 VSS input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4336 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4337 a_242396_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_241938_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4338 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4339 vrefA VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4340 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4341 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4342 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4343 peak_detector_0/vpeak peak_detector_0/verr VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4344 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4345 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4346 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4347 a_275374_n146348# sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4348 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4349 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4350 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4351 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4352 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4353 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4354 vampm input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4355 dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4356 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4357 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4358 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4359 VDD a_242951_n121443# a_242867_n121345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4360 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4361 biquad_gm_c_filter_0/gm_c_stage_1/vtail_diff vintm vintm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4362 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4363 input_amplifier_0/diff_fold_casc_ota_0/vfoldm VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4364 VSS input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4365 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4366 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4367 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4368 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4369 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4370 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X4371 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X4372 vpeak vpeak vpeak VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4373 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4374 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4375 vpeak_sampled vpeak_sampled vpeak_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4376 vampp VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X4377 a_223872_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_224330_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X4378 sample_and_hold_0/vholdm vcp_sampled sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X4379 a_242526_n123369# a_242358_n123343# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X4380 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4381 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4382 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4383 a_356329_n164260# dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4384 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4385 vintm vampm biquad_gm_c_filter_0/gm_c_stage_0/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4386 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/vcom_buf VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4387 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4388 VDD low_freq_pll_0/cs_ring_osc_0/vosc2 low_freq_pll_0/freq_div_0/vin VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4389 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4390 dac_8bit_0/c7m dac_8bit_0/amux_2to1_0/SELB vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4391 dac_8bit_1/c1m sample dac_8bit_1/amux_2to1_7/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4392 a_242783_n123343# a_242085_n123337# a_242526_n123369# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4393 dac_8bit_0/c1m dac_8bit_0/amux_2to1_7/SELB vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4394 a_163060_n102324# input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4395 a_239330_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X4396 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4397 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4398 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4399 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4400 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4401 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X4402 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4403 VDD a_239883_n115151# a_239870_n114759# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4404 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4405 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4406 VSS VSS vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4407 a_236632_n119618# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout a_236174_n119618# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4408 VSS vcp_sampled sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X4409 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4410 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4411 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4412 a_383050_n152139# dac_8bit_1/latched_comparator_folded_0/vcompm_buf VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4413 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4414 VDD a_245481_n123343# a_245649_n123369# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4415 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4416 input_amplifier_0/vop1 input_amplifier_0/rst input_amplifier_0/vim2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4417 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4418 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 vcp_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4419 a_242526_n121599# a_242358_n121345# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X4420 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4421 VSS vcp a_238770_n150168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4422 a_239143_n115125# a_238627_n115125# a_239048_n115125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4423 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4424 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4425 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4426 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4427 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4428 input_amplifier_0/vim1 input_amplifier_0/txgate_4/txb vincm VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4429 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4430 a_245565_n123343# a_244783_n123337# a_245481_n123343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4431 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4432 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4433 VDD vbiasp biquad_gm_c_filter_0/ibiasn1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X4434 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4435 input_amplifier_0/diff_fold_casc_ota_1/vcascnp input_amplifier_0/diff_fold_casc_ota_1/vbias3 vampp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4436 input_amplifier_0/vim2 input_amplifier_0/txgate_1/txb input_amplifier_0/venp1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4437 dac_8bit_1/c3m sample dac_8bit_1/amux_2to1_4/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4438 dac_8bit_0/c3m dac_8bit_0/amux_2to1_4/SELB vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4439 VSS VSS biquad_gm_c_filter_0/ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4440 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4441 biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail1 vintm biquad_gm_c_filter_0/gm_c_stage_0/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4442 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4443 a_243138_n114759# a_242380_n114857# a_242575_n114888# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4444 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4445 dac_8bit_0/amux_2to1_8/SELB sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4446 a_244971_n122255# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4447 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4448 vcp_sampled vcp_sampled vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4449 vlowB q1B dac_8bit_1/amux_2to1_7/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4450 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4451 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4452 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4453 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4454 dac_8bit_1/latched_comparator_folded_0/vlatchm vlowB dac_8bit_1/latched_comparator_folded_0/vtailp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4455 VSS vpeak_sampled sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X4456 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4457 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4458 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4459 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4460 vampm input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4461 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4462 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4463 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4464 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4465 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4466 adc_vcaparrayB dac_8bit_1/adc_run vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4467 a_242867_n120257# a_242085_n120623# a_242783_n120257# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4468 input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4469 input_amplifier_0/vip1 input_amplifier_0/rst vincm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4470 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4471 VDD VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4472 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4473 vampp VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X4474 adc_vcaparrayA dac_8bit_0/adc_run vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4475 dac_8bit_1/c6m sample dac_8bit_1/amux_2to1_1/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4476 a_245151_n121167# a_244617_n121161# a_245056_n121167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4477 dac_8bit_0/c6m dac_8bit_0/amux_2to1_1/SELB vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4478 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4479 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4480 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4481 vcp_sampled vcp_sampled vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4482 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4483 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4484 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4485 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4486 vampm input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vfoldm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4487 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4488 vlowA VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4489 VSS a_242526_n123369# a_242484_n122965# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4490 dac_8bit_1/amux_2to1_9/SELB q0B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4491 vlowB VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4492 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp vse peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4493 a_242506_n114759# a_242419_n114983# a_242102_n114873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4494 vlowB q3B dac_8bit_1/amux_2to1_4/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4495 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4496 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4497 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4498 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4499 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4500 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4501 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 a_275374_n146348# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4502 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/vom1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4503 input_amplifier_0/diff_fold_casc_ota_0/vcascnp input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/vop1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4504 vrefB VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4505 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4506 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/vip2 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X4507 sample_and_hold_0/vholdm vcp_sampled sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X4508 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4509 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4510 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4511 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4512 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4513 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4514 diff_to_se_converter_0/vip diff_to_se_converter_0/txgate_0/txb vfiltp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4515 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4516 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4517 a_227412_n122869# low_freq_pll_0/cs_ring_osc_0/vpbias a_226954_n122869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X4518 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4519 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4520 VSS VSS low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4521 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4522 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q a_241919_n122799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4523 VSS a_242783_n121167# a_242951_n121193# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4524 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4525 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4526 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X4527 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X4528 VDD vbiasp vcp_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X4529 vlowA VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4530 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4531 vlowB q6B dac_8bit_1/amux_2to1_1/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4532 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4533 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4534 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/vip2 input_amplifier_0/diff_fold_casc_ota_1/vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X4535 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X4536 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4537 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn2 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4538 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X4539 vrefB VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4540 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4541 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 a_356329_n164260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4542 dac_8bit_1/ibiasn dac_8bit_1/ibiasn dac_8bit_1/ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4543 vampm input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4544 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4545 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4546 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 input_amplifier_0/ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4547 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4548 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4549 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X4550 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4551 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4552 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4553 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4554 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q a_242951_n123369# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4555 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X4556 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp vse peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4557 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4558 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 vocm input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X4559 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4560 a_336955_n185409# a_336401_n185569# a_336608_n185510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4561 vcp_sampled vcp_sampled vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4562 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4563 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4564 dac_8bit_0/latched_comparator_folded_0/vcompm_buf dac_8bit_0/latched_comparator_folded_0/vcompmb VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4565 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X4566 VSS VSS dac_8bit_0/amux_2to1_9/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4567 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4568 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4569 VSS a_338149_n185569# a_338156_n185665# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4570 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4571 adc_vcaparrayB dac_8bit_1/c2m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4572 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4573 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4574 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X4575 a_228328_n122869# low_freq_pll_0/cs_ring_osc_0/vpbias low_freq_pll_0/cs_ring_osc_0/vpbias VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X4576 a_163060_n102324# input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4577 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4578 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4579 a_275374_n180872# sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4580 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4581 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4582 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn biquad_gm_c_filter_0/gm_c_stage_2/vcmcn VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4583 input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4584 VDD VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4585 VDD input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X4586 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4587 a_241188_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_241646_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X4588 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4589 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4590 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4591 biquad_gm_c_filter_0/ibiasn2 biquad_gm_c_filter_0/ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4592 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X4593 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4594 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4595 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X4596 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4597 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4598 dac_8bit_1/latched_comparator_folded_0/vlatchp adc_clk dac_8bit_1/latched_comparator_folded_0/vlatchm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X4599 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4600 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4601 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4602 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4603 a_241938_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_241480_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4604 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4605 vampp input_amplifier_0/txgate_3/txb input_amplifier_0/venp2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4606 dac_8bit_1/ibiasn dac_8bit_1/ibiasn dac_8bit_1/ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4607 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4608 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_243770_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4609 VSS VSS dac_8bit_0/amux_2to1_5/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4610 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4611 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X4612 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4613 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4614 dac_8bit_0/amux_2to1_9/Y q0A vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4615 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4616 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X4617 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4618 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4619 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4620 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4621 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4622 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4623 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4624 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4625 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_8/A a_246080_n122255# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4626 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4627 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn vintp biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4628 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4629 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X4630 vse diff_to_se_converter_0/vim sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X4631 a_275374_n146348# sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4632 dac_8bit_1/cdumm dac_8bit_1/amux_2to1_6/SELB vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4633 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4634 a_336955_n185409# a_336408_n185665# a_336608_n185510# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4635 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4636 VDD VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4637 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4638 VSS VSS input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4639 dac_8bit_0/latched_comparator_folded_0/vtailp dac_8bit_0/vcom_buf dac_8bit_0/latched_comparator_folded_0/vlatchp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4640 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4641 input_amplifier_0/venm2 input_amplifier_0/vip2 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X4642 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4643 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4644 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4645 VDD vbiasp biquad_gm_c_filter_0/ibiasn4 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X4646 vampm input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4647 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4648 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4649 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4650 input_amplifier_0/vip2 VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4651 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4652 input_amplifier_0/diff_fold_casc_ota_0/vcascnm input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4653 VDD input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X4654 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4655 vampp gain_ctrl_1 input_amplifier_0/venp2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4656 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn biquad_gm_c_filter_0/gm_c_stage_3/vcmcn VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4657 vrefB dac_8bit_1/amux_2to1_12/SELB dac_8bit_1/amux_2to1_5/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4658 vpeak_sampled vpeak_sampled VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4659 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4660 dac_8bit_1/c4m dac_8bit_1/amux_2to1_3/SELB vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4661 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 a_356329_n164260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4662 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4663 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4664 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4665 dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4666 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4667 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4668 VDD low_freq_pll_0/pfd_cp_lpf_0/vQA low_freq_pll_0/pfd_cp_lpf_0/vQAb VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4669 vlowB VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4670 dac_8bit_1/latched_comparator_folded_0/vlatchm vlowB dac_8bit_1/latched_comparator_folded_0/vtailp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4671 dac_8bit_0/vcom_buf dac_8bit_0/vcom_buf dac_8bit_0/vcom_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4672 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4673 comparator_0/vcompp comparator_0/vcompp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4674 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4675 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4676 sample_and_hold_1/vhold sample vpeak VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4677 comparator_0/ibiasn comparator_0/ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4678 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4679 VSS dac_8bit_0/latched_comparator_folded_0/vcomppb dac_8bit_0/latched_comparator_folded_0/vcompp_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4680 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 vpeak VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4681 a_230869_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin a_230411_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X4682 VDD input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X4683 a_275374_n146348# sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4684 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4685 adc_vcaparrayB dac_8bit_1/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4686 input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4687 a_237498_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_237956_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X4688 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4689 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4690 VDD vbiasp diff_to_se_converter_0/ibiasn VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X4691 VSS biquad_gm_c_filter_0/ibiasn2 biquad_gm_c_filter_0/ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4692 dac_8bit_0/amux_2to1_12/SELB q2A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4693 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4694 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4695 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4696 a_221582_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_222040_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X4697 VDD input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X4698 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4699 input_amplifier_0/diff_fold_casc_ota_1/M1d input_amplifier_0/diff_fold_casc_ota_1/M1d input_amplifier_0/diff_fold_casc_ota_1/M1d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4700 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4701 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4702 vrefB dac_8bit_1/amux_2to1_15/SELB dac_8bit_1/amux_2to1_2/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4703 input_amplifier_0/diff_fold_casc_ota_1/vcascnp input_amplifier_0/diff_fold_casc_ota_1/vbias3 vampp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4704 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4705 VSS a_245481_n121345# a_245649_n121443# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4706 input_amplifier_0/vop1 VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X4707 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4708 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4709 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 a_275374_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4710 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4711 vlowB VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4712 VSS dac_8bit_1/vcom_buf sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X4713 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4714 a_245565_n122433# a_244783_n122799# a_245481_n122433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4715 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4716 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4717 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4718 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4719 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4720 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4721 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4722 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4723 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4724 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4725 a_356329_n164260# dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4726 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/M2d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4727 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 a_189446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4728 dac_8bit_0/amux_2to1_15/SELB q5A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4729 input_amplifier_0/diff_fold_casc_ota_1/vcascnm input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4730 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4731 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_0/A a_243382_n120301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4732 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4733 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4734 a_239883_n115151# a_239708_n115125# a_240062_n115125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4735 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4736 a_236480_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_236022_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4737 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4738 input_amplifier_0/venp2 input_amplifier_0/txgate_3/txb vampp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4739 a_238770_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin a_238312_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4740 biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail2 vfiltm biquad_gm_c_filter_0/gm_c_stage_3/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4741 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4742 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4743 VSS biquad_gm_c_filter_0/ibiasn3 biquad_gm_c_filter_0/ibiasn3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4744 input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc vocm input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X4745 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4746 vlowB VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4747 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X4748 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4749 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4750 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4751 VSS vse sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X4752 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4753 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4754 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4755 VDD input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X4756 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X4757 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4758 low_freq_pll_0/cs_ring_osc_0/vosc2 low_freq_pll_0/cs_ring_osc_0/vosc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4759 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4760 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4761 a_221481_n130007# low_freq_pll_0/cs_ring_osc_0/vosc a_221023_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X4762 input_amplifier_0/diff_fold_casc_ota_0/vcascnp input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/vop1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4763 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4764 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vfoldm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4765 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4766 VDD a_242526_n123369# a_242453_n123343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4767 VSS a_337592_n185460# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_2/Q VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4768 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4769 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4770 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4771 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4772 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4773 VDD input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X4774 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4775 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4776 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4777 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4778 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4779 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4780 VSS VSS dac_8bit_0/ibiasp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=2e+06u
X4781 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4782 sample_and_hold_1/vhold VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X4783 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4784 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X4785 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn vfiltm biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4786 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4787 a_241328_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_240870_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4788 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q a_241919_n122249# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4789 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4790 VDD input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X4791 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4792 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4793 biquad_gm_c_filter_0/gm_c_stage_3/vtail_diff vintm vfiltm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4794 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4795 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4796 input_amplifier_0/vop1 VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X4797 a_223770_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin a_223312_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4798 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4799 vcp_sampled sample dac_8bit_0/cdumm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4800 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4801 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/vip2 input_amplifier_0/diff_fold_casc_ota_1/vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X4802 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4803 a_230412_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin a_229954_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4804 low_freq_pll_0/ibiasn low_freq_pll_0/ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4805 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4806 a_242358_n123343# a_241919_n123337# a_242273_n123343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4807 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_245649_n122281# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4808 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4809 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4810 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4811 dac_8bit_0/latched_comparator_folded_0/vcompp dac_8bit_0/latched_comparator_folded_0/vcompm VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4812 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4813 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4814 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X4815 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4816 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4817 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X4818 a_244954_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4819 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4820 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4821 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4822 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4823 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4824 VSS dac_8bit_1/ibiasn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4825 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4826 a_241634_n115151# a_241731_n115151# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4827 input_amplifier_0/diff_fold_casc_ota_1/vcascnp input_amplifier_0/diff_fold_casc_ota_1/vbias3 vampp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4828 adc_vcaparrayB dac_8bit_1/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4829 VDD input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vfoldm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4830 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4831 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4832 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4833 dac_8bit_0/amux_2to1_6/B dac_8bit_0/amux_2to1_11/SELB vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4834 vcp_sampled sample dac_8bit_0/c4m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4835 VDD VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4836 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4837 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4838 input_amplifier_0/diff_fold_casc_ota_1/vcascnp input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4839 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4840 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 a_356329_n164260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4841 VSS low_freq_pll_0/ibiasn low_freq_pll_0/ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4842 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4843 dac_8bit_1/latched_comparator_folded_0/vtailp vlowB dac_8bit_1/latched_comparator_folded_0/vlatchm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4844 VSS VSS input_amplifier_0/vim2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4845 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn1 vocm_filt biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4846 vampm input_amplifier_0/vip2 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X4847 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4848 dac_8bit_0/amux_2to1_7/SELB sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4849 VSS a_335749_n185813# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/Q_N VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4850 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q a_242951_n121443# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4851 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4852 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4853 biquad_gm_c_filter_0/gm_c_stage_1/vtail_diff VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4854 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4855 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X4856 a_242783_n122433# a_242085_n122799# a_242526_n122687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4857 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4858 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4859 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4860 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4861 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4862 VDD input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X4863 a_241023_n130007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X4864 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4865 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4866 a_226496_n122869# low_freq_pll_0/cs_ring_osc_0/vpbias a_226954_n122869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X4867 VSS diff_to_se_converter_0/ibiasn diff_to_se_converter_0/ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4868 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4869 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4870 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4871 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4872 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4873 dac_8bit_0/amux_2to1_3/B dac_8bit_0/amux_2to1_14/SELB vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4874 biquad_gm_c_filter_0/ibiasn1 biquad_gm_c_filter_0/ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4875 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4876 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4877 adc_vcaparrayB dac_8bit_1/c2m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4878 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4879 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4880 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4881 adc_vcaparrayA dac_8bit_0/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4882 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4883 VSS VSS sample_and_hold_0/vholdm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4884 a_232244_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin a_231786_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4885 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4886 low_freq_pll_0/pfd_cp_lpf_0/vRSTN low_freq_pll_0/pfd_cp_lpf_0/vQA a_241105_n115125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4887 a_241327_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_240869_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X4888 VDD VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4889 dac_8bit_0/amux_2to1_4/SELB sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4890 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4891 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4892 dac_8bit_1/amux_2to1_10/SELB q1B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4893 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4894 VSS VSS vlowA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4895 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/M6d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4896 VSS VSS low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4897 VDD a_335844_n185460# pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4898 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4899 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4900 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4901 a_242484_n121877# a_242085_n122249# a_242358_n122255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4902 input_amplifier_0/diff_fold_casc_ota_0/M6d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4903 vrefB VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4904 a_243312_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_242854_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4905 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4906 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4907 a_230411_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin a_229953_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X4908 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4909 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4910 a_237956_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_238414_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X4911 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4912 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4913 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4914 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4915 a_336955_n185243# a_336408_n184969# a_336608_n185269# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4916 diff_to_se_converter_0/vim vfiltm sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X4917 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4918 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4919 a_244953_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X4920 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4921 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4922 dac_8bit_0/amux_2to1_1/SELB sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4923 dac_8bit_1/amux_2to1_13/SELB q3B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4924 VSS VSS vlowA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4925 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4926 VDD a_242951_n121193# a_243382_n121167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4927 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4928 input_amplifier_0/vop1 input_amplifier_0/vop1 input_amplifier_0/vop1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4929 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4930 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/diff_fold_casc_ota_0/vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X4931 vrefB VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4932 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4933 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4934 input_amplifier_0/venm2 gain_ctrl_1 vampm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4935 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4936 input_amplifier_0/diff_fold_casc_ota_1/M2d input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/M3d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4937 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4938 VDD vbiasp peak_detector_0/ibiasn1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X4939 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4940 dac_8bit_0/latched_comparator_folded_0/vlatchp adc_clk dac_8bit_0/latched_comparator_folded_0/vlatchm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X4941 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4942 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4943 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4944 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4945 a_228478_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_228020_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X4946 vintp VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4947 VDD VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4948 VDD input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/M6d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4949 dac_8bit_1/amux_2to1_16/SELB q6B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4950 a_246328_n134960# vcp a_245870_n134960# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4951 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4952 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4953 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4954 a_242104_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_241646_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X4955 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4956 input_amplifier_0/diff_fold_casc_ota_1/M6d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4957 a_337592_n185460# a_337864_n185555# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4958 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4959 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4960 VSS input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4961 comparator_0/vo1 comparator_0/vcompp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4962 dac_8bit_0/amux_2to1_11/SELB VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4963 dac_8bit_1/amux_2to1_0/SELB sample VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4964 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4965 VSS VSS dac_8bit_0/amux_2to1_7/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4966 a_336537_n185409# a_336408_n185665# a_336116_n185555# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4967 sample_and_hold_1/vholdm sample vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4968 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4969 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4970 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X4971 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4972 a_232243_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin a_231785_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X4973 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q a_241919_n122799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4974 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 vampp input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X4975 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4976 VSS peak_detector_0/ibiasn1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4977 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4978 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4979 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4980 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4981 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4982 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4983 a_275374_n146348# sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4984 vpeak_sampled sample dac_8bit_1/c0m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4985 a_221582_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X4986 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4987 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4988 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4989 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X4990 VSS VSS biquad_gm_c_filter_0/gm_c_stage_3/vtail_diff VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4991 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4992 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4993 dac_8bit_0/amux_2to1_0/B VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4994 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4995 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4996 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4997 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 a_230446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4998 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4999 dac_8bit_0/amux_2to1_14/SELB q4A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5000 vampp input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5001 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5002 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5003 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5004 VSS VSS dac_8bit_0/amux_2to1_4/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5005 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X5006 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/csinvn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X5007 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/diff_fold_casc_ota_1/vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X5008 adc_vcaparrayA dac_8bit_0/c3m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5009 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5010 dac_8bit_0/amux_2to1_7/B q1A vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5011 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5012 input_amplifier_0/diff_fold_casc_ota_1/M2d input_amplifier_0/diff_fold_casc_ota_1/M2d input_amplifier_0/diff_fold_casc_ota_1/M2d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5013 comparator_0/ibiasn comparator_0/ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X5014 dac_8bit_1/latched_comparator_folded_0/vlatchp VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5015 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5016 a_238465_n122049# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout a_238007_n122049# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X5017 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5018 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5019 a_335749_n185269# a_335844_n185269# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5020 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5021 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 a_275374_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5022 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5023 vampm VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X5024 diff_to_se_converter_0/vim vfiltm sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X5025 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5026 input_amplifier_0/vip2 input_amplifier_0/txgate_0/txb input_amplifier_0/venm1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5027 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X5028 dac_8bit_1/amux_2to1_9/Y dac_8bit_1/amux_2to1_9/SELB vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5029 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5030 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5031 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5032 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5033 dac_8bit_1/c2m dac_8bit_1/amux_2to1_5/SELB vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5034 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5035 vcp_sampled VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5036 a_356329_n164260# dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5037 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5038 adc_vcaparrayA VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5039 VSS input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5040 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5041 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5042 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5043 VDD a_242526_n122687# a_242453_n122433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5044 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5045 input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5046 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5047 a_356329_n113250# dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5048 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/csinvp VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X5049 VSS VSS dac_8bit_0/amux_2to1_1/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5050 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5051 a_237855_n130007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin a_237397_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X5052 comparator_0/vcompm comparator_0/vcompm VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5053 a_336608_n185269# a_336408_n184969# a_336757_n185243# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5054 dac_8bit_0/amux_2to1_4/B q3A vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5055 VDD vbiasp comparator_0/ibiasn VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X5056 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5057 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5058 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5059 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5060 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5061 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn vfiltp biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5062 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5063 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5064 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5065 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5066 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5067 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5068 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5069 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5070 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5071 dac_8bit_1/c5m dac_8bit_1/amux_2to1_2/SELB vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5072 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5073 vlowB dac_8bit_1/adc_run adc_vcaparrayB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5074 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5075 input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc vocm input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X5076 a_162668_n147576# diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5077 dac_8bit_1/amux_2to1_6/SELB sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5078 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5079 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5080 VDD VDD dac_8bit_0/latched_comparator_folded_0/vlatchp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5081 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5082 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5083 dac_8bit_0/amux_2to1_1/B q6A vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5084 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5085 a_222396_n150168# vcp a_221938_n150168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X5086 a_162668_n147576# diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5087 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 vse VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5088 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5089 adc_vcaparrayB dac_8bit_1/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5090 VSS input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5091 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5092 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5093 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5094 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5095 a_230446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5096 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5097 a_222855_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin a_222397_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X5098 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn2 vocm_filt biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5099 vrefA VSS dac_8bit_0/amux_2to1_6/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5100 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 vse VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5101 dac_8bit_1/amux_2to1_3/SELB sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5102 vincm input_amplifier_0/rst input_amplifier_0/vim1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5103 vampp input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5104 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5105 VDD dac_8bit_1/latched_comparator_folded_0/vcompp dac_8bit_1/latched_comparator_folded_0/vcomppb VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5106 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5107 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5108 peak_detector_0/vpeak peak_detector_rst VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5109 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 a_189446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5110 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5111 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5112 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5113 adc_vcaparrayA dac_8bit_0/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5114 a_237397_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_236939_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X5115 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X5116 dac_8bit_1/ibiasp VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=2e+06u
X5117 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5118 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5119 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5120 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5121 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5122 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5123 dac_8bit_1/latched_comparator_folded_0/vlatchp adc_clk dac_8bit_1/latched_comparator_folded_0/vlatchm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X5124 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5125 a_189446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5126 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X5127 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5128 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5129 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 vpeak VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5130 dac_8bit_0/c0m sample vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5131 input_amplifier_0/diff_fold_casc_ota_0/M1d input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5132 VSS a_242419_n114983# a_242380_n114857# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5133 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5134 VDD dac_8bit_1/comp_outm adc_compB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5135 a_242783_n121167# a_241919_n121161# a_242526_n121193# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5136 a_226481_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_226023_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X5137 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X5138 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5139 a_228771_n130007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_228313_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X5140 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5141 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5142 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5143 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5144 vrefA q4A dac_8bit_0/amux_2to1_3/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5145 a_242909_n120789# a_241919_n121161# a_242783_n121167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5146 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5147 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5148 biquad_gm_c_filter_0/gm_c_stage_2/vcmc VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5149 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5150 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5151 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X5152 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5153 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5154 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5155 dac_8bit_1/amux_2to1_9/SELB q0B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5156 VSS pulse_generator_0/sky130_fd_sc_hd__inv_1_0/Y a_338703_n185243# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5157 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5158 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 vampm input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X5159 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5160 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5161 a_356329_n164260# dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5162 VSS vcp_sampled sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X5163 dac_8bit_0/amux_2to1_6/B dac_8bit_0/amux_2to1_6/SELB dac_8bit_0/cdumm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5164 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5165 VDD VDD vpeak VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5166 a_338703_n185243# a_338149_n185269# a_338356_n185269# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5167 dac_8bit_1/vcom_buf dac_8bit_1/vcom_buf dac_8bit_1/vcom_buf VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5168 VSS VSS biquad_gm_c_filter_0/gm_c_stage_3/vbiasp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X5169 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5170 VDD a_245649_n123369# a_246080_n123343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5171 a_239405_n115125# a_239361_n114883# a_239239_n115125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5172 input_amplifier_0/diff_fold_casc_ota_1/vcascnp input_amplifier_0/diff_fold_casc_ota_1/vbias3 vampp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5173 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5174 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5175 dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5176 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 a_356329_n164260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5177 input_amplifier_0/diff_fold_casc_ota_0/vcascnm input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/vom1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5178 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5179 a_242273_n121167# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5180 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5181 dac_8bit_0/latched_comparator_folded_0/vcompm dac_8bit_0/latched_comparator_folded_0/vcompp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5182 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5183 dac_8bit_1/latched_comparator_folded_0/vcompp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5184 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5185 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5186 vpeak_sampled dac_8bit_1/amux_2to1_0/SELB dac_8bit_1/c7m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5187 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5188 dac_8bit_0/amux_2to1_0/B sample dac_8bit_0/c7m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5189 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5190 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5191 VSS biquad_gm_c_filter_0/gm_c_stage_1/vcmc biquad_gm_c_filter_0/gm_c_stage_1/vcmc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X5192 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5193 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5194 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5195 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5196 vcp_sampled sample dac_8bit_0/c2m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5197 VDD vbiasp peak_detector_0/ibiasn2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X5198 VDD a_337497_n185813# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/D VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5199 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5200 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5201 VSS VSS dac_8bit_1/amux_2to1_6/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5202 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 a_162668_n147576# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5203 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X5204 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5205 diff_to_se_converter_0/ibiasn diff_to_se_converter_0/ibiasn diff_to_se_converter_0/ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5206 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5207 dac_8bit_0/amux_2to1_3/B dac_8bit_0/amux_2to1_3/SELB dac_8bit_0/c4m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5208 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5209 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5210 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5211 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5212 VDD adc_clk dac_8bit_1/latched_comparator_folded_0/vcompm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5213 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5214 dac_8bit_1/c7m sample dac_8bit_1/amux_2to1_0/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5215 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5216 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5217 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5218 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 a_162668_n147576# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5219 VDD vbiasp vpeak_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X5220 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/vcom_buf VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5221 VDD dac_8bit_0/latched_comparator_folded_0/vcompm dac_8bit_0/latched_comparator_folded_0/vcompp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5222 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5223 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5224 biquad_gm_c_filter_0/gm_c_stage_3/vcmc VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5225 VDD VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5226 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5227 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5228 dac_8bit_0/amux_2to1_5/B dac_8bit_0/amux_2to1_12/SELB vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5229 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5230 vcp_sampled sample dac_8bit_0/c5m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5231 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5232 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5233 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5234 VSS VSS dac_8bit_1/amux_2to1_3/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5235 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5236 a_336757_n185421# a_336537_n185409# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5237 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5238 VDD VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5239 dac_8bit_1/amux_2to1_6/B VSS vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5240 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5241 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5242 a_228020_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_228478_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X5243 dac_8bit_0/amux_2to1_0/B dac_8bit_0/amux_2to1_0/SELB dac_8bit_0/c7m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5244 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5245 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5246 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5247 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/vip2 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X5248 dac_8bit_0/latched_comparator_folded_0/vlatchm dac_8bit_0/latched_comparator_folded_0/vlatchp VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X5249 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5250 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5251 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5252 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5253 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5254 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5255 a_356329_n113250# dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5256 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5257 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5258 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5259 a_242358_n122433# a_241919_n122799# a_242273_n122799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5260 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5261 a_223414_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_222956_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X5262 comparator_0/vcompm comparator_0/vcompm comparator_0/vcompm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5263 VDD VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5264 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5265 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X5266 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5267 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5268 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5269 a_242273_n122799# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5270 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5271 dac_8bit_0/amux_2to1_2/B dac_8bit_0/amux_2to1_15/SELB vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5272 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 vampp input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X5273 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5274 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5275 VSS VSS dac_8bit_1/amux_2to1_0/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5276 diff_to_se_converter_0/ibiasn diff_to_se_converter_0/ibiasn diff_to_se_converter_0/ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5277 a_336336_n185243# a_335844_n185269# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5278 dac_8bit_1/amux_2to1_3/B q4B vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5279 low_freq_pll_0/ibiasn vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X5280 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5281 a_237956_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_237498_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X5282 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5283 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5284 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_5/A a_243382_n123343# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5285 VSS VSS vlowA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5286 VSS VSS input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5287 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5288 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5289 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5290 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5291 vampm input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vfoldm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5292 input_amplifier_0/txgate_2/txb gain_ctrl_1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5293 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5294 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X5295 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 a_230446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5296 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5297 vcp VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5298 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5299 VDD dac_8bit_0/latched_comparator_folded_0/vcompm dac_8bit_0/latched_comparator_folded_0/vcompp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5300 vincm VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5301 a_236938_n150168# vcp a_236480_n150168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X5302 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5303 vrefB q0B dac_8bit_1/amux_2to1_9/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5304 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5305 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X5306 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5307 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5308 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5309 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5310 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5311 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5312 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X5313 vcp sample sample_and_hold_0/vhold VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5314 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X5315 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5316 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5317 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5318 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5319 VSS peak_detector_0/ibiasn1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5320 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5321 input_amplifier_0/ibiasn1 input_amplifier_0/ibiasn1 input_amplifier_0/ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5322 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5323 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5324 VSS VSS vlowA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5325 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5326 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5327 VDD biquad_gm_c_filter_0/gm_c_stage_0/vcmcn biquad_gm_c_filter_0/gm_c_stage_0/vcmc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5328 VSS vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5329 biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail1 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X5330 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_10/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5331 a_224330_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X5332 a_242453_n123343# a_241919_n123337# a_242358_n123343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5333 VSS VSS vincm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5334 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X5335 biquad_gm_c_filter_0/gm_c_stage_2/vbiasp biquad_gm_c_filter_0/ibiasn4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X5336 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vfoldp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5337 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5338 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn2 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5339 input_amplifier_0/vom1 VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X5340 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5341 low_freq_pll_0/freq_div_0/vin low_freq_pll_0/cs_ring_osc_0/vosc2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5342 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5343 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5344 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_6/A a_246080_n121167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5345 VSS vcp a_223770_n150168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X5346 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5347 VDD a_338149_n185569# a_338156_n185665# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5348 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5349 VSS VSS vlowA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5350 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5351 dac_8bit_1/amux_2to1_9/Y dac_8bit_1/amux_2to1_8/SELB dac_8bit_1/c0m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5352 a_239870_n114759# a_238793_n115125# a_239708_n115125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5353 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5354 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5355 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X5356 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5357 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5358 a_236174_n119618# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X5359 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5360 dac_8bit_0/amux_2to1_12/SELB q2A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5361 VDD VDD dac_8bit_1/vcom_buf VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5362 VDD low_freq_pll_0/pfd_cp_lpf_0/vpdiode low_freq_pll_0/pfd_cp_lpf_0/vpdiode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5363 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5364 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5365 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X5366 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5367 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5368 adc_vcaparrayB dac_8bit_1/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5369 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 a_189446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5370 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5371 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5372 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5373 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5374 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1.2e+07u w=2e+06u
X5375 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5376 input_amplifier_0/diff_fold_casc_ota_1/vcascnm input_amplifier_0/diff_fold_casc_ota_1/vbias3 vampm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5377 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5378 a_245481_n123343# a_244617_n123337# a_245224_n123369# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5379 vpeak_sampled sample dac_8bit_1/c1m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5380 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5381 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5382 input_amplifier_0/diff_fold_casc_ota_1/vcascnm input_amplifier_0/diff_fold_casc_ota_1/vbias3 vampm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5383 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5384 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_238771_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X5385 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5386 input_amplifier_0/txgate_2/txb gain_ctrl_1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5387 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5388 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5389 dac_8bit_1/amux_2to1_5/B dac_8bit_1/amux_2to1_5/SELB dac_8bit_1/c2m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5390 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5391 a_245607_n122965# a_244617_n123337# a_245481_n123343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5392 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5393 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5394 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5395 input_amplifier_0/vom1 input_amplifier_0/vom1 input_amplifier_0/vom1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5396 VDD biquad_gm_c_filter_0/gm_c_stage_1/vcmcn biquad_gm_c_filter_0/gm_c_stage_1/vcmc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5397 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5398 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/vim2 input_amplifier_0/diff_fold_casc_ota_1/vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X5399 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5400 a_230446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5401 VSS peak_detector_0/ibiasn2 peak_detector_0/ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5402 dac_8bit_0/amux_2to1_15/SELB q5A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5403 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5404 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5405 VDD input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vfoldp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5406 a_230446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5407 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5408 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5409 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5410 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X5411 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5412 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5413 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5414 a_242783_n120257# a_241919_n120623# a_242526_n120511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5415 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5416 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5417 dac_8bit_0/amux_2to1_0/B q7A vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5418 VSS biquad_gm_c_filter_0/ibiasn3 biquad_gm_c_filter_0/ibiasn3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X5419 dac_8bit_1/amux_2to1_7/B dac_8bit_1/amux_2to1_10/SELB vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5420 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5421 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5422 vpeak_sampled sample dac_8bit_1/c3m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5423 dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5424 dac_8bit_1/latched_comparator_folded_0/vtailp dac_8bit_1/vcom_buf dac_8bit_1/latched_comparator_folded_0/vlatchp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5425 a_275374_n180872# sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5426 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X5427 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5428 VSS VSS input_amplifier_0/vip2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5429 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5430 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5431 VSS VSS vfiltm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5432 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5433 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5434 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5435 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5436 dac_8bit_0/vcom_buf VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X5437 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5438 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5439 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_9/A a_246080_n122477# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5440 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5441 VSS vbiasn dac_8bit_0/ibiasp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=2e+06u
X5442 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5443 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5444 dac_8bit_1/latched_comparator_folded_0/vlatchp dac_8bit_1/latched_comparator_folded_0/vlatchm VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X5445 dac_8bit_0/amux_2to1_9/Y q0A vrefA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5446 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5447 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5448 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5449 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5450 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5451 adc_vcaparrayB dac_8bit_1/c2m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5452 a_226954_n122869# low_freq_pll_0/cs_ring_osc_0/vpbias a_226496_n122869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X5453 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5454 peak_detector_0/verr peak_detector_0/verr peak_detector_0/verr VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5455 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5456 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5457 VDD comparator_0/vcompm comparator_0/vcompm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5458 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X5459 a_242273_n120623# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5460 VSS a_245649_n121443# a_246080_n121389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5461 dac_8bit_1/amux_2to1_4/B dac_8bit_1/amux_2to1_13/SELB vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5462 vpeak_sampled sample dac_8bit_1/c6m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5463 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5464 input_amplifier_0/diff_fold_casc_ota_1/vcascnp input_amplifier_0/diff_fold_casc_ota_1/vbias3 vampp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5465 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5466 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5467 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5468 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5469 vcp_sampled vcp_sampled VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5470 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/M1d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5471 VSS dac_8bit_1/vcom_buf sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X5472 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5473 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 a_217060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5474 VDD a_335749_n185269# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5475 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5476 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5477 VSS biquad_gm_c_filter_0/ibiasn1 biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X5478 dac_8bit_1/amux_2to1_5/SELB sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5479 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5480 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5481 input_amplifier_0/vim1 vincm sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X5482 VSS sample dac_8bit_1/adc_run VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5483 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5484 vlowA dac_8bit_0/amux_2to1_11/SELB dac_8bit_0/amux_2to1_6/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5485 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5486 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5487 a_275374_n146348# sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5488 input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vfoldp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5489 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5490 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5491 a_241938_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_241480_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X5492 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5493 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5494 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5495 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5496 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5497 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5498 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5499 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5500 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5501 dac_8bit_1/amux_2to1_1/B dac_8bit_1/amux_2to1_16/SELB vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5502 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5503 input_amplifier_0/diff_fold_casc_ota_0/vcascnp input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/vop1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5504 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5505 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5506 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5507 a_244783_n121711# a_244617_n121711# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5508 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/vip2 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X5509 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5510 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5511 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5512 vrefA q2A dac_8bit_0/amux_2to1_5/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5513 dac_8bit_1/amux_2to1_2/SELB sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5514 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 a_356329_n113250# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5515 input_amplifier_0/diff_fold_casc_ota_1/vcascnm input_amplifier_0/diff_fold_casc_ota_1/vbias3 vampm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5516 VDD a_242783_n123343# a_242951_n123369# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5517 a_244783_n121711# a_244617_n121711# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5518 VSS VSS vlowB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5519 VDD vbiasp peak_detector_0/ibiasn2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X5520 vlowA dac_8bit_0/amux_2to1_14/SELB dac_8bit_0/amux_2to1_3/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5521 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5522 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5523 vcp_sampled sample sample_and_hold_0/vholdm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5524 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5525 sample_and_hold_1/vhold VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X5526 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5527 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 vpeak_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5528 input_amplifier_0/diff_fold_casc_ota_1/M2d input_amplifier_0/diff_fold_casc_ota_1/M2d input_amplifier_0/diff_fold_casc_ota_1/M2d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5529 input_amplifier_0/vip1 input_amplifier_0/txgate_5/txb vincm VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5530 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5531 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5532 input_amplifier_0/venp2 gain_ctrl_1 vampp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5533 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5534 a_226188_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_226646_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X5535 a_239361_n114883# a_239143_n115125# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5536 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5537 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5538 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5539 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5540 dac_8bit_0/c1m sample vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5541 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5542 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5543 VDD input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/M1d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5544 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X5545 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5546 a_356329_n113250# dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5547 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5548 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 a_163060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5549 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5550 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_9/A a_246080_n122477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5551 input_amplifier_0/venm1 input_amplifier_0/vom1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X5552 a_242273_n122255# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5553 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5554 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5555 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5556 vrefA q5A dac_8bit_0/amux_2to1_2/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5557 VDD low_freq_pll_0/pfd_cp_lpf_0/vpbias low_freq_pll_0/pfd_cp_lpf_0/vswitchh VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X5558 VSS VSS vlowB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5559 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5560 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5561 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5562 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5563 a_242506_n114759# a_242380_n114857# a_242102_n114873# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5564 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5565 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5566 vlowA dac_8bit_0/amux_2to1_17/SELB dac_8bit_0/amux_2to1_0/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5567 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5568 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5569 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5570 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5571 a_356329_n113250# dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5572 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5573 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5574 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5575 dac_8bit_1/amux_2to1_10/SELB q1B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5576 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5577 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5578 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5579 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5580 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5581 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5582 input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vbias3 a_163060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5583 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X5584 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5585 VSS input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5586 a_239330_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_238872_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X5587 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5588 dac_8bit_0/c3m sample vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5589 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5590 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5591 a_275374_n146348# sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5592 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5593 a_338285_n185243# a_338156_n184969# a_337864_n185269# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5594 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5595 a_189446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5596 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5597 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5598 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5599 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5600 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 vse VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5601 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5602 a_338084_n185421# a_337592_n185460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5603 VSS VSS vlowB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5604 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5605 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5606 a_238312_n150168# vcp a_237854_n150168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X5607 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5608 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5609 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5610 adc_vcaparrayA dac_8bit_0/c3m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5611 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5612 vintp vampp biquad_gm_c_filter_0/gm_c_stage_0/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5613 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5614 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X5615 VSS a_242951_n121443# a_242909_n121711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5616 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5617 dac_8bit_1/amux_2to1_13/SELB q3B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5618 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 a_230446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5619 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5620 biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail1 vocm_filt biquad_gm_c_filter_0/gm_c_stage_1/vcmcn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5621 vampm VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X5622 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5623 dac_8bit_0/amux_2to1_2/B dac_8bit_0/amux_2to1_2/SELB dac_8bit_0/c5m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5624 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5625 input_amplifier_0/diff_fold_casc_ota_0/vfoldp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5626 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X5627 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn vse peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5628 a_356329_n164260# dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5629 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5630 dac_8bit_0/c6m sample vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5631 VDD VDD input_amplifier_0/diff_fold_casc_ota_0/vfoldp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5632 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5633 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5634 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5635 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5636 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X5637 VSS VSS low_freq_pll_0/ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X5638 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5639 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5640 dac_8bit_0/latched_comparator_folded_0/vlatchp dac_8bit_0/vcom_buf dac_8bit_0/latched_comparator_folded_0/vtailp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5641 a_236480_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin a_236022_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X5642 a_242453_n122433# a_241919_n122799# a_242358_n122433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5643 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_245649_n122531# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5644 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5645 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5646 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5647 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5648 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5649 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5650 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5651 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5652 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5653 dac_8bit_1/amux_2to1_16/SELB q6B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5654 a_238006_n119618# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout a_237548_n119618# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X5655 VSS VSS dac_8bit_1/amux_2to1_2/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5656 VDD input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X5657 dac_8bit_1/amux_2to1_5/B q2B vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5658 VDD VDD input_amplifier_0/vop1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5659 dac_8bit_0/latched_comparator_folded_0/vtailp vlowA dac_8bit_0/latched_comparator_folded_0/vlatchm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5660 vse diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5661 comparator_0/ibiasn comparator_0/ibiasn comparator_0/ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X5662 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5663 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5664 input_amplifier_0/venp2 input_amplifier_0/vim2 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X5665 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5666 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5667 a_217060_n102324# input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5668 VSS a_245649_n123369# a_245607_n122965# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5669 input_amplifier_0/venp2 input_amplifier_0/vim2 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X5670 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5671 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5672 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5673 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5674 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5675 biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail1 vfiltp biquad_gm_c_filter_0/gm_c_stage_3/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5676 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5677 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5678 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5679 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_7/A a_246080_n121389# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5680 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5681 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5682 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X5683 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5684 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5685 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5686 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5687 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X5688 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5689 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5690 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5691 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5692 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5693 a_245481_n122433# a_244617_n122799# a_245224_n122687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5694 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5695 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5696 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/verr VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5697 vlowB dac_8bit_1/amux_2to1_9/SELB dac_8bit_1/amux_2to1_9/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5698 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5699 dac_8bit_1/latched_comparator_folded_0/vlatchp dac_8bit_1/vcom_buf dac_8bit_1/latched_comparator_folded_0/vtailp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5700 a_221480_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin a_221022_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X5701 adc_vcaparrayB dac_8bit_1/c2m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5702 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 a_275374_n146348# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5703 a_223770_n131500# low_freq_pll_0/cs_ring_osc_0/vosc a_223312_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X5704 VSS input_amplifier_0/ibiasn2 input_amplifier_0/ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5705 dac_8bit_1/amux_2to1_2/B q5B vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5706 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5707 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5708 a_230446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5709 VSS a_245224_n122687# a_245182_n122799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5710 input_amplifier_0/diff_fold_casc_ota_0/M1d input_amplifier_0/diff_fold_casc_ota_0/M1d input_amplifier_0/diff_fold_casc_ota_0/M1d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5711 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5712 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5713 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5714 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5715 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5716 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5717 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5718 dac_8bit_0/latched_comparator_folded_0/vlatchm adc_clk dac_8bit_0/latched_comparator_folded_0/vlatchp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X5719 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5720 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5721 VDD VDD biquad_gm_c_filter_0/gm_c_stage_0/vcmcn VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5722 a_275374_n180872# sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5723 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5724 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5725 vrefB q1B dac_8bit_1/amux_2to1_7/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5726 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5727 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5728 adc_vcaparrayA dac_8bit_0/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5729 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5730 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5731 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5732 VDD input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X5733 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5734 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5735 vlowB dac_8bit_1/amux_2to1_12/SELB dac_8bit_1/amux_2to1_5/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5736 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5737 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5738 VDD sample pulse_generator_0/sky130_fd_sc_hd__inv_1_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5739 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5740 a_162668_n147576# diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5741 biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail2 vocm_filt biquad_gm_c_filter_0/gm_c_stage_1/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5742 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5743 VDD VDD low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X5744 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5745 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5746 VDD VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5747 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn vse peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5748 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5749 a_163060_n102324# input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5750 biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail2 biquad_gm_c_filter_0/ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X5751 vampp input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vfoldp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5752 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5753 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5754 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/vim2 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X5755 input_amplifier_0/txgate_6/txb input_amplifier_0/rst VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5756 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5757 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/vim1 input_amplifier_0/diff_fold_casc_ota_0/vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X5758 dac_8bit_0/ibiasp vbiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=2e+06u
X5759 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/vop1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5760 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5761 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5762 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5763 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5764 sample_and_hold_0/vhold VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X5765 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5766 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X5767 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5768 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5769 vrefB q3B dac_8bit_1/amux_2to1_4/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5770 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5771 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 vpeak_sampled VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5772 dac_8bit_0/amux_2to1_9/Y VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5773 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5774 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5775 VSS a_245649_n121193# a_246080_n121167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5776 VDD input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X5777 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5778 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5779 a_230446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5780 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5781 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5782 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X5783 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X5784 vampp VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X5785 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5786 VDD VDD vintm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5787 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X5788 a_275374_n180872# sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5789 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5790 biquad_gm_c_filter_0/gm_c_stage_2/vcmc VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X5791 dac_8bit_1/amux_2to1_7/B dac_8bit_1/amux_2to1_7/SELB dac_8bit_1/c1m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5792 VSS a_245481_n122255# a_245649_n122281# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5793 a_242526_n122281# a_242358_n122255# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5794 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5795 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5796 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5797 low_freq_pll_0/ibiasn low_freq_pll_0/ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X5798 dac_8bit_1/cdumm sample vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5799 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5800 VSS VSS low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X5801 vfiltm VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5802 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5803 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5804 dac_8bit_0/cdumm dac_8bit_0/amux_2to1_6/SELB dac_8bit_0/amux_2to1_6/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5805 VDD VDD biquad_gm_c_filter_0/gm_c_stage_1/vcmcn VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5806 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5807 a_217060_n102324# input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5808 vrefB q6B dac_8bit_1/amux_2to1_1/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5809 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 vcp_sampled VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5810 a_241022_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X5811 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X5812 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5813 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5814 a_243312_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_242854_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X5815 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn vse peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5816 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5817 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5818 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5819 vpeak_sampled VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X5820 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5821 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5822 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_1/A a_243382_n121167# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5823 VDD dac_8bit_0/latched_comparator_folded_0/vcompp dac_8bit_0/latched_comparator_folded_0/vcompm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5824 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5825 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5826 a_244783_n121161# a_244617_n121161# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5827 input_amplifier_0/vom1 VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5828 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5829 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 a_163060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5830 dac_8bit_1/amux_2to1_4/B dac_8bit_1/amux_2to1_4/SELB dac_8bit_1/c3m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5831 VSS VSS input_amplifier_0/vom1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5832 vrefA dac_8bit_0/amux_2to1_17/SELB dac_8bit_0/amux_2to1_0/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5833 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5834 dac_8bit_1/c4m sample vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5835 VSS a_242783_n121345# a_242951_n121443# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5836 low_freq_pll_0/pfd_cp_lpf_0/VQBb low_freq_pll_0/pfd_cp_lpf_0/vQB VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5837 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5838 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5839 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5840 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5841 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5842 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5843 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5844 dac_8bit_0/c4m dac_8bit_0/amux_2to1_3/SELB dac_8bit_0/amux_2to1_3/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5845 VDD input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X5846 VDD low_freq_pll_0/pfd_cp_lpf_0/vpbias low_freq_pll_0/pfd_cp_lpf_0/vpbias VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X5847 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 vpeak_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5848 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5849 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5850 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X5851 a_242358_n122255# a_242085_n122249# a_242273_n122255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5852 input_amplifier_0/diff_fold_casc_ota_1/vcascnm input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5853 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5854 input_amplifier_0/vim2 gain_ctrl_0 input_amplifier_0/venp1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5855 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5856 vpeak_sampled VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5857 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5858 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5859 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5860 a_242484_n121711# a_242085_n121711# a_242358_n121345# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5861 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/vcom_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5862 a_336401_n185269# adc_clk VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5863 input_amplifier_0/txgate_4/txb input_amplifier_0/rst VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5864 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5865 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5866 a_238770_n132168# vcp a_238312_n132168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X5867 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5868 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5869 dac_8bit_1/amux_2to1_0/B dac_8bit_1/amux_2to1_17/SELB vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5870 VSS input_amplifier_0/diff_fold_casc_ota_0/M13d input_amplifier_0/diff_fold_casc_ota_0/M13d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5871 VDD comparator_0/vcompp comparator_0/vcompp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5872 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5873 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X5874 VDD VDD vfiltm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5875 VDD low_freq_pll_0/pfd_cp_lpf_0/vRSTN a_241731_n115151# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5876 dac_8bit_1/amux_2to1_1/B dac_8bit_1/amux_2to1_1/SELB dac_8bit_1/c6m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5877 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5878 a_189446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5879 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5880 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5881 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5882 a_241105_n115125# low_freq_pll_0/pfd_cp_lpf_0/vQB VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5883 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_6/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5884 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn vse peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5885 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5886 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5887 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X5888 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5889 a_222040_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_222498_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X5890 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5891 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5892 dac_8bit_0/amux_2to1_7/B q1A vrefA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5893 VDD input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X5894 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5895 a_245607_n122799# a_244617_n122799# a_245481_n122433# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5896 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5897 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5898 a_338703_n185409# a_338156_n185665# a_338356_n185510# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5899 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5900 sample_and_hold_0/vholdm sample vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5901 a_238414_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_238872_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X5902 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5903 comparator_0/vcompm comparator_0/vcompm comparator_0/vcompm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5904 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5905 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5906 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X5907 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5908 VSS dac_8bit_0/vcom_buf sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X5909 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5910 a_245224_n122281# a_245056_n122255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X5911 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5912 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5913 biquad_gm_c_filter_0/ibiasn4 biquad_gm_c_filter_0/ibiasn4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X5914 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5915 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5916 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5917 VSS a_242951_n121193# a_242909_n120789# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5918 input_amplifier_0/txgate_3/txb gain_ctrl_1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5919 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5920 dac_8bit_1/comp_outm adc_compB VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5921 a_245224_n121599# a_245056_n121345# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5922 a_245481_n122255# a_244783_n122249# a_245224_n122281# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5923 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5924 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5925 dac_8bit_0/amux_2to1_4/B q3A vrefA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5926 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 a_162668_n147576# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5927 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5928 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X5929 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 a_230446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5930 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5931 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5932 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5933 VSS VSS sample_and_hold_0/vholdm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5934 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5935 adc_vcaparrayA dac_8bit_0/cdumm sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5936 peak_detector_0/vpeak VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X5937 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5938 a_231328_n134960# vcp a_230870_n134960# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X5939 a_356329_n113250# dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5940 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5941 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5942 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5943 a_217060_n102324# input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5944 peak_detector_0/verr peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5945 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q a_242951_n122281# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5946 VSS VSS biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X5947 VDD vbiasp low_freq_pll_0/ibiasn VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X5948 dac_8bit_1/latched_comparator_folded_0/vcompmb dac_8bit_1/latched_comparator_folded_0/vcompm VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5949 a_275374_n146348# sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5950 VSS low_freq_pll_0/pfd_cp_lpf_0/vRSTN a_239405_n115125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5951 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5952 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X5953 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5954 VSS a_242526_n120511# a_242484_n120623# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5955 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5956 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5957 a_356329_n164260# dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5958 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5959 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5960 vlowA dac_8bit_0/amux_2to1_15/SELB dac_8bit_0/amux_2to1_2/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5961 VDD input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X5962 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5963 diff_to_se_converter_0/txgate_0/txb diff_to_se_converter_0/rst VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5964 a_338149_n185269# adc_clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5965 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5966 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5967 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5968 dac_8bit_0/amux_2to1_1/B q6A vrefA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5969 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5970 VDD a_337592_n185460# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_2/Q VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5971 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/csinvp VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X5972 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5973 VDD VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5974 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5975 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5976 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5977 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5978 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5979 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5980 vfiltm diff_to_se_converter_0/rst diff_to_se_converter_0/vim VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5981 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5982 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5983 input_amplifier_0/diff_fold_casc_ota_0/M1d input_amplifier_0/diff_fold_casc_ota_0/M1d input_amplifier_0/diff_fold_casc_ota_0/M1d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5984 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn vse peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5985 a_226786_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_226328_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X5986 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X5987 VDD comparator_0/vcompm comparator_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5988 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5989 a_356329_n164260# dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5990 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5991 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5992 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5993 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X5994 vampm input_amplifier_0/txgate_2/txb input_amplifier_0/venm2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5995 input_amplifier_0/diff_fold_casc_ota_1/vcascnm input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5996 VSS VSS vlowB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5997 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5998 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5999 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/vim2 input_amplifier_0/diff_fold_casc_ota_1/vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X6000 VDD VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6001 VDD input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X6002 comparator_0/vo1 comparator_0/vo1 comparator_0/vo1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6003 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6004 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6005 VSS biquad_gm_c_filter_0/gm_c_stage_3/vcmc biquad_gm_c_filter_0/gm_c_stage_3/vtail_diff VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X6006 vpeak_sampled vpeak_sampled vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6007 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6008 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6009 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6010 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6011 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6012 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6013 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6014 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6015 a_237854_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_237396_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6016 adc_vcaparrayB dac_8bit_1/c1m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6017 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6018 dac_8bit_1/c0m dac_8bit_1/amux_2to1_8/SELB dac_8bit_1/amux_2to1_9/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6019 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 a_275374_n146348# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6020 VSS input_amplifier_0/ibiasn2 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6021 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6022 VSS a_245224_n122281# a_245182_n121877# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6023 VDD VDD vpeak_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6024 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn vintm biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6025 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6026 a_238793_n115125# a_238627_n115125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6027 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6028 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6029 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1.2e+07u w=2e+06u
X6030 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6031 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6032 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn1 vocm_filt biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6033 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X6034 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6035 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/csinvp VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X6036 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X6037 a_222855_n130007# low_freq_pll_0/cs_ring_osc_0/vosc a_222397_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X6038 input_amplifier_0/txgate_3/txb gain_ctrl_1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6039 input_amplifier_0/diff_fold_casc_ota_0/vcascnm input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6040 low_freq_pll_0/pfd_cp_lpf_0/vpdiode low_freq_pll_0/pfd_cp_lpf_0/VQBb low_freq_pll_0/pfd_cp_lpf_0/vswitchl VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6041 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6042 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6043 biquad_gm_c_filter_0/ibiasn2 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X6044 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6045 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6046 a_239361_n114883# a_239143_n115125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X6047 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6048 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6049 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6050 VSS input_amplifier_0/ibiasn1 input_amplifier_0/ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6051 a_237397_n130007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin a_236939_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X6052 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6053 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6054 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6055 a_226954_n122869# low_freq_pll_0/cs_ring_osc_0/vpbias a_227412_n122869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X6056 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6057 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6058 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6059 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6060 biquad_gm_c_filter_0/ibiasn3 biquad_gm_c_filter_0/ibiasn3 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X6061 a_226481_n130007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_226023_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X6062 vintm vfiltp biquad_gm_c_filter_0/gm_c_stage_2/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6063 a_275374_n180872# sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6064 diff_to_se_converter_0/txgate_0/txb diff_to_se_converter_0/rst VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6065 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6066 VDD input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X6067 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6068 vrefA VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6069 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6070 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6071 VDD low_freq_pll_0/cs_ring_osc_0/vpbias a_240730_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X6072 VDD VDD dac_8bit_0/amux_2to1_6/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6073 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6074 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X6075 sample_and_hold_0/vholdm vcp_sampled sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X6076 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6077 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6078 VSS dac_8bit_0/latched_comparator_folded_0/vcompp_buf a_383508_n101129# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6079 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X6080 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6081 a_226785_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_226327_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X6082 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6083 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X6084 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6085 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6086 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6087 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6088 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6089 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6090 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6091 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6092 a_246328_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin a_245870_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6093 vpeak_sampled vpeak_sampled vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6094 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6095 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/vim1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X6096 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6097 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6098 vlowA VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6099 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6100 a_228770_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_228312_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6101 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/M1d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6102 a_222397_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin a_221939_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X6103 input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6104 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6105 biquad_gm_c_filter_0/ibiasn1 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X6106 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6107 VDD VDD dac_8bit_0/amux_2to1_3/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6108 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6109 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6110 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6111 vlowB dac_8bit_1/amux_2to1_10/SELB dac_8bit_1/amux_2to1_7/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6112 VDD peak_detector_0/verr peak_detector_0/vpeak VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6113 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6114 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6115 dac_8bit_1/amux_2to1_6/B VSS vrefB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6116 pulse_generator_0/sky130_fd_sc_hd__inv_1_1/A pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A a_335507_n185243# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6117 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6118 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6119 a_242909_n120623# a_241919_n120623# a_242783_n120257# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X6120 vpeak_sampled sample sample_and_hold_1/vholdm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6121 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6122 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6123 VSS input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6124 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6125 a_230446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6126 dac_8bit_0/amux_2to1_6/B dac_8bit_0/amux_2to1_11/SELB vlowA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6127 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6128 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 vpeak VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6129 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6130 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6131 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6132 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6133 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6134 adc_compB dac_8bit_1/latched_comparator_folded_0/vcompm_buf VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6135 VDD a_338356_n185510# a_338285_n185409# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X6136 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6137 dac_8bit_1/latched_comparator_folded_0/vlatchm adc_clk dac_8bit_1/latched_comparator_folded_0/vcompm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X6138 a_242358_n121345# a_242085_n121711# a_242273_n121711# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6139 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_242951_n120355# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6140 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6141 input_amplifier_0/vop1 input_amplifier_0/vim1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X6142 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6143 a_275374_n180872# sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6144 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6145 VDD VDD dac_8bit_0/amux_2to1_0/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6146 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6147 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6148 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6149 vlowB dac_8bit_1/amux_2to1_13/SELB dac_8bit_1/amux_2to1_4/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6150 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6151 adc_vcaparrayA dac_8bit_0/c2m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6152 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/vim2 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X6153 dac_8bit_1/amux_2to1_3/B q4B vrefB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6154 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6155 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6156 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6157 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6158 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6159 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6160 a_227562_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_227104_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X6161 VDD VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6162 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6163 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6164 dac_8bit_1/ibiasn dac_8bit_1/ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6165 dac_8bit_0/amux_2to1_3/B dac_8bit_0/amux_2to1_14/SELB vlowA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6166 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6167 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6168 VDD VDD vintp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6169 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6170 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6171 VSS a_242951_n123369# a_243382_n123343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6172 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/vcom_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6173 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X6174 a_338703_n185243# a_338156_n184969# a_338356_n185269# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6175 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 a_162668_n147576# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6176 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X6177 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6178 input_amplifier_0/vip1 vhpf sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X6179 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6180 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6181 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6182 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X6183 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6184 dac_8bit_0/amux_2to1_7/B VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6185 VSS input_amplifier_0/ibiasn2 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6186 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6187 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6188 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6189 a_246327_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin a_245869_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X6190 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6191 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6192 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6193 vlowB dac_8bit_1/amux_2to1_16/SELB dac_8bit_1/amux_2to1_1/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6194 biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail2 vintp biquad_gm_c_filter_0/gm_c_stage_0/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6195 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6196 VSS input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6197 adc_vcaparrayB dac_8bit_1/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6198 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6199 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6200 VSS biquad_gm_c_filter_0/ibiasn1 biquad_gm_c_filter_0/ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X6201 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 a_356329_n164260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6202 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6203 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6204 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6205 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6206 dac_8bit_1/c7m sample dac_8bit_1/amux_2to1_0/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6207 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6208 dac_8bit_0/c7m dac_8bit_0/amux_2to1_0/SELB vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6209 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6210 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6211 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6212 dac_8bit_1/c2m sample vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6213 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6214 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vfoldp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6215 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6216 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6217 vlowB sample adc_vcaparrayB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6218 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6219 VDD dac_8bit_0/latched_comparator_folded_0/vcompp dac_8bit_0/latched_comparator_folded_0/vcompm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6220 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6221 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6222 dac_8bit_0/c2m dac_8bit_0/amux_2to1_5/SELB dac_8bit_0/amux_2to1_5/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6223 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6224 input_amplifier_0/vip1 vhpf sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X6225 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6226 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn vse peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6227 dac_8bit_0/amux_2to1_4/B VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6228 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6229 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 vpeak VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6230 dac_8bit_0/latched_comparator_folded_0/vlatchm VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6231 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X6232 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6233 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_5/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6234 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6235 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6236 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn vintp biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6237 dac_8bit_0/amux_2to1_9/Y sample dac_8bit_0/c0m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6238 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6239 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6240 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6241 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6242 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 a_163060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6243 a_228478_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X6244 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6245 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6246 dac_8bit_1/c5m sample vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6247 VDD VDD vfiltp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6248 input_amplifier_0/venp1 input_amplifier_0/vop1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X6249 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6250 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6251 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6252 vlowB q7B dac_8bit_1/amux_2to1_0/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6253 dac_8bit_0/c5m dac_8bit_0/amux_2to1_2/SELB dac_8bit_0/amux_2to1_2/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6254 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6255 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 a_356329_n164260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6256 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6257 VSS vpeak_sampled sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X6258 dac_8bit_0/amux_2to1_1/B VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6259 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/vim2 input_amplifier_0/diff_fold_casc_ota_1/vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X6260 VSS biquad_gm_c_filter_0/ibiasn4 biquad_gm_c_filter_0/ibiasn4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X6261 a_222956_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_222498_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X6262 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6263 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6264 input_amplifier_0/txgate_7/txb input_amplifier_0/rst VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6265 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 vse VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6266 VDD VDD dac_8bit_1/amux_2to1_9/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6267 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.4e+07u
X6268 VDD VDD vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6269 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6270 vampp input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6271 VDD VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6272 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6273 input_amplifier_0/ibiasn1 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X6274 dac_8bit_0/latched_comparator_folded_0/vlatchm adc_clk dac_8bit_0/latched_comparator_folded_0/vlatchp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X6275 dac_8bit_0/amux_2to1_5/B sample dac_8bit_0/c2m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6276 VSS VSS input_amplifier_0/vop1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6277 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6278 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6279 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6280 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6281 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6282 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6283 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6284 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6285 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6286 a_221938_n150168# vcp a_221480_n150168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6287 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6288 VSS low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_227702_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6289 VDD input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vfoldp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6290 input_amplifier_0/venp1 input_amplifier_0/vop1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X6291 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 a_275374_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6292 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6293 VDD VDD low_freq_pll_0/cs_ring_osc_0/vosc VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X6294 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6295 VDD VDD input_amplifier_0/vim2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6296 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/vip2 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X6297 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6298 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X6299 VDD a_245224_n122281# a_245151_n122255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6300 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6301 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6302 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6303 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6304 dac_8bit_0/latched_comparator_folded_0/vcompm_buf dac_8bit_0/latched_comparator_folded_0/vcompmb VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6305 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6306 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6307 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6308 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6309 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6310 a_356329_n164260# dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6311 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6312 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6313 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6314 VDD VDD dac_8bit_1/amux_2to1_5/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6315 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6316 VDD VDD vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6317 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6318 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6319 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6320 low_freq_pll_0/cs_ring_osc_0/vosc low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout a_238923_n122049# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X6321 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6322 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6323 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6324 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6325 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6326 VDD input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/M6d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6327 a_236939_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_236481_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X6328 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6329 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin a_238771_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X6330 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6331 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6332 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X6333 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/vim1 input_amplifier_0/diff_fold_casc_ota_0/vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X6334 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6335 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6336 dac_8bit_1/amux_2to1_9/Y dac_8bit_1/amux_2to1_9/SELB vlowB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6337 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6338 sample_and_hold_0/vhold VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6339 input_amplifier_0/diff_fold_casc_ota_1/vcascnm input_amplifier_0/diff_fold_casc_ota_1/vbias3 vampm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6340 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/vcom_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6341 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6342 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6343 a_245056_n122255# a_244617_n122249# a_244971_n122255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X6344 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6345 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6346 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6347 a_242526_n122687# a_242358_n122433# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X6348 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/M2d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6349 input_amplifier_0/vop1 input_amplifier_0/vop1 input_amplifier_0/vop1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6350 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6351 adc_vcaparrayA dac_8bit_0/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6352 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6353 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6354 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X6355 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6356 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6357 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6358 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6359 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
X6360 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6361 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X6362 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6363 adc_vcaparrayA sample vlowA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6364 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6365 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 a_275374_n146348# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6366 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6367 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6368 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6369 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6370 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6371 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6372 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin a_223771_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X6373 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6374 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X6375 input_amplifier_0/txgate_1/txb gain_ctrl_0 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6376 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6377 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6378 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 input_amplifier_0/ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6379 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6380 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6381 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6382 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6383 a_356329_n113250# dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6384 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6385 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6386 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6387 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6388 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6389 VSS VSS biquad_gm_c_filter_0/gm_c_stage_1/vtail_diff VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X6390 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6391 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6392 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6393 vse VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X6394 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6395 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q a_241919_n123337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6396 low_freq_pll_0/pfd_cp_lpf_0/vpdiode VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6397 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6398 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6399 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6400 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6401 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6402 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6403 VSS dac_8bit_0/latched_comparator_folded_0/vlatchp dac_8bit_0/latched_comparator_folded_0/vlatchm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X6404 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6405 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6406 dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6407 VDD input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/M2d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6408 VDD dac_8bit_0/latched_comparator_folded_0/vcomppb dac_8bit_0/latched_comparator_folded_0/vcompp_buf VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6409 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X6410 VDD low_freq_pll_0/cs_ring_osc_0/vpbias a_236582_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X6411 a_336359_n185787# a_335844_n185460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6412 dac_8bit_1/c1m dac_8bit_1/amux_2to1_7/SELB dac_8bit_1/amux_2to1_7/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6413 a_227855_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_227397_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X6414 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X6415 comparator_0/vmirror comparator_0/vcompm VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6416 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6417 dac_8bit_1/amux_2to1_6/B VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6418 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6419 dac_8bit_1/ibiasp dac_8bit_1/ibiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6420 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6421 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6422 vpeak sample sample_and_hold_1/vhold VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6423 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6424 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6425 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6426 input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc vocm input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X6427 a_245182_n120789# a_244783_n121161# a_245056_n121167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X6428 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X6429 peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6430 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6431 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6432 input_amplifier_0/diff_fold_casc_ota_1/vcascnm input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6433 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn vse peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6434 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6435 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6436 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6437 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6438 vintp vfiltm biquad_gm_c_filter_0/gm_c_stage_2/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6439 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6440 low_freq_pll_0/ibiasn low_freq_pll_0/ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X6441 VDD input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vfoldm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6442 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6443 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6444 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6445 peak_detector_0/vpeak VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X6446 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6447 adc_vcaparrayA dac_8bit_0/c0m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6448 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6449 dac_8bit_1/c3m dac_8bit_1/amux_2to1_4/SELB dac_8bit_1/amux_2to1_4/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6450 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 a_230446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6451 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X6452 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6453 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6454 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/diff_fold_casc_ota_1/vbias2 vampp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6455 dac_8bit_1/amux_2to1_3/B VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6456 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6457 input_amplifier_0/vip2 gain_ctrl_0 input_amplifier_0/venm1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6458 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6459 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6460 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6461 dac_8bit_0/latched_comparator_folded_0/vlatchp adc_clk dac_8bit_0/latched_comparator_folded_0/vlatchm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X6462 vfiltm vintm biquad_gm_c_filter_0/gm_c_stage_3/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6463 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6464 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6465 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/vim2 input_amplifier_0/diff_fold_casc_ota_1/vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X6466 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6467 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6468 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6469 input_amplifier_0/diff_fold_casc_ota_0/vcascnm input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/vom1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6470 VSS VSS biquad_gm_c_filter_0/gm_c_stage_0/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6471 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6472 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6473 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X6474 a_337864_n185555# a_338149_n185569# a_338084_n185421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X6475 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6476 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6477 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6478 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6479 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6480 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6481 a_244971_n122255# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6482 VSS input_amplifier_0/ibiasn2 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6483 VDD a_242951_n123369# a_242867_n123343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6484 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6485 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6486 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X6487 vlowB VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6488 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6489 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6490 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6491 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/vim1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X6492 dac_8bit_1/c6m dac_8bit_1/amux_2to1_1/SELB dac_8bit_1/amux_2to1_1/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6493 input_amplifier_0/diff_fold_casc_ota_0/vcascnp input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/vop1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6494 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6495 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6496 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6497 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6498 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6499 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6500 a_237040_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_236582_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X6501 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6502 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X6503 vlowA VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6504 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6505 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6506 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6507 a_356329_n164260# dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6508 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6509 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6510 VSS VDD a_243138_n114759# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6511 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X6512 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 a_356329_n164260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6513 comparator_0/vcompp vfiltm comparator_0/vtail VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6514 VSS input_amplifier_0/ibiasn1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6515 VDD VDD dac_8bit_0/amux_2to1_2/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6516 a_236022_n150168# vcp low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/csinvn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6517 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X6518 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6519 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6520 dac_8bit_1/amux_2to1_5/B q2B vrefB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6521 VDD low_freq_pll_0/cs_ring_osc_0/vosc2 low_freq_pll_0/freq_div_0/vin VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6522 input_amplifier_0/ibiasn2 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X6523 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6524 dac_8bit_0/latched_comparator_folded_0/vtailp dac_8bit_0/latched_comparator_folded_0/vtailp dac_8bit_0/latched_comparator_folded_0/vtailp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6525 input_amplifier_0/diff_fold_casc_ota_1/M1d input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6526 dac_8bit_0/amux_2to1_5/B dac_8bit_0/amux_2to1_12/SELB vlowA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6527 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 a_217060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6528 input_amplifier_0/vip1 vhpf sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X6529 vlowA VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6530 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6531 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6532 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6533 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6534 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6535 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/M1d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6536 sample_and_hold_0/vholdm VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6537 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6538 vfiltm diff_to_se_converter_0/rst diff_to_se_converter_0/vim VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6539 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6540 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_2/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6541 VDD a_245649_n121193# a_245565_n121167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6542 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6543 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X6544 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6545 a_163060_n102324# input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6546 a_224330_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_223872_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X6547 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6548 input_amplifier_0/ibiasn2 input_amplifier_0/ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6549 VSS a_338356_n185269# a_338285_n185243# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6550 input_amplifier_0/diff_fold_casc_ota_1/vcascnp input_amplifier_0/diff_fold_casc_ota_1/vbias3 vampp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6551 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6552 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6553 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6554 dac_8bit_1/amux_2to1_2/B q5B vrefB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6555 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6556 a_228786_n119618# vcp a_228328_n119618# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6557 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6558 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6559 peak_detector_0/ibiasn2 peak_detector_0/ibiasn2 peak_detector_0/ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6560 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6561 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/vip2 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X6562 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6563 VSS VSS biquad_gm_c_filter_0/gm_c_stage_0/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6564 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6565 VDD input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vfoldp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6566 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6567 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6568 dac_8bit_0/amux_2to1_2/B dac_8bit_0/amux_2to1_15/SELB vlowA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6569 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6570 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6571 a_223312_n150168# vcp a_222854_n150168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6572 input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X6573 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6574 vlowA VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6575 VDD a_245224_n121599# a_245151_n121345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6576 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6577 vampp input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vfoldp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6578 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 a_356329_n113250# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6579 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6580 a_242867_n122255# a_242085_n122249# a_242783_n122255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6581 vincm input_amplifier_0/txgate_5/txb input_amplifier_0/vip1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6582 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6583 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn2 vocm_filt biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6584 VDD a_245649_n122531# a_246080_n122477# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6585 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6586 input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X6587 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6588 VSS VSS adc_vcaparrayB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6589 vampp input_amplifier_0/txgate_3/txb input_amplifier_0/venp2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6590 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6591 dac_8bit_0/amux_2to1_8/SELB sample VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6592 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/vim1 input_amplifier_0/diff_fold_casc_ota_0/vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X6593 diff_to_se_converter_0/vim VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6594 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6595 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6596 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6597 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6598 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6599 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6600 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6601 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6602 a_221480_n131500# low_freq_pll_0/cs_ring_osc_0/vosc a_221022_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6603 biquad_gm_c_filter_0/gm_c_stage_2/vtail_diff biquad_gm_c_filter_0/ibiasn4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X6604 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6605 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6606 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6607 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6608 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6609 VDD low_freq_pll_0/pfd_cp_lpf_0/vQA low_freq_pll_0/pfd_cp_lpf_0/vRSTN VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6610 a_238313_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_237855_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X6611 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6612 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 a_275374_n146348# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6613 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X6614 comparator_0/vtail comparator_0/vtail comparator_0/vtail VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X6615 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6616 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6617 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6618 biquad_gm_c_filter_0/gm_c_stage_0/vtail_diff vampm vintm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6619 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X6620 VDD low_freq_pll_0/freq_div_0/vin a_241919_n120623# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6621 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X6622 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6623 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6624 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/vcom_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6625 input_amplifier_0/diff_fold_casc_ota_1/vcascnm input_amplifier_0/diff_fold_casc_ota_1/vbias3 vampm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6626 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6627 VSS a_245481_n122433# a_245649_n122531# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6628 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6629 diff_to_se_converter_0/vip vocm_filt sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X6630 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6631 adc_vcaparrayA dac_8bit_0/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6632 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6633 dac_8bit_0/amux_2to1_7/B sample dac_8bit_0/c1m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6634 biquad_gm_c_filter_0/ibiasn1 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X6635 a_356329_n164260# dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6636 dac_8bit_0/cdumm dac_8bit_0/amux_2to1_6/SELB vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6637 dac_8bit_0/latched_comparator_folded_0/vtailp vlowA dac_8bit_0/latched_comparator_folded_0/vlatchm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6638 VSS biquad_gm_c_filter_0/ibiasn2 biquad_gm_c_filter_0/ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X6639 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6640 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/verr VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6641 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6642 input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X6643 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6644 VDD VDD low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X6645 peak_detector_0/ibiasn1 peak_detector_0/ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6646 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6647 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6648 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6649 VDD a_242575_n114888# a_242506_n114759# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X6650 dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6651 a_242085_n121711# a_241919_n121711# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6652 VSS input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6653 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6654 dac_8bit_0/amux_2to1_0/SELB sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6655 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6656 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X6657 a_242085_n121711# a_241919_n121711# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6658 input_amplifier_0/diff_fold_casc_ota_0/vcascnm input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/vom1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6659 biquad_gm_c_filter_0/ibiasn1 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X6660 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6661 dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6662 dac_8bit_0/latched_comparator_folded_0/vlatchm vlowA dac_8bit_0/latched_comparator_folded_0/vtailp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6663 input_amplifier_0/vop1 input_amplifier_0/txgate_6/txb input_amplifier_0/vim2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6664 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6665 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6666 vcp_sampled vcp_sampled vcp_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6667 VDD vbiasp biquad_gm_c_filter_0/ibiasn2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X6668 VDD VDD dac_8bit_1/amux_2to1_7/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6669 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6670 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6671 VDD VDD vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6672 dac_8bit_0/amux_2to1_4/B sample dac_8bit_0/c3m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6673 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X6674 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6675 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6676 dac_8bit_0/ibiasn dac_8bit_0/ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6677 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6678 dac_8bit_0/c4m dac_8bit_0/amux_2to1_3/SELB vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6679 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6680 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6681 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6682 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X6683 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6684 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6685 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6686 VSS a_239883_n115151# a_239817_n115125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6687 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6688 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6689 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6690 dac_8bit_1/amux_2to1_17/SELB q7B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6691 a_336359_n184877# a_335844_n185269# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6692 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6693 a_189446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6694 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6695 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6696 a_241022_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6697 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6698 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6699 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X6700 VDD VDD dac_8bit_1/amux_2to1_4/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6701 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6702 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6703 VDD VDD vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6704 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6705 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 a_356329_n113250# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6706 dac_8bit_0/amux_2to1_1/B sample dac_8bit_0/c6m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6707 low_freq_pll_0/pfd_cp_lpf_0/vswitchh VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X6708 VDD a_239708_n115125# a_239883_n115151# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6709 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6710 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6711 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6712 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6713 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6714 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6715 dac_8bit_1/amux_2to1_7/B dac_8bit_1/amux_2to1_10/SELB vlowB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6716 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6717 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6718 a_228328_n122869# low_freq_pll_0/cs_ring_osc_0/vpbias a_227870_n122869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X6719 vlowB VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6720 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6721 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6722 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6723 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6724 input_amplifier_0/vop1 input_amplifier_0/vim1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X6725 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6726 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6727 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6728 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6729 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6730 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6731 adc_vcaparrayA dac_8bit_0/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6732 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6733 VDD VDD dac_8bit_1/amux_2to1_1/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6734 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6735 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6736 a_242104_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_242562_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X6737 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6738 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6739 VDD VDD vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6740 input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vbias3 a_163060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6741 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6742 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6743 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6744 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6745 a_236480_n132168# vcp a_236022_n132168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6746 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6747 a_244971_n121711# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6748 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6749 VDD a_242951_n122531# a_242867_n122433# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6750 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6751 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6752 dac_8bit_1/amux_2to1_4/B dac_8bit_1/amux_2to1_13/SELB vlowB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6753 VDD VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6754 VDD VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6755 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6756 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6757 vlowB VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6758 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q a_242951_n122531# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6759 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6760 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6761 input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vfoldm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6762 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6763 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6764 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6765 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X6766 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6767 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6768 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6769 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6770 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6771 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6772 VDD VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6773 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6774 vintm biquad_gm_c_filter_0/gm_c_stage_2/vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6775 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6776 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6777 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/vim2 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X6778 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X6779 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6780 vampm VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6781 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/vim1 input_amplifier_0/diff_fold_casc_ota_0/vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X6782 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6783 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6784 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/csinvp low_freq_pll_0/cs_ring_osc_0/vpbias a_239330_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X6785 input_amplifier_0/vop1 input_amplifier_0/vop1 input_amplifier_0/vop1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6786 biquad_gm_c_filter_0/ibiasn1 biquad_gm_c_filter_0/ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X6787 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6788 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6789 dac_8bit_1/amux_2to1_1/B dac_8bit_1/amux_2to1_16/SELB vlowB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6790 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X6791 vcp_sampled dac_8bit_0/amux_2to1_8/SELB dac_8bit_0/c0m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6792 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 a_275374_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6793 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6794 peak_detector_0/ibiasn2 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X6795 VSS pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/D a_336955_n185409# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6796 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6797 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6798 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6799 VDD a_242951_n120355# a_243382_n120301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6800 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 a_163060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6801 dac_8bit_0/latched_comparator_folded_0/vcompm VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6802 a_223770_n132168# vcp a_223312_n132168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6803 a_356329_n164260# dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6804 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6805 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6806 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6807 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6808 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6809 dac_8bit_1/amux_2to1_5/B VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6810 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6811 VDD VDD biquad_gm_c_filter_0/gm_c_stage_2/vcmcn2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6812 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6813 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6814 dac_8bit_0/amux_2to1_0/B q7A vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6815 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6816 VSS VSS vintm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6817 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6818 VDD a_336401_n185269# a_336408_n184969# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6819 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6820 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6821 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6822 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X6823 dac_8bit_1/c0m dac_8bit_1/amux_2to1_8/SELB vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6824 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6825 dac_8bit_0/c0m sample dac_8bit_0/amux_2to1_9/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6826 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6827 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6828 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6829 a_162668_n147576# diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6830 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6831 diff_to_se_converter_0/ibiasn diff_to_se_converter_0/ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6832 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6833 biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail1 vintp biquad_gm_c_filter_0/gm_c_stage_1/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6834 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6835 input_amplifier_0/venp1 gain_ctrl_0 input_amplifier_0/vim2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6836 a_244971_n123343# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6837 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6838 input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6839 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6840 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 input_amplifier_0/ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6841 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6842 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6843 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6844 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6845 a_222498_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_222956_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X6846 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6847 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6848 a_230160_n119618# vcp a_229702_n119618# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6849 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6850 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6851 dac_8bit_1/amux_2to1_2/B VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6852 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X6853 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X6854 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6855 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6856 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 vpeak VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6857 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6858 vfiltm biquad_gm_c_filter_0/gm_c_stage_3/vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6859 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6860 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6861 a_242867_n121345# a_242085_n121711# a_242783_n121345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6862 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6863 a_245481_n121345# a_244783_n121711# a_245224_n121599# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X6864 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6865 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6866 input_amplifier_0/venm2 input_amplifier_0/txgate_2/txb vampm VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6867 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6868 dac_8bit_1/amux_2to1_6/B sample dac_8bit_1/cdumm VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6869 vcp_sampled dac_8bit_0/amux_2to1_6/SELB dac_8bit_0/cdumm VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6870 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6871 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6872 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6873 vse VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6874 a_245151_n122255# a_244617_n122249# a_245056_n122255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6875 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6876 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6877 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6878 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_0/A a_243382_n120301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6879 VSS peak_detector_0/vpeak sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X6880 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6881 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6882 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6883 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6884 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6885 input_amplifier_0/ibiasn1 input_amplifier_0/ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6886 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6887 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6888 VDD VDD input_amplifier_0/vip2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6889 VDD VDD vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6890 comparator_0/vcompm vfiltp comparator_0/vtail VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6891 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6892 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 a_356329_n113250# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6893 dac_8bit_0/latched_comparator_folded_0/vlatchm vlowA dac_8bit_0/latched_comparator_folded_0/vtailp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6894 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/csinvn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6895 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6896 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X6897 a_237854_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin a_237396_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6898 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X6899 VDD VDD biquad_gm_c_filter_0/gm_c_stage_3/vcmcn2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6900 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6901 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6902 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6903 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6904 VDD VDD input_amplifier_0/diff_fold_casc_ota_0/vfoldm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6905 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6906 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6907 VDD input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/M2d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6908 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X6909 VDD VDD vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6910 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6911 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6912 dac_8bit_1/amux_2to1_3/B sample dac_8bit_1/c4m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6913 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6914 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6915 vcp_sampled dac_8bit_0/amux_2to1_3/SELB dac_8bit_0/c4m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6916 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6917 VDD comparator_0/vcompm comparator_0/vcompp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6918 VSS a_242783_n122255# a_242951_n122281# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6919 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6920 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/csinvp VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X6921 dac_8bit_1/latched_comparator_folded_0/vlatchm VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X6922 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/M1d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6923 sample_and_hold_0/vholdm sample vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6924 a_217060_n102324# input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6925 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6926 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6927 VDD VDD vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6928 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6929 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6930 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6931 a_244783_n122249# a_244617_n122249# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6932 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6933 VSS vbiasn dac_8bit_1/ibiasp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=2e+06u
X6934 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6935 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6936 a_230446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6937 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6938 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6939 a_242377_n115125# a_241731_n115151# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6940 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6941 a_243771_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_243313_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X6942 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6943 VDD VDD vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6944 input_amplifier_0/diff_fold_casc_ota_0/vcascnp input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6945 dac_8bit_1/amux_2to1_0/B sample dac_8bit_1/c7m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6946 a_242085_n121161# a_241919_n121161# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6947 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6948 vcp_sampled dac_8bit_0/amux_2to1_0/SELB dac_8bit_0/c7m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6949 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6950 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6951 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/verr VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6952 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/vip2 input_amplifier_0/diff_fold_casc_ota_1/vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X6953 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 a_189446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6954 a_222854_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin a_222396_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6955 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6956 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6957 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6958 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6959 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6960 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6961 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6962 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6963 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6964 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6965 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6966 vampm input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6967 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6968 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X6969 diff_to_se_converter_0/vim diff_to_se_converter_0/rst vfiltm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6970 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6971 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6972 low_freq_pll_0/pfd_cp_lpf_0/vndiode low_freq_pll_0/pfd_cp_lpf_0/vQA low_freq_pll_0/pfd_cp_lpf_0/vswitchh VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6973 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6974 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X6975 input_amplifier_0/vim1 input_amplifier_0/rst vincm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6976 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6977 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6978 a_237396_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_236938_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6979 input_amplifier_0/txgate_0/txb gain_ctrl_0 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6980 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X6981 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6982 vlowA sample adc_vcaparrayA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6983 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn2 vocm_filt biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6984 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X6985 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6986 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6987 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6988 VDD VDD vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6989 a_337497_n185269# a_337592_n185269# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6990 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6991 a_230446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6992 comparator_0/vo1 comparator_0/vmirror VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6993 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X6994 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6995 biquad_gm_c_filter_0/ibiasn2 biquad_gm_c_filter_0/ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X6996 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6997 a_226480_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_226022_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X6998 a_163060_n102324# input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6999 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7000 a_228770_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_228312_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X7001 input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X7002 dac_8bit_0/amux_2to1_7/SELB sample VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7003 a_222397_n130007# low_freq_pll_0/cs_ring_osc_0/vosc a_221939_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X7004 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7005 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7006 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7007 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7008 a_275374_n180872# sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7009 biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail2 vocm_filt biquad_gm_c_filter_0/gm_c_stage_2/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7010 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7011 adc_vcaparrayB dac_8bit_1/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7012 vpeak_sampled vpeak_sampled VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7013 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7014 a_242102_n114873# a_242380_n114857# a_242336_n114759# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7015 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/verr VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7016 input_amplifier_0/rst rst_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7017 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7018 low_freq_pll_0/pfd_cp_lpf_0/vswitchh VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7019 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7020 VDD VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7021 diff_to_se_converter_0/vip vocm_filt sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X7022 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 a_356329_n164260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7023 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7024 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7025 vcomp comparator_0/vo1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7026 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7027 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X7028 biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail2 vfiltm biquad_gm_c_filter_0/gm_c_stage_3/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7029 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7030 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7031 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7032 VDD low_freq_pll_0/cs_ring_osc_0/vpbias a_225730_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X7033 low_freq_pll_0/pfd_cp_lpf_0/vswitchl VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7034 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7035 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7036 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7037 input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vbias3 a_217060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7038 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7039 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 a_356329_n113250# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7040 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7041 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7042 VSS dac_8bit_1/latched_comparator_folded_0/vlatchm dac_8bit_1/latched_comparator_folded_0/vlatchp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X7043 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7044 input_amplifier_0/venp2 input_amplifier_0/vim2 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X7045 dac_8bit_0/amux_2to1_4/SELB sample VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7046 VDD input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vfoldp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7047 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7048 vampp VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X7049 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7050 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7051 adc_vcaparrayA dac_8bit_0/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7052 a_231328_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin a_230870_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X7053 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7054 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7055 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X7056 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7057 dac_8bit_0/latched_comparator_folded_0/vtailp dac_8bit_0/ibiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X7058 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7059 a_240730_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_241188_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X7060 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7061 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7062 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7063 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7064 a_244783_n121161# a_244617_n121161# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7065 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7066 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7067 dac_8bit_0/c2m dac_8bit_0/amux_2to1_5/SELB vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7068 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7069 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7070 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X7071 biquad_gm_c_filter_0/gm_c_stage_2/vtail_diff vfiltm vintp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7072 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7073 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7074 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/vim2 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X7075 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7076 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7077 VDD VDD low_freq_pll_0/pfd_cp_lpf_0/vswitchh VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X7078 sample_and_hold_1/vhold VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X7079 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7080 a_238872_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_239330_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X7081 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7082 input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X7083 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X7084 biquad_gm_c_filter_0/ibiasn1 biquad_gm_c_filter_0/ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X7085 vpeak_sampled dac_8bit_1/amux_2to1_8/SELB dac_8bit_1/c0m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7086 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7087 dac_8bit_0/amux_2to1_1/SELB sample VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7088 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7089 a_222956_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_223414_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X7090 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7091 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7092 peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7093 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 a_230446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7094 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7095 biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail1 vocm_filt biquad_gm_c_filter_0/gm_c_stage_2/vcmcn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7096 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7097 dac_8bit_0/c5m dac_8bit_0/amux_2to1_2/SELB vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7098 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7099 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7100 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7101 input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vbias3 a_163060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7102 vpeak vpeak vpeak VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7103 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7104 a_189446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7105 low_freq_pll_0/freq_div_0/vout a_245649_n121193# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7106 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7107 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7108 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/vcom_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7109 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7110 vincm input_amplifier_0/rst input_amplifier_0/vim1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7111 vpeak_sampled dac_8bit_1/amux_2to1_5/SELB dac_8bit_1/c2m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7112 input_amplifier_0/diff_fold_casc_ota_0/M6d input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7113 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7114 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X7115 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7116 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X7117 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7118 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7119 VDD VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7120 VDD a_242783_n120257# a_242951_n120355# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7121 VDD VDD vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7122 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7123 sample_and_hold_1/vholdm VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7124 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 a_189446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7125 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7126 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/vim1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X7127 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X7128 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X7129 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7130 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7131 VDD VDD dac_8bit_1/latched_comparator_folded_0/vlatchm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7132 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7133 VDD VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7134 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7135 input_amplifier_0/venm2 input_amplifier_0/vip2 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X7136 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7137 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7138 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7139 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7140 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 a_230446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7141 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7142 a_231327_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin a_230869_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X7143 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7144 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_3/A a_243382_n121389# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7145 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7146 vlowB VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7147 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7148 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7149 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7150 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7151 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X7152 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7153 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 a_217060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7154 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7155 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7156 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7157 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7158 VSS biquad_gm_c_filter_0/gm_c_stage_1/vcmc biquad_gm_c_filter_0/gm_c_stage_1/vtail_diff VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X7159 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7160 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7161 VDD VDD vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7162 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X7163 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7164 dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7165 dac_8bit_0/latched_comparator_folded_0/vcompp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7166 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7167 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/vcom_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7168 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7169 a_245151_n121345# a_244617_n121711# a_245056_n121345# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7170 VDD input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vfoldm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7171 a_217060_n102324# input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7172 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7173 vcomp comparator_0/vo1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7174 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7175 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7176 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7177 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7178 a_225870_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_225412_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X7179 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7180 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7181 input_amplifier_0/diff_fold_casc_ota_1/M6d input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7182 vlowB VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7183 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7184 a_237549_n122049# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout a_237091_n122049# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X7185 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7186 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7187 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/vim2 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X7188 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7189 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7190 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7191 diff_to_se_converter_0/ibiasn diff_to_se_converter_0/ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7192 a_162668_n147576# diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7193 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7194 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7195 VDD VDD vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7196 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_7/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7197 biquad_gm_c_filter_0/gm_c_stage_0/vtail_diff vampp vintp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7198 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7199 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7200 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7201 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7202 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7203 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q a_241919_n123337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7204 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7205 vfiltp diff_to_se_converter_0/rst diff_to_se_converter_0/vip VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7206 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7207 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X7208 a_237091_n122049# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout a_236633_n122049# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X7209 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7210 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7211 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7212 a_162668_n147576# diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7213 adc_vcaparrayB sample vlowB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7214 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7215 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7216 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7217 vpeak_sampled sample dac_8bit_1/c7m VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7218 a_236939_n130007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin a_236481_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X7219 vcp_sampled dac_8bit_0/amux_2to1_7/SELB dac_8bit_0/c1m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7220 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7221 dac_8bit_1/latched_comparator_folded_0/vlatchm VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X7222 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7223 VSS biquad_gm_c_filter_0/ibiasn4 biquad_gm_c_filter_0/ibiasn4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X7224 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7225 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7226 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7227 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7228 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7229 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7230 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7231 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7232 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7233 VSS dac_8bit_0/latched_comparator_folded_0/vcompp dac_8bit_0/latched_comparator_folded_0/vcomppb VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7234 biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail1 vocm_filt biquad_gm_c_filter_0/gm_c_stage_1/vcmcn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7235 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7236 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7237 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7238 VDD VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7239 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7240 dac_8bit_1/amux_2to1_6/SELB sample VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7241 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7242 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7243 adc_vcaparrayA dac_8bit_0/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7244 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7245 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7246 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7247 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7248 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7249 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7250 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 a_356329_n113250# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7251 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7252 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7253 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7254 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7255 diff_to_se_converter_0/vip VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7256 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7257 dac_8bit_1/c1m dac_8bit_1/amux_2to1_7/SELB vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7258 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7259 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7260 dac_8bit_0/c1m sample dac_8bit_0/amux_2to1_7/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7261 dac_8bit_1/amux_2to1_0/B dac_8bit_1/amux_2to1_17/SELB vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7262 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_238770_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X7263 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7264 a_230446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7265 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp vse peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7266 adc_compA dac_8bit_0/comp_outm a_383050_n101129# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7267 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7268 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X7269 vcp_sampled dac_8bit_0/amux_2to1_4/SELB dac_8bit_0/c3m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7270 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7271 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7272 dac_8bit_0/amux_2to1_6/B VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7273 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7274 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7275 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/verr VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7276 input_amplifier_0/vop1 input_amplifier_0/rst input_amplifier_0/vim2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7277 dac_8bit_0/latched_comparator_folded_0/vtailp vlowA dac_8bit_0/latched_comparator_folded_0/vlatchm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7278 dac_8bit_1/amux_2to1_3/SELB sample VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7279 a_221939_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin a_221481_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X7280 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs low_freq_pll_0/cs_ring_osc_0/vosc a_223771_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X7281 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7282 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7283 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7284 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7285 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X7286 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/diff_fold_casc_ota_1/vbias2 vampp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7287 vampm input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7288 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7289 a_230446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7290 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7291 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X7292 vrefA dac_8bit_0/amux_2to1_9/SELB dac_8bit_0/amux_2to1_9/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7293 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7294 a_245056_n121345# a_244617_n121711# a_244971_n121711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X7295 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7296 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7297 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7298 input_amplifier_0/vim2 input_amplifier_0/txgate_1/txb input_amplifier_0/venp1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7299 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7300 dac_8bit_1/c3m dac_8bit_1/amux_2to1_4/SELB vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7301 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X7302 dac_8bit_0/c3m sample dac_8bit_0/amux_2to1_4/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7303 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7304 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7305 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7306 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7307 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/vim2 input_amplifier_0/diff_fold_casc_ota_1/vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X7308 vcp_sampled dac_8bit_0/amux_2to1_1/SELB dac_8bit_0/c6m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7309 dac_8bit_1/ibiasn vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X7310 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7311 VDD comparator_0/vcompp comparator_0/vcompm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7312 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7313 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7314 a_275374_n180872# sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7315 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7316 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7317 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 a_275374_n146348# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7318 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_245649_n122531# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7319 VSS VSS biquad_gm_c_filter_0/gm_c_stage_3/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7320 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7321 VDD VDD vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7322 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7323 dac_8bit_0/amux_2to1_3/B VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7324 dac_8bit_1/latched_comparator_folded_0/vlatchp dac_8bit_1/vcom_buf dac_8bit_1/latched_comparator_folded_0/vtailp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7325 biquad_gm_c_filter_0/ibiasn3 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X7326 VSS vse sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X7327 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7328 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7329 a_242484_n122965# a_242085_n123337# a_242358_n123343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X7330 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X7331 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7332 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7333 input_amplifier_0/diff_fold_casc_ota_0/M3d VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7334 biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail2 biquad_gm_c_filter_0/ibiasn4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X7335 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7336 a_227855_n130007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_227397_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X7337 a_245224_n121193# a_245056_n121167# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7338 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7339 VDD VDD vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7340 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7341 biquad_gm_c_filter_0/ibiasn3 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X7342 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7343 a_239048_n115125# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7344 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7345 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7346 vrefA dac_8bit_0/amux_2to1_12/SELB dac_8bit_0/amux_2to1_5/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7347 dac_8bit_1/amux_2to1_2/B sample dac_8bit_1/c5m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7348 vcp_sampled dac_8bit_0/amux_2to1_2/SELB dac_8bit_0/c5m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7349 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 vpeak_sampled VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7350 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7351 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7352 VSS VSS dac_8bit_0/latched_comparator_folded_0/vlatchp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X7353 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7354 dac_8bit_1/c6m dac_8bit_1/amux_2to1_1/SELB vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7355 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7356 dac_8bit_0/c6m sample dac_8bit_0/amux_2to1_1/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7357 vcp_sampled vcp_sampled vcp_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7358 vincm VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7359 biquad_gm_c_filter_0/gm_c_stage_0/vtail_diff VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X7360 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7361 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7362 VDD low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_227701_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X7363 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7364 VDD a_242951_n122281# a_243382_n122255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7365 VDD VDD vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7366 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7367 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X7368 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7369 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7370 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7371 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7372 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7373 VDD VDD vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7374 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7375 VDD low_freq_pll_0/cs_ring_osc_0/vpbias a_221582_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X7376 a_163060_n102324# input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7377 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X7378 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7379 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7380 VDD VDD vpeak_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7381 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7382 input_amplifier_0/diff_fold_casc_ota_1/M1d input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7383 dac_8bit_0/latched_comparator_folded_0/vcompp adc_clk dac_8bit_0/latched_comparator_folded_0/vlatchp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X7384 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7385 a_189446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7386 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7387 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7388 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7389 input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vbias3 a_217060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7390 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7391 dac_8bit_0/c7m sample vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7392 biquad_gm_c_filter_0/gm_c_stage_2/vbiasp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7393 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7394 a_245056_n121167# a_244783_n121161# a_244971_n121167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7395 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7396 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X7397 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp vse peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7398 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7399 VDD VDD vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7400 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7401 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7402 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7403 a_227397_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_226939_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X7404 a_236582_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_237040_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X7405 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X7406 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7407 dac_8bit_1/amux_2to1_17/SELB q7B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7408 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7409 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/vim1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X7410 VDD VDD low_freq_pll_0/pfd_cp_lpf_0/vndiode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7411 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7412 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7413 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7414 vampp VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7415 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7416 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1.2e+07u w=2e+06u
X7417 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 a_230446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7418 peak_detector_0/ibiasn2 peak_detector_0/ibiasn2 peak_detector_0/ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7419 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7420 VSS a_245649_n122531# a_246080_n122477# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7421 VDD biquad_gm_c_filter_0/gm_c_stage_2/vcmcn1 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7422 VSS VSS biquad_gm_c_filter_0/gm_c_stage_3/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7423 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7424 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7425 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7426 low_freq_pll_0/ibiasn low_freq_pll_0/ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X7427 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X7428 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7429 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7430 input_amplifier_0/diff_fold_casc_ota_0/vcascnm input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7431 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7432 VDD comparator_0/vcompp comparator_0/vo1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7433 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7434 VDD VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7435 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7436 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/csinvp low_freq_pll_0/cs_ring_osc_0/vpbias a_228478_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X7437 VSS dac_8bit_0/ibiasn dac_8bit_0/ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7438 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7439 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7440 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q a_245649_n121443# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7441 input_amplifier_0/diff_fold_casc_ota_0/vcascnm input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/vom1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7442 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7443 VSS dac_8bit_0/vcom_buf sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X7444 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7445 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7446 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7447 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X7448 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 a_275374_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7449 sample_and_hold_1/vhold VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7450 input_amplifier_0/venp1 gain_ctrl_0 input_amplifier_0/vim2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7451 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7452 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7453 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7454 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7455 VDD adc_clk dac_8bit_1/latched_comparator_folded_0/vcompp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7456 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X7457 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7458 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7459 biquad_gm_c_filter_0/gm_c_stage_3/vbiasp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7460 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7461 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 a_275374_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7462 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7463 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7464 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7465 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7466 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7467 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7468 vpeak_sampled dac_8bit_1/amux_2to1_6/SELB dac_8bit_1/cdumm VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7469 dac_8bit_0/amux_2to1_6/B sample dac_8bit_0/cdumm VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7470 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7471 a_227702_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_227244_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X7472 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_10/A a_246080_n123343# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7473 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7474 input_amplifier_0/venm1 gain_ctrl_0 input_amplifier_0/vip2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7475 a_222040_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_221582_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X7476 a_244783_n122799# a_244617_n122799# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7477 biquad_gm_c_filter_0/gm_c_stage_3/vtail_diff vintp vfiltp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7478 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7479 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7480 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7481 dac_8bit_1/amux_2to1_9/Y VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7482 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7483 vcp_sampled VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7484 dac_8bit_1/latched_comparator_folded_0/vlatchm adc_clk dac_8bit_1/latched_comparator_folded_0/vlatchp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X7485 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn vintm biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7486 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_244617_n121711# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7487 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7488 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X7489 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7490 input_amplifier_0/diff_fold_casc_ota_0/M6d input_amplifier_0/diff_fold_casc_ota_0/M6d input_amplifier_0/diff_fold_casc_ota_0/M6d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7491 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7492 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7493 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7494 dac_8bit_0/amux_2to1_9/Y dac_8bit_0/amux_2to1_9/SELB vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7495 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_244617_n121711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7496 VSS vcp_sampled sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X7497 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7498 a_221022_n150168# vcp low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/csinvn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X7499 dac_8bit_1/latched_comparator_folded_0/vtailp dac_8bit_1/vcom_buf dac_8bit_1/latched_comparator_folded_0/vlatchp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7500 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7501 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7502 input_amplifier_0/venp2 input_amplifier_0/txgate_3/txb vampp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7503 VDD biquad_gm_c_filter_0/gm_c_stage_3/vcmcn1 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7504 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 a_275374_n146348# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7505 VSS VSS biquad_gm_c_filter_0/gm_c_stage_2/vtail_diff VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X7506 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7507 a_238923_n122049# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout a_238465_n122049# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X7508 input_amplifier_0/diff_fold_casc_ota_1/vcascnm input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7509 vpeak_sampled dac_8bit_1/amux_2to1_7/SELB dac_8bit_1/c1m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7510 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7511 VSS input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7512 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7513 VSS pulse_generator_0/sky130_fd_sc_hd__inv_1_1/A peak_detector_rst VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7514 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7515 input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/M3d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7516 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 a_356329_n113250# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7517 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7518 dac_8bit_1/cdumm sample dac_8bit_1/amux_2to1_6/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7519 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7520 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7521 input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc vocm input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X7522 vpeak_sampled dac_8bit_1/amux_2to1_3/SELB dac_8bit_1/c4m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7523 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7524 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7525 dac_8bit_0/amux_2to1_3/B sample dac_8bit_0/c4m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7526 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X7527 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7528 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7529 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7530 low_freq_pll_0/cs_ring_osc_0/vosc2 low_freq_pll_0/cs_ring_osc_0/vosc VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7531 input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7532 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7533 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7534 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7535 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7536 a_217060_n102324# input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7537 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7538 vlowA VSS dac_8bit_0/amux_2to1_6/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7539 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7540 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X7541 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7542 a_162668_n147576# diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7543 peak_detector_0/ibiasn1 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X7544 a_236023_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X7545 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7546 comparator_0/vtail vfiltp comparator_0/vcompm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7547 a_238313_n130007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin a_237855_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X7548 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7549 VDD VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7550 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7551 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7552 vpeak_sampled dac_8bit_1/amux_2to1_4/SELB dac_8bit_1/c3m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7553 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7554 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/vim1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X7555 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7556 dac_8bit_1/c4m sample dac_8bit_1/amux_2to1_3/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7557 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7558 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7559 a_336608_n185510# a_336401_n185569# a_336784_n185787# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7560 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/vcom_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7561 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7562 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7563 VDD VDD vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7564 vrefB q7B dac_8bit_1/amux_2to1_0/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7565 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7566 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7567 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7568 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7569 vlowA q4A dac_8bit_0/amux_2to1_3/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7570 peak_detector_0/verr peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7571 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7572 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7573 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7574 VSS a_242951_n122531# a_242909_n122799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7575 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7576 VSS VSS vcp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7577 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7578 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7579 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7580 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7581 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7582 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7583 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7584 VDD sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7585 dac_8bit_0/vcom_buf VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X7586 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7587 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X7588 a_227701_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_227243_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X7589 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7590 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7591 vpeak_sampled dac_8bit_1/amux_2to1_1/SELB dac_8bit_1/c6m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7592 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7593 input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/M3d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7594 low_freq_pll_0/pfd_cp_lpf_0/VQBb low_freq_pll_0/pfd_cp_lpf_0/vQB VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7595 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7596 a_336955_n185243# a_336401_n185269# a_336608_n185269# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X7597 a_242783_n122255# a_241919_n122249# a_242526_n122281# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7598 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7599 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7600 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X7601 vcp_sampled sample sample_and_hold_0/vholdm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7602 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7603 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7604 VDD VDD vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7605 a_163060_n102324# input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7606 dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7607 a_356329_n164260# dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7608 a_223313_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin a_222855_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X7609 a_242909_n121877# a_241919_n122249# a_242783_n122255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X7610 a_163060_n102324# input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7611 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7612 VDD VDD vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7613 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7614 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7615 vlowA q7A dac_8bit_0/amux_2to1_0/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7616 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7617 vse diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7618 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X7619 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7620 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7621 biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail2 vintm biquad_gm_c_filter_0/gm_c_stage_2/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7622 VSS comparator_0/ibiasn comparator_0/vtail VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X7623 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7624 VSS VSS low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X7625 VDD input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vfoldp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7626 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7627 VDD a_335749_n185813# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7628 low_freq_pll_0/pfd_cp_lpf_0/vRSTN low_freq_pll_0/pfd_cp_lpf_0/vQB VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7629 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7630 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7631 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7632 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7633 VDD dac_8bit_1/ibiasp dac_8bit_1/latched_comparator_folded_0/vtailp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X7634 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X7635 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7636 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7637 peak_detector_0/ibiasn1 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X7638 a_242273_n122255# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7639 adc_vcaparrayB dac_8bit_1/c2m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7640 low_freq_pll_0/pfd_cp_lpf_0/vndiode low_freq_pll_0/pfd_cp_lpf_0/vndiode VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7641 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7642 input_amplifier_0/vom1 input_amplifier_0/vom1 input_amplifier_0/vom1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7643 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp vse peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7644 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7645 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7646 VSS biquad_gm_c_filter_0/ibiasn2 biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X7647 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7648 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7649 VDD VDD vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7650 a_275374_n180872# sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7651 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7652 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7653 VDD VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7654 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/vim1 input_amplifier_0/diff_fold_casc_ota_0/vfoldp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X7655 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn vintm biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7656 input_amplifier_0/diff_fold_casc_ota_0/vcascnp input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7657 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7658 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7659 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7660 a_217060_n102324# input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7661 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7662 peak_detector_0/verr VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X7663 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7664 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7665 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7666 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7667 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7668 a_226038_n122869# low_freq_pll_0/cs_ring_osc_0/vpbias a_225580_n122869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X7669 VSS a_242951_n120355# a_243382_n120301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7670 biquad_gm_c_filter_0/gm_c_stage_2/vtail_diff vfiltp vintm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7671 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 vampm input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X7672 vse vse vse VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7673 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q a_245649_n123369# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7674 input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X7675 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7676 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7677 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7678 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7679 VSS input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7680 dac_8bit_1/amux_2to1_5/SELB sample VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7681 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7682 dac_8bit_1/amux_2to1_9/Y sample dac_8bit_1/c0m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7683 VDD sample dac_8bit_1/adc_run VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7684 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7685 a_243478_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_243020_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X7686 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7687 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7688 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7689 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7690 VSS VSS biquad_gm_c_filter_0/gm_c_stage_2/vbiasp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X7691 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7692 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7693 vse diff_to_se_converter_0/vim sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X7694 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7695 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7696 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7697 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7698 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_228771_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X7699 low_freq_pll_0/ibiasn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X7700 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7701 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7702 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7703 VSS VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7704 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 a_162668_n147576# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7705 input_amplifier_0/vim2 input_amplifier_0/txgate_6/txb input_amplifier_0/vop1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7706 vpeak VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X7707 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7708 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7709 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X7710 peak_detector_0/verr peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7711 input_amplifier_0/vom1 input_amplifier_0/rst input_amplifier_0/vip2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7712 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7713 dac_8bit_0/amux_2to1_5/B VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7714 a_275374_n146348# sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7715 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7716 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7717 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7718 dac_8bit_1/amux_2to1_2/SELB sample VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7719 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7720 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X7721 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7722 dac_8bit_0/amux_2to1_0/B q7A vrefA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7723 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 a_230446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7724 VDD VDD input_amplifier_0/diff_fold_casc_ota_0/M3d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7725 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7726 a_242813_n115125# low_freq_pll_0/pfd_cp_lpf_0/vRSTN VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7727 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7728 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7729 VSS a_245649_n122281# a_246080_n122255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7730 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7731 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7732 vrefA dac_8bit_0/amux_2to1_10/SELB dac_8bit_0/amux_2to1_7/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7733 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.4e+07u
X7734 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7735 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X7736 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X7737 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7738 dac_8bit_0/amux_2to1_6/B VSS vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7739 a_239883_n115151# low_freq_pll_0/pfd_cp_lpf_0/vRSTN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7740 a_237498_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_237040_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X7741 input_amplifier_0/diff_fold_casc_ota_1/vcascnp input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7742 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7743 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7744 vlowB q0B dac_8bit_1/amux_2to1_9/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7745 biquad_gm_c_filter_0/gm_c_stage_1/vbiasp biquad_gm_c_filter_0/ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X7746 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 a_275374_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7747 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7748 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7749 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X7750 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7751 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7752 dac_8bit_1/latched_comparator_folded_0/vtailp dac_8bit_1/vcom_buf dac_8bit_1/latched_comparator_folded_0/vlatchp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7753 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7754 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7755 a_227104_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_227562_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X7756 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7757 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7758 input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X7759 sample_and_hold_0/vhold VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X7760 dac_8bit_0/amux_2to1_2/B VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7761 a_227562_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_228020_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X7762 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7763 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7764 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X7765 adc_vcaparrayB dac_8bit_1/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7766 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7767 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7768 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X7769 a_221480_n132168# vcp a_221022_n132168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X7770 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7771 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp vse peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7772 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/vbias2 vampm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7773 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7774 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7775 VDD VDD vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7776 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7777 vrefA dac_8bit_0/amux_2to1_13/SELB dac_8bit_0/amux_2to1_4/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7778 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7779 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7780 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7781 dac_8bit_0/amux_2to1_3/B q4A vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7782 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7783 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7784 vlowB q2B dac_8bit_1/amux_2to1_5/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7785 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7786 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7787 a_244783_n122249# a_244617_n122249# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7788 VDD biquad_gm_c_filter_0/gm_c_stage_0/vbiasp biquad_gm_c_filter_0/gm_c_stage_0/vbiasp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7789 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7790 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7791 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7792 dac_8bit_0/vcom_buf VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X7793 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7794 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7795 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7796 VSS a_242783_n122433# a_242951_n122531# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7797 VDD VDD input_amplifier_0/vom1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7798 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7799 VDD input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/M1d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7800 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7801 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/csinvp low_freq_pll_0/cs_ring_osc_0/vpbias a_224330_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X7802 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7803 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7804 a_217060_n102324# input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7805 a_227870_n119618# vcp a_227412_n119618# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X7806 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7807 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 a_275374_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7808 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7809 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7810 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q a_244617_n121161# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7811 VDD VDD vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7812 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7813 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7814 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7815 vrefA dac_8bit_0/amux_2to1_16/SELB dac_8bit_0/amux_2to1_1/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7816 input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X7817 dac_8bit_0/latched_comparator_folded_0/vlatchp VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X7818 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7819 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7820 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7821 a_242484_n122799# a_242085_n122799# a_242358_n122433# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X7822 VSS vcp_sampled vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7823 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7824 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_8/A a_246080_n122255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7825 input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X7826 input_amplifier_0/vom1 input_amplifier_0/vip1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X7827 VSS dac_8bit_1/vcom_buf sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X7828 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7829 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7830 adc_vcaparrayB VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7831 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/vfoldm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X7832 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7833 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7834 VSS input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7835 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 a_275374_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7836 VDD dac_8bit_0/latched_comparator_folded_0/vcompp_buf dac_8bit_0/comp_outm VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7837 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 a_356329_n113250# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7838 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/csinvn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X7839 VDD VDD vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7840 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7841 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7842 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7843 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7844 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7845 dac_8bit_0/c0m sample dac_8bit_0/amux_2to1_9/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7846 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7847 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7848 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7849 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7850 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7851 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7852 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7853 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7854 VDD biquad_gm_c_filter_0/gm_c_stage_1/vbiasp biquad_gm_c_filter_0/gm_c_stage_1/vbiasp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7855 a_336608_n185269# a_336401_n185269# a_336784_n184877# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7856 VSS dac_8bit_1/ibiasn dac_8bit_1/ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7857 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7858 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7859 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7860 diff_to_se_converter_0/rst rst_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7861 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn2 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn2 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7862 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7863 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7864 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7865 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7866 VSS a_242951_n122281# a_242909_n121877# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7867 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7868 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7869 a_245224_n122687# a_245056_n122433# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7870 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7871 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7872 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7873 VDD pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A pulse_generator_0/sky130_fd_sc_hd__inv_1_1/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7874 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7875 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7876 input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X7877 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7878 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X7879 input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vfoldm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7880 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7881 a_241481_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_241023_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X7882 a_243771_n130007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_243313_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X7883 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp vse peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7884 a_242783_n121345# a_241919_n121711# a_242526_n121599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7885 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7886 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X7887 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7888 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7889 sample_and_hold_1/vhold VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X7890 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7891 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7892 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7893 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7894 biquad_gm_c_filter_0/ibiasn4 biquad_gm_c_filter_0/ibiasn4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X7895 vse VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X7896 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/csinvn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X7897 vlowA q0A dac_8bit_0/amux_2to1_9/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7898 a_222854_n131500# low_freq_pll_0/cs_ring_osc_0/vosc a_222396_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X7899 vpeak_sampled dac_8bit_1/amux_2to1_5/SELB dac_8bit_1/c2m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7900 dac_8bit_0/amux_2to1_5/B sample dac_8bit_0/c2m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7901 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7902 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X7903 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7904 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7905 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7906 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7907 dac_8bit_1/amux_2to1_7/B VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7908 vcp_sampled VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7909 VSS pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A a_338703_n185409# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7910 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7911 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7912 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X7913 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7914 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7915 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7916 dac_8bit_0/amux_2to1_7/B dac_8bit_0/amux_2to1_10/SELB vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7917 a_237396_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin a_236938_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X7918 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7919 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7920 VDD input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vfoldp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7921 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/vcom_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7922 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7923 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7924 dac_8bit_1/latched_comparator_folded_0/vtailp dac_8bit_1/latched_comparator_folded_0/vtailp dac_8bit_1/latched_comparator_folded_0/vtailp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X7925 a_336116_n185555# a_336401_n185569# a_336336_n185421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X7926 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7927 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7928 a_242273_n121711# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7929 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7930 input_amplifier_0/vip2 input_amplifier_0/txgate_0/txb input_amplifier_0/venm1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7931 a_162668_n147576# diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7932 dac_8bit_1/amux_2to1_9/Y q0B vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7933 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7934 vfiltm diff_to_se_converter_0/txgate_1/txb diff_to_se_converter_0/vim VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7935 VDD a_338149_n185269# a_338156_n184969# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7936 dac_8bit_1/c2m sample dac_8bit_1/amux_2to1_5/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7937 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7938 a_226480_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_226022_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X7939 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7940 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7941 vpeak_sampled dac_8bit_1/amux_2to1_2/SELB dac_8bit_1/c5m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7942 input_amplifier_0/txgate_6/txb input_amplifier_0/rst VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7943 dac_8bit_0/amux_2to1_2/B sample dac_8bit_0/c5m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7944 biquad_gm_c_filter_0/gm_c_stage_3/vcmc VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X7945 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn2 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn2 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7946 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 a_356329_n113250# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7947 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn vintp biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7948 VSS input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7949 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7950 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7951 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7952 dac_8bit_1/amux_2to1_4/B VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7953 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7954 adc_vcaparrayB dac_8bit_1/c1m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7955 vcp_sampled VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7956 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7957 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 a_275374_n146348# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7958 dac_8bit_1/ibiasp vbiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=2e+06u
X7959 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7960 dac_8bit_0/amux_2to1_4/B dac_8bit_0/amux_2to1_13/SELB vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7961 VSS biquad_gm_c_filter_0/ibiasn4 biquad_gm_c_filter_0/ibiasn4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X7962 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7963 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn1 vocm_filt biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7964 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7965 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7966 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7967 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7968 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7969 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7970 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7971 vrefB dac_8bit_1/amux_2to1_11/SELB dac_8bit_1/amux_2to1_6/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7972 sample_and_hold_1/vholdm vpeak_sampled sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X7973 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7974 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X7975 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7976 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7977 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7978 diff_to_se_converter_0/rst rst_n VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7979 VDD pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/D a_336955_n185409# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7980 dac_8bit_1/c5m sample dac_8bit_1/amux_2to1_2/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7981 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X7982 a_222396_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin a_221938_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X7983 a_244783_n122799# a_244617_n122799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7984 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X7985 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7986 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7987 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7988 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7989 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7990 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7991 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7992 input_amplifier_0/diff_fold_casc_ota_0/M6d input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7993 input_amplifier_0/diff_fold_casc_ota_0/vcascnp input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7994 vcp_sampled sample sample_and_hold_0/vholdm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7995 VDD low_freq_pll_0/freq_div_0/vout a_238627_n115125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7996 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/vcom_buf VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7997 dac_8bit_1/amux_2to1_1/B VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7998 a_243020_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_243478_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X7999 vcp_sampled VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8000 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8001 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8002 vlowA q5A dac_8bit_0/amux_2to1_2/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8003 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8004 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 a_356329_n164260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8005 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8006 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8007 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8008 dac_8bit_0/amux_2to1_1/B dac_8bit_0/amux_2to1_16/SELB vrefA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8009 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8010 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8011 peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8012 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn2 vocm_filt biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8013 vrefB dac_8bit_1/amux_2to1_14/SELB dac_8bit_1/amux_2to1_3/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8014 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8015 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8016 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8017 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8018 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8019 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8020 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8021 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X8022 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8023 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8024 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X8025 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8026 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8027 a_336537_n185243# a_336408_n184969# a_336116_n185269# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8028 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8029 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8030 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8031 a_242273_n123343# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8032 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn vintm biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8033 input_amplifier_0/txgate_7/txb input_amplifier_0/rst VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8034 input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vbias3 a_163060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8035 VDD VDD vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8036 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8037 adc_vcaparrayA dac_8bit_0/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8038 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8039 dac_8bit_0/amux_2to1_0/B VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8040 a_336336_n185421# a_335844_n185460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8041 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8042 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8043 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8044 VSS comparator_0/vmirror comparator_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8045 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8046 input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8047 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8048 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X8049 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8050 a_238872_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_238414_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X8051 input_amplifier_0/diff_fold_casc_ota_1/M6d input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8052 VSS VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8053 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8054 low_freq_pll_0/pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/Q_N a_240447_n115125# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8055 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8056 vrefB dac_8bit_1/amux_2to1_17/SELB dac_8bit_1/amux_2to1_0/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8057 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 a_230446_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8058 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8059 biquad_gm_c_filter_0/ibiasn3 biquad_gm_c_filter_0/ibiasn3 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X8060 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8061 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X8062 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1.2e+07u w=2e+06u
X8063 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8064 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8065 comparator_0/vmirror comparator_0/vmirror comparator_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8066 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8067 a_225730_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_226188_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X8068 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1.2e+07u w=2e+06u
X8069 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8070 input_amplifier_0/ibiasn1 input_amplifier_0/ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8071 VDD input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vfoldm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8072 input_amplifier_0/diff_fold_casc_ota_1/M6d input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8073 input_amplifier_0/diff_fold_casc_ota_1/vcascnp input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8074 input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8075 a_383508_n101129# adc_compA dac_8bit_0/comp_outm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8076 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8077 a_237854_n132168# vcp a_237396_n132168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X8078 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8079 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8080 VDD vbiasp biquad_gm_c_filter_0/ibiasn4 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X8081 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8082 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X8083 VDD VDD vcp_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8084 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8085 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8086 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8087 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8088 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8089 VSS VSS low_freq_pll_0/pfd_cp_lpf_0/vndiode VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8090 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8091 VDD low_freq_pll_0/pfd_cp_lpf_0/vpbias low_freq_pll_0/pfd_cp_lpf_0/vswitchh VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X8092 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8093 input_amplifier_0/venm1 gain_ctrl_0 input_amplifier_0/vip2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8094 vintm vintm biquad_gm_c_filter_0/gm_c_stage_1/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8095 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8096 biquad_gm_c_filter_0/gm_c_stage_3/vtail_diff vintm vfiltm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8097 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8098 a_229702_n119618# vcp a_229244_n119618# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X8099 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8100 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8101 dac_8bit_0/latched_comparator_folded_0/vcompmb dac_8bit_0/latched_comparator_folded_0/vcompm VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8102 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8103 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8104 VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8105 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X8106 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8107 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X8108 VSS VSS biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X8109 adc_vcaparrayA dac_8bit_0/c2m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8110 comparator_0/ibiasn vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X8111 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8112 VSS input_amplifier_0/ibiasn2 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8113 a_335507_n185243# pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8114 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X8115 a_239708_n115125# a_238793_n115125# a_239361_n114883# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8116 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8117 a_242526_n121193# a_242358_n121167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X8118 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8119 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8120 biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail1 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X8121 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8122 a_223414_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_223872_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X8123 VDD VDD input_amplifier_0/diff_fold_casc_ota_1/M6d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8124 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8125 a_242085_n122249# a_241919_n122249# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8126 dac_8bit_1/amux_2to1_7/B sample dac_8bit_1/c1m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8127 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8128 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8129 input_amplifier_0/diff_fold_casc_ota_0/M1d input_amplifier_0/diff_fold_casc_ota_0/M1d input_amplifier_0/diff_fold_casc_ota_0/M1d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8130 vpeak_sampled vpeak_sampled vpeak_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8131 a_242526_n120511# a_242358_n120257# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8132 input_amplifier_0/venm2 input_amplifier_0/vip2 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X8133 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8134 a_242783_n121167# a_242085_n121161# a_242526_n121193# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8135 input_amplifier_0/diff_fold_casc_ota_0/vcascnp input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/vop1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8136 VSS peak_detector_0/verr sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X8137 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8138 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X8139 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X8140 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8141 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8142 VSS a_242575_n114888# a_242506_n114759# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8143 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8144 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8145 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X8146 vrefA dac_8bit_0/amux_2to1_11/SELB dac_8bit_0/amux_2to1_6/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8147 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8148 vampm input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8149 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8150 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X8151 VDD a_245481_n121167# a_245649_n121193# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8152 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8153 comparator_0/vtail vfiltm comparator_0/vcompp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8154 vlowA VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8155 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8156 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8157 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8158 input_amplifier_0/txgate_1/txb gain_ctrl_0 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8159 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8160 dac_8bit_1/amux_2to1_4/B sample dac_8bit_1/c3m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8161 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8162 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8163 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8164 a_245565_n121167# a_244783_n121161# a_245481_n121167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8165 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8166 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8167 low_freq_pll_0/pfd_cp_lpf_0/vpbias low_freq_pll_0/ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X8168 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8169 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8170 dac_8bit_0/amux_2to1_5/B q2A vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8171 vpeak_sampled VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8172 vlowB q1B dac_8bit_1/amux_2to1_7/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8173 VSS vpeak sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X8174 vcp_sampled vcp_sampled VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8175 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X8176 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 a_275374_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8177 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 a_163060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8178 dac_8bit_1/amux_2to1_6/B dac_8bit_1/amux_2to1_11/SELB vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8179 vrefA dac_8bit_0/amux_2to1_14/SELB dac_8bit_0/amux_2to1_3/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8180 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X8181 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8182 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8183 a_336784_n185787# a_336537_n185409# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8184 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8185 sample_and_hold_0/vhold sample vcp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8186 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8187 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8188 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8189 vlowB dac_8bit_1/adc_run adc_vcaparrayB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8190 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8191 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8192 adc_vcaparrayB dac_8bit_1/c3m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8193 dac_8bit_1/amux_2to1_1/B sample dac_8bit_1/c6m VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8194 VSS dac_8bit_1/ibiasn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8195 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8196 VDD peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8197 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8198 dac_8bit_0/amux_2to1_2/B q5A vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8199 dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8200 vpeak_sampled VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8201 vlowB q3B dac_8bit_1/amux_2to1_4/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8202 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc vampm input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X8203 a_162668_n147576# diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8204 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8205 VSS VSS dac_8bit_0/latched_comparator_folded_0/vlatchm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X8206 dac_8bit_1/amux_2to1_3/B dac_8bit_1/amux_2to1_14/SELB vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8207 VDD diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8208 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8209 a_236938_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_236480_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X8210 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin a_238770_n131500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X8211 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8212 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 a_275374_n146348# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8213 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X8214 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8215 adc_vcaparrayA dac_8bit_0/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8216 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8217 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8218 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8219 a_356329_n164260# dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8220 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 a_217060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8221 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8222 adc_vcaparrayB dac_8bit_1/c4m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8223 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8224 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8225 adc_vcaparrayA dac_8bit_0/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8226 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/vcom_buf VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8227 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X8228 a_221939_n130007# low_freq_pll_0/cs_ring_osc_0/vosc a_221481_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X8229 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8230 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8231 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8232 a_242085_n121161# a_241919_n121161# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8233 dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8234 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X8235 VDD input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vfoldm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8236 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8237 a_338356_n185510# a_338156_n185665# a_338505_n185421# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8238 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8239 vlowB q6B dac_8bit_1/amux_2to1_1/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8240 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8241 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8242 VSS dac_8bit_0/vcom_buf sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X8243 input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X8244 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/diff_fold_casc_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8245 vpeak vpeak vpeak VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8246 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8247 input_amplifier_0/vom1 input_amplifier_0/vip1 sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X8248 input_amplifier_0/diff_fold_casc_ota_0/vcascnp input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/vop1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8249 low_freq_pll_0/ibiasn low_freq_pll_0/ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X8250 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8251 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8252 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8253 VDD VDD vincm VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8254 VDD dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8255 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8256 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn2 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8257 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8258 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8259 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8260 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8261 a_356329_n113250# dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8262 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8263 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin a_223770_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X8264 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X8265 input_amplifier_0/ibiasn2 input_amplifier_0/ibiasn2 input_amplifier_0/ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8266 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8267 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8268 dac_8bit_1/c7m dac_8bit_1/amux_2to1_0/SELB dac_8bit_1/amux_2to1_0/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8269 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8270 dac_8bit_0/c1m sample dac_8bit_0/amux_2to1_7/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8271 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=2e+06u
X8272 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8273 VDD pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/D a_336955_n185243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8274 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/vim2 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X8275 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_2/A a_243382_n122255# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8276 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8277 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8278 a_356329_n164260# dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8279 vincm input_amplifier_0/rst input_amplifier_0/vip1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8280 input_amplifier_0/vip1 vhpf sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X8281 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8282 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q a_242951_n121193# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8283 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8284 vse diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8285 a_225869_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_225411_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X8286 a_383050_n101129# dac_8bit_0/latched_comparator_folded_0/vcompm_buf VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8287 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8288 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8289 VSS input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8290 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8291 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 a_163060_n102324# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8292 VDD vbiasp biquad_gm_c_filter_0/ibiasn1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X8293 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8294 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8295 input_amplifier_0/vim2 input_amplifier_0/txgate_6/txb input_amplifier_0/vop1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8296 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8297 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8298 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8299 a_227854_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_227396_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X8300 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8301 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 a_356329_n164260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8302 dac_8bit_0/c3m sample dac_8bit_0/amux_2to1_4/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8303 a_242358_n123343# a_242085_n123337# a_242273_n123343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8304 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8305 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8306 input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X8307 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8308 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8309 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8310 vlowA q1A dac_8bit_0/amux_2to1_7/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8311 VSS dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8312 input_amplifier_0/vim2 input_amplifier_0/rst input_amplifier_0/vop1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8313 dac_8bit_0/latched_comparator_folded_0/vlatchm vlowA dac_8bit_0/latched_comparator_folded_0/vtailp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8314 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X8315 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X8316 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8317 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8318 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8319 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8320 vrefB dac_8bit_1/amux_2to1_9/SELB dac_8bit_1/amux_2to1_9/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8321 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8322 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_8/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8323 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8324 VDD a_245481_n122433# a_245649_n122531# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8325 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8326 VSS comparator_0/ibiasn comparator_0/ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X8327 VSS sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8328 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8329 adc_vcaparrayA dac_8bit_0/adc_run vlowA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8330 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8331 input_amplifier_0/venp1 input_amplifier_0/txgate_1/txb input_amplifier_0/vim2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8332 VDD low_freq_pll_0/pfd_cp_lpf_0/vpbias low_freq_pll_0/pfd_cp_lpf_0/vpbias VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X8333 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8334 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8335 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8336 a_227397_n130007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_226939_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X8337 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8338 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X8339 dac_8bit_0/c6m sample dac_8bit_0/amux_2to1_1/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8340 VSS VSS vintm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8341 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X8342 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8343 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8344 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8345 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8346 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8347 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8348 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn vfiltp biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8349 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8350 dac_8bit_1/amux_2to1_7/B q1B vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8351 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8352 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X8353 dac_8bit_0/amux_2to1_9/SELB q0A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8354 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8355 vlowA VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8356 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8357 vlowA q3A dac_8bit_0/amux_2to1_4/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8358 VSS biquad_gm_c_filter_0/ibiasn2 biquad_gm_c_filter_0/ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X8359 a_245224_n123369# a_245056_n123343# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X8360 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8361 input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/M3d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8362 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8363 a_226646_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias a_226188_n140786# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X8364 adc_vcaparrayB dac_8bit_1/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8365 vrefA VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8366 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8367 peak_detector_0/verr peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8368 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 vpeak_sampled VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8369 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8370 a_245481_n123343# a_244783_n123337# a_245224_n123369# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8371 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8372 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X8373 a_336401_n185269# adc_clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8374 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8375 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8376 a_275374_n146348# sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8377 a_221582_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias a_222040_n145742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X8378 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8379 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8380 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8381 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8382 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X8383 dac_8bit_1/amux_2to1_4/B q3B vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8384 peak_detector_0/ibiasn2 peak_detector_0/ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8385 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8386 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8387 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X8388 a_245224_n121599# a_245056_n121345# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X8389 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8390 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X8391 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8392 vlowA q6A dac_8bit_0/amux_2to1_1/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8393 VSS input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8394 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8395 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8396 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8397 VSS input_amplifier_0/ibiasn2 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8398 VSS peak_detector_0/vpeak sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X8399 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8400 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8401 a_225412_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_224954_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X8402 vpeak sample sample_and_hold_1/vhold VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8403 peak_detector_0/verr peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8404 vrefA VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8405 VSS a_242526_n121599# a_242484_n121711# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8406 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 a_356329_n113250# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8407 adc_vcaparrayA dac_8bit_0/c2m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8408 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8409 dac_8bit_0/ibiasn dac_8bit_0/ibiasn dac_8bit_0/ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8410 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8411 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8412 adc_vcaparrayB adc_vcaparrayB sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8413 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn2 vocm_filt biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8414 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8415 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8416 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8417 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8418 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8419 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 a_275374_n180872# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8420 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8421 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8422 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8423 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8424 VSS biquad_gm_c_filter_0/ibiasn3 biquad_gm_c_filter_0/ibiasn3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X8425 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X8426 VSS peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8427 vrefB dac_8bit_1/amux_2to1_15/SELB dac_8bit_1/amux_2to1_2/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8428 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8429 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8430 a_239954_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X8431 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8432 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8433 dac_8bit_1/amux_2to1_1/B q6B vlowB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8434 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8435 input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8436 VSS low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8437 a_236633_n122049# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout a_236175_n122049# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X8438 input_amplifier_0/diff_fold_casc_ota_0/M13d input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/M6d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8439 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8440 VSS input_amplifier_0/ibiasn1 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8441 input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/diff_fold_casc_ota_0/M2d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8442 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 vocm input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X8443 diff_to_se_converter_0/vim vfiltm sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=8e+06u
X8444 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8445 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8446 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8447 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8448 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8449 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8450 VDD VDD peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8451 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8452 VDD a_245481_n121345# a_245649_n121443# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8453 VSS input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8454 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8455 low_freq_pll_0/pfd_cp_lpf_0/vpbias VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X8456 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8457 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8458 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8459 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8460 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8461 a_336784_n184877# a_336537_n185243# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8462 VSS a_245224_n123369# a_245182_n122965# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8463 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8464 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8465 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X8466 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8467 VDD input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/M6d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8468 vintp vintp biquad_gm_c_filter_0/gm_c_stage_1/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8469 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8470 a_236023_n130007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X8471 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8472 peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8473 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8474 a_230446_n180872# peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8475 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8476 dac_8bit_0/latched_comparator_folded_0/vlatchp adc_clk dac_8bit_0/latched_comparator_folded_0/vlatchm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X8477 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8478 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8479 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8480 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q a_242951_n122531# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8481 input_amplifier_0/vip1 input_amplifier_0/txgate_5/txb vincm VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8482 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8483 input_amplifier_0/diff_fold_casc_ota_1/M2d input_amplifier_0/diff_fold_casc_ota_1/M2d input_amplifier_0/diff_fold_casc_ota_1/M2d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8484 adc_vcaparrayB dac_8bit_1/c2m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8485 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8486 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8487 dac_8bit_0/ibiasn dac_8bit_0/ibiasn dac_8bit_0/ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8488 a_227244_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_226786_n135628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X8489 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X8490 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8491 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8492 input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8493 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8494 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1.2e+07u
X8495 a_275374_n180872# sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8496 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8497 VDD a_242526_n121193# a_242453_n121167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8498 a_242885_n115125# a_242506_n114759# a_242813_n115125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8499 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8500 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8501 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8502 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8503 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8504 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 vse VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8505 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8506 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8507 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8508 a_238312_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_237854_n149500# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X8509 dac_8bit_1/cdumm sample dac_8bit_1/amux_2to1_6/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8510 a_225411_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_224953_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X8511 input_amplifier_0/diff_fold_casc_ota_1/M13d input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/M6d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8512 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8513 dac_8bit_0/cdumm dac_8bit_0/amux_2to1_6/SELB vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8514 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8515 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8516 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8517 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8518 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8519 adc_vcaparrayB dac_8bit_1/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8520 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8521 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8522 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8523 adc_vcaparrayA dac_8bit_0/c5m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8524 biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail1 vocm_filt biquad_gm_c_filter_0/gm_c_stage_0/vcmcn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8525 VSS biquad_gm_c_filter_0/gm_c_stage_2/vcmc biquad_gm_c_filter_0/gm_c_stage_2/vtail_diff VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X8526 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8527 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8528 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8529 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8530 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8531 a_221023_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X8532 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X8533 vfiltm diff_to_se_converter_0/txgate_1/txb diff_to_se_converter_0/vim VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8534 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8535 a_239953_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X8536 a_223313_n130007# low_freq_pll_0/cs_ring_osc_0/vosc a_222855_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X8537 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8538 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8539 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8540 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8541 a_238793_n115125# a_238627_n115125# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8542 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X8543 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X8544 a_242358_n121167# a_241919_n121161# a_242273_n121167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8545 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8546 a_356329_n164260# dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8547 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8548 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 vpeak VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8549 VSS VSS low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X8550 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8551 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8552 dac_8bit_1/c4m sample dac_8bit_1/amux_2to1_3/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8553 vrefA dac_8bit_0/amux_2to1_12/SELB dac_8bit_0/amux_2to1_5/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8554 VSS dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8555 dac_8bit_0/c4m dac_8bit_0/amux_2to1_3/SELB vcp_sampled VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8556 dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8557 vlowA VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8558 dac_8bit_0/latched_comparator_folded_0/vlatchm vlowA dac_8bit_0/latched_comparator_folded_0/vtailp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8559 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8560 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/M2d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8561 vlowB VSS dac_8bit_1/amux_2to1_6/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8562 VDD sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8563 VSS input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8564 VDD a_336608_n185510# a_336537_n185409# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X8565 adc_vcaparrayA dac_8bit_0/c7m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8566 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2e+06u
X8567 VSS sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8568 vrefB VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8569 VDD VDD adc_vcaparrayB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8570 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8571 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8572 diff_to_se_converter_0/vim VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8573 vpeak_sampled VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8574 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8575 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8576 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=8e+06u
X8577 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 a_162668_n147576# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8578 dac_8bit_1/amux_2to1_5/B dac_8bit_1/amux_2to1_12/SELB vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8579 a_242909_n121711# a_241919_n121711# a_242783_n121345# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8580 biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail1 vintp biquad_gm_c_filter_0/gm_c_stage_2/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8581 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8582 vrefA dac_8bit_0/amux_2to1_15/SELB dac_8bit_0/amux_2to1_2/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8583 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8584 VSS input_amplifier_0/ibiasn2 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8585 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8586 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8587 a_227243_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_226785_n138121# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X8588 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M3d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8589 peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8590 dac_8bit_1/amux_2to1_0/B dac_8bit_1/amux_2to1_17/SELB vlowB VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8591 dac_8bit_0/ibiasn vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=4e+06u
X8592 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8593 vlowA VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8594 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8595 vlowB q4B dac_8bit_1/amux_2to1_3/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8596 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8597 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8598 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=800000u
X8599 a_242358_n122433# a_242085_n122799# a_242273_n122799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8600 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q a_242951_n121443# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8601 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8602 adc_vcaparrayA adc_vcaparrayA sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8603 input_amplifier_0/ibiasn1 input_amplifier_0/ibiasn1 input_amplifier_0/ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8604 VSS input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8605 vse vse vse VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8606 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8607 dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8608 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8609 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8610 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/vbias2 vampm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8611 a_356329_n113250# dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8612 vpeak_sampled VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8613 biquad_gm_c_filter_0/ibiasn4 biquad_gm_c_filter_0/ibiasn4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X8614 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/vim1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=1.2e+06u
X8615 vampm VSS sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X8616 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8617 a_217060_n102324# input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8618 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8619 dac_8bit_1/amux_2to1_2/B dac_8bit_1/amux_2to1_15/SELB vrefB VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8620 VSS peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8621 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8622 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8623 VDD dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8624 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8625 sample_and_hold_0/vholdm sample vcp_sampled VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8626 a_237040_n127742# low_freq_pll_0/cs_ring_osc_0/vpbias a_237498_n127742# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X8627 adc_vcaparrayB dac_8bit_1/c6m sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
X8628 a_226939_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_226481_n148007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X8629 VSS diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8630 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_228771_n130007# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
C0 vpeak_sampled dac_8bit_1/c5m 1.94fF
C1 sample dac_8bit_1/amux_2to1_9/Y 2.66fF
C2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/vholdm 10.10fF
C3 low_freq_pll_0/pfd_cp_lpf_0/vQAb low_freq_pll_0/pfd_cp_lpf_0/vQB 0.05fF
C4 diff_to_se_converter_0/ibiasn rst_n 6.55fF
C5 dac_8bit_1/amux_2to1_0/SELB VDD 1.15fF
C6 a_337592_n185269# a_338356_n185269# 0.02fF
C7 a_337864_n185269# a_338149_n185269# 0.09fF
C8 sample dac_8bit_0/amux_2to1_0/B 2.60fF
C9 a_242783_n123343# a_242085_n122799# 0.01fF
C10 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d 15.11fF
C11 a_231328_n134960# vcp 0.03fF
C12 vampp input_amplifier_0/venp2 7.13fF
C13 comparator_0/ibiasn comparator_0/vtail 4.69fF
C14 biquad_gm_c_filter_0/gm_c_stage_0/vbiasp biquad_gm_c_filter_0/gm_c_stage_0/vcmcn 0.53fF
C15 a_243382_n121167# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/A 0.05fF
C16 low_freq_pll_0/cs_ring_osc_0/vpbias a_236582_n145742# 0.51fF
C17 a_242336_n114759# a_242102_n114873# 0.04fF
C18 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample 12.70fF
C19 vintm biquad_gm_c_filter_0/gm_c_stage_3/vcmcn 0.19fF
C20 dac_8bit_0/amux_2to1_5/SELB dac_8bit_0/c2m 1.59fF
C21 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/vholdm 19.15fF
C22 dac_8bit_0/amux_2to1_9/SELB VDD 1.15fF
C23 a_242358_n122255# a_242484_n121877# 0.02fF
C24 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_245649_n122281# 0.02fF
C25 a_338149_n185569# VDD 0.87fF
C26 dac_8bit_1/ibiasp dac_8bit_1/latched_comparator_folded_0/vlatchm 0.04fF
C27 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vbias1 0.55fF
C28 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d 1.74fF
C29 sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp 0.28fF
C30 a_222498_n145742# VDD 0.40fF
C31 a_242380_n114857# a_242506_n114759# 0.41fF
C32 gain_ctrl_1 VDD 0.48fF
C33 a_242419_n114983# a_242575_n114888# 0.42fF
C34 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 13.36fF
C35 a_242358_n121345# a_242951_n121443# 0.02fF
C36 a_242526_n121599# a_242783_n121345# 0.11fF
C37 vampm VDD 5.50fF
C38 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 0.04fF
C39 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 32.00fF
C40 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/vcom_buf 9.19fF
C41 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_239954_n135628# 0.03fF
C42 a_245056_n121345# a_244617_n122249# 0.01fF
C43 a_244617_n121711# a_245056_n122255# 0.01fF
C44 a_236582_n145742# a_238414_n145742# 0.65fF
C45 a_237040_n145742# a_237956_n145742# 2.26fF
C46 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d VDD 9.36fF
C47 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y a_242085_n123337# 0.61fF
C48 a_241919_n123337# a_242526_n123369# 0.37fF
C49 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc input_amplifier_0/vim1 8.59fF
C50 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/ibiasn1 1.61fF
C51 VDD a_241919_n123337# 0.79fF
C52 peak_detector_rst pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A 0.01fF
C53 input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vfoldm 3.26fF
C54 comparator_0/ibiasn vcp_sampled 0.55fF
C55 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d 6.93fF
C56 vrefA dac_8bit_0/amux_2to1_3/B 2.44fF
C57 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp 19.65fF
C58 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d 3.28fF
C59 low_freq_pll_0/cs_ring_osc_0/vosc low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/csinvn 0.09fF
C60 dac_8bit_0/ibiasn vbiasp 4.26fF
C61 vfiltm biquad_gm_c_filter_0/gm_c_stage_2/vtail_diff 0.33fF
C62 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/csinvn low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.09fF
C63 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VDD 2.04fF
C64 a_336784_n185787# a_336608_n185510# 0.04fF
C65 dac_8bit_0/amux_2to1_11/SELB VDD 1.15fF
C66 a_242783_n123343# a_242909_n122965# 0.04fF
C67 a_244617_n123337# a_245056_n122433# 0.01fF
C68 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/A 0.10fF
C69 input_amplifier_0/txgate_4/txb input_amplifier_0/vim1 0.35fF
C70 a_245056_n123343# a_244617_n122799# 0.01fF
C71 a_336784_n184877# VDD 0.02fF
C72 a_244617_n121161# a_244783_n121711# 0.09fF
C73 a_337497_n185813# a_336401_n185569# 0.07fF
C74 a_244783_n121161# a_244617_n121711# 0.09fF
C75 a_242085_n122799# VDD 0.43fF
C76 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp 12.50fF
C77 dac_8bit_0/c1m dac_8bit_0/c7m 2.24fF
C78 dac_8bit_0/c2m dac_8bit_0/c5m 1.02fF
C79 dac_8bit_0/cdumm dac_8bit_0/c6m 0.86fF
C80 sample dac_8bit_1/c1m 2.36fF
C81 a_242783_n123343# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q 0.04fF
C82 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout a_237090_n119618# 0.03fF
C83 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.02fF
C84 VDD input_amplifier_0/vop1 7.32fF
C85 a_238007_n122049# VDD 0.01fF
C86 dac_8bit_0/amux_2to1_17/SELB q7A 2.36fF
C87 vpeak vse 15.31fF
C88 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror 0.69fF
C89 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn1 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn2 0.17fF
C90 peak_detector_0/ibiasn1 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d 0.40fF
C91 vlowA dac_8bit_0/latched_comparator_folded_0/vlatchm 4.52fF
C92 gain_ctrl_0 input_amplifier_0/venp1 0.55fF
C93 dac_8bit_1/ibiasp adc_clk 3.87fF
C94 dac_8bit_1/latched_comparator_folded_0/vlatchm VDD 6.80fF
C95 input_amplifier_0/diff_fold_casc_ota_1/M2d vampp 14.54fF
C96 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm vpeak 24.37fF
C97 input_amplifier_0/vip2 input_amplifier_0/txgate_7/txb 0.59fF
C98 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 21.43fF
C99 input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vcascnm 16.60fF
C100 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vbias2 0.10fF
C101 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn 9.20fF
C102 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vcascnp 18.64fF
C103 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d 0.56fF
C104 biquad_gm_c_filter_0/gm_c_stage_0/vbiasp vintp 0.44fF
C105 VDD input_amplifier_0/txgate_5/txb 3.26fF
C106 input_amplifier_0/ibiasn1 low_freq_pll_0/ibiasn 0.22fF
C107 dac_8bit_0/amux_2to1_2/B VDD 4.57fF
C108 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn a_356329_n113250# 0.11fF
C109 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp 1.94fF
C110 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn biquad_gm_c_filter_0/gm_c_stage_2/vcmcn1 1.18fF
C111 biquad_gm_c_filter_0/gm_c_stage_2/vbiasp biquad_gm_c_filter_0/gm_c_stage_2/vcmcn2 0.88fF
C112 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/vcom_buf 16.56fF
C113 vcp a_247244_n134960# 0.03fF
C114 peak_detector_0/verr a_230446_n180872# 19.89fF
C115 a_225580_n122869# a_227412_n122869# 0.67fF
C116 a_226038_n122869# a_226954_n122869# 2.26fF
C117 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/B a_335749_n185269# 0.02fF
C118 low_freq_pll_0/pfd_cp_lpf_0/vRSTN a_242102_n114873# 0.57fF
C119 a_239708_n115125# low_freq_pll_0/pfd_cp_lpf_0/vQB 0.02fF
C120 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VDD 12.54fF
C121 a_241919_n121711# VDD 0.79fF
C122 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q a_242951_n122281# 0.02fF
C123 a_245056_n121345# a_245182_n121711# 0.02fF
C124 adc_vcaparrayB dac_8bit_1/ibiasp 35.67fF
C125 a_242484_n122965# a_242358_n123343# 0.02fF
C126 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc vocm 0.07fF
C127 a_242951_n120355# a_243382_n120301# 0.31fF
C128 biquad_gm_c_filter_0/ibiasn1 biquad_gm_c_filter_0/gm_c_stage_0/vbiasp 1.23fF
C129 dac_8bit_1/latched_comparator_folded_0/vcompp adc_compB 0.70fF
C130 peak_detector_0/ibiasn2 vfiltm 0.18fF
C131 input_amplifier_0/rst input_amplifier_0/diff_fold_casc_ota_0/vbias2 0.11fF
C132 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d 0.70fF
C133 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp 0.28fF
C134 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q a_242951_n123369# 0.02fF
C135 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q VDD 1.02fF
C136 a_245056_n122433# a_245151_n122433# 0.04fF
C137 a_238872_n127742# VDD 0.09fF
C138 a_237396_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.03fF
C139 a_242336_n114759# VDD 0.01fF
C140 vcp a_237396_n132168# 0.03fF
C141 a_338149_n185569# a_338703_n185409# 0.21fF
C142 a_337864_n185555# a_338107_n185787# 0.05fF
C143 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 input_amplifier_0/ibiasn1 3.91fF
C144 peak_detector_0/ibiasn1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp 0.16fF
C145 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d 1.84fF
C146 a_275374_n146348# sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp 10.36fF
C147 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d 1.13fF
C148 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q VDD 2.18fF
C149 a_337592_n185460# a_337864_n185555# 0.67fF
C150 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin a_223312_n149500# 0.03fF
C151 vintp biquad_gm_c_filter_0/gm_c_stage_2/vcmcn 1.12fF
C152 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 adc_vcaparrayA 0.08fF
C153 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/A VDD 0.62fF
C154 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_226023_n130007# 0.03fF
C155 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm 0.08fF
C156 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror 4.50fF
C157 input_amplifier_0/venp2 input_amplifier_0/vim2 43.85fF
C158 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y a_243382_n122477# 0.11fF
C159 a_245151_n121345# VDD 0.02fF
C160 adc_clk VDD 7.70fF
C161 dac_8bit_1/c7m dac_8bit_1/c5m 1.37fF
C162 input_amplifier_0/rst vocm 0.65fF
C163 low_freq_pll_0/cs_ring_osc_0/vpbias a_227104_n140786# 0.83fF
C164 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/A 1.66fF
C165 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp 11.53fF
C166 a_242358_n121167# a_242783_n121167# 0.03fF
C167 input_amplifier_0/diff_fold_casc_ota_1/vfoldp vampp 0.18fF
C168 dac_8bit_0/c3m dac_8bit_0/ibiasn 0.19fF
C169 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp 19.65fF
C170 input_amplifier_0/diff_fold_casc_ota_1/vcascnm a_163060_n102324# 9.83fF
C171 diff_to_se_converter_0/ibiasn diff_to_se_converter_0/vim 3.75fF
C172 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d 3.28fF
C173 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/vom1 5.16fF
C174 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc 6.63fF
C175 dac_8bit_0/c1m adc_vcaparrayA 18.08fF
C176 dac_8bit_0/c3m dac_8bit_0/ibiasp 0.26fF
C177 a_245056_n121167# a_245182_n120789# 0.02fF
C178 biquad_gm_c_filter_0/ibiasn3 diff_to_se_converter_0/ibiasn 19.23fF
C179 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d 10.82fF
C180 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/A VDD 0.62fF
C181 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d vpeak 15.32fF
C182 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d 2.62fF
C183 vintm biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail1 0.07fF
C184 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_243313_n148007# 0.03fF
C185 dac_8bit_0/c6m VDD 2.50fF
C186 a_241919_n121711# a_242526_n121599# 0.37fF
C187 comparator_0/vcompp comparator_0/vtail 0.30fF
C188 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y a_242085_n121711# 0.61fF
C189 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn 0.61fF
C190 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 12.94fF
C191 dac_8bit_1/amux_2to1_0/B q7B 1.99fF
C192 dac_8bit_1/ibiasn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 0.18fF
C193 adc_vcaparrayB VDD 3.82fF
C194 a_336116_n185269# a_336336_n185243# 0.04fF
C195 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A a_336401_n185269# 0.03fF
C196 sample sample_and_hold_0/vholdm 0.82fF
C197 vampp input_amplifier_0/txgate_3/txb 0.36fF
C198 a_238627_n115125# a_238793_n115125# 1.60fF
C199 vampp vocm 1.32fF
C200 vfiltp biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail1 2.83fF
C201 input_amplifier_0/rst input_amplifier_0/vom1 11.10fF
C202 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_2/Q VDD 0.28fF
C203 dac_8bit_1/amux_2to1_1/B q6B 1.99fF
C204 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y a_244971_n123343# 0.38fF
C205 biquad_gm_c_filter_0/ibiasn3 vbiasp 3.72fF
C206 biquad_gm_c_filter_0/ibiasn2 input_amplifier_0/ibiasn1 0.18fF
C207 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias3 0.02fF
C208 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d 0.12fF
C209 a_239251_n114759# VDD 0.27fF
C210 a_242867_n122255# VDD 0.02fF
C211 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vcascnp 18.64fF
C212 input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vcascnm 16.60fF
C213 dac_8bit_1/c1m dac_8bit_1/amux_2to1_7/B 1.72fF
C214 q7A vrefA 0.88fF
C215 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_240869_n138121# 0.03fF
C216 a_226038_n122869# low_freq_pll_0/cs_ring_osc_0/vpbias 0.66fF
C217 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp 0.81fF
C218 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp 13.60fF
C219 low_freq_pll_0/pfd_cp_lpf_0/vRSTN VDD 2.28fF
C220 a_244617_n121711# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y 0.04fF
C221 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d 3.07fF
C222 vampp input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc 4.23fF
C223 dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 8.87fF
C224 a_241022_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs 0.03fF
C225 vpeak_sampled VDD 20.42fF
C226 a_225730_n140786# VDD 0.73fF
C227 input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc vampp 0.86fF
C228 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp 6.59fF
C229 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d 5.99fF
C230 a_245224_n122281# a_244971_n122255# 0.04fF
C231 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d 14.22fF
C232 vse diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d 9.65fF
C233 vintm biquad_gm_c_filter_0/gm_c_stage_1/vcmcn 1.20fF
C234 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_3/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/A 0.35fF
C235 vpeak_sampled dac_8bit_1/amux_2to1_3/SELB 2.07fF
C236 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin a_247702_n135628# 0.03fF
C237 low_freq_pll_0/pfd_cp_lpf_0/vQAb a_241634_n115151# 0.04fF
C238 low_freq_pll_0/cs_ring_osc_0/vpbias a_224330_n127742# 0.77fF
C239 low_freq_pll_0/cs_ring_osc_0/vosc a_222397_n130007# 0.03fF
C240 diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 2.30fF
C241 a_338285_n185409# pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A 0.05fF
C242 a_245481_n121345# a_245481_n122255# 0.07fF
C243 vlowB q0B 2.75fF
C244 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_243382_n120301# 0.37fF
C245 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror 1.41fF
C246 biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail1 biquad_gm_c_filter_0/gm_c_stage_1/vtail_diff 0.49fF
C247 gain_ctrl_0 input_amplifier_0/txgate_1/txb 0.48fF
C248 peak_detector_0/ibiasn1 vcp_sampled 3.90fF
C249 vfiltm biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail2 0.32fF
C250 a_338703_n185409# adc_clk 0.05fF
C251 rst_n input_amplifier_0/vop1 3.30fF
C252 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y a_242951_n120355# 0.17fF
C253 a_241919_n120623# a_242783_n120257# 0.09fF
C254 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_244617_n121711# 0.49fF
C255 a_337497_n185813# adc_clk 0.12fF
C256 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/vtail_casc 10.25fF
C257 diff_to_se_converter_0/ibiasn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 0.18fF
C258 a_245481_n123343# a_245481_n122433# 0.07fF
C259 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y 0.01fF
C260 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/A 0.01fF
C261 a_245649_n121193# a_245649_n121443# 0.09fF
C262 vpeak_sampled dac_8bit_1/amux_2to1_5/B 0.38fF
C263 low_freq_pll_0/pfd_cp_lpf_0/VQBb low_freq_pll_0/pfd_cp_lpf_0/vpdiode 0.10fF
C264 a_245870_n134960# vcp 0.03fF
C265 input_amplifier_0/diff_fold_casc_ota_0/vcascnm a_217060_n102324# 9.83fF
C266 a_245649_n122281# VDD 0.45fF
C267 vcp low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin 4.16fF
C268 dac_8bit_0/c4m dac_8bit_0/amux_2to1_3/B 1.72fF
C269 sample_and_hold_1/vhold VDD 0.64fF
C270 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A a_337592_n185269# 0.03fF
C271 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y a_246080_n121167# 0.11fF
C272 dac_8bit_1/c2m dac_8bit_1/c0m 0.39fF
C273 dac_8bit_1/cdumm dac_8bit_1/c1m 1.32fF
C274 a_242358_n122433# a_242453_n122433# 0.04fF
C275 a_242526_n122281# VDD 0.23fF
C276 a_242273_n120623# a_242273_n121167# 0.02fF
C277 a_242273_n120623# VDD 0.15fF
C278 peak_detector_0/verr VDD 6.63fF
C279 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/csinvp a_242562_n140786# 0.10fF
C280 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y a_242526_n121193# 0.15fF
C281 a_242085_n120623# VDD 0.43fF
C282 a_336608_n185510# VDD 0.36fF
C283 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/vim2 3.57fF
C284 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD 1.49fF
C285 adc_vcaparrayB dac_8bit_1/c3m 29.30fF
C286 a_244783_n122249# a_245224_n122281# 0.28fF
C287 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm 23.84fF
C288 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d 1.84fF
C289 low_freq_pll_0/pfd_cp_lpf_0/vQA a_242102_n114873# 0.02fF
C290 a_245224_n121193# VDD 0.23fF
C291 input_amplifier_0/txgate_6/txb input_amplifier_0/rst 0.36fF
C292 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/csinvp low_freq_pll_0/cs_ring_osc_0/vpbias 0.31fF
C293 dac_8bit_1/amux_2to1_1/B VDD 4.57fF
C294 sample vlowB 4.89fF
C295 a_222956_n127742# VDD 0.69fF
C296 a_337497_n185813# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_2/Q 0.37fF
C297 sample dac_8bit_1/amux_2to1_8/SELB 2.36fF
C298 sample pulse_generator_0/sky130_fd_sc_hd__inv_1_0/Y 0.16fF
C299 a_336408_n184969# VDD 0.45fF
C300 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 21.43fF
C301 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/Q_N pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/B 0.24fF
C302 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d 16.02fF
C303 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y a_243382_n122255# 0.11fF
C304 q6A vlowA 2.75fF
C305 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VDD 11.66fF
C306 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q a_242951_n121443# 0.02fF
C307 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm 0.08fF
C308 input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/diff_fold_casc_ota_0/M1d 8.30fF
C309 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_3/A VDD 0.48fF
C310 sample dac_8bit_0/amux_2to1_0/SELB 2.37fF
C311 input_amplifier_0/vip2 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc 3.62fF
C312 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d 0.04fF
C313 dac_8bit_1/amux_2to1_2/SELB dac_8bit_1/amux_2to1_2/B 1.51fF
C314 low_freq_pll_0/cs_ring_osc_0/vosc vcp 5.08fF
C315 dac_8bit_0/latched_comparator_folded_0/vcompp VDD 6.16fF
C316 a_227562_n140786# a_228478_n140786# 0.79fF
C317 input_amplifier_0/venm1 VDD 1.10fF
C318 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 0.08fF
C319 biquad_gm_c_filter_0/ibiasn3 biquad_gm_c_filter_0/gm_c_stage_3/vtail_diff 0.06fF
C320 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vbias4 36.08fF
C321 input_amplifier_0/rst input_amplifier_0/diff_fold_casc_ota_0/M13d 0.11fF
C322 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias3 60.63fF
C323 vocm input_amplifier_0/vim2 0.14fF
C324 input_amplifier_0/diff_fold_casc_ota_1/M13d input_amplifier_0/diff_fold_casc_ota_1/vtail_casc 0.04fF
C325 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vbias3 0.04fF
C326 VDD a_245056_n122433# 0.36fF
C327 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vtail_casc 1.56fF
C328 a_336116_n185555# a_336401_n185569# 0.09fF
C329 biquad_gm_c_filter_0/gm_c_stage_2/vbiasp VDD 3.04fF
C330 a_335844_n185460# a_336408_n185665# 0.11fF
C331 a_243382_n123343# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y 0.11fF
C332 a_245224_n123369# a_245649_n123369# 0.04fF
C333 a_241919_n121161# a_242358_n121345# 0.02fF
C334 a_244783_n123337# a_245481_n123343# 0.44fF
C335 biquad_gm_c_filter_0/ibiasn2 vfiltp 0.19fF
C336 q0A dac_8bit_1/ibiasp 0.02fF
C337 vpeak_sampled dac_8bit_1/c3m 1.94fF
C338 a_242526_n122281# a_242526_n121599# 0.05fF
C339 a_236582_n127742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/csinvp 0.08fF
C340 a_237956_n127742# a_238414_n127742# 0.02fF
C341 a_242085_n122249# a_242358_n122255# 0.38fF
C342 a_338156_n184969# a_338356_n185269# 0.38fF
C343 a_337864_n185269# a_338285_n185243# 0.11fF
C344 a_232244_n134960# vcp 0.03fF
C345 dac_8bit_1/amux_2to1_0/B dac_8bit_1/amux_2to1_17/SELB 1.59fF
C346 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y 0.03fF
C347 dac_8bit_0/c5m dac_8bit_0/c4m 1.41fF
C348 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD 7.64fF
C349 a_383508_n152139# dac_8bit_1/comp_outm 0.05fF
C350 q6B dac_8bit_1/amux_2to1_16/SELB 2.36fF
C351 a_244783_n122249# a_244783_n122799# 0.05fF
C352 input_amplifier_0/diff_fold_casc_ota_0/vbias4 vocm 0.69fF
C353 low_freq_pll_0/cs_ring_osc_0/vpbias a_237498_n145742# 0.63fF
C354 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn2 VDD 1.51fF
C355 a_240730_n140786# a_241646_n140786# 2.99fF
C356 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 33.98fF
C357 a_242720_n114759# a_242102_n114873# 0.01fF
C358 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d 2.72fF
C359 dac_8bit_0/comp_outm a_383508_n101129# 0.05fF
C360 adc_clk pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.19fF
C361 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VDD 12.54fF
C362 input_amplifier_0/vom1 input_amplifier_0/vim2 4.56fF
C363 a_338356_n185510# VDD 0.36fF
C364 a_242085_n121161# a_242085_n121711# 0.05fF
C365 a_223414_n145742# VDD 0.14fF
C366 input_amplifier_0/diff_fold_casc_ota_1/M2d input_amplifier_0/diff_fold_casc_ota_1/M1d 8.30fF
C367 a_242575_n114888# a_242506_n114759# 0.50fF
C368 a_242951_n121443# a_242783_n121345# 0.67fF
C369 dac_8bit_0/ibiasn dac_8bit_0/c6m 0.19fF
C370 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_240870_n135628# 0.03fF
C371 dac_8bit_1/c7m VDD 2.60fF
C372 dac_8bit_0/ibiasp dac_8bit_0/c6m 0.26fF
C373 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A a_335844_n185269# 0.44fF
C374 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/M6d 1.84fF
C375 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD 19.81fF
C376 input_amplifier_0/diff_fold_casc_ota_0/M1d input_amplifier_0/diff_fold_casc_ota_0/vfoldp 6.26fF
C377 input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/diff_fold_casc_ota_0/vbias2 1.06fF
C378 dac_8bit_0/amux_2to1_17/SELB vrefA 2.12fF
C379 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD 19.81fF
C380 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y 0.42fF
C381 a_236582_n145742# a_239330_n145742# 0.14fF
C382 a_237040_n145742# a_238872_n145742# 0.43fF
C383 a_237498_n145742# a_238414_n145742# 1.92fF
C384 dac_8bit_0/amux_2to1_6/B vrefA 2.44fF
C385 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn biquad_gm_c_filter_0/gm_c_stage_1/vcmcn2 1.28fF
C386 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y a_242358_n123343# 0.16fF
C387 a_241919_n123337# a_242951_n123369# 0.11fF
C388 a_242273_n120623# low_freq_pll_0/freq_div_0/vin 0.02fF
C389 input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vbias4 28.62fF
C390 a_244783_n121711# a_245056_n121345# 0.38fF
C391 vampm input_amplifier_0/diff_fold_casc_ota_1/vcascnm 18.97fF
C392 biquad_gm_c_filter_0/gm_c_stage_2/vcmc VDD 2.70fF
C393 q0A VDD 3.81fF
C394 diff_to_se_converter_0/ibiasn low_freq_pll_0/ibiasn 8.26fF
C395 low_freq_pll_0/freq_div_0/vin a_242085_n120623# 0.06fF
C396 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin 0.40fF
C397 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 3.02fF
C398 a_337497_n185269# VDD 0.35fF
C399 dac_8bit_0/amux_2to1_2/SELB VDD 1.15fF
C400 a_245056_n121167# a_244617_n121711# 0.02fF
C401 a_242358_n122433# VDD 0.36fF
C402 a_244617_n121161# a_245056_n121345# 0.02fF
C403 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout a_238006_n119618# 0.03fF
C404 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_5/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q 0.15fF
C405 low_freq_pll_0/pfd_cp_lpf_0/vQA VDD 3.16fF
C406 a_238923_n122049# VDD 0.01fF
C407 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/A 0.09fF
C408 gain_ctrl_1 input_amplifier_0/venp2 0.79fF
C409 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/csinvn low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin 0.09fF
C410 a_217060_n102324# vocm 0.12fF
C411 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_245481_n122433# 0.05fF
C412 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d VDD 7.37fF
C413 vampm input_amplifier_0/venp2 2.93fF
C414 dac_8bit_0/ibiasn vpeak_sampled 5.00fF
C415 dac_8bit_0/amux_2to1_5/B VDD 4.57fF
C416 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/A 0.09fF
C417 input_amplifier_0/diff_fold_casc_ota_1/M1d input_amplifier_0/diff_fold_casc_ota_1/vfoldp 6.26fF
C418 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/M6d 1.84fF
C419 input_amplifier_0/diff_fold_casc_ota_1/M2d input_amplifier_0/diff_fold_casc_ota_1/vbias2 1.06fF
C420 input_amplifier_0/ibiasn1 biquad_gm_c_filter_0/ibiasn4 0.19fF
C421 m1_326207_n110098# adc_vcaparrayA 0.06fF
C422 dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d 9.79fF
C423 vbiasp low_freq_pll_0/ibiasn 2.19fF
C424 a_275374_n146348# sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror 8.05fF
C425 biquad_gm_c_filter_0/ibiasn2 vintm 0.15fF
C426 vcp low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/csinvn 0.08fF
C427 vlowB dac_8bit_1/amux_2to1_7/B 1.86fF
C428 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp 0.28fF
C429 q5A vlowA 2.75fF
C430 a_337864_n185269# a_338084_n185243# 0.04fF
C431 a_338156_n184969# a_338703_n185243# 0.26fF
C432 diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 10.10fF
C433 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/diff_fold_casc_ota_0/M3d 0.12fF
C434 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp a_162668_n147576# 10.36fF
C435 low_freq_pll_0/pfd_cp_lpf_0/vRSTN a_242419_n114983# 0.86fF
C436 a_225580_n122869# a_228328_n122869# 0.14fF
C437 input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/vom1 0.38fF
C438 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/diff_fold_casc_ota_0/vbias2 2.32fF
C439 a_226496_n122869# a_227412_n122869# 1.98fF
C440 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc 0.08fF
C441 a_226038_n122869# a_227870_n122869# 0.43fF
C442 vampp vocm_filt 0.28fF
C443 a_239143_n115125# VDD 0.33fF
C444 input_amplifier_0/vom1 a_217060_n102324# 8.05fF
C445 VDD dac_8bit_1/amux_2to1_16/SELB 1.15fF
C446 dac_8bit_0/c3m dac_8bit_0/c1m 0.07fF
C447 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm 23.84fF
C448 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/vhold 28.95fF
C449 dac_8bit_0/amux_2to1_9/Y dac_8bit_0/amux_2to1_9/SELB 1.59fF
C450 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q a_242951_n123369# 0.38fF
C451 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.40fF
C452 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn 2.30fF
C453 a_238312_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.03fF
C454 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/csinvp VDD 0.48fF
C455 a_242720_n114759# VDD 0.27fF
C456 vcp a_238312_n132168# 0.03fF
C457 vocm_filt vfiltp 2.96fF
C458 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VDD 6.84fF
C459 a_338356_n185510# a_338703_n185409# 0.11fF
C460 a_244617_n123337# a_244783_n123337# 2.23fF
C461 input_amplifier_0/diff_fold_casc_ota_0/vfoldp vocm 0.14fF
C462 input_amplifier_0/txgate_6/txb input_amplifier_0/vim2 0.60fF
C463 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q a_245649_n122531# 0.02fF
C464 a_337592_n185460# a_338156_n185665# 0.11fF
C465 a_337864_n185555# a_338149_n185569# 0.09fF
C466 dac_8bit_0/amux_2to1_16/SELB vlowA 1.62fF
C467 peak_detector_0/ibiasn2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm 0.08fF
C468 dac_8bit_1/amux_2to1_0/B vrefB 2.44fF
C469 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_226939_n130007# 0.03fF
C470 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/vip2 3.11fF
C471 diff_to_se_converter_0/rst vfiltp 0.55fF
C472 a_245565_n121345# VDD 0.02fF
C473 a_242854_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs 0.03fF
C474 input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vcascnm 11.77fF
C475 dac_8bit_0/latched_comparator_folded_0/vcompm VDD 5.25fF
C476 a_242951_n121193# a_243382_n121167# 0.31fF
C477 low_freq_pll_0/pfd_cp_lpf_0/vpdiode VDD 1.10fF
C478 low_freq_pll_0/cs_ring_osc_0/vpbias a_228020_n140786# 0.92fF
C479 dac_8bit_1/c7m dac_8bit_1/c3m 1.31fF
C480 input_amplifier_0/txgate_0/txb VDD 3.08fF
C481 vampp input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 0.69fF
C482 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc 0.55fF
C483 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/M13d 6.93fF
C484 biquad_gm_c_filter_0/ibiasn2 diff_to_se_converter_0/ibiasn 0.36fF
C485 input_amplifier_0/diff_fold_casc_ota_1/M2d vampm 0.38fF
C486 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc 0.08fF
C487 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/diff_fold_casc_ota_1/vbias2 2.32fF
C488 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/M3d 0.12fF
C489 a_335749_n185269# VDD 0.38fF
C490 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 a_230446_n180872# 8.05fF
C491 input_amplifier_0/ibiasn2 input_amplifier_0/ibiasn1 6.32fF
C492 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/vip 1.41fF
C493 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y 0.30fF
C494 a_239048_n115125# a_238793_n115125# 0.22fF
C495 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/A VDD 0.62fF
C496 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d 0.75fF
C497 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp 0.08fF
C498 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 44.84fF
C499 a_241188_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias 0.66fF
C500 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/csinvp VDD 0.48fF
C501 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d VDD 11.46fF
C502 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/vom1 2.90fF
C503 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc 0.96fF
C504 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y a_242358_n121345# 0.16fF
C505 a_241919_n121711# a_242951_n121443# 0.11fF
C506 dac_8bit_1/amux_2to1_7/SELB dac_8bit_1/c1m 1.59fF
C507 a_337497_n185813# a_337497_n185269# 0.04fF
C508 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp diff_to_se_converter_0/vip 0.86fF
C509 a_244617_n121711# a_244617_n122249# 0.08fF
C510 a_336408_n184969# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.06fF
C511 biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail1 biquad_gm_c_filter_0/gm_c_stage_3/vtail_diff 0.49fF
C512 a_238793_n115125# a_239361_n114883# 0.41fF
C513 a_238627_n115125# low_freq_pll_0/pfd_cp_lpf_0/vRSTN 0.86fF
C514 low_freq_pll_0/cs_ring_osc_0/vosc2 VDD 0.58fF
C515 dac_8bit_1/ibiasn vlowA 0.28fF
C516 input_amplifier_0/diff_fold_casc_ota_0/M13d input_amplifier_0/diff_fold_casc_ota_0/vbias4 0.04fF
C517 adc_compB VDD 2.44fF
C518 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_224954_n135628# 0.03fF
C519 vocm_filt biquad_gm_c_filter_0/gm_c_stage_3/vcmcn2 0.38fF
C520 a_229954_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.03fF
C521 dac_8bit_0/latched_comparator_folded_0/vtailp VDD 1.69fF
C522 biquad_gm_c_filter_0/ibiasn2 biquad_gm_c_filter_0/gm_c_stage_1/vtail_diff 0.06fF
C523 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm 0.51fF
C524 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 1.65fF
C525 a_246080_n123343# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/A 0.05fF
C526 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm 0.08fF
C527 input_amplifier_0/diff_fold_casc_ota_1/vbias2 vocm 0.49fF
C528 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 6.00fF
C529 low_freq_pll_0/pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/Q_N a_240447_n115125# 0.14fF
C530 dac_8bit_0/latched_comparator_folded_0/vcompmb dac_8bit_0/latched_comparator_folded_0/vcompm_buf 0.31fF
C531 biquad_gm_c_filter_0/ibiasn1 input_amplifier_0/ibiasn1 0.19fF
C532 biquad_gm_c_filter_0/ibiasn2 vbiasp 2.86fF
C533 input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc vocm 2.51fF
C534 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn vampp 0.49fF
C535 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d VDD 9.36fF
C536 a_244617_n123337# a_244617_n122799# 0.08fF
C537 a_335749_n185269# a_335749_n185813# 0.04fF
C538 input_amplifier_0/diff_fold_casc_ota_0/M1d input_amplifier_0/vop1 0.54fF
C539 a_245151_n122255# VDD 0.02fF
C540 vse diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 13.30fF
C541 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 1.13fF
C542 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 0.61fF
C543 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_241785_n138121# 0.03fF
C544 a_226954_n122869# low_freq_pll_0/cs_ring_osc_0/vpbias 0.83fF
C545 dac_8bit_0/c0m dac_8bit_1/ibiasn 0.20fF
C546 comparator_0/vcompm VDD 5.99fF
C547 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_244617_n122799# 0.03fF
C548 a_241938_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs 0.03fF
C549 low_freq_pll_0/cs_ring_osc_0/vosc a_221022_n131500# 0.03fF
C550 a_226646_n140786# VDD 0.40fF
C551 a_236175_n122049# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout 0.03fF
C552 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc 0.10fF
C553 dac_8bit_0/amux_2to1_6/SELB dac_8bit_0/amux_2to1_6/B 1.51fF
C554 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/M13d 0.18fF
C555 adc_vcaparrayB dac_8bit_1/c4m 111.85fF
C556 dac_8bit_1/ibiasn sample 4.69fF
C557 biquad_gm_c_filter_0/ibiasn3 vpeak_sampled 0.42fF
C558 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc 0.96fF
C559 input_amplifier_0/diff_fold_casc_ota_1/vfoldp vampm 2.90fF
C560 a_245056_n122255# a_245182_n121877# 0.02fF
C561 a_336757_n185421# a_336608_n185510# 0.02fF
C562 a_336955_n185409# a_336408_n185665# 0.26fF
C563 vfiltp biquad_gm_c_filter_0/ibiasn4 0.17fF
C564 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y a_242273_n122255# 0.38fF
C565 vintm vocm_filt 6.20fF
C566 vpeak_sampled dac_8bit_1/amux_2to1_5/SELB 2.07fF
C567 input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc input_amplifier_0/vom1 2.27fF
C568 vlowA dac_8bit_0/amux_2to1_1/B 1.86fF
C569 vcp_sampled dac_8bit_0/amux_2to1_0/B 0.38fF
C570 q4A vlowA 2.75fF
C571 a_246080_n121389# a_246080_n122255# 0.04fF
C572 low_freq_pll_0/cs_ring_osc_0/vosc a_223313_n130007# 0.03fF
C573 input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/diff_fold_casc_ota_0/M13d 0.70fF
C574 comparator_0/vmirror comparator_0/vo1 1.16fF
C575 dac_8bit_0/amux_2to1_3/SELB dac_8bit_0/c4m 1.59fF
C576 input_amplifier_0/vip2 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 0.15fF
C577 gain_ctrl_1 input_amplifier_0/txgate_3/txb 0.36fF
C578 pulse_generator_0/sky130_fd_sc_hd__inv_1_1/A pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/Q_N 0.21fF
C579 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 8.90fF
C580 input_amplifier_0/diff_fold_casc_ota_0/M13d a_217060_n102324# 1.44fF
C581 dac_8bit_0/latched_comparator_folded_0/vcomppb VDD 0.47fF
C582 a_242273_n123343# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y 0.38fF
C583 vampm vocm 4.93fF
C584 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y a_243382_n120301# 0.11fF
C585 a_337864_n185555# adc_clk 0.05fF
C586 vocm_filt biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail2 2.82fF
C587 a_246080_n123343# a_246080_n122477# 0.04fF
C588 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y 0.42fF
C589 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y a_244971_n122799# 0.38fF
C590 a_245481_n121167# a_245481_n121345# 0.05fF
C591 vpeak_sampled dac_8bit_1/c4m 1.94fF
C592 a_246786_n134960# vcp 0.03fF
C593 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/vop1 1.24fF
C594 dac_8bit_1/amux_2to1_1/SELB VDD 1.15fF
C595 a_241919_n121161# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q 0.03fF
C596 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD 1.49fF
C597 dac_8bit_0/amux_2to1_15/SELB vlowA 1.62fF
C598 a_246080_n122255# VDD 0.37fF
C599 vampp input_amplifier_0/ibiasn2 0.16fF
C600 a_337497_n185269# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.21fF
C601 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 4.16fF
C602 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A a_338156_n184969# 0.02fF
C603 sample dac_8bit_0/amux_2to1_1/B 2.66fF
C604 a_242358_n122433# a_242484_n122799# 0.02fF
C605 a_242951_n122281# VDD 0.45fF
C606 a_225580_n122869# VDD 4.03fF
C607 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q 0.02fF
C608 vampp vintp 0.87fF
C609 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 9.20fF
C610 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 21.43fF
C611 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/csinvp a_243478_n140786# 0.16fF
C612 input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc 6.63fF
C613 vampm input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc 5.06fF
C614 a_242358_n120257# VDD 0.36fF
C615 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 input_amplifier_0/vim2 1.29fF
C616 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/D VDD 0.40fF
C617 low_freq_pll_0/cs_ring_osc_0/vosc2 low_freq_pll_0/freq_div_0/vin 1.01fF
C618 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y a_242951_n121193# 0.17fF
C619 input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc vampm 2.27fF
C620 a_244783_n122249# a_245649_n122281# 0.11fF
C621 a_245224_n122281# a_245056_n122255# 0.59fF
C622 diff_to_se_converter_0/ibiasn vocm_filt 3.00fF
C623 input_amplifier_0/vop1 vocm 1.39fF
C624 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y a_244971_n121167# 0.38fF
C625 a_245649_n121193# VDD 0.45fF
C626 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 16.73fF
C627 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 28.69fF
C628 a_242085_n121711# a_242273_n121711# 0.26fF
C629 a_223872_n127742# VDD 0.09fF
C630 a_336608_n185269# VDD 0.36fF
C631 a_337864_n185555# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_2/Q 0.04fF
C632 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/diff_fold_casc_ota_0/M13d 1.62fF
C633 a_242526_n121193# a_242273_n121167# 0.04fF
C634 a_242526_n121193# VDD 0.23fF
C635 vintp vfiltp 1.72fF
C636 vpeak_sampled a_275374_n180872# 21.33fF
C637 diff_to_se_converter_0/ibiasn diff_to_se_converter_0/rst 0.36fF
C638 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_236481_n148007# 0.03fF
C639 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm 12.61fF
C640 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d 10.82fF
C641 dac_8bit_0/latched_comparator_folded_0/vlatchp adc_clk 0.39fF
C642 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y 0.42fF
C643 VDD a_245481_n122433# 0.22fF
C644 vocm_filt biquad_gm_c_filter_0/gm_c_stage_1/vtail_diff 1.19fF
C645 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d 2.62fF
C646 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp 0.73fF
C647 a_336116_n185555# a_336608_n185510# 0.03fF
C648 a_336401_n185569# a_336408_n185665# 2.23fF
C649 a_335844_n185460# a_336537_n185409# 0.04fF
C650 a_245056_n123343# a_245481_n123343# 0.03fF
C651 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn vintm 0.42fF
C652 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/A 1.64fF
C653 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn2 vfiltm 0.19fF
C654 input_amplifier_0/vom1 input_amplifier_0/vop1 55.78fF
C655 dac_8bit_0/c0m dac_8bit_0/c7m 0.85fF
C656 dac_8bit_0/c1m dac_8bit_0/c6m 2.24fF
C657 dac_8bit_0/c2m dac_8bit_0/c4m 1.04fF
C658 dac_8bit_0/cdumm dac_8bit_0/c5m 0.43fF
C659 sample dac_8bit_1/c0m 2.36fF
C660 a_242783_n122255# a_242085_n121711# 0.01fF
C661 peak_detector_0/vpeak peak_detector_0/verr 1.01fF
C662 a_242358_n122255# a_242358_n121345# 0.05fF
C663 a_242085_n122249# a_242783_n122255# 0.44fF
C664 a_336955_n185409# a_336955_n185243# 0.02fF
C665 a_237956_n127742# a_239330_n127742# 0.01fF
C666 a_237498_n127742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/csinvp 0.09fF
C667 a_238414_n127742# a_238872_n127742# 0.01fF
C668 a_338149_n185269# a_338285_n185243# 0.37fF
C669 a_336408_n184969# a_336116_n185555# 0.01fF
C670 a_338156_n184969# pulse_generator_0/sky130_fd_sc_hd__inv_1_0/Y 0.61fF
C671 low_freq_pll_0/pfd_cp_lpf_0/vQAb VDD 3.39fF
C672 a_242783_n123343# a_242783_n122433# 0.07fF
C673 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/csinvn vcp 0.08fF
C674 sample dac_8bit_0/c7m 2.10fF
C675 a_245224_n122281# a_245224_n122687# 0.03fF
C676 dac_8bit_1/c5m dac_8bit_1/amux_2to1_2/B 2.37fF
C677 low_freq_pll_0/cs_ring_osc_0/vpbias a_238414_n145742# 0.76fF
C678 input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 0.69fF
C679 a_241188_n140786# a_242104_n140786# 2.26fF
C680 a_240730_n140786# a_242562_n140786# 0.65fF
C681 a_243138_n114759# a_242380_n114857# 0.22fF
C682 biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail2 biquad_gm_c_filter_0/ibiasn4 0.19fF
C683 vcp a_221022_n150168# 0.03fF
C684 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/Q_N VDD 0.47fF
C685 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/vpeak 0.71fF
C686 dac_8bit_0/amux_2to1_3/B VDD 4.57fF
C687 a_242526_n121193# a_242526_n121599# 0.03fF
C688 a_224330_n145742# VDD 0.06fF
C689 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/vim 4.81fF
C690 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/vhold 6.29fF
C691 q3A vlowA 2.75fF
C692 a_242951_n121443# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_3/A 0.04fF
C693 a_242783_n121345# a_243382_n121389# 0.02fF
C694 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm 2.00fF
C695 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_241786_n135628# 0.03fF
C696 vcomp low_freq_pll_0/pfd_cp_lpf_0/vQAb 0.04fF
C697 vintm biquad_gm_c_filter_0/gm_c_stage_2/vcmcn1 0.12fF
C698 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q a_242273_n122255# 0.02fF
C699 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp 1.03fF
C700 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror 14.22fF
C701 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d 1.91fF
C702 a_237498_n145742# a_239330_n145742# 0.24fF
C703 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp diff_to_se_converter_0/vim 0.86fF
C704 a_237956_n145742# a_238872_n145742# 1.33fF
C705 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d 16.02fF
C706 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp 19.65fF
C707 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/verr 3.16fF
C708 dac_8bit_1/comp_outm adc_clk 0.04fF
C709 a_244783_n121711# a_245481_n121345# 0.44fF
C710 a_245224_n121599# a_245649_n121443# 0.04fF
C711 adc_compA a_383050_n101129# 0.05fF
C712 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm vse 2.13fF
C713 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp 1.94fF
C714 vocm_filt biquad_gm_c_filter_0/gm_c_stage_1/vcmcn2 0.28fF
C715 dac_8bit_0/amux_2to1_5/SELB VDD 1.15fF
C716 a_244783_n123337# VDD 0.43fF
C717 dac_8bit_0/latched_comparator_folded_0/vtailp dac_8bit_0/ibiasp 1.91fF
C718 diff_to_se_converter_0/ibiasn biquad_gm_c_filter_0/ibiasn4 0.38fF
C719 a_242783_n123343# a_242867_n123343# 0.05fF
C720 biquad_gm_c_filter_0/gm_c_stage_2/vcmc biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail1 0.15fF
C721 vcp a_221022_n132168# 0.03fF
C722 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_226939_n148007# 0.03fF
C723 adc_vcaparrayA vlowA 1.95fF
C724 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d vse 4.90fF
C725 a_337864_n185269# VDD 0.22fF
C726 a_244783_n122799# a_245224_n122687# 0.28fF
C727 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/Q_N a_335749_n185813# 0.21fF
C728 a_337497_n185813# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/D 0.22fF
C729 a_242783_n122433# VDD 0.22fF
C730 vintm biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail1 2.84fF
C731 gain_ctrl_0 input_amplifier_0/rst 1.43fF
C732 dac_8bit_0/amux_2to1_14/SELB vlowA 1.62fF
C733 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout a_238922_n119618# 0.03fF
C734 a_236582_n127742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin 0.90fF
C735 vcp_sampled sample_and_hold_0/vholdm 44.74fF
C736 input_amplifier_0/ibiasn2 input_amplifier_0/vim2 0.61fF
C737 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y VDD 0.93fF
C738 vintp vintm 13.75fF
C739 a_238627_n115125# a_239143_n115125# 0.42fF
C740 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q a_245649_n121193# 0.02fF
C741 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_9/A 0.07fF
C742 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y a_242273_n122799# 0.38fF
C743 dac_8bit_1/c6m dac_8bit_1/c5m 1.39fF
C744 a_237040_n145742# VDD 1.55fF
C745 dac_8bit_1/c7m dac_8bit_1/c4m 1.44fF
C746 dac_8bit_0/c0m adc_vcaparrayA 15.13fF
C747 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn a_275374_n180872# 0.11fF
C748 a_240062_n115125# low_freq_pll_0/pfd_cp_lpf_0/vRSTN 0.01fF
C749 VDD input_amplifier_0/vip1 0.62fF
C750 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 3.47fF
C751 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm 16.88fF
C752 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp peak_detector_0/vpeak 0.86fF
C753 vbiasp biquad_gm_c_filter_0/ibiasn4 1.75fF
C754 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD 7.64fF
C755 vlowB dac_8bit_1/latched_comparator_folded_0/vlatchp 0.16fF
C756 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn 16.73fF
C757 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 28.69fF
C758 dac_8bit_1/latched_comparator_folded_0/vtailp dac_8bit_1/latched_comparator_folded_0/vlatchm 1.85fF
C759 dac_8bit_0/c5m VDD 2.56fF
C760 a_245411_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.03fF
C761 biquad_gm_c_filter_0/ibiasn1 vintm 0.98fF
C762 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm 0.08fF
C763 adc_vcaparrayA sample 0.40fF
C764 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm 20.84fF
C765 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 1.35fF
C766 a_226954_n122869# a_227870_n122869# 1.33fF
C767 peak_detector_0/ibiasn2 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d 0.38fF
C768 a_338356_n185269# a_338703_n185243# 0.11fF
C769 a_226496_n122869# a_228328_n122869# 0.24fF
C770 low_freq_pll_0/pfd_cp_lpf_0/vRSTN a_242506_n114759# 0.37fF
C771 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp 0.73fF
C772 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 1.65fF
C773 input_amplifier_0/txgate_6/txb input_amplifier_0/vop1 0.36fF
C774 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm 0.08fF
C775 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror 4.50fF
C776 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm 0.51fF
C777 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y 0.30fF
C778 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/Q_N 0.24fF
C779 a_239708_n115125# VDD 0.39fF
C780 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 1.13fF
C781 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn 0.21fF
C782 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp a_356329_n164260# 10.36fF
C783 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn a_275374_n146348# 0.11fF
C784 a_242453_n123343# a_242358_n123343# 0.04fF
C785 a_242867_n123343# VDD 0.02fF
C786 a_229702_n119618# vcp 0.03fF
C787 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d 6.93fF
C788 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp 19.65fF
C789 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d 3.28fF
C790 vocm_filt biquad_gm_c_filter_0/gm_c_stage_3/vtail_diff 1.19fF
C791 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp 0.28fF
C792 diff_to_se_converter_0/ibiasn input_amplifier_0/ibiasn2 0.63fF
C793 vpeak_sampled low_freq_pll_0/ibiasn 0.48fF
C794 a_245481_n122433# a_245565_n122433# 0.05fF
C795 VDD a_244617_n122799# 0.78fF
C796 input_amplifier_0/venm2 VDD 2.02fF
C797 a_221023_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin 0.03fF
C798 q1A vlowA 2.75fF
C799 a_338356_n185510# a_338532_n185787# 0.04fF
C800 a_244617_n123337# a_245056_n123343# 0.63fF
C801 input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/M13d 9.82fF
C802 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y a_245224_n123369# 0.15fF
C803 a_241919_n121161# a_241919_n121711# 0.20fF
C804 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d vse 0.58fF
C805 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 6.88fF
C806 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs 0.40fF
C807 a_337592_n185460# a_338285_n185409# 0.04fF
C808 a_337864_n185555# a_338356_n185510# 0.03fF
C809 a_338149_n185569# a_338156_n185665# 2.23fF
C810 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm 32.00fF
C811 sample_and_hold_0/vhold VDD 0.64fF
C812 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_227855_n130007# 0.03fF
C813 sample dac_8bit_1/amux_2to1_0/B 2.60fF
C814 a_236022_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin 0.03fF
C815 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 vse 7.98fF
C816 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d 2.62fF
C817 vlowB dac_8bit_1/adc_run 0.35fF
C818 a_243770_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs 0.03fF
C819 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_226022_n149500# 0.03fF
C820 dac_8bit_0/latched_comparator_folded_0/vlatchp dac_8bit_0/latched_comparator_folded_0/vcompp 0.36fF
C821 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/A a_243382_n120301# 0.05fF
C822 a_239048_n115125# a_239251_n114759# 0.02fF
C823 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/A 0.09fF
C824 dac_8bit_0/comp_outm VDD 0.67fF
C825 dac_8bit_0/amux_2to1_9/Y q0A 1.99fF
C826 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 33.98fF
C827 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 2.21fF
C828 a_245056_n121167# a_245151_n121167# 0.04fF
C829 biquad_gm_c_filter_0/ibiasn1 diff_to_se_converter_0/ibiasn 0.37fF
C830 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD 1.46fF
C831 input_amplifier_0/ibiasn2 vbiasp 0.77fF
C832 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_0/Q_N pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/D 0.02fF
C833 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 28.69fF
C834 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/vholdm 2.13fF
C835 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn 16.73fF
C836 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror 2.23fF
C837 vintp biquad_gm_c_filter_0/gm_c_stage_1/vtail_diff 3.07fF
C838 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 8.42fF
C839 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm 4.75fF
C840 a_239251_n114759# a_239361_n114883# 0.23fF
C841 q2A vlowA 2.75fF
C842 a_242104_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias 0.83fF
C843 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y a_242783_n121345# 0.14fF
C844 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm 5.03fF
C845 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 6.88fF
C846 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d 7.88fF
C847 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror 0.69fF
C848 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm 0.19fF
C849 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp 3.66fF
C850 a_337592_n185460# a_337592_n185269# 0.09fF
C851 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y 0.13fF
C852 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp 13.60fF
C853 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d 2.72fF
C854 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d 0.12fF
C855 a_239361_n114883# low_freq_pll_0/pfd_cp_lpf_0/vRSTN 0.37fF
C856 q7A VDD 6.38fF
C857 adc_compB dac_8bit_1/latched_comparator_folded_0/vcomppb 0.03fF
C858 a_241919_n123337# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y 0.35fF
C859 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_225870_n135628# 0.03fF
C860 adc_clk a_336408_n185665# 0.06fF
C861 low_freq_pll_0/cs_ring_osc_0/vosc2 low_freq_pll_0/cs_ring_osc_0/vosc 0.27fF
C862 a_230870_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.03fF
C863 a_244617_n121711# a_244783_n121711# 2.23fF
C864 a_241022_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs 0.03fF
C865 peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d a_189446_n180872# 1.44fF
C866 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin VDD 4.26fF
C867 biquad_gm_c_filter_0/ibiasn1 vbiasp 3.10fF
C868 comparator_0/ibiasn input_amplifier_0/ibiasn1 0.27fF
C869 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_241023_n130007# 0.03fF
C870 vpeak_sampled dac_8bit_1/amux_2to1_6/B 0.38fF
C871 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y 0.13fF
C872 a_335844_n185269# a_335844_n185460# 0.09fF
C873 a_239870_n114759# VDD 0.01fF
C874 dac_8bit_0/amux_2to1_13/SELB vlowA 1.62fF
C875 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp 11.53fF
C876 a_244617_n121161# a_244617_n121711# 0.20fF
C877 a_241919_n122799# VDD 0.79fF
C878 vcp_sampled dac_8bit_0/amux_2to1_0/SELB 2.07fF
C879 a_241919_n122249# a_242085_n121711# 0.02fF
C880 a_242909_n121711# a_242783_n121345# 0.04fF
C881 a_241919_n122249# a_242085_n122249# 2.23fF
C882 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_242701_n138121# 0.03fF
C883 a_227870_n122869# low_freq_pll_0/cs_ring_osc_0/vpbias 0.93fF
C884 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror 2.23fF
C885 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn1 VDD 3.44fF
C886 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d 5.99fF
C887 a_242085_n122799# a_242526_n122687# 0.28fF
C888 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp 1.03fF
C889 a_242854_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs 0.03fF
C890 peak_detector_0/ibiasn1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp 0.13fF
C891 low_freq_pll_0/cs_ring_osc_0/vosc a_221938_n131500# 0.03fF
C892 a_237091_n122049# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout 0.03fF
C893 a_227562_n140786# VDD 0.14fF
C894 vampm input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 0.45fF
C895 vfiltm VDD 2.98fF
C896 adc_vcaparrayB dac_8bit_1/c2m 57.70fF
C897 biquad_gm_c_filter_0/ibiasn2 vpeak_sampled 0.41fF
C898 dac_8bit_0/amux_2to1_4/B vlowA 1.86fF
C899 a_336955_n185409# a_336537_n185409# 0.04fF
C900 low_freq_pll_0/pfd_cp_lpf_0/VQBb low_freq_pll_0/pfd_cp_lpf_0/vQB 1.54fF
C901 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp 13.60fF
C902 vpeak a_189446_n180872# 19.89fF
C903 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm 23.84fF
C904 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d 13.66fF
C905 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm a_356329_n164260# 10.16fF
C906 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 3.45fF
C907 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d peak_detector_0/verr 0.58fF
C908 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp 1.94fF
C909 vintp biquad_gm_c_filter_0/gm_c_stage_1/vcmcn2 0.10fF
C910 dac_8bit_1/amux_2to1_2/B VDD 4.57fF
C911 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp 7.95fF
C912 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d 15.11fF
C913 input_amplifier_0/txgate_7/txb input_amplifier_0/rst 0.36fF
C914 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_7/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_8/A 0.04fF
C915 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q 0.02fF
C916 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 adc_vcaparrayB 0.71fF
C917 a_240730_n140786# VDD 0.73fF
C918 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp vse 5.59fF
C919 gain_ctrl_0 input_amplifier_0/vim2 0.52fF
C920 a_242453_n121345# VDD 0.02fF
C921 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d 4.98fF
C922 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d 10.82fF
C923 sample dac_8bit_0/amux_2to1_1/SELB 2.36fF
C924 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm 3.14fF
C925 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp 11.53fF
C926 input_amplifier_0/venm1 input_amplifier_0/vom1 29.19fF
C927 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc 6.12fF
C928 a_246080_n121389# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/A 0.05fF
C929 dac_8bit_0/latched_comparator_folded_0/vcompp_buf dac_8bit_0/latched_comparator_folded_0/vcompp 0.02fF
C930 dac_8bit_0/cdumm dac_8bit_0/amux_2to1_6/B 1.72fF
C931 dac_8bit_1/amux_2to1_2/B q5B 1.99fF
C932 low_freq_pll_0/pfd_cp_lpf_0/vswitchl vcp 0.07fF
C933 a_338156_n185665# adc_clk 0.73fF
C934 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y 0.66fF
C935 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_10/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_9/A 0.04fF
C936 a_246080_n121167# a_246080_n121389# 0.04fF
C937 dac_8bit_0/amux_2to1_4/B sample 2.66fF
C938 vpeak_sampled dac_8bit_1/c2m 1.94fF
C939 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y 0.42fF
C940 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn vampm 0.51fF
C941 vpeak_sampled vpeak 0.12fF
C942 a_242951_n122531# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q 0.39fF
C943 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/ibiasn2 1.60fF
C944 rst_n input_amplifier_0/vip1 0.23fF
C945 a_243382_n122255# VDD 0.37fF
C946 a_226496_n122869# VDD 1.24fF
C947 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/rst 0.11fF
C948 input_amplifier_0/ibiasn1 input_amplifier_0/vim1 0.17fF
C949 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/A VDD 0.62fF
C950 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y 1.64fF
C951 a_242783_n120257# VDD 0.22fF
C952 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y a_243382_n121167# 0.11fF
C953 a_242867_n121345# VDD 0.02fF
C954 a_245056_n122255# a_245649_n122281# 0.02fF
C955 a_245224_n122281# a_245481_n122255# 0.11fF
C956 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/vholdm 2.37fF
C957 vintp biquad_gm_c_filter_0/gm_c_stage_3/vtail_diff 0.33fF
C958 adc_clk a_336955_n185243# 0.02fF
C959 a_246080_n121167# VDD 0.37fF
C960 input_amplifier_0/txgate_2/txb VDD 3.08fF
C961 dac_8bit_0/amux_2to1_10/SELB vlowA 1.62fF
C962 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/ibiasn 0.03fF
C963 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 1.65fF
C964 a_242358_n121345# a_242273_n121711# 0.11fF
C965 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm 0.51fF
C966 dac_8bit_0/ibiasn dac_8bit_0/c5m 0.19fF
C967 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/csinvp VDD 0.48fF
C968 a_338156_n185665# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_2/Q 0.01fF
C969 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/D VDD 0.41fF
C970 dac_8bit_0/ibiasp dac_8bit_0/c5m 0.26fF
C971 dac_8bit_1/c6m VDD 2.50fF
C972 a_242358_n121167# a_242484_n120789# 0.02fF
C973 a_242085_n121161# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q 0.03fF
C974 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 0.21fF
C975 a_242951_n121193# VDD 0.45fF
C976 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm a_162668_n147576# 10.16fF
C977 a_241919_n121711# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y 0.35fF
C978 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm 16.88fF
C979 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp adc_vcaparrayA 0.86fF
C980 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 3.47fF
C981 a_241919_n121161# a_242085_n120623# 0.02fF
C982 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_237397_n148007# 0.03fF
C983 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d 0.16fF
C984 dac_8bit_0/amux_2to1_7/B vrefA 2.44fF
C985 low_freq_pll_0/freq_div_0/vout a_238793_n115125# 0.04fF
C986 dac_8bit_1/amux_2to1_2/SELB dac_8bit_1/c5m 1.59fF
C987 dac_8bit_0/latched_comparator_folded_0/vlatchp dac_8bit_0/latched_comparator_folded_0/vcompm 1.33fF
C988 dac_8bit_1/amux_2to1_4/SELB dac_8bit_1/amux_2to1_4/B 1.51fF
C989 peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp 12.69fF
C990 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_9/A 0.48fF
C991 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d 1.74fF
C992 dac_8bit_0/c2m dac_8bit_0/cdumm 10.49fF
C993 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d 0.82fF
C994 dac_8bit_1/latched_comparator_folded_0/vcompm dac_8bit_1/latched_comparator_folded_0/vcompmb 0.23fF
C995 a_336401_n185569# a_336537_n185409# 0.37fF
C996 a_336408_n185665# a_336608_n185510# 0.38fF
C997 a_245649_n123369# a_246080_n123343# 0.31fF
C998 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q a_244971_n123343# 0.02fF
C999 vpeak sample_and_hold_1/vhold 1.71fF
C1000 dac_8bit_0/amux_2to1_3/SELB VDD 1.15fF
C1001 dac_8bit_0/amux_2to1_12/SELB vlowA 1.62fF
C1002 vpeak peak_detector_0/verr 0.05fF
C1003 a_242951_n122281# a_242951_n121443# 0.09fF
C1004 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y 0.03fF
C1005 a_238872_n127742# a_239330_n127742# 0.02fF
C1006 a_238414_n127742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/csinvp 0.10fF
C1007 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/vcom_buf 8.06fF
C1008 a_338356_n185269# pulse_generator_0/sky130_fd_sc_hd__inv_1_0/Y 0.04fF
C1009 a_336401_n185269# a_336401_n185569# 0.08fF
C1010 a_336408_n184969# a_336408_n185665# 0.06fF
C1011 vampm input_amplifier_0/ibiasn2 0.16fF
C1012 pulse_generator_0/sky130_fd_sc_hd__inv_1_1/A pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A 0.26fF
C1013 a_243382_n123343# a_243382_n122477# 0.04fF
C1014 low_freq_pll_0/pfd_cp_lpf_0/vpbias VDD 5.78fF
C1015 diff_to_se_converter_0/txgate_0/txb vfiltp 0.35fF
C1016 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.04fF
C1017 a_244783_n121161# a_245224_n121193# 0.28fF
C1018 a_245056_n122255# a_245056_n122433# 0.08fF
C1019 dac_8bit_0/amux_2to1_17/SELB VDD 1.15fF
C1020 low_freq_pll_0/cs_ring_osc_0/vpbias a_239330_n145742# 0.77fF
C1021 a_241646_n140786# a_242562_n140786# 1.92fF
C1022 a_240730_n140786# a_243478_n140786# 0.14fF
C1023 peak_detector_0/ibiasn1 peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d 0.13fF
C1024 vampm vintp 2.82fF
C1025 a_241188_n140786# a_243020_n140786# 0.43fF
C1026 input_amplifier_0/txgate_1/txb input_amplifier_0/venp1 0.35fF
C1027 dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp 23.02fF
C1028 a_243138_n114759# a_242575_n114888# 0.13fF
C1029 a_242720_n114759# a_242506_n114759# 0.23fF
C1030 dac_8bit_0/amux_2to1_6/B VDD 4.57fF
C1031 peak_detector_0/ibiasn2 VDD 5.62fF
C1032 a_336116_n185269# a_336408_n184969# 0.44fF
C1033 input_amplifier_0/rst input_amplifier_0/vim1 0.81fF
C1034 dac_8bit_0/latched_comparator_folded_0/vtailp dac_8bit_0/latched_comparator_folded_0/vlatchp 2.00fF
C1035 vcp a_221938_n150168# 0.03fF
C1036 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 vpeak 5.84fF
C1037 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn 8.02fF
C1038 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y a_244971_n122255# 0.38fF
C1039 diff_to_se_converter_0/vip vfiltm 1.07fF
C1040 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 58.37fF
C1041 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d 1.84fF
C1042 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d 1.51fF
C1043 a_242358_n121167# a_242358_n121345# 0.08fF
C1044 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp 4.15fF
C1045 a_243382_n121389# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_3/A 0.25fF
C1046 vlowB dac_8bit_1/amux_2to1_9/Y 1.90fF
C1047 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_242702_n135628# 0.03fF
C1048 dac_8bit_1/amux_2to1_8/SELB dac_8bit_1/amux_2to1_9/Y 1.51fF
C1049 vcomp low_freq_pll_0/pfd_cp_lpf_0/vpbias 0.10fF
C1050 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm adc_vcaparrayA 6.31fF
C1051 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm 2.00fF
C1052 a_238414_n145742# a_239330_n145742# 0.79fF
C1053 dac_8bit_0/amux_2to1_0/SELB dac_8bit_0/amux_2to1_0/B 1.51fF
C1054 a_245056_n121345# a_245481_n121345# 0.03fF
C1055 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/A 1.64fF
C1056 dac_8bit_0/c3m dac_8bit_0/c0m 0.07fF
C1057 a_245056_n123343# VDD 0.36fF
C1058 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp 1.94fF
C1059 dac_8bit_0/vcom_buf VDD 5.69fF
C1060 peak_detector_0/ibiasn1 input_amplifier_0/ibiasn1 0.76fF
C1061 vcp a_221938_n132168# 0.03fF
C1062 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_227855_n148007# 0.03fF
C1063 a_338149_n185269# VDD 0.81fF
C1064 dac_8bit_0/c3m sample 2.36fF
C1065 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_4/A VDD 0.48fF
C1066 a_239048_n115125# a_239143_n115125# 0.13fF
C1067 a_245224_n122687# a_245056_n122433# 0.59fF
C1068 a_244783_n122799# a_245649_n122531# 0.11fF
C1069 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 input_amplifier_0/ibiasn1 1.79fF
C1070 peak_detector_0/ibiasn1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror 0.40fF
C1071 a_275374_n146348# sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d 0.79fF
C1072 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/A 0.03fF
C1073 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/vcom_buf 9.19fF
C1074 a_237498_n127742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin 0.25fF
C1075 vfiltm rst_n 0.48fF
C1076 dac_8bit_1/amux_2to1_1/B vrefB 2.44fF
C1077 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VDD 23.91fF
C1078 a_239361_n114883# a_239143_n115125# 0.50fF
C1079 a_238627_n115125# a_239708_n115125# 0.27fF
C1080 a_238793_n115125# a_239883_n115151# 0.10fF
C1081 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror 17.44fF
C1082 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm 2.41fF
C1083 VDD input_amplifier_0/diff_fold_casc_ota_0/vfoldm 20.43fF
C1084 a_237956_n145742# VDD 0.69fF
C1085 sample vcp 0.90fF
C1086 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn1 VDD 3.44fF
C1087 dac_8bit_1/c7m dac_8bit_1/c2m 2.04fF
C1088 dac_8bit_1/c6m dac_8bit_1/c3m 1.31fF
C1089 dac_8bit_1/comp_outm adc_compB 1.08fF
C1090 a_245224_n121599# VDD 0.23fF
C1091 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror 4.50fF
C1092 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 6.00fF
C1093 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 2.79fF
C1094 dac_8bit_1/amux_2to1_2/B dac_8bit_1/amux_2to1_15/SELB 1.59fF
C1095 dac_8bit_0/c2m VDD 2.47fF
C1096 a_241919_n120623# VDD 0.79fF
C1097 sample_and_hold_0/vhold sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp 0.28fF
C1098 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d 1.74fF
C1099 a_242526_n122281# a_242526_n122687# 0.03fF
C1100 a_241105_n115125# low_freq_pll_0/pfd_cp_lpf_0/vRSTN 0.05fF
C1101 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y a_244783_n122249# 0.61fF
C1102 a_244617_n122249# a_245224_n122281# 0.37fF
C1103 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp vpeak 0.86fF
C1104 dac_8bit_0/amux_2to1_9/SELB vlowA 1.62fF
C1105 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d 5.21fF
C1106 a_246327_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.03fF
C1107 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y VDD 0.93fF
C1108 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp 0.73fF
C1109 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d 2.62fF
C1110 a_338356_n185269# a_338505_n185243# 0.02fF
C1111 a_227412_n122869# a_228328_n122869# 0.79fF
C1112 pulse_generator_0/sky130_fd_sc_hd__inv_1_0/Y a_338703_n185243# 0.35fF
C1113 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 24.81fF
C1114 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn 32.00fF
C1115 a_245056_n123343# a_245151_n123343# 0.04fF
C1116 sample dac_8bit_1/amux_2to1_0/SELB 2.46fF
C1117 low_freq_pll_0/pfd_cp_lpf_0/vQB VDD 0.49fF
C1118 a_336408_n184969# a_336955_n185243# 0.26fF
C1119 a_226480_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.03fF
C1120 vpeak_sampled biquad_gm_c_filter_0/ibiasn4 0.43fF
C1121 a_245481_n122433# a_245607_n122799# 0.04fF
C1122 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm 19.65fF
C1123 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_225411_n138121# 0.03fF
C1124 a_221939_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin 0.03fF
C1125 dac_8bit_1/vcom_buf a_356329_n164260# 19.89fF
C1126 a_230411_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.03fF
C1127 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y a_245649_n123369# 0.17fF
C1128 a_244617_n123337# a_245481_n123343# 0.09fF
C1129 dac_8bit_0/amux_2to1_11/SELB vlowA 1.62fF
C1130 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/vcom_buf 16.56fF
C1131 peak_detector_0/ibiasn1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 0.26fF
C1132 a_338156_n185665# a_338356_n185510# 0.38fF
C1133 a_338149_n185569# a_338285_n185409# 0.37fF
C1134 a_242358_n122255# a_241919_n121711# 0.01fF
C1135 input_amplifier_0/diff_fold_casc_ota_1/M6d VDD 11.14fF
C1136 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_228771_n130007# 0.03fF
C1137 a_222956_n145742# a_223414_n145742# 0.02fF
C1138 a_221582_n145742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/csinvp 0.08fF
C1139 a_236938_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin 0.03fF
C1140 VDD input_amplifier_0/diff_fold_casc_ota_0/M3d 1.56fF
C1141 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc 23.17fF
C1142 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn biquad_gm_c_filter_0/gm_c_stage_3/vcmcn1 1.18fF
C1143 vrefA VDD 29.33fF
C1144 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y VDD 0.91fF
C1145 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror 14.22fF
C1146 a_244783_n122249# a_244617_n122799# 0.09fF
C1147 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_226938_n149500# 0.03fF
C1148 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d 1.91fF
C1149 a_244617_n122249# a_244783_n122799# 0.09fF
C1150 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp 1.03fF
C1151 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 32.00fF
C1152 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn vfiltm 1.20fF
C1153 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn2 vocm_filt 0.28fF
C1154 comparator_0/vcompp vfiltp 0.57fF
C1155 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_8/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/A 0.35fF
C1156 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp 0.81fF
C1157 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d 3.07fF
C1158 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp 13.60fF
C1159 vampp input_amplifier_0/diff_fold_casc_ota_1/vtail_casc 1.62fF
C1160 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d VDD 1.27fF
C1161 comparator_0/ibiasn diff_to_se_converter_0/ibiasn 0.28fF
C1162 a_338532_n184877# VDD 0.02fF
C1163 dac_8bit_1/latched_comparator_folded_0/vcompm dac_8bit_1/latched_comparator_folded_0/vcompp 1.51fF
C1164 a_242783_n121167# a_242867_n121167# 0.05fF
C1165 a_242085_n121161# a_241919_n121711# 0.09fF
C1166 vcp_sampled dac_8bit_0/amux_2to1_1/B 0.38fF
C1167 vlowA dac_8bit_0/amux_2to1_2/B 1.86fF
C1168 vpeak_sampled dac_8bit_1/amux_2to1_6/SELB 2.07fF
C1169 a_243020_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias 0.92fF
C1170 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_3/A 0.27fF
C1171 input_amplifier_0/venp2 input_amplifier_0/venm2 9.34fF
C1172 a_337864_n185555# a_337864_n185269# 0.07fF
C1173 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_245649_n122281# 0.39fF
C1174 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/D pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.17fF
C1175 a_236022_n150168# vcp 0.03fF
C1176 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm 6.29fF
C1177 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_226786_n135628# 0.03fF
C1178 a_231786_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.03fF
C1179 dac_8bit_0/latched_comparator_folded_0/vcompp_buf dac_8bit_0/latched_comparator_folded_0/vcomppb 0.32fF
C1180 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y a_245224_n121599# 0.15fF
C1181 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD 1.49fF
C1182 input_amplifier_0/rst input_amplifier_0/txgate_4/txb 0.36fF
C1183 a_244617_n121711# a_245056_n121345# 0.63fF
C1184 a_241938_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs 0.03fF
C1185 vpeak_sampled input_amplifier_0/ibiasn2 0.44fF
C1186 vcp_sampled input_amplifier_0/ibiasn1 0.83fF
C1187 comparator_0/ibiasn vbiasp 7.29fF
C1188 low_freq_pll_0/freq_div_0/vin a_241919_n120623# 0.41fF
C1189 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_241939_n130007# 0.03fF
C1190 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vbias1 2.10fF
C1191 biquad_gm_c_filter_0/gm_c_stage_2/vcmc vocm_filt 0.24fF
C1192 a_245649_n123369# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.39fF
C1193 adc_clk a_336401_n185269# 0.45fF
C1194 a_221582_n145742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin 0.90fF
C1195 dac_8bit_1/amux_2to1_2/SELB VDD 1.15fF
C1196 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VDD 15.85fF
C1197 peak_detector_0/ibiasn2 rst_n 9.31fF
C1198 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin a_236023_n130007# 0.03fF
C1199 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y 0.06fF
C1200 a_242273_n122255# VDD 0.15fF
C1201 a_243382_n123343# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/A 0.05fF
C1202 input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc VDD 5.35fF
C1203 a_241919_n122249# a_242358_n121345# 0.01fF
C1204 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_0/vcom_buf 0.58fF
C1205 sample dac_8bit_0/amux_2to1_2/B 2.66fF
C1206 vcp a_227870_n119618# 0.03fF
C1207 a_335749_n185269# a_336116_n185269# 0.02fF
C1208 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y 0.30fF
C1209 a_242085_n122799# a_242951_n122531# 0.11fF
C1210 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD 25.41fF
C1211 a_242526_n122687# a_242358_n122433# 0.59fF
C1212 a_243770_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs 0.03fF
C1213 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 13.66fF
C1214 low_freq_pll_0/cs_ring_osc_0/vosc a_222854_n131500# 0.03fF
C1215 vlowA adc_clk 0.47fF
C1216 a_228478_n140786# VDD 0.06fF
C1217 a_238007_n122049# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout 0.03fF
C1218 dac_8bit_1/latched_comparator_folded_0/vcompmb VDD 0.47fF
C1219 dac_8bit_0/amux_2to1_6/SELB dac_8bit_0/cdumm 1.59fF
C1220 a_245056_n122255# a_245151_n122255# 0.04fF
C1221 biquad_gm_c_filter_0/ibiasn1 vpeak_sampled 0.42fF
C1222 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn1 biquad_gm_c_filter_0/gm_c_stage_0/vcmc 2.37fF
C1223 vocm_filt biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail2 4.74fF
C1224 input_amplifier_0/rst input_amplifier_0/diff_fold_casc_ota_0/vbias1 0.14fF
C1225 diff_to_se_converter_0/vim vfiltm 36.96fF
C1226 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VDD 1.49fF
C1227 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d 3.60fF
C1228 vrefB dac_8bit_1/amux_2to1_16/SELB 2.12fF
C1229 biquad_gm_c_filter_0/ibiasn3 vfiltm 0.17fF
C1230 biquad_gm_c_filter_0/gm_c_stage_2/vbiasp biquad_gm_c_filter_0/ibiasn4 0.04fF
C1231 VDD dac_8bit_1/amux_2to1_4/B 4.57fF
C1232 a_241646_n140786# VDD 0.40fF
C1233 vcp low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin 3.55fF
C1234 vcp_sampled dac_8bit_0/c7m 1.94fF
C1235 peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 0.56fF
C1236 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn 8.02fF
C1237 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q a_242273_n121711# 0.02fF
C1238 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD 1.45fF
C1239 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp 1.03fF
C1240 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn biquad_gm_c_filter_0/gm_c_stage_0/vcmcn2 1.28fF
C1241 sample adc_clk 0.58fF
C1242 a_338285_n185409# adc_clk 0.05fF
C1243 input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc 28.15fF
C1244 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_6/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_7/A 0.04fF
C1245 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vfoldp 0.12fF
C1246 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vcascnm 10.63fF
C1247 dac_8bit_0/vcom_buf dac_8bit_0/ibiasp 0.20fF
C1248 dac_8bit_0/cdumm dac_8bit_0/c4m 0.43fF
C1249 dac_8bit_0/c1m dac_8bit_0/c5m 1.12fF
C1250 low_freq_pll_0/cs_ring_osc_0/vpbias a_237040_n127742# 0.66fF
C1251 dac_8bit_0/c0m dac_8bit_0/c6m 0.85fF
C1252 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 44.84fF
C1253 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 a_356329_n113250# 8.26fF
C1254 biquad_gm_c_filter_0/gm_c_stage_2/vbiasp biquad_gm_c_filter_0/gm_c_stage_2/vcmcn1 0.19fF
C1255 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q 0.21fF
C1256 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/vcom_buf 5.70fF
C1257 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A pulse_generator_0/sky130_fd_sc_hd__inv_1_0/Y 0.04fF
C1258 sample dac_8bit_0/c6m 2.17fF
C1259 a_243382_n122477# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q 0.37fF
C1260 peak_detector_0/ibiasn1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn 0.15fF
C1261 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VDD 12.54fF
C1262 a_227412_n122869# VDD 0.52fF
C1263 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VDD 7.64fF
C1264 comparator_0/vtail vfiltp 0.28fF
C1265 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 3.02fF
C1266 adc_vcaparrayB sample 1.26fF
C1267 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q a_242951_n122531# 0.02fF
C1268 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_0/A VDD 0.48fF
C1269 input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 0.59fF
C1270 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn 2.79fF
C1271 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 6.00fF
C1272 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc input_amplifier_0/vim2 8.59fF
C1273 dac_8bit_0/c2m dac_8bit_0/ibiasn 0.19fF
C1274 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q VDD 0.38fF
C1275 dac_8bit_0/c2m dac_8bit_0/ibiasp 0.26fF
C1276 a_245649_n122281# a_245481_n122255# 0.67fF
C1277 biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail1 biquad_gm_c_filter_0/gm_c_stage_2/vtail_diff 0.49fF
C1278 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD 6.84fF
C1279 adc_clk a_337592_n185269# 0.21fF
C1280 biquad_gm_c_filter_0/gm_c_stage_2/vcmc biquad_gm_c_filter_0/ibiasn4 0.11fF
C1281 biquad_gm_c_filter_0/gm_c_stage_0/vcmc biquad_gm_c_filter_0/gm_c_stage_0/vtail_diff 0.03fF
C1282 a_243382_n121167# VDD 0.37fF
C1283 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d 0.56fF
C1284 a_242526_n122281# a_242358_n122255# 0.59fF
C1285 low_freq_pll_0/cs_ring_osc_0/vosc low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/csinvp 1.18fF
C1286 a_241919_n121161# a_242358_n120257# 0.01fF
C1287 vintp biquad_gm_c_filter_0/gm_c_stage_2/vbiasp 0.32fF
C1288 comparator_0/vcompm comparator_0/vmirror 1.29fF
C1289 comparator_0/vcompp comparator_0/vo1 1.27fF
C1290 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_238313_n148007# 0.03fF
C1291 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm 0.51fF
C1292 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d VDD 11.46fF
C1293 a_244971_n121167# VDD 0.15fF
C1294 a_242273_n120623# a_242526_n120511# 0.04fF
C1295 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail2 0.58fF
C1296 dac_8bit_0/amux_2to1_6/SELB VDD 1.15fF
C1297 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_225730_n140786# 0.82fF
C1298 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp 23.52fF
C1299 dac_8bit_0/latched_comparator_folded_0/vcompm_buf dac_8bit_0/latched_comparator_folded_0/vcompm 0.02fF
C1300 a_241919_n121161# a_242526_n121193# 0.37fF
C1301 input_amplifier_0/diff_fold_casc_ota_1/vfoldm vampp 5.90fF
C1302 a_336408_n185665# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/D 0.61fF
C1303 a_336608_n185510# a_336537_n185409# 0.59fF
C1304 a_242085_n120623# a_242526_n120511# 0.28fF
C1305 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc 16.79fF
C1306 input_amplifier_0/diff_fold_casc_ota_1/vcascnm input_amplifier_0/diff_fold_casc_ota_1/vcascnp 12.37fF
C1307 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/vip 0.28fF
C1308 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc 0.16fF
C1309 vpeak_sampled sample 14.19fF
C1310 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 33.98fF
C1311 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn2 vintp 2.15fF
C1312 vintm biquad_gm_c_filter_0/gm_c_stage_1/vcmc 0.10fF
C1313 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn1 biquad_gm_c_filter_0/gm_c_stage_2/vcmc 2.37fF
C1314 a_242783_n122255# a_242783_n121345# 0.07fF
C1315 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/vim1 3.14fF
C1316 input_amplifier_0/vip2 input_amplifier_0/rst 0.93fF
C1317 a_239330_n127742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/csinvp 0.16fF
C1318 a_336401_n185269# a_336608_n185510# 0.01fF
C1319 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_5/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_4/A 0.04fF
C1320 a_242085_n120623# a_242085_n121161# 0.06fF
C1321 a_244783_n121161# a_245649_n121193# 0.11fF
C1322 a_245224_n121193# a_245056_n121167# 0.59fF
C1323 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/A 0.01fF
C1324 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VDD 1.46fF
C1325 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y 0.01fF
C1326 a_241634_n115151# VDD 0.29fF
C1327 a_245649_n122281# a_245649_n122531# 0.09fF
C1328 dac_8bit_1/c6m dac_8bit_1/c4m 1.44fF
C1329 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VDD 25.41fF
C1330 a_242484_n121711# a_242358_n121345# 0.02fF
C1331 a_242104_n140786# a_243020_n140786# 1.33fF
C1332 a_241646_n140786# a_243478_n140786# 0.24fF
C1333 a_222956_n127742# a_223414_n127742# 0.02fF
C1334 a_221582_n127742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/csinvp 0.08fF
C1335 dac_8bit_1/c3m dac_8bit_1/amux_2to1_4/B 1.72fF
C1336 a_336116_n185269# a_336608_n185269# 0.03fF
C1337 input_amplifier_0/vip1 input_amplifier_0/vom1 29.62fF
C1338 vincm input_amplifier_0/vim1 39.51fF
C1339 a_336408_n184969# a_336401_n185269# 2.23fF
C1340 input_amplifier_0/rst input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc 0.11fF
C1341 diff_to_se_converter_0/ibiasn peak_detector_0/ibiasn1 0.76fF
C1342 vcp a_222854_n150168# 0.03fF
C1343 biquad_gm_c_filter_0/ibiasn3 peak_detector_0/ibiasn2 0.41fF
C1344 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/A 0.01fF
C1345 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y 0.01fF
C1346 a_242951_n121193# a_242951_n121443# 0.09fF
C1347 dac_8bit_0/c4m VDD 2.41fF
C1348 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d 0.82fF
C1349 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs VDD 4.44fF
C1350 input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 0.12fF
C1351 input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc 28.15fF
C1352 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vcascnm 10.63fF
C1353 vintp biquad_gm_c_filter_0/gm_c_stage_2/vcmc 0.10fF
C1354 vampp input_amplifier_0/vip2 0.80fF
C1355 sample sample_and_hold_1/vhold 4.50fF
C1356 dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 14.42fF
C1357 vampp input_amplifier_0/diff_fold_casc_ota_1/M13d 9.72fF
C1358 a_245649_n121443# a_246080_n121389# 0.31fF
C1359 dac_8bit_1/latched_comparator_folded_0/vcompp VDD 6.16fF
C1360 input_amplifier_0/diff_fold_casc_ota_1/M3d vampp 0.98fF
C1361 a_245481_n123343# VDD 0.22fF
C1362 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/vhold 1.41fF
C1363 peak_detector_0/ibiasn1 vbiasp 4.09fF
C1364 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 10.85fF
C1365 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d 0.81fF
C1366 vcp a_222854_n132168# 0.03fF
C1367 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_228771_n148007# 0.03fF
C1368 vintm biquad_gm_c_filter_0/gm_c_stage_1/vbiasp 0.61fF
C1369 a_338285_n185243# VDD 0.23fF
C1370 a_245056_n122433# a_245649_n122531# 0.02fF
C1371 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q a_244971_n122799# 0.02fF
C1372 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/B VDD 0.43fF
C1373 a_245224_n122687# a_245481_n122433# 0.11fF
C1374 vintp biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail2 0.32fF
C1375 dac_8bit_1/c0m dac_8bit_1/amux_2to1_9/Y 1.72fF
C1376 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q 0.07fF
C1377 sample dac_8bit_1/amux_2to1_1/B 2.66fF
C1378 a_239361_n114883# a_239708_n115125# 0.13fF
C1379 low_freq_pll_0/pfd_cp_lpf_0/vRSTN a_239883_n115151# 0.70fF
C1380 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q 0.42fF
C1381 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail2 0.58fF
C1382 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn1 biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail1 0.58fF
C1383 a_238872_n145742# VDD 0.09fF
C1384 dac_8bit_0/c7m dac_8bit_0/amux_2to1_0/B 2.37fF
C1385 vampp input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 2.44fF
C1386 a_245649_n121443# VDD 0.45fF
C1387 biquad_gm_c_filter_0/gm_c_stage_1/vcmc biquad_gm_c_filter_0/gm_c_stage_1/vtail_diff 0.03fF
C1388 vfiltp biquad_gm_c_filter_0/gm_c_stage_3/vbiasp 0.68fF
C1389 dac_8bit_0/comp_outm dac_8bit_0/latched_comparator_folded_0/vcompp_buf 0.21fF
C1390 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/vop1 4.72fF
C1391 biquad_gm_c_filter_0/ibiasn1 biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail2 0.15fF
C1392 a_242358_n122255# a_242358_n122433# 0.08fF
C1393 a_244617_n122249# a_245649_n122281# 0.11fF
C1394 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y a_245056_n122255# 0.16fF
C1395 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/vip 6.29fF
C1396 a_247243_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.03fF
C1397 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q a_244971_n121167# 0.02fF
C1398 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn a_189446_n180872# 0.11fF
C1399 low_freq_pll_0/pfd_cp_lpf_0/vswitchl low_freq_pll_0/pfd_cp_lpf_0/vpdiode 0.08fF
C1400 a_241919_n121711# a_242273_n121711# 0.21fF
C1401 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD 7.64fF
C1402 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/B a_335749_n185813# 0.45fF
C1403 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y a_242273_n121167# 0.38fF
C1404 input_amplifier_0/diff_fold_casc_ota_0/vcascnm input_amplifier_0/diff_fold_casc_ota_0/vcascnp 12.37fF
C1405 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y VDD 0.91fF
C1406 a_336401_n185269# a_337497_n185269# 0.07fF
C1407 a_336608_n185269# a_336955_n185243# 0.11fF
C1408 gain_ctrl_0 input_amplifier_0/venm1 0.55fF
C1409 a_227396_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.03fF
C1410 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/vim2 7.34fF
C1411 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/vhold 0.08fF
C1412 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm 2.41fF
C1413 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_226327_n138121# 0.03fF
C1414 a_222855_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin 0.03fF
C1415 dac_8bit_0/adc_run VDD 3.10fF
C1416 vintm biquad_gm_c_filter_0/gm_c_stage_3/vcmc 0.10fF
C1417 vpeak_sampled dac_8bit_1/amux_2to1_7/B 0.38fF
C1418 q0A vlowA 2.75fF
C1419 a_231327_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.03fF
C1420 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y a_246080_n123343# 0.11fF
C1421 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp VDD 19.81fF
C1422 vcp_sampled dac_8bit_0/amux_2to1_1/SELB 2.07fF
C1423 a_338356_n185510# a_338285_n185409# 0.59fF
C1424 dac_8bit_1/c1m dac_8bit_1/c0m 12.39fF
C1425 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin vcp 3.55fF
C1426 vse diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 9.01fF
C1427 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 8.02fF
C1428 a_223414_n145742# a_223872_n145742# 0.01fF
C1429 a_222956_n145742# a_224330_n145742# 0.01fF
C1430 input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/diff_fold_casc_ota_0/vbias1 11.84fF
C1431 a_237854_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin 0.03fF
C1432 a_222498_n145742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/csinvp 0.09fF
C1433 peak_detector_0/ibiasn2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp 0.16fF
C1434 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn2 biquad_gm_c_filter_0/gm_c_stage_3/vbiasp 0.88fF
C1435 sample dac_8bit_1/c7m 2.10fF
C1436 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d 0.21fF
C1437 a_244617_n122249# a_245056_n122433# 0.02fF
C1438 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_227854_n149500# 0.03fF
C1439 a_245056_n122255# a_244617_n122799# 0.02fF
C1440 biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail1 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn1 0.58fF
C1441 biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail2 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn 0.58fF
C1442 biquad_gm_c_filter_0/ibiasn3 biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail2 0.19fF
C1443 diff_to_se_converter_0/ibiasn vcp_sampled 0.51fF
C1444 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vbias3 1.29fF
C1445 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/diff_fold_casc_ota_0/vtail_casc 8.06fF
C1446 input_amplifier_0/diff_fold_casc_ota_1/M13d input_amplifier_0/diff_fold_casc_ota_1/vbias4 0.04fF
C1447 dac_8bit_0/amux_2to1_5/B vlowA 1.86fF
C1448 adc_vcaparrayB dac_8bit_1/cdumm 11.56fF
C1449 dac_8bit_0/amux_2to1_4/B vcp_sampled 0.38fF
C1450 input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_1/vbias3 0.02fF
C1451 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias4 1.53fF
C1452 biquad_gm_c_filter_0/gm_c_stage_0/vcmc VDD 2.70fF
C1453 a_242358_n121167# a_241919_n121711# 0.02fF
C1454 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn 3.02fF
C1455 dac_8bit_1/amux_2to1_3/B VDD 4.57fF
C1456 input_amplifier_0/vop1 input_amplifier_0/vim1 30.73fF
C1457 a_242783_n122255# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q 0.05fF
C1458 a_221582_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias 0.51fF
C1459 q0A sample 0.07fF
C1460 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d VDD 7.37fF
C1461 a_338149_n185569# a_338156_n184969# 0.02fF
C1462 a_338156_n185665# a_337864_n185269# 0.01fF
C1463 sample dac_8bit_0/amux_2to1_2/SELB 2.36fF
C1464 input_amplifier_0/vip2 input_amplifier_0/vim2 23.69fF
C1465 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_246080_n122255# 0.37fF
C1466 dac_8bit_1/amux_2to1_3/SELB dac_8bit_1/amux_2to1_3/B 1.51fF
C1467 a_236938_n150168# vcp 0.03fF
C1468 peak_detector_0/ibiasn1 vcp 0.21fF
C1469 dac_8bit_1/vcom_buf dac_8bit_1/ibiasp 0.02fF
C1470 input_amplifier_0/diff_fold_casc_ota_0/vbias3 vocm 12.04fF
C1471 vcp_sampled a_275374_n146348# 21.33fF
C1472 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn1 VDD 3.44fF
C1473 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_227702_n135628# 0.03fF
C1474 input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 0.36fF
C1475 q3B dac_8bit_1/amux_2to1_4/B 1.99fF
C1476 a_232702_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.03fF
C1477 vincm input_amplifier_0/txgate_4/txb 0.36fF
C1478 a_244617_n121711# a_245481_n121345# 0.09fF
C1479 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y a_245649_n121443# 0.17fF
C1480 vcp_sampled vbiasp 11.70fF
C1481 a_244617_n123337# VDD 0.78fF
C1482 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/vim 1.42fF
C1483 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_242855_n130007# 0.03fF
C1484 dac_8bit_0/amux_2to1_5/B sample 2.66fF
C1485 a_222498_n145742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin 0.25fF
C1486 vpeak_sampled dac_8bit_1/cdumm 1.94fF
C1487 input_amplifier_0/diff_fold_casc_ota_1/M2d input_amplifier_0/diff_fold_casc_ota_1/vbias1 11.84fF
C1488 a_246080_n123343# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.37fF
C1489 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin a_236939_n130007# 0.03fF
C1490 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y a_244783_n122799# 0.61fF
C1491 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q a_245649_n121443# 0.39fF
C1492 a_244617_n122799# a_245224_n122687# 0.37fF
C1493 VDD dac_8bit_1/amux_2to1_4/SELB 1.15fF
C1494 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VDD 2.04fF
C1495 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/vcom_buf 8.06fF
C1496 vcp a_228786_n119618# 0.03fF
C1497 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm 13.76fF
C1498 input_amplifier_0/diff_fold_casc_ota_0/M1d input_amplifier_0/diff_fold_casc_ota_0/vfoldm 13.09fF
C1499 input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/diff_fold_casc_ota_0/M6d 2.00fF
C1500 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vfoldp 6.84fF
C1501 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VDD 1.49fF
C1502 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q VDD 2.23fF
C1503 a_221582_n145742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs 0.82fF
C1504 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 6.00fF
C1505 a_337497_n185269# a_337592_n185269# 0.31fF
C1506 a_335844_n185269# a_336408_n184969# 0.11fF
C1507 a_242526_n122687# a_242783_n122433# 0.11fF
C1508 a_242358_n122433# a_242951_n122531# 0.02fF
C1509 low_freq_pll_0/cs_ring_osc_0/vosc a_223770_n131500# 0.03fF
C1510 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn biquad_gm_c_filter_0/gm_c_stage_1/vcmcn1 1.18fF
C1511 biquad_gm_c_filter_0/gm_c_stage_1/vbiasp biquad_gm_c_filter_0/gm_c_stage_1/vcmcn2 0.88fF
C1512 a_238923_n122049# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout 0.03fF
C1513 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q 0.02fF
C1514 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vcascnm 0.69fF
C1515 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 input_amplifier_0/vim2 0.10fF
C1516 input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vbias3 5.67fF
C1517 a_238770_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin 0.03fF
C1518 input_amplifier_0/diff_fold_casc_ota_1/M13d a_163060_n102324# 1.44fF
C1519 q6A q5A 9.23fF
C1520 comparator_0/ibiasn vpeak_sampled 0.57fF
C1521 dac_8bit_1/latched_comparator_folded_0/vcompm VDD 5.25fF
C1522 a_336784_n185787# VDD 0.02fF
C1523 vampm input_amplifier_0/diff_fold_casc_ota_1/vtail_casc 1.58fF
C1524 dac_8bit_0/vcom_buf dac_8bit_0/latched_comparator_folded_0/vlatchp 3.59fF
C1525 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn2 VDD 1.51fF
C1526 biquad_gm_c_filter_0/ibiasn2 vfiltm 0.16fF
C1527 a_242783_n122255# a_242867_n122255# 0.05fF
C1528 dac_8bit_0/ibiasn dac_8bit_0/c4m 0.19fF
C1529 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror a_189446_n180872# 8.05fF
C1530 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 0.61fF
C1531 dac_8bit_1/c5m VDD 2.56fF
C1532 dac_8bit_0/ibiasp dac_8bit_0/c4m 0.26fF
C1533 a_242562_n140786# VDD 0.14fF
C1534 a_241731_n115151# a_242380_n114857# 0.10fF
C1535 low_freq_pll_0/pfd_cp_lpf_0/VQBb VDD 0.42fF
C1536 a_242085_n122249# a_242085_n121711# 0.06fF
C1537 dac_8bit_0/amux_2to1_9/Y vrefA 1.93fF
C1538 dac_8bit_1/vcom_buf VDD 5.69fF
C1539 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 4.16fF
C1540 input_amplifier_0/diff_fold_casc_ota_0/vcascnp vocm 0.19fF
C1541 low_freq_pll_0/pfd_cp_lpf_0/vpbias low_freq_pll_0/ibiasn 0.05fF
C1542 dac_8bit_0/c2m dac_8bit_0/c1m 1.20fF
C1543 VDD a_245151_n122433# 0.02fF
C1544 dac_8bit_0/amux_2to1_16/SELB q6A 2.36fF
C1545 dac_8bit_0/latched_comparator_folded_0/vtailp vlowA 1.83fF
C1546 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_0/vholdm 0.86fF
C1547 peak_detector_0/ibiasn2 low_freq_pll_0/ibiasn 0.70fF
C1548 a_244783_n123337# a_244971_n123343# 0.26fF
C1549 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_9/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/A 0.35fF
C1550 dac_8bit_0/amux_2to1_4/SELB VDD 1.15fF
C1551 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vfoldp 6.84fF
C1552 input_amplifier_0/diff_fold_casc_ota_1/M1d input_amplifier_0/diff_fold_casc_ota_1/vfoldm 13.09fF
C1553 input_amplifier_0/diff_fold_casc_ota_1/M2d input_amplifier_0/diff_fold_casc_ota_1/M6d 2.00fF
C1554 low_freq_pll_0/cs_ring_osc_0/vpbias a_237956_n127742# 0.83fF
C1555 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/csinvn low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.09fF
C1556 a_236582_n127742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs 0.82fF
C1557 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp 0.08fF
C1558 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d 1.26fF
C1559 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/diff_fold_casc_ota_0/M6d 18.03fF
C1560 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc 0.09fF
C1561 input_amplifier_0/diff_fold_casc_ota_0/M1d input_amplifier_0/diff_fold_casc_ota_0/M3d 2.62fF
C1562 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/diff_fold_casc_ota_0/vbias2 1.45fF
C1563 a_228328_n122869# VDD 0.06fF
C1564 input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 2.44fF
C1565 dac_8bit_0/amux_2to1_7/B VDD 4.57fF
C1566 input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vcascnp 3.37fF
C1567 gain_ctrl_0 input_amplifier_0/txgate_0/txb 0.36fF
C1568 low_freq_pll_0/cs_ring_osc_0/vpbias low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/csinvp 0.31fF
C1569 dac_8bit_0/c3m vcp_sampled 1.94fF
C1570 a_245481_n122255# a_246080_n122255# 0.02fF
C1571 a_245649_n122281# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_8/A 0.04fF
C1572 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/vpeak 0.75fF
C1573 adc_clk a_338156_n184969# 0.23fF
C1574 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/vim 19.24fF
C1575 a_241919_n122249# a_242085_n122799# 0.09fF
C1576 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp 0.08fF
C1577 input_amplifier_0/diff_fold_casc_ota_0/vfoldm vocm 0.16fF
C1578 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/vhold 0.71fF
C1579 a_242783_n121167# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q 0.05fF
C1580 q6A dac_8bit_1/ibiasn 0.20fF
C1581 a_242358_n122255# a_242951_n122281# 0.02fF
C1582 a_242526_n122281# a_242783_n122255# 0.11fF
C1583 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/csinvn 0.09fF
C1584 a_239143_n115125# a_239883_n115151# 0.02fF
C1585 vcp_sampled vcp 0.12fF
C1586 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y 0.41fF
C1587 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/verr 13.64fF
C1588 a_242453_n121167# VDD 0.02fF
C1589 a_242453_n120257# a_242358_n120257# 0.04fF
C1590 dac_8bit_1/amux_2to1_3/B q4B 1.99fF
C1591 input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc 1.62fF
C1592 a_245224_n121599# a_244971_n121711# 0.04fF
C1593 dac_8bit_1/amux_2to1_4/SELB dac_8bit_1/c3m 1.59fF
C1594 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_226646_n140786# 0.22fF
C1595 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp vse 1.42fF
C1596 a_241919_n121161# a_242951_n121193# 0.11fF
C1597 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc 2.10fF
C1598 a_242085_n120623# a_242951_n120355# 0.11fF
C1599 a_242526_n120511# a_242358_n120257# 0.59fF
C1600 a_336537_n185409# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/D 0.04fF
C1601 dac_8bit_0/latched_comparator_folded_0/vcompm_buf dac_8bit_0/comp_outm 0.12fF
C1602 input_amplifier_0/diff_fold_casc_ota_1/M1d input_amplifier_0/diff_fold_casc_ota_1/M3d 2.62fF
C1603 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/vbias2 1.45fF
C1604 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/diff_fold_casc_ota_1/M6d 18.03fF
C1605 dac_8bit_1/latched_comparator_folded_0/vlatchp dac_8bit_1/latched_comparator_folded_0/vlatchm 3.86fF
C1606 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc 0.09fF
C1607 a_242453_n122433# VDD 0.02fF
C1608 a_236582_n127742# VDD 0.73fF
C1609 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.42fF
C1610 a_243382_n122255# a_243382_n121389# 0.04fF
C1611 input_amplifier_0/venp1 input_amplifier_0/vim2 2.01fF
C1612 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d 1.51fF
C1613 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/M3d 0.61fF
C1614 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc 2.70fF
C1615 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/vom1 2.33fF
C1616 dac_8bit_1/amux_2to1_2/B vrefB 2.44fF
C1617 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/D a_336408_n185665# 0.02fF
C1618 a_242526_n120511# a_242526_n121193# 0.05fF
C1619 a_242720_n114759# a_243138_n114759# 0.02fF
C1620 a_245056_n121167# a_245649_n121193# 0.02fF
C1621 a_241919_n122249# a_241919_n121711# 0.08fF
C1622 a_245224_n121193# a_245481_n121167# 0.11fF
C1623 q6B VDD 3.49fF
C1624 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin a_221022_n149500# 0.03fF
C1625 a_245481_n122255# a_245481_n122433# 0.05fF
C1626 a_242102_n114873# VDD 0.39fF
C1627 biquad_gm_c_filter_0/gm_c_stage_3/vcmc biquad_gm_c_filter_0/gm_c_stage_3/vtail_diff 0.03fF
C1628 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q a_242951_n121443# 0.39fF
C1629 a_242562_n140786# a_243478_n140786# 0.79fF
C1630 a_223414_n127742# a_223872_n127742# 0.01fF
C1631 dac_8bit_1/c7m dac_8bit_1/cdumm 0.86fF
C1632 a_222956_n127742# a_224330_n127742# 0.01fF
C1633 dac_8bit_1/c6m dac_8bit_1/c2m 2.04fF
C1634 dac_8bit_1/c5m dac_8bit_1/c3m 0.66fF
C1635 a_222498_n127742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/csinvp 0.09fF
C1636 a_241919_n122799# a_242526_n122687# 0.37fF
C1637 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y a_242085_n122799# 0.61fF
C1638 a_242885_n115125# a_242575_n114888# 0.07fF
C1639 q6A q4A 0.10fF
C1640 q6A dac_8bit_0/amux_2to1_1/B 1.99fF
C1641 a_336408_n184969# a_336537_n185243# 0.28fF
C1642 input_amplifier_0/diff_fold_casc_ota_0/M13d input_amplifier_0/diff_fold_casc_ota_0/vbias3 0.48fF
C1643 a_336401_n185269# a_336608_n185269# 0.63fF
C1644 vocm_filt biquad_gm_c_filter_0/gm_c_stage_3/vcmcn1 1.07fF
C1645 dac_8bit_0/cdumm VDD 2.41fF
C1646 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 0.03fF
C1647 dac_8bit_1/amux_2to1_13/SELB dac_8bit_1/amux_2to1_4/B 1.59fF
C1648 a_242085_n121161# a_242526_n121193# 0.28fF
C1649 vcp a_223770_n150168# 0.03fF
C1650 dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d 0.73fF
C1651 biquad_gm_c_filter_0/ibiasn2 biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail2 0.13fF
C1652 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 a_275374_n180872# 8.05fF
C1653 biquad_gm_c_filter_0/ibiasn2 peak_detector_0/ibiasn2 0.40fF
C1654 a_242783_n121167# a_242783_n121345# 0.05fF
C1655 vocm_filt vfiltm 0.78fF
C1656 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm 0.19fF
C1657 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 6.88fF
C1658 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn 0.61fF
C1659 input_amplifier_0/diff_fold_casc_ota_0/M3d vocm 0.07fF
C1660 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 12.94fF
C1661 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror a_275374_n180872# 8.05fF
C1662 q6B q5B 9.23fF
C1663 a_241919_n122249# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q 0.03fF
C1664 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A a_335844_n185460# 0.02fF
C1665 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm 16.88fF
C1666 dac_8bit_1/amux_2to1_8/SELB dac_8bit_1/c0m 1.59fF
C1667 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_241023_n148007# 0.03fF
C1668 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_1/vhold 0.86fF
C1669 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 3.47fF
C1670 peak_detector_0/ibiasn2 peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d 0.13fF
C1671 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/vop1 2.63fF
C1672 low_freq_pll_0/cs_ring_osc_0/vosc low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.40fF
C1673 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/A VDD 0.62fF
C1674 vpeak_sampled sample_and_hold_1/vholdm 44.75fF
C1675 sample dac_8bit_1/amux_2to1_1/SELB 2.36fF
C1676 diff_to_se_converter_0/rst vfiltm 0.65fF
C1677 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/vip2 2.97fF
C1678 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 a_275374_n146348# 8.05fF
C1679 dac_8bit_1/latched_comparator_folded_0/vcompp dac_8bit_1/latched_comparator_folded_0/vcomppb 0.23fF
C1680 dac_8bit_0/amux_2to1_0/SELB dac_8bit_0/c7m 1.59fF
C1681 dac_8bit_1/latched_comparator_folded_0/vlatchp adc_clk 0.39fF
C1682 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc 0.12fF
C1683 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp 1.94fF
C1684 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD 1.46fF
C1685 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin 0.38fF
C1686 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/M13d 1.61fF
C1687 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_10/A VDD 0.48fF
C1688 dac_8bit_1/ibiasp VDD 4.58fF
C1689 input_amplifier_0/diff_fold_casc_ota_1/vfoldm vampm 2.33fF
C1690 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc 2.70fF
C1691 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/M3d 0.61fF
C1692 vcp a_223770_n132168# 0.03fF
C1693 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs VDD 4.44fF
C1694 a_242783_n123343# a_242526_n123369# 0.11fF
C1695 a_245649_n121193# low_freq_pll_0/freq_div_0/vout 0.38fF
C1696 a_242783_n123343# VDD 0.22fF
C1697 a_245649_n122531# a_245481_n122433# 0.67fF
C1698 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d 1.51fF
C1699 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp vse 3.50fF
C1700 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 3.45fF
C1701 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/vom1 3.33fF
C1702 input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc 13.41fF
C1703 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/vhold 2.30fF
C1704 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm 28.76fF
C1705 a_335749_n185269# a_335844_n185269# 0.31fF
C1706 peak_detector_0/ibiasn2 vpeak 9.74fF
C1707 low_freq_pll_0/pfd_cp_lpf_0/vRSTN a_240447_n115125# 0.10fF
C1708 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_4/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/A 0.35fF
C1709 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d vse 0.73fF
C1710 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/csinvp VDD 0.48fF
C1711 dac_8bit_0/amux_2to1_7/SELB dac_8bit_0/amux_2to1_7/B 1.51fF
C1712 a_221582_n127742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.82fF
C1713 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc vocm 1.38fF
C1714 a_246080_n121389# VDD 0.37fF
C1715 peak_detector_0/ibiasn1 vpeak_sampled 10.65fF
C1716 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y 0.30fF
C1717 input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc vocm 1.38fF
C1718 vcp a_229954_n134960# 0.03fF
C1719 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 5.47fF
C1720 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y 0.01fF
C1721 a_242951_n122281# a_242951_n122531# 0.09fF
C1722 vocm_filt biquad_gm_c_filter_0/gm_c_stage_2/vtail_diff 1.19fF
C1723 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/vhold 6.29fF
C1724 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y a_245481_n122255# 0.14fF
C1725 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm 2.00fF
C1726 a_240730_n140786# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs 0.82fF
C1727 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/csinvp low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.10fF
C1728 vpeak_sampled dac_8bit_1/amux_2to1_7/SELB 2.07fF
C1729 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp 11.53fF
C1730 vlowA dac_8bit_0/amux_2to1_3/B 1.86fF
C1731 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm 3.14fF
C1732 vcp_sampled dac_8bit_0/amux_2to1_2/B 0.38fF
C1733 sample_and_hold_1/vhold sample_and_hold_1/vholdm 21.72fF
C1734 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 13.36fF
C1735 q5A dac_8bit_1/ibiasn 0.20fF
C1736 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin a_245412_n135628# 0.03fF
C1737 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/B a_336116_n185555# 0.04fF
C1738 input_amplifier_0/diff_fold_casc_ota_0/M6d input_amplifier_0/vop1 0.31fF
C1739 low_freq_pll_0/cs_ring_osc_0/vpbias a_222040_n127742# 0.66fF
C1740 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 8.42fF
C1741 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm 4.75fF
C1742 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror 2.23fF
C1743 a_337592_n185460# pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A 0.03fF
C1744 vampm input_amplifier_0/vip2 16.51fF
C1745 vcp low_freq_pll_0/cs_ring_osc_0/vpbias 13.40fF
C1746 a_241919_n121161# a_241919_n120623# 0.08fF
C1747 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_242085_n120623# 0.03fF
C1748 peak_detector_0/verr peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d 4.82fF
C1749 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc 6.12fF
C1750 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/D a_336955_n185243# 0.35fF
C1751 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 24.81fF
C1752 a_242085_n123337# a_242358_n123343# 0.38fF
C1753 VDD a_242526_n123369# 0.23fF
C1754 a_242273_n121167# VDD 0.15fF
C1755 vampm input_amplifier_0/diff_fold_casc_ota_1/M13d 3.51fF
C1756 input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc 0.16fF
C1757 input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc 16.79fF
C1758 a_228312_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.03fF
C1759 dac_8bit_1/latched_comparator_folded_0/vcompmb dac_8bit_1/comp_outm 0.03fF
C1760 input_amplifier_0/diff_fold_casc_ota_1/M3d vampm 3.23fF
C1761 input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc 13.41fF
C1762 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_227243_n138121# 0.03fF
C1763 a_223771_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin 0.03fF
C1764 vfiltm biquad_gm_c_filter_0/ibiasn4 0.17fF
C1765 a_232243_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.03fF
C1766 adc_vcaparrayB dac_8bit_1/adc_run 0.36fF
C1767 dac_8bit_1/amux_2to1_3/SELB VDD 1.15fF
C1768 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q 0.14fF
C1769 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/diff_fold_casc_ota_0/M13d 6.93fF
C1770 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror 4.50fF
C1771 sample dac_8bit_0/amux_2to1_3/B 2.66fF
C1772 q5B VDD 3.49fF
C1773 a_223414_n145742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/csinvp 0.10fF
C1774 a_223872_n145742# a_224330_n145742# 0.02fF
C1775 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y a_244783_n121161# 0.61fF
C1776 a_244617_n121161# a_245224_n121193# 0.37fF
C1777 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 13.66fF
C1778 vcomp VDD 10.91fF
C1779 input_amplifier_0/vip2 input_amplifier_0/vop1 0.79fF
C1780 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_228770_n149500# 0.03fF
C1781 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror 0.69fF
C1782 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm 3.14fF
C1783 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp 0.81fF
C1784 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d 7.88fF
C1785 peak_detector_0/ibiasn1 peak_detector_0/verr 0.51fF
C1786 q6A q3A 0.10fF
C1787 q5A q4A 9.15fF
C1788 dac_8bit_1/amux_2to1_3/B dac_8bit_1/amux_2to1_14/SELB 1.59fF
C1789 biquad_gm_c_filter_0/ibiasn2 biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail2 0.79fF
C1790 vampm input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 0.10fF
C1791 a_335749_n185813# VDD 0.38fF
C1792 vocm_filt biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail2 4.74fF
C1793 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/A 0.01fF
C1794 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_244971_n122255# 0.02fF
C1795 sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn 10.10fF
C1796 biquad_gm_c_filter_0/gm_c_stage_0/vbiasp vintm 0.51fF
C1797 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp 6.59fF
C1798 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/verr 3.50fF
C1799 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp 4.15fF
C1800 dac_8bit_0/amux_2to1_5/SELB sample 2.36fF
C1801 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_2/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q 0.07fF
C1802 q6B q4B 0.10fF
C1803 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_2/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/A 0.35fF
C1804 a_222498_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias 0.63fF
C1805 VDD dac_8bit_1/amux_2to1_5/B 4.57fF
C1806 input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc input_amplifier_0/vop1 0.70fF
C1807 vcp_sampled dac_8bit_0/c6m 1.94fF
C1808 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp 6.59fF
C1809 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/vholdm 5.59fF
C1810 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d 5.99fF
C1811 input_amplifier_0/txgate_1/txb input_amplifier_0/vim2 0.53fF
C1812 a_245151_n123343# VDD 0.02fF
C1813 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror vse 4.81fF
C1814 a_338149_n185569# a_338356_n185269# 0.01fF
C1815 a_338156_n185665# a_338149_n185269# 0.02fF
C1816 a_241919_n122249# a_242526_n122281# 0.37fF
C1817 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d 15.11fF
C1818 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp 7.95fF
C1819 a_237854_n150168# vcp 0.03fF
C1820 vlowB dac_8bit_1/amux_2to1_0/B 1.86fF
C1821 a_242526_n121599# VDD 0.23fF
C1822 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d a_356329_n113250# 0.79fF
C1823 dac_8bit_0/amux_2to1_15/SELB q5A 2.36fF
C1824 dac_8bit_0/amux_2to1_16/SELB dac_8bit_0/amux_2to1_1/B 1.59fF
C1825 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y a_246080_n121389# 0.11fF
C1826 diff_to_se_converter_0/vip diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm 0.75fF
C1827 biquad_gm_c_filter_0/gm_c_stage_2/vtail_diff biquad_gm_c_filter_0/ibiasn4 0.06fF
C1828 vintp biquad_gm_c_filter_0/gm_c_stage_3/vcmcn1 0.78fF
C1829 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_243771_n130007# 0.03fF
C1830 dac_8bit_0/c0m dac_8bit_0/c5m 0.43fF
C1831 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 9.20fF
C1832 dac_8bit_0/c1m dac_8bit_0/c4m 1.12fF
C1833 a_242273_n123343# a_242273_n122799# 0.02fF
C1834 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin a_237855_n130007# 0.03fF
C1835 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/M13d 0.18fF
C1836 a_244617_n122799# a_245649_n122531# 0.11fF
C1837 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y a_245056_n122433# 0.16fF
C1838 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q a_246080_n121389# 0.37fF
C1839 vintp vfiltm 3.06fF
C1840 vintm biquad_gm_c_filter_0/gm_c_stage_2/vcmcn 2.62fF
C1841 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_6/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/A 0.35fF
C1842 sample dac_8bit_0/c5m 2.16fF
C1843 a_236582_n127742# a_237498_n127742# 2.99fF
C1844 a_222498_n145742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs 0.22fF
C1845 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d 3.07fF
C1846 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp 13.60fF
C1847 dac_8bit_1/c4m dac_8bit_1/amux_2to1_3/B 1.72fF
C1848 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp 0.81fF
C1849 a_337592_n185269# a_337864_n185269# 0.67fF
C1850 a_335844_n185269# a_336608_n185269# 0.02fF
C1851 a_244971_n121711# a_244971_n121167# 0.02fF
C1852 a_242951_n122531# a_242783_n122433# 0.67fF
C1853 vcp_sampled vpeak_sampled 4.14fF
C1854 dac_8bit_0/cdumm dac_8bit_0/ibiasn 0.19fF
C1855 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y VDD 0.93fF
C1856 vocm_filt biquad_gm_c_filter_0/gm_c_stage_1/vcmcn1 1.07fF
C1857 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp 0.28fF
C1858 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d 0.70fF
C1859 a_338703_n185409# VDD 0.16fF
C1860 dac_8bit_0/cdumm dac_8bit_0/ibiasp 0.42fF
C1861 low_freq_pll_0/freq_div_0/vin VDD 1.03fF
C1862 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/vholdm 2.13fF
C1863 a_242358_n122255# a_241919_n122799# 0.02fF
C1864 a_244617_n122249# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y 0.35fF
C1865 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_244783_n122249# 0.09fF
C1866 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail2 0.58fF
C1867 a_337497_n185813# VDD 0.35fF
C1868 q4A dac_8bit_1/ibiasn 0.20fF
C1869 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp 0.73fF
C1870 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/verr 0.73fF
C1871 a_242102_n114873# a_242419_n114983# 0.27fF
C1872 a_243478_n140786# VDD 0.06fF
C1873 a_241731_n115151# a_242575_n114888# 0.02fF
C1874 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q VDD 2.23fF
C1875 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d a_162668_n147576# 1.44fF
C1876 VDD dac_8bit_1/c3m 2.41fF
C1877 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d 0.16fF
C1878 a_242085_n121711# a_242358_n121345# 0.38fF
C1879 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 vse 0.08fF
C1880 q6A q1A 0.10fF
C1881 sample sample_and_hold_0/vhold 4.52fF
C1882 q7A vlowA 2.75fF
C1883 dac_8bit_0/amux_2to1_7/SELB VDD 1.15fF
C1884 VDD a_245565_n122433# 0.02fF
C1885 diff_to_se_converter_0/vip VDD 1.80fF
C1886 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d 0.12fF
C1887 a_245056_n123343# a_244971_n123343# 0.11fF
C1888 peak_detector_0/ibiasn2 biquad_gm_c_filter_0/ibiasn4 0.42fF
C1889 dac_8bit_1/ibiasp dac_8bit_0/ibiasp 5.08fF
C1890 low_freq_pll_0/cs_ring_osc_0/vpbias a_238872_n127742# 0.92fF
C1891 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d VDD 11.46fF
C1892 vintp biquad_gm_c_filter_0/gm_c_stage_2/vtail_diff 2.75fF
C1893 a_237498_n127742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs 0.22fF
C1894 q4B VDD 3.49fF
C1895 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm 3.14fF
C1896 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 13.36fF
C1897 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp 11.53fF
C1898 a_236633_n122049# VDD 0.01fF
C1899 dac_8bit_1/c5m dac_8bit_1/c4m 1.41fF
C1900 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn 8.02fF
C1901 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 0.56fF
C1902 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 58.37fF
C1903 q5A q3A 0.10fF
C1904 q6A q2A 0.10fF
C1905 a_244617_n122249# a_244617_n122799# 0.20fF
C1906 vocm_filt biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail2 2.82fF
C1907 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp 0.08fF
C1908 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d 0.75fF
C1909 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d 3.60fF
C1910 a_246080_n122255# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_8/A 0.25fF
C1911 dac_8bit_1/latched_comparator_folded_0/vcompp dac_8bit_1/comp_outm 0.08fF
C1912 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm vpeak 16.67fF
C1913 adc_clk a_338356_n185269# 0.04fF
C1914 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp a_275374_n180872# 10.36fF
C1915 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 1.13fF
C1916 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d 0.75fF
C1917 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d 3.60fF
C1918 a_241919_n122249# a_242358_n122433# 0.02fF
C1919 q5B q4B 9.15fF
C1920 q6B q3B 0.10fF
C1921 vse vfiltp 0.29fF
C1922 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d 1.51fF
C1923 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_1/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q 0.07fF
C1924 VDD rst_n 2.71fF
C1925 dac_8bit_1/ibiasn dac_8bit_0/c7m 0.20fF
C1926 a_242951_n122281# a_242783_n122255# 0.67fF
C1927 input_amplifier_0/venp1 input_amplifier_0/vop1 29.41fF
C1928 a_239883_n115151# a_239708_n115125# 0.62fF
C1929 dac_8bit_1/amux_2to1_15/SELB VDD 1.15fF
C1930 a_245056_n121345# a_245151_n121345# 0.04fF
C1931 a_242273_n123343# a_242085_n123337# 0.26fF
C1932 dac_8bit_0/ibiasn VDD 2.20fF
C1933 dac_8bit_0/ibiasp VDD 2.69fF
C1934 a_242526_n120511# a_242783_n120257# 0.11fF
C1935 peak_detector_0/ibiasn2 input_amplifier_0/ibiasn2 2.51fF
C1936 a_242358_n120257# a_242951_n120355# 0.02fF
C1937 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn 3.02fF
C1938 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp 4.15fF
C1939 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d 0.56fF
C1940 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_0/Q_N VDD 0.31fF
C1941 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q a_242085_n123337# 0.08fF
C1942 a_244783_n122799# a_244971_n122799# 0.26fF
C1943 vcp sample_and_hold_0/vholdm 8.80fF
C1944 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VDD 11.66fF
C1945 a_237498_n127742# VDD 0.40fF
C1946 a_236022_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.03fF
C1947 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn 5.68fF
C1948 vcp a_236022_n132168# 0.03fF
C1949 dac_8bit_1/amux_2to1_15/SELB q5B 2.36fF
C1950 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_2/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_3/A 0.04fF
C1951 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y 0.29fF
C1952 a_242783_n120257# a_242085_n121161# 0.01fF
C1953 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp adc_vcaparrayB 0.86fF
C1954 a_242358_n120257# a_242358_n121167# 0.05fF
C1955 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm 16.88fF
C1956 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 3.47fF
C1957 a_242085_n120623# a_242783_n121167# 0.01fF
C1958 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y 0.13fF
C1959 sample dac_8bit_1/amux_2to1_2/B 2.66fF
C1960 dac_8bit_1/amux_2to1_4/B vrefB 2.44fF
C1961 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin a_221938_n149500# 0.03fF
C1962 a_245649_n121193# a_245481_n121167# 0.67fF
C1963 a_242419_n114983# VDD 0.89fF
C1964 a_246080_n122255# a_246080_n122477# 0.04fF
C1965 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm 20.84fF
C1966 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q a_243382_n121389# 0.37fF
C1967 a_223872_n127742# a_224330_n127742# 0.02fF
C1968 a_223414_n127742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/csinvp 0.10fF
C1969 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y a_242358_n122433# 0.16fF
C1970 a_241919_n122799# a_242951_n122531# 0.11fF
C1971 a_336608_n185269# a_336537_n185243# 0.59fF
C1972 a_336401_n185269# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/D 0.42fF
C1973 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror 17.44fF
C1974 a_242526_n121193# a_242358_n121167# 0.59fF
C1975 low_freq_pll_0/cs_ring_osc_0/vpbias a_225730_n140786# 0.51fF
C1976 a_242085_n121161# a_242951_n121193# 0.11fF
C1977 biquad_gm_c_filter_0/ibiasn1 peak_detector_0/ibiasn2 0.40fF
C1978 a_243382_n121167# a_243382_n121389# 0.04fF
C1979 a_244783_n121161# a_244971_n121167# 0.26fF
C1980 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d vpeak 0.58fF
C1981 q3A dac_8bit_1/ibiasn 0.20fF
C1982 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d 1.26fF
C1983 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A a_336401_n185569# 0.03fF
C1984 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d 5.21fF
C1985 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_241939_n148007# 0.03fF
C1986 vcomp a_242419_n114983# 0.51fF
C1987 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 28.76fF
C1988 peak_detector_0/verr peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 12.80fF
C1989 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn 9.20fF
C1990 comparator_0/vcompp comparator_0/vcompm 7.44fF
C1991 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/csinvp 0.10fF
C1992 q5A q1A 0.10fF
C1993 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn vse 10.10fF
C1994 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn VDD 4.05fF
C1995 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 1.11fF
C1996 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 a_356329_n164260# 8.05fF
C1997 adc_clk a_338703_n185243# 0.05fF
C1998 input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 0.37fF
C1999 input_amplifier_0/vip2 input_amplifier_0/venm1 2.01fF
C2000 q6B q1B 0.10fF
C2001 diff_to_se_converter_0/vim diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm 2.13fF
C2002 vpeak_sampled dac_8bit_1/amux_2to1_9/Y 0.38fF
C2003 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp 0.73fF
C2004 a_242783_n123343# a_242951_n123369# 0.67fF
C2005 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d 2.62fF
C2006 a_245649_n122531# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_9/A 0.04fF
C2007 low_freq_pll_0/pfd_cp_lpf_0/vswitchl low_freq_pll_0/pfd_cp_lpf_0/vQB 0.44fF
C2008 a_245481_n122433# a_246080_n122477# 0.02fF
C2009 a_246080_n121167# low_freq_pll_0/freq_div_0/vout 0.37fF
C2010 a_239239_n115125# a_239143_n115125# 0.07fF
C2011 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_5/A VDD 0.48fF
C2012 adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn 2.30fF
C2013 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 28.76fF
C2014 vintp biquad_gm_c_filter_0/gm_c_stage_1/vcmcn1 0.15fF
C2015 vcp_sampled dac_8bit_0/amux_2to1_2/SELB 2.07fF
C2016 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm adc_vcaparrayB 6.31fF
C2017 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm 2.00fF
C2018 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp 24.81fF
C2019 q3B VDD 3.49fF
C2020 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VDD 1.49fF
C2021 a_244971_n122255# VDD 0.15fF
C2022 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror 2.23fF
C2023 sample dac_8bit_1/c6m 2.17fF
C2024 q5A q2A 0.10fF
C2025 q4A q3A 7.24fF
C2026 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d 7.88fF
C2027 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp 3.66fF
C2028 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm 5.03fF
C2029 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror 0.69fF
C2030 a_238627_n115125# VDD 0.90fF
C2031 a_222498_n127742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.22fF
C2032 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin VDD 4.26fF
C2033 dac_8bit_0/amux_2to1_17/SELB vlowA 1.62fF
C2034 adc_compA adc_clk 0.05fF
C2035 adc_vcaparrayB dac_8bit_1/c1m 18.08fF
C2036 dac_8bit_0/amux_2to1_5/B vcp_sampled 0.38fF
C2037 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d 1.91fF
C2038 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror 14.22fF
C2039 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp 1.03fF
C2040 dac_8bit_0/amux_2to1_6/B vlowA 1.86fF
C2041 a_242783_n122255# a_242783_n122433# 0.05fF
C2042 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_8/A 0.27fF
C2043 q6B q2B 0.10fF
C2044 q5B q3B 0.10fF
C2045 a_241646_n140786# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs 0.22fF
C2046 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin a_246328_n135628# 0.03fF
C2047 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/B a_336408_n185665# 0.01fF
C2048 low_freq_pll_0/cs_ring_osc_0/vpbias a_222956_n127742# 0.83fF
C2049 biquad_gm_c_filter_0/gm_c_stage_0/vbiasp vampm 0.12fF
C2050 sample dac_8bit_0/amux_2to1_3/SELB 2.36fF
C2051 low_freq_pll_0/cs_ring_osc_0/vosc a_221023_n130007# 0.03fF
C2052 a_338149_n185569# pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A 0.25fF
C2053 dac_8bit_1/amux_2to1_14/SELB VDD 1.15fF
C2054 a_242867_n120257# a_242783_n120257# 0.05fF
C2055 low_freq_pll_0/pfd_cp_lpf_0/vswitchh low_freq_pll_0/pfd_cp_lpf_0/vndiode 0.15fF
C2056 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/D a_337592_n185269# 0.37fF
C2057 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/rst 0.14fF
C2058 a_242526_n123369# a_242951_n123369# 0.04fF
C2059 dac_8bit_0/latched_comparator_folded_0/vlatchm adc_clk 0.68fF
C2060 dac_8bit_0/c1m dac_8bit_0/amux_2to1_7/B 1.72fF
C2061 dac_8bit_1/latched_comparator_folded_0/vcomppb VDD 0.47fF
C2062 dac_8bit_0/amux_2to1_14/SELB q4A 2.36fF
C2063 VDD a_242951_n123369# 0.45fF
C2064 a_242273_n120623# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y 0.38fF
C2065 diff_to_se_converter_0/vim VDD 1.92fF
C2066 a_241919_n121161# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y 0.35fF
C2067 biquad_gm_c_filter_0/ibiasn3 VDD 2.91fF
C2068 a_241919_n120623# a_242526_n120511# 0.37fF
C2069 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y a_242085_n120623# 0.61fF
C2070 low_freq_pll_0/cs_ring_osc_0/vosc VDD 8.63fF
C2071 q1A dac_8bit_1/ibiasn 0.20fF
C2072 diff_to_se_converter_0/ibiasn vse 1.71fF
C2073 dac_8bit_0/amux_2to1_6/B sample 2.66fF
C2074 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/csinvp low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.10fF
C2075 dac_8bit_0/vcom_buf vlowA 1.79fF
C2076 vpeak_sampled dac_8bit_1/c1m 1.94fF
C2077 VDD dac_8bit_1/amux_2to1_5/SELB 1.15fF
C2078 a_244783_n122249# VDD 0.43fF
C2079 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm 20.84fF
C2080 a_224330_n145742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/csinvp 0.16fF
C2081 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm 0.08fF
C2082 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 1.35fF
C2083 a_241919_n120623# a_242085_n121161# 0.02fF
C2084 a_335749_n185269# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/Q_N 0.21fF
C2085 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y a_245056_n121167# 0.16fF
C2086 a_244617_n121161# a_245649_n121193# 0.11fF
C2087 a_242085_n122799# a_242273_n122799# 0.26fF
C2088 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs VDD 4.44fF
C2089 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d 10.82fF
C2090 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y 0.41fF
C2091 q6B q7B 11.40fF
C2092 a_336116_n185555# VDD 0.22fF
C2093 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 13.66fF
C2094 q2A dac_8bit_1/ibiasn 0.20fF
C2095 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d 6.93fF
C2096 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm 2.00fF
C2097 low_freq_pll_0/pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/Q_N low_freq_pll_0/pfd_cp_lpf_0/vRSTN 0.08fF
C2098 a_240730_n140786# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.90fF
C2099 input_amplifier_0/venp2 VDD 3.10fF
C2100 dac_8bit_1/c4m VDD 2.41fF
C2101 a_223414_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias 0.76fF
C2102 q1B VDD 3.49fF
C2103 peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn 0.21fF
C2104 a_221582_n127742# VDD 0.73fF
C2105 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d 1.15fF
C2106 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 1.13fF
C2107 comparator_0/vcompm comparator_0/vtail 0.31fF
C2108 sample a_338149_n185269# 0.02fF
C2109 peak_detector_0/vpeak VDD 1.89fF
C2110 a_338356_n185510# a_338356_n185269# 0.05fF
C2111 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/vcom_buf 0.73fF
C2112 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y a_242358_n122255# 0.16fF
C2113 a_241919_n122249# a_242951_n122281# 0.11fF
C2114 a_238770_n150168# vcp 0.03fF
C2115 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q a_242085_n121711# 0.09fF
C2116 a_242951_n121443# VDD 0.45fF
C2117 q4A q1A 0.10fF
C2118 dac_8bit_1/amux_2to1_3/SELB dac_8bit_1/c4m 1.59fF
C2119 adc_vcaparrayA dac_8bit_0/c7m 854.85fF
C2120 dac_8bit_1/amux_2to1_5/SELB dac_8bit_1/amux_2to1_5/B 1.51fF
C2121 input_amplifier_0/vip1 input_amplifier_0/vim1 16.87fF
C2122 a_227104_n140786# a_227562_n140786# 0.02fF
C2123 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp 0.86fF
C2124 dac_8bit_0/cdumm dac_8bit_0/c1m 1.32fF
C2125 dac_8bit_0/c2m dac_8bit_0/c0m 0.39fF
C2126 q5B q1B 0.10fF
C2127 dac_8bit_0/ibiasn dac_8bit_0/ibiasp 8.77fF
C2128 diff_to_se_converter_0/ibiasn diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp 0.03fF
C2129 dac_8bit_0/c2m sample 2.36fF
C2130 a_335749_n185813# a_336116_n185555# 0.02fF
C2131 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y low_freq_pll_0/freq_div_0/vout 0.10fF
C2132 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/ibiasn 0.18fF
C2133 a_244783_n123337# a_245224_n123369# 0.28fF
C2134 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y a_245481_n122433# 0.14fF
C2135 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin a_238771_n130007# 0.03fF
C2136 q2B VDD 3.49fF
C2137 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror adc_vcaparrayA 1.41fF
C2138 a_236582_n127742# a_238414_n127742# 0.65fF
C2139 a_237040_n127742# a_237956_n127742# 2.26fF
C2140 a_337864_n185269# a_338156_n184969# 0.44fF
C2141 a_337592_n185269# a_338149_n185269# 0.11fF
C2142 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD 6.84fF
C2143 low_freq_pll_0/freq_div_0/vout low_freq_pll_0/pfd_cp_lpf_0/vQB 0.12fF
C2144 a_230870_n134960# vcp 0.03fF
C2145 a_242951_n122531# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_4/A 0.04fF
C2146 a_242783_n122433# a_243382_n122477# 0.02fF
C2147 q4A q2A 0.10fF
C2148 vrefA vlowA 9.06fF
C2149 dac_8bit_0/amux_2to1_9/Y VDD 4.57fF
C2150 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q a_242273_n122799# 0.02fF
C2151 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VDD 11.66fF
C2152 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 44.84fF
C2153 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 a_162668_n147576# 8.26fF
C2154 input_amplifier_0/venm1 input_amplifier_0/venp1 6.43fF
C2155 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d 0.16fF
C2156 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn 5.68fF
C2157 a_338532_n185787# VDD 0.02fF
C2158 input_amplifier_0/vip2 input_amplifier_0/txgate_0/txb 0.53fF
C2159 q5B q2B 0.10fF
C2160 q4B q3B 7.24fF
C2161 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VDD 11.66fF
C2162 adc_clk pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A 0.79fF
C2163 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d 2.72fF
C2164 a_337864_n185555# VDD 0.22fF
C2165 a_242358_n122255# a_242273_n122255# 0.11fF
C2166 vlowB dac_8bit_1/latched_comparator_folded_0/vlatchm 4.52fF
C2167 a_222040_n145742# VDD 1.55fF
C2168 a_242380_n114857# a_242575_n114888# 0.49fF
C2169 a_242102_n114873# a_242506_n114759# 0.13fF
C2170 a_242085_n121711# a_242783_n121345# 0.44fF
C2171 a_242526_n121599# a_242951_n121443# 0.04fF
C2172 a_242085_n122249# a_242783_n121345# 0.01fF
C2173 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_1/vcom_buf 0.58fF
C2174 dac_8bit_1/amux_2to1_13/SELB VDD 1.15fF
C2175 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD 7.64fF
C2176 input_amplifier_0/diff_fold_casc_ota_1/M2d VDD 9.25fF
C2177 VDD input_amplifier_0/diff_fold_casc_ota_0/M1d 10.42fF
C2178 dac_8bit_0/amux_2to1_1/SELB dac_8bit_0/amux_2to1_1/B 1.51fF
C2179 q2B dac_8bit_1/amux_2to1_5/B 1.99fF
C2180 dac_8bit_1/vcom_buf dac_8bit_1/latched_comparator_folded_0/vtailp 2.62fF
C2181 a_241919_n123337# a_242085_n123337# 2.23fF
C2182 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn VDD 4.05fF
C2183 adc_compA dac_8bit_0/latched_comparator_folded_0/vcompp 0.70fF
C2184 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d 5.48fF
C2185 dac_8bit_1/ibiasn vbiasp 2.20fF
C2186 VDD q7B 3.29fF
C2187 diff_to_se_converter_0/vim diff_to_se_converter_0/vip 22.65fF
C2188 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 a_189446_n180872# 8.26fF
C2189 dac_8bit_1/amux_2to1_14/SELB q4B 2.36fF
C2190 low_freq_pll_0/cs_ring_osc_0/vpbias low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/csinvp 0.31fF
C2191 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD 25.41fF
C2192 a_336359_n184877# VDD 0.02fF
C2193 a_242085_n122799# a_242085_n123337# 0.06fF
C2194 dac_8bit_1/amux_2to1_3/B vrefB 2.44fF
C2195 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout a_236632_n119618# 0.03fF
C2196 a_237549_n122049# VDD 0.01fF
C2197 peak_detector_0/ibiasn2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 0.13fF
C2198 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d VDD 9.36fF
C2199 dac_8bit_1/c5m dac_8bit_1/c2m 1.02fF
C2200 dac_8bit_1/c4m dac_8bit_1/c3m 1.18fF
C2201 dac_8bit_1/c6m dac_8bit_1/cdumm 0.86fF
C2202 dac_8bit_1/c7m dac_8bit_1/c1m 2.24fF
C2203 q5B q7B 0.10fF
C2204 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y 0.06fF
C2205 vcp low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin 4.28fF
C2206 dac_8bit_0/latched_comparator_folded_0/vlatchp VDD 4.86fF
C2207 dac_8bit_0/c1m VDD 2.47fF
C2208 vlowB adc_clk 0.47fF
C2209 adc_clk pulse_generator_0/sky130_fd_sc_hd__inv_1_0/Y 0.41fF
C2210 dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 8.87fF
C2211 diff_to_se_converter_0/ibiasn input_amplifier_0/ibiasn1 0.26fF
C2212 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y 0.06fF
C2213 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/vcom_buf 5.70fF
C2214 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y a_244617_n122249# 0.04fF
C2215 a_242783_n122255# a_243382_n122255# 0.02fF
C2216 input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 0.13fF
C2217 a_242951_n122281# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_2/A 0.04fF
C2218 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/csinvp low_freq_pll_0/cs_ring_osc_0/vpbias 0.31fF
C2219 a_337864_n185269# a_338107_n184877# 0.05fF
C2220 biquad_gm_c_filter_0/ibiasn3 rst_n 0.19fF
C2221 input_amplifier_0/diff_fold_casc_ota_1/vfoldp VDD 17.12fF
C2222 low_freq_pll_0/pfd_cp_lpf_0/vRSTN a_241731_n115151# 0.70fF
C2223 a_239883_n115151# low_freq_pll_0/pfd_cp_lpf_0/vQB 0.39fF
C2224 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d VDD 9.36fF
C2225 sample dac_8bit_1/amux_2to1_2/SELB 2.36fF
C2226 q3A q1A 0.10fF
C2227 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d VDD 7.37fF
C2228 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vbias4 36.08fF
C2229 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vbias3 0.04fF
C2230 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias2 14.23fF
C2231 a_245565_n121167# VDD 0.02fF
C2232 input_amplifier_0/rst input_amplifier_0/vim2 2.20fF
C2233 adc_vcaparrayB vlowB 1.95fF
C2234 a_242273_n123343# a_242358_n123343# 0.11fF
C2235 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 12.94fF
C2236 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror a_356329_n113250# 8.05fF
C2237 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 0.61fF
C2238 q4B q1B 0.10fF
C2239 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn1 vocm_filt 1.07fF
C2240 peak_detector_rst pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/B 0.03fF
C2241 a_242951_n120355# a_242783_n120257# 0.67fF
C2242 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_245649_n121443# 0.02fF
C2243 vampp input_amplifier_0/diff_fold_casc_ota_1/vbias4 14.85fF
C2244 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q a_242085_n123337# 0.01fF
C2245 a_244617_n123337# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y 0.04fF
C2246 a_242085_n122249# a_242085_n122799# 0.05fF
C2247 a_245056_n122433# a_244971_n122799# 0.11fF
C2248 a_238414_n127742# VDD 0.14fF
C2249 a_236938_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.03fF
C2250 vcp a_236938_n132168# 0.03fF
C2251 input_amplifier_0/txgate_3/txb VDD 3.08fF
C2252 input_amplifier_0/ibiasn1 vbiasp 1.06fF
C2253 dac_8bit_1/amux_2to1_10/SELB VDD 1.15fF
C2254 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q a_244783_n122799# 0.08fF
C2255 a_244617_n122799# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y 0.35fF
C2256 input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc 3.62fF
C2257 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/A 0.03fF
C2258 VDD vocm 0.07fF
C2259 a_242951_n120355# a_242951_n121193# 0.09fF
C2260 a_337497_n185813# a_337864_n185555# 0.02fF
C2261 a_245481_n121167# a_246080_n121167# 0.02fF
C2262 a_245649_n121193# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_6/A 0.04fF
C2263 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin a_222854_n149500# 0.03fF
C2264 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_8/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_9/A 0.04fF
C2265 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/Q_N pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/Q_N 0.02fF
C2266 a_242506_n114759# VDD 0.32fF
C2267 sample dac_8bit_1/amux_2to1_4/B 2.66fF
C2268 q3A q2A 6.48fF
C2269 vampp vintm 0.44fF
C2270 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y a_242783_n122433# 0.14fF
C2271 a_224330_n127742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/csinvp 0.16fF
C2272 a_244971_n121711# VDD 0.15fF
C2273 a_336537_n185243# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/D 0.04fF
C2274 vampp input_amplifier_0/vim2 14.59fF
C2275 dac_8bit_1/comp_outm VDD 0.67fF
C2276 low_freq_pll_0/cs_ring_osc_0/vpbias a_226646_n140786# 0.63fF
C2277 a_242358_n121167# a_242951_n121193# 0.02fF
C2278 a_242526_n121193# a_242783_n121167# 0.11fF
C2279 dac_8bit_0/c3m dac_8bit_1/ibiasn 0.20fF
C2280 q4B q2B 0.10fF
C2281 comparator_0/ibiasn peak_detector_0/ibiasn2 8.91fF
C2282 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_1/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_3/A 0.04fF
C2283 VDD low_freq_pll_0/ibiasn 2.04fF
C2284 a_245056_n121167# a_244971_n121167# 0.11fF
C2285 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/vip 0.71fF
C2286 vpeak_sampled dac_8bit_1/amux_2to1_8/SELB 2.07fF
C2287 vcp_sampled dac_8bit_0/amux_2to1_3/B 0.38fF
C2288 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn2 vocm_filt 0.28fF
C2289 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d 2.72fF
C2290 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp 2.79fF
C2291 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror 6.00fF
C2292 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 a_189446_n180872# 8.05fF
C2293 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VDD 5.18fF
C2294 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_242855_n148007# 0.03fF
C2295 vintm vfiltp 0.71fF
C2296 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VDD 12.54fF
C2297 dac_8bit_1/amux_2to1_12/SELB VDD 1.15fF
C2298 a_241919_n121711# a_242085_n121711# 2.23fF
C2299 input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc VDD 8.68fF
C2300 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_0/vcom_buf 0.86fF
C2301 a_242085_n122249# a_241919_n121711# 0.02fF
C2302 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 24.81fF
C2303 pulse_generator_0/sky130_fd_sc_hd__inv_1_1/A a_335749_n185269# 0.05fF
C2304 VDD input_amplifier_0/vom1 5.57fF
C2305 sample sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 12.79fF
C2306 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A a_336408_n184969# 0.03fF
C2307 dac_8bit_0/amux_2to1_13/SELB q3A 2.36fF
C2308 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d VDD 7.37fF
C2309 comparator_0/vcompp vfiltm 0.28fF
C2310 dac_8bit_0/latched_comparator_folded_0/vcompp_buf VDD 0.53fF
C2311 vampp a_163060_n102324# 19.89fF
C2312 dac_8bit_0/amux_2to1_5/SELB vcp_sampled 2.07fF
C2313 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/A 0.62fF
C2314 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 1.35fF
C2315 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm 20.84fF
C2316 a_336359_n185787# VDD 0.02fF
C2317 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm 0.08fF
C2318 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn biquad_gm_c_filter_0/gm_c_stage_0/vcmc 0.05fF
C2319 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_5/A a_242951_n123369# 0.04fF
C2320 a_244617_n123337# a_244971_n123343# 0.21fF
C2321 vocm_filt biquad_gm_c_filter_0/gm_c_stage_0/vtail_diff 1.19fF
C2322 vfiltp biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail2 0.07fF
C2323 a_246080_n122477# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_9/A 0.25fF
C2324 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_226481_n148007# 0.03fF
C2325 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d VDD 11.46fF
C2326 a_242085_n122249# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q 0.03fF
C2327 dac_8bit_1/ibiasp dac_8bit_1/latched_comparator_folded_0/vtailp 1.91fF
C2328 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y 0.08fF
C2329 dac_8bit_0/amux_2to1_4/B q3A 1.99fF
C2330 a_239048_n115125# VDD 0.60fF
C2331 vincm input_amplifier_0/ibiasn1 0.20fF
C2332 a_242453_n122255# VDD 0.02fF
C2333 vse diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 3.47fF
C2334 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d a_162668_n147576# 0.79fF
C2335 peak_detector_0/ibiasn2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror 3.13fF
C2336 diff_to_se_converter_0/txgate_1/txb vfiltm 0.35fF
C2337 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y a_244617_n122799# 0.04fF
C2338 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d 3.07fF
C2339 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_240411_n138121# 0.03fF
C2340 q4B q7B 0.10fF
C2341 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn biquad_gm_c_filter_0/gm_c_stage_0/vcmcn1 1.18fF
C2342 a_225580_n122869# low_freq_pll_0/cs_ring_osc_0/vpbias 0.60fF
C2343 biquad_gm_c_filter_0/gm_c_stage_0/vbiasp biquad_gm_c_filter_0/gm_c_stage_0/vcmcn2 0.88fF
C2344 q5A dac_8bit_0/amux_2to1_2/B 1.99fF
C2345 a_239361_n114883# VDD 0.32fF
C2346 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d VDD 7.37fF
C2347 dac_8bit_1/amux_2to1_12/SELB dac_8bit_1/amux_2to1_5/B 1.59fF
C2348 dac_8bit_0/amux_2to1_7/SELB dac_8bit_0/c1m 1.59fF
C2349 a_243382_n122255# a_243382_n122477# 0.04fF
C2350 VDD dac_8bit_1/amux_2to1_17/SELB 1.15fF
C2351 a_244783_n122249# a_244971_n122255# 0.26fF
C2352 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc 2.12fF
C2353 diff_to_se_converter_0/ibiasn vfiltp 0.49fF
C2354 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vfoldm 0.12fF
C2355 dac_8bit_0/amux_2to1_6/SELB sample 2.36fF
C2356 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 33.98fF
C2357 VDD dac_8bit_1/amux_2to1_6/B 4.57fF
C2358 a_241919_n122249# a_241919_n122799# 0.20fF
C2359 vcp_sampled dac_8bit_0/c5m 1.94fF
C2360 a_243382_n121389# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/A 0.05fF
C2361 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin a_247244_n135628# 0.03fF
C2362 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 33.98fF
C2363 low_freq_pll_0/cs_ring_osc_0/vpbias a_223872_n127742# 0.92fF
C2364 biquad_gm_c_filter_0/gm_c_stage_2/vbiasp biquad_gm_c_filter_0/gm_c_stage_2/vcmcn 0.53fF
C2365 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/vcom_buf 24.36fF
C2366 low_freq_pll_0/cs_ring_osc_0/vosc a_221939_n130007# 0.03fF
C2367 a_338356_n185510# pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A 0.05fF
C2368 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD 25.41fF
C2369 q2A q1A 3.80fF
C2370 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_242783_n120257# 0.05fF
C2371 vlowB dac_8bit_1/amux_2to1_1/B 1.86fF
C2372 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs 0.40fF
C2373 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q 0.08fF
C2374 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/D a_338156_n184969# 0.01fF
C2375 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d VDD 11.46fF
C2376 q6B vrefB 0.88fF
C2377 dac_8bit_0/latched_comparator_folded_0/vlatchm dac_8bit_0/latched_comparator_folded_0/vcompm 0.54fF
C2378 q3B q1B 0.10fF
C2379 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y a_244971_n121711# 0.38fF
C2380 biquad_gm_c_filter_0/ibiasn2 VDD 1.26fF
C2381 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_242951_n121193# 0.02fF
C2382 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y a_242358_n120257# 0.16fF
C2383 a_241919_n120623# a_242951_n120355# 0.11fF
C2384 dac_8bit_1/latched_comparator_folded_0/vtailp VDD 1.69fF
C2385 input_amplifier_0/rst input_amplifier_0/diff_fold_casc_ota_0/vfoldp 0.11fF
C2386 dac_8bit_0/c0m dac_8bit_0/c4m 0.43fF
C2387 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm 5.03fF
C2388 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/A VDD 0.62fF
C2389 biquad_gm_c_filter_0/gm_c_stage_0/vcmc biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail1 0.15fF
C2390 dac_8bit_1/amux_2to1_9/SELB VDD 1.15fF
C2391 peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d VDD 1.27fF
C2392 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.06fF
C2393 a_245412_n134960# vcp 0.03fF
C2394 sample dac_8bit_0/c4m 2.36fF
C2395 a_241919_n121161# a_242273_n121167# 0.21fF
C2396 a_241919_n121161# VDD 0.79fF
C2397 a_245056_n122255# VDD 0.36fF
C2398 vcp_sampled sample_and_hold_0/vhold 4.88fF
C2399 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VDD 2.04fF
C2400 dac_8bit_0/c3m dac_8bit_0/c7m 1.31fF
C2401 a_241919_n120623# a_242358_n121167# 0.01fF
C2402 vintp biquad_gm_c_filter_0/gm_c_stage_0/vcmc 0.10fF
C2403 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 13.36fF
C2404 input_amplifier_0/rst vincm 0.92fF
C2405 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 28.69fF
C2406 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y a_245481_n121167# 0.14fF
C2407 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 2.79fF
C2408 peak_detector_0/ibiasn2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 0.21fF
C2409 a_242358_n122433# a_242273_n122799# 0.11fF
C2410 input_amplifier_0/txgate_6/txb VDD 3.08fF
C2411 a_241919_n122799# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y 0.35fF
C2412 dac_8bit_0/c1m dac_8bit_0/ibiasn 0.19fF
C2413 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn1 biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail1 0.58fF
C2414 biquad_gm_c_filter_0/gm_c_stage_0/vbiasp biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail2 0.90fF
C2415 dac_8bit_0/c1m dac_8bit_0/ibiasp 0.26fF
C2416 q3B q2B 6.48fF
C2417 dac_8bit_0/latched_comparator_folded_0/vtailp dac_8bit_0/latched_comparator_folded_0/vlatchm 1.85fF
C2418 a_336408_n185665# VDD 0.45fF
C2419 input_amplifier_0/diff_fold_casc_ota_1/M1d vampp 0.54fF
C2420 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y a_242085_n121161# 0.61fF
C2421 input_amplifier_0/diff_fold_casc_ota_1/vbias4 a_163060_n102324# 14.02fF
C2422 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc 0.86fF
C2423 a_241646_n140786# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.25fF
C2424 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn1 vintp 0.91fF
C2425 a_244783_n121161# VDD 0.43fF
C2426 a_224330_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias 0.77fF
C2427 low_freq_pll_0/pfd_cp_lpf_0/vQA a_241731_n115151# 0.39fF
C2428 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 32.00fF
C2429 vintm biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail2 0.32fF
C2430 biquad_gm_c_filter_0/ibiasn1 biquad_gm_c_filter_0/gm_c_stage_0/vcmc 0.11fF
C2431 VDD dac_8bit_1/c2m 2.47fF
C2432 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn1 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn2 0.17fF
C2433 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn biquad_gm_c_filter_0/gm_c_stage_2/vcmc 0.05fF
C2434 a_222498_n127742# VDD 0.40fF
C2435 dac_8bit_1/amux_2to1_11/SELB VDD 1.15fF
C2436 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/vim1 7.75fF
C2437 a_336116_n185269# VDD 0.22fF
C2438 a_338285_n185409# a_338285_n185243# 0.05fF
C2439 vpeak VDD 5.79fF
C2440 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y a_242783_n122255# 0.14fF
C2441 VDD input_amplifier_0/diff_fold_casc_ota_0/M13d 1.24fF
C2442 low_freq_pll_0/cs_ring_osc_0/vosc a_221582_n127742# 2.75fF
C2443 a_243382_n121389# VDD 0.37fF
C2444 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm 13.76fF
C2445 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VDD 11.66fF
C2446 comparator_0/vtail vfiltm 2.70fF
C2447 dac_8bit_0/amux_2to1_8/SELB VDD 1.15fF
C2448 low_freq_pll_0/pfd_cp_lpf_0/vswitchl low_freq_pll_0/pfd_cp_lpf_0/VQBb 0.28fF
C2449 a_227562_n140786# a_228020_n140786# 0.01fF
C2450 a_227104_n140786# a_228478_n140786# 0.01fF
C2451 input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc 0.22fF
C2452 adc_compA dac_8bit_0/latched_comparator_folded_0/vcomppb 0.03fF
C2453 input_amplifier_0/rst input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc 0.11fF
C2454 a_242273_n122255# a_242273_n121711# 0.02fF
C2455 dac_8bit_1/amux_2to1_13/SELB q3B 2.36fF
C2456 VDD a_245224_n122687# 0.23fF
C2457 a_225730_n140786# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.90fF
C2458 a_335844_n185460# a_336401_n185569# 0.11fF
C2459 a_242783_n123343# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y 0.14fF
C2460 dac_8bit_0/adc_run vlowA 0.35fF
C2461 a_244783_n123337# a_245649_n123369# 0.11fF
C2462 a_242273_n123343# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q 0.02fF
C2463 a_245224_n123369# a_245056_n123343# 0.59fF
C2464 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_9/A 0.27fF
C2465 input_amplifier_0/venm2 input_amplifier_0/vip2 44.02fF
C2466 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d 6.93fF
C2467 rst_n low_freq_pll_0/ibiasn 0.51fF
C2468 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc 2.12fF
C2469 a_242085_n122249# a_242526_n122281# 0.28fF
C2470 a_237498_n127742# a_238414_n127742# 1.92fF
C2471 a_237040_n127742# a_238872_n127742# 0.43fF
C2472 a_236582_n127742# a_239330_n127742# 0.14fF
C2473 a_338156_n184969# a_338149_n185269# 2.23fF
C2474 a_337592_n185269# a_338285_n185243# 0.04fF
C2475 a_337864_n185269# a_338356_n185269# 0.03fF
C2476 q3B q7B 0.10fF
C2477 a_243382_n122477# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_4/A 0.25fF
C2478 a_231786_n134960# vcp 0.03fF
C2479 comparator_0/vmirror VDD 2.51fF
C2480 dac_8bit_1/c2m dac_8bit_1/amux_2to1_5/B 1.72fF
C2481 dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 13.20fF
C2482 low_freq_pll_0/cs_ring_osc_0/vpbias a_237040_n145742# 0.66fF
C2483 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_1/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/A 0.35fF
C2484 input_amplifier_0/diff_fold_casc_ota_1/vbias2 vampp 1.14fF
C2485 peak_detector_0/ibiasn1 peak_detector_0/ibiasn2 5.18fF
C2486 VDD vrefB 29.33fF
C2487 rst_n input_amplifier_0/vom1 0.16fF
C2488 biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail1 biquad_gm_c_filter_0/gm_c_stage_0/vtail_diff 0.49fF
C2489 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d 5.99fF
C2490 a_338156_n185665# VDD 0.46fF
C2491 low_freq_pll_0/pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/Q_N low_freq_pll_0/pfd_cp_lpf_0/vRSTN 0.09fF
C2492 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/vim 2.37fF
C2493 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp 2.72fF
C2494 vintm biquad_gm_c_filter_0/gm_c_stage_1/vtail_diff 4.99fF
C2495 a_222956_n145742# VDD 0.69fF
C2496 dac_8bit_1/ibiasn dac_8bit_0/c6m 0.20fF
C2497 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/A 0.10fF
C2498 dac_8bit_0/c3m adc_vcaparrayA 29.30fF
C2499 a_242419_n114983# a_242506_n114759# 0.16fF
C2500 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/vhold 0.75fF
C2501 vintp biquad_gm_c_filter_0/gm_c_stage_0/vtail_diff 0.58fF
C2502 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/A 1.64fF
C2503 a_242358_n121345# a_242783_n121345# 0.03fF
C2504 dac_8bit_0/adc_run sample 0.38fF
C2505 dac_8bit_0/amux_2to1_4/B dac_8bit_0/amux_2to1_13/SELB 1.59fF
C2506 dac_8bit_0/amux_2to1_10/SELB q1A 2.36fF
C2507 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_240412_n135628# 0.03fF
C2508 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A a_335749_n185269# 0.50fF
C2509 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 13.36fF
C2510 dac_8bit_1/ibiasn adc_vcaparrayB 1.12fF
C2511 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_241919_n120623# 0.03fF
C2512 q6A q0A 0.10fF
C2513 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail1 0.58fF
C2514 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn1 biquad_gm_c_filter_0/gm_c_stage_3/vcmc 2.37fF
C2515 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d 1.15fF
C2516 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/verr 21.50fF
C2517 q5B vrefB 0.88fF
C2518 dac_8bit_0/amux_2to1_15/SELB dac_8bit_0/amux_2to1_2/B 1.59fF
C2519 a_241919_n123337# a_242358_n123343# 0.63fF
C2520 q2B q1B 3.80fF
C2521 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y a_242526_n123369# 0.15fF
C2522 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y 0.91fF
C2523 peak_detector_0/verr vse 1.09fF
C2524 vfiltp biquad_gm_c_filter_0/gm_c_stage_3/vtail_diff 2.76fF
C2525 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d 0.12fF
C2526 a_244783_n121711# a_245224_n121599# 0.28fF
C2527 vocm_filt VDD 1.73fF
C2528 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/vop1 4.33fF
C2529 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias3 0.02fF
C2530 biquad_gm_c_filter_0/ibiasn1 biquad_gm_c_filter_0/gm_c_stage_0/vtail_diff 0.06fF
C2531 vlowB dac_8bit_1/amux_2to1_16/SELB 1.62fF
C2532 a_242526_n122687# a_242526_n123369# 0.05fF
C2533 a_336955_n185243# VDD 0.15fF
C2534 a_337592_n185460# a_336401_n185569# 0.02fF
C2535 peak_detector_rst q6B 0.12fF
C2536 a_242526_n122687# VDD 0.23fF
C2537 input_amplifier_0/diff_fold_casc_ota_0/vbias4 a_217060_n102324# 14.02fF
C2538 a_243382_n123343# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q 0.45fF
C2539 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout a_237548_n119618# 0.03fF
C2540 sample dac_8bit_1/amux_2to1_3/B 2.66fF
C2541 dac_8bit_1/amux_2to1_5/B vrefB 2.44fF
C2542 diff_to_se_converter_0/rst VDD 0.64fF
C2543 a_238465_n122049# VDD 0.01fF
C2544 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q a_244783_n121161# 0.09fF
C2545 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/A 0.02fF
C2546 a_244617_n121161# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y 0.35fF
C2547 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_245649_n122531# 0.39fF
C2548 vampp gain_ctrl_1 0.45fF
C2549 dac_8bit_0/c6m dac_8bit_0/amux_2to1_1/B 2.37fF
C2550 dac_8bit_1/c3m dac_8bit_1/c2m 0.16fF
C2551 vampm vampp 31.15fF
C2552 input_amplifier_0/rst input_amplifier_0/vop1 9.48fF
C2553 dac_8bit_0/latched_comparator_folded_0/vcompm_buf VDD 0.53fF
C2554 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d 8.42fF
C2555 diff_to_se_converter_0/ibiasn vbiasp 3.91fF
C2556 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm 23.84fF
C2557 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/vpeak 28.95fF
C2558 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 3.45fF
C2559 vintm biquad_gm_c_filter_0/gm_c_stage_1/vcmcn2 2.12fF
C2560 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn 32.00fF
C2561 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp 0.28fF
C2562 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm 0.19fF
C2563 a_243382_n122255# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_2/A 0.25fF
C2564 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 6.88fF
C2565 vcp a_247702_n134960# 0.03fF
C2566 a_244971_n121711# a_244971_n122255# 0.02fF
C2567 biquad_gm_c_filter_0/ibiasn2 rst_n 0.18fF
C2568 q1B q7B 0.10fF
C2569 low_freq_pll_0/pfd_cp_lpf_0/vRSTN a_242380_n114857# 0.33fF
C2570 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/B a_335844_n185269# 0.01fF
C2571 a_240447_n115125# low_freq_pll_0/pfd_cp_lpf_0/vQB 0.59fF
C2572 vcp low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/csinvn 0.08fF
C2573 dac_8bit_0/amux_2to1_12/SELB q2A 2.36fF
C2574 sample dac_8bit_1/amux_2to1_4/SELB 2.36fF
C2575 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn1 biquad_gm_c_filter_0/gm_c_stage_3/vbiasp 0.19fF
C2576 input_amplifier_0/rst input_amplifier_0/txgate_5/txb 0.36fF
C2577 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y VDD 0.91fF
C2578 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs VDD 4.44fF
C2579 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp 0.73fF
C2580 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d 0.56fF
C2581 adc_compB dac_8bit_1/latched_comparator_folded_0/vcompp_buf 0.12fF
C2582 a_245481_n121345# a_245565_n121345# 0.05fF
C2583 vfiltm biquad_gm_c_filter_0/gm_c_stage_3/vbiasp 0.44fF
C2584 biquad_gm_c_filter_0/gm_c_stage_1/vcmc biquad_gm_c_filter_0/gm_c_stage_1/vcmcn1 2.37fF
C2585 biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail2 biquad_gm_c_filter_0/gm_c_stage_1/vbiasp 0.90fF
C2586 a_244971_n123343# VDD 0.15fF
C2587 biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail1 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn 0.58fF
C2588 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d VDD 1.27fF
C2589 biquad_gm_c_filter_0/ibiasn3 biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail1 0.07fF
C2590 dac_8bit_1/amux_2to1_0/SELB dac_8bit_1/amux_2to1_0/B 1.51fF
C2591 a_242783_n120257# a_243382_n120301# 0.02fF
C2592 a_242951_n120355# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_0/A 0.04fF
C2593 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp 4.15fF
C2594 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/diff_fold_casc_ota_0/vtail_casc 10.25fF
C2595 input_amplifier_0/diff_fold_casc_ota_1/M13d input_amplifier_0/diff_fold_casc_ota_1/vbias3 0.48fF
C2596 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vbias3 60.63fF
C2597 a_237854_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.03fF
C2598 a_239330_n127742# VDD 0.06fF
C2599 vcp a_237854_n132168# 0.03fF
C2600 vcp_sampled dac_8bit_0/amux_2to1_3/SELB 2.07fF
C2601 a_338356_n185510# a_338505_n185421# 0.02fF
C2602 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror vse 15.92fF
C2603 a_338156_n185665# a_338703_n185409# 0.26fF
C2604 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d 0.75fF
C2605 low_freq_pll_0/pfd_cp_lpf_0/VQBb low_freq_pll_0/freq_div_0/vout 0.10fF
C2606 a_275374_n146348# sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm 10.16fF
C2607 a_242783_n120257# a_242783_n121167# 0.07fF
C2608 a_337592_n185460# a_338149_n185569# 0.11fF
C2609 low_freq_pll_0/pfd_cp_lpf_0/vQA low_freq_pll_0/pfd_cp_lpf_0/vndiode 0.13fF
C2610 a_246080_n121167# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_6/A 0.25fF
C2611 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin a_223770_n149500# 0.03fF
C2612 sample dac_8bit_1/c5m 2.16fF
C2613 q2B q7B 0.10fF
C2614 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_226481_n130007# 0.03fF
C2615 a_221582_n145742# a_222498_n145742# 2.99fF
C2616 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_4/A 0.27fF
C2617 a_242396_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs 0.03fF
C2618 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn VDD 4.05fF
C2619 dac_8bit_0/c7m dac_8bit_0/c6m 2.04fF
C2620 dac_8bit_0/amux_2to1_7/B vlowA 1.86fF
C2621 adc_vcaparrayB dac_8bit_1/c0m 15.13fF
C2622 a_242951_n121193# a_242783_n121167# 0.67fF
C2623 dac_8bit_0/amux_2to1_6/B vcp_sampled 0.38fF
C2624 peak_detector_0/ibiasn2 vcp_sampled 6.54fF
C2625 low_freq_pll_0/cs_ring_osc_0/vpbias a_227562_n140786# 0.76fF
C2626 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 24.81fF
C2627 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/vim2 0.07fF
C2628 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q VDD 0.38fF
C2629 VDD biquad_gm_c_filter_0/ibiasn4 1.72fF
C2630 vintm biquad_gm_c_filter_0/gm_c_stage_3/vtail_diff 2.72fF
C2631 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn 3.02fF
C2632 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/vhold 0.71fF
C2633 biquad_gm_c_filter_0/ibiasn3 low_freq_pll_0/ibiasn 2.19fF
C2634 q7A dac_8bit_0/amux_2to1_0/B 1.99fF
C2635 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm 0.08fF
C2636 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror 4.50fF
C2637 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_244617_n122249# 0.51fF
C2638 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm 0.51fF
C2639 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 1.65fF
C2640 a_239048_n115125# a_238627_n115125# 0.23fF
C2641 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_243771_n148007# 0.03fF
C2642 sample dac_8bit_0/amux_2to1_4/SELB 2.36fF
C2643 a_240730_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias 0.51fF
C2644 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 13.36fF
C2645 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y a_242526_n121599# 0.15fF
C2646 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm 3.14fF
C2647 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp 11.53fF
C2648 a_241919_n121711# a_242358_n121345# 0.63fF
C2649 input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/diff_fold_casc_ota_0/vfoldp 1.90fF
C2650 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vfoldm 2.33fF
C2651 input_amplifier_0/txgate_3/txb input_amplifier_0/venp2 0.58fF
C2652 peak_detector_rst VDD 2.90fF
C2653 a_241919_n122249# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y 0.35fF
C2654 q5A q0A 0.10fF
C2655 peak_detector_0/verr peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d 9.65fF
C2656 q4B vrefB 0.88fF
C2657 a_238627_n115125# a_239361_n114883# 0.16fF
C2658 dac_8bit_1/amux_2to1_10/SELB q1B 2.36fF
C2659 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 3.02fF
C2660 biquad_gm_c_filter_0/gm_c_stage_1/vbiasp biquad_gm_c_filter_0/gm_c_stage_1/vcmcn1 0.19fF
C2661 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vtail_casc 1.56fF
C2662 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc 0.01fF
C2663 q6B q0B 0.10fF
C2664 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp 0.73fF
C2665 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d 2.62fF
C2666 vampm input_amplifier_0/diff_fold_casc_ota_1/vbias4 28.62fF
C2667 dac_8bit_0/amux_2to1_7/B sample 2.66fF
C2668 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn1 VDD 3.44fF
C2669 vocm_filt diff_to_se_converter_0/vip 30.61fF
C2670 vpeak_sampled dac_8bit_1/c0m 1.85fF
C2671 dac_8bit_0/c3m dac_8bit_0/amux_2to1_4/B 1.72fF
C2672 peak_detector_rst q5B 0.12fF
C2673 VDD dac_8bit_1/amux_2to1_6/SELB 1.15fF
C2674 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror 17.44fF
C2675 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm 2.41fF
C2676 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD 6.84fF
C2677 diff_to_se_converter_0/vip diff_to_se_converter_0/rst 0.40fF
C2678 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_241327_n138121# 0.03fF
C2679 a_226496_n122869# low_freq_pll_0/cs_ring_osc_0/vpbias 0.73fF
C2680 input_amplifier_0/diff_fold_casc_ota_0/vcascnm vocm 0.06fF
C2681 dac_8bit_1/amux_2to1_15/SELB vrefB 2.12fF
C2682 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm 4.75fF
C2683 vampm vintm 1.21fF
C2684 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 1.65fF
C2685 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror 14.22fF
C2686 a_241480_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs 0.03fF
C2687 low_freq_pll_0/pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/Q_N low_freq_pll_0/pfd_cp_lpf_0/vQA 0.13fF
C2688 vampm input_amplifier_0/vim2 1.34fF
C2689 a_226188_n140786# VDD 1.55fF
C2690 dac_8bit_0/c2m vcp_sampled 1.94fF
C2691 input_amplifier_0/ibiasn2 VDD 1.86fF
C2692 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_2/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_4/A 0.04fF
C2693 dac_8bit_0/comp_outm adc_compA 1.08fF
C2694 a_245056_n122255# a_244971_n122255# 0.11fF
C2695 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp 7.95fF
C2696 a_336359_n185787# a_336116_n185555# 0.05fF
C2697 a_336955_n185409# a_336401_n185569# 0.21fF
C2698 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/verr 15.92fF
C2699 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y 0.06fF
C2700 input_amplifier_0/diff_fold_casc_ota_1/M2d input_amplifier_0/diff_fold_casc_ota_1/vfoldp 1.90fF
C2701 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vfoldm 2.33fF
C2702 a_241919_n122249# a_242273_n122255# 0.21fF
C2703 vintp VDD 2.28fF
C2704 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/vholdm 4.81fF
C2705 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp 13.60fF
C2706 low_freq_pll_0/pfd_cp_lpf_0/vswitchh vcp 0.15fF
C2707 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d 3.07fF
C2708 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp 0.81fF
C2709 low_freq_pll_0/cs_ring_osc_0/vpbias low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/csinvp 0.31fF
C2710 low_freq_pll_0/cs_ring_osc_0/vosc a_222855_n130007# 0.03fF
C2711 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm vse 19.24fF
C2712 vocm_filt rst_n 0.22fF
C2713 input_amplifier_0/diff_fold_casc_ota_0/M1d input_amplifier_0/diff_fold_casc_ota_0/vbias2 6.85fF
C2714 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/diff_fold_casc_ota_0/M6d 10.15fF
C2715 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/M3d 5.14fF
C2716 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp 6.59fF
C2717 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d 5.99fF
C2718 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_0/A 0.07fF
C2719 adc_vcaparrayA dac_8bit_0/c6m 427.49fF
C2720 input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vcascnm 18.97fF
C2721 diff_to_se_converter_0/rst rst_n 0.23fF
C2722 a_242273_n123343# a_241919_n123337# 0.21fF
C2723 dac_8bit_1/amux_2to1_12/SELB q2B 2.36fF
C2724 q0A dac_8bit_1/ibiasn 0.20fF
C2725 vampm a_163060_n102324# 8.05fF
C2726 biquad_gm_c_filter_0/ibiasn1 VDD 7.42fF
C2727 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y a_242783_n120257# 0.14fF
C2728 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y 0.42fF
C2729 input_amplifier_0/vop1 input_amplifier_0/vim2 35.47fF
C2730 a_337592_n185460# adc_clk 0.20fF
C2731 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 8.02fF
C2732 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 58.37fF
C2733 dac_8bit_0/cdumm sample 2.36fF
C2734 biquad_gm_c_filter_0/ibiasn3 biquad_gm_c_filter_0/ibiasn2 24.60fF
C2735 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q a_241919_n123337# 0.49fF
C2736 a_244617_n122799# a_244971_n122799# 0.21fF
C2737 a_246328_n134960# vcp 0.03fF
C2738 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q 0.08fF
C2739 a_245481_n122255# VDD 0.22fF
C2740 a_336955_n185243# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.04fF
C2741 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_6/A 0.27fF
C2742 a_242085_n122799# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q 0.03fF
C2743 a_242358_n122255# VDD 0.36fF
C2744 a_242453_n120257# VDD 0.02fF
C2745 input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vbias4 14.85fF
C2746 a_242526_n120511# VDD 0.23fF
C2747 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y a_242358_n121167# 0.16fF
C2748 a_336537_n185409# VDD 0.23fF
C2749 sample_and_hold_0/vhold sample_and_hold_0/vholdm 21.72fF
C2750 a_244783_n122249# a_245056_n122255# 0.38fF
C2751 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/M3d 5.14fF
C2752 input_amplifier_0/diff_fold_casc_ota_1/M1d input_amplifier_0/diff_fold_casc_ota_1/vbias2 6.85fF
C2753 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/M6d 10.15fF
C2754 a_244617_n121161# a_244971_n121167# 0.21fF
C2755 a_245056_n121167# VDD 0.36fF
C2756 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm 0.08fF
C2757 q0B VDD 3.49fF
C2758 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 1.35fF
C2759 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/verr 7.98fF
C2760 dac_8bit_1/ibiasp sample 0.46fF
C2761 a_337592_n185460# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_2/Q 0.33fF
C2762 a_336401_n185269# VDD 0.81fF
C2763 a_223414_n127742# VDD 0.14fF
C2764 a_242085_n121161# a_242273_n121167# 0.26fF
C2765 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp 4.15fF
C2766 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/vholdm 0.08fF
C2767 input_amplifier_0/diff_fold_casc_ota_0/M1d input_amplifier_0/vom1 14.05fF
C2768 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc 0.08fF
C2769 a_242085_n121161# VDD 0.43fF
C2770 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc 0.15fF
C2771 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_2/A 0.27fF
C2772 low_freq_pll_0/cs_ring_osc_0/vosc a_222498_n127742# 0.25fF
C2773 q4A q0A 0.10fF
C2774 q3B vrefB 0.88fF
C2775 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_236023_n148007# 0.03fF
C2776 dac_8bit_1/amux_2to1_5/SELB dac_8bit_1/c2m 1.59fF
C2777 a_228020_n140786# a_228478_n140786# 0.02fF
C2778 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q a_241919_n122249# 0.49fF
C2779 vocm_filt biquad_gm_c_filter_0/gm_c_stage_3/vcmcn 2.51fF
C2780 vlowA VDD 44.16fF
C2781 q5B q0B 0.10fF
C2782 VDD a_245649_n122531# 0.45fF
C2783 biquad_gm_c_filter_0/ibiasn2 biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail1 0.07fF
C2784 a_336116_n185555# a_336408_n185665# 0.44fF
C2785 a_335844_n185460# a_336608_n185510# 0.02fF
C2786 a_226646_n140786# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.25fF
C2787 a_245224_n123369# a_245481_n123343# 0.11fF
C2788 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_5/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y 0.27fF
C2789 a_245056_n123343# a_245649_n123369# 0.02fF
C2790 peak_detector_rst q4B 0.12fF
C2791 input_amplifier_0/diff_fold_casc_ota_0/vbias2 vocm 0.42fF
C2792 dac_8bit_0/amux_2to1_17/SELB dac_8bit_0/amux_2to1_0/B 1.59fF
C2793 vpeak_sampled dac_8bit_1/amux_2to1_0/B 0.38fF
C2794 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs 0.38fF
C2795 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q 0.04fF
C2796 input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/vop1 14.54fF
C2797 a_237956_n127742# a_238872_n127742# 1.33fF
C2798 a_242085_n122249# a_242951_n122281# 0.11fF
C2799 rst_n biquad_gm_c_filter_0/ibiasn4 0.19fF
C2800 a_237498_n127742# a_239330_n127742# 0.24fF
C2801 a_338149_n185269# a_338356_n185269# 0.63fF
C2802 a_338156_n184969# a_338285_n185243# 0.28fF
C2803 a_336116_n185269# a_336116_n185555# 0.07fF
C2804 a_232702_n134960# vcp 0.03fF
C2805 dac_8bit_1/c7m dac_8bit_1/c0m 0.85fF
C2806 dac_8bit_1/c4m dac_8bit_1/c2m 1.04fF
C2807 dac_8bit_1/c5m dac_8bit_1/cdumm 0.43fF
C2808 dac_8bit_1/c6m dac_8bit_1/c1m 2.24fF
C2809 dac_8bit_1/amux_2to1_14/SELB vrefB 2.12fF
C2810 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q 0.08fF
C2811 dac_8bit_0/c0m VDD 2.48fF
C2812 low_freq_pll_0/cs_ring_osc_0/vpbias a_237956_n145742# 0.83fF
C2813 input_amplifier_0/vop1 a_217060_n102324# 19.89fF
C2814 low_freq_pll_0/freq_div_0/vout VDD 0.55fF
C2815 a_221582_n127742# a_222498_n127742# 2.99fF
C2816 dac_8bit_1/latched_comparator_folded_0/vcompm_buf adc_compB 0.20fF
C2817 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs VDD 4.44fF
C2818 a_242720_n114759# a_242380_n114857# 0.12fF
C2819 a_242137_n115125# a_241731_n115151# 0.04fF
C2820 input_amplifier_0/diff_fold_casc_ota_1/M6d input_amplifier_0/diff_fold_casc_ota_1/M13d 0.56fF
C2821 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc 0.12fF
C2822 peak_detector_0/vpeak vpeak 16.10fF
C2823 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d a_275374_n180872# 0.79fF
C2824 sample VDD 81.17fF
C2825 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc 0.15fF
C2826 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc 0.08fF
C2827 input_amplifier_0/diff_fold_casc_ota_1/M1d vampm 14.05fF
C2828 a_242783_n122255# a_242909_n121877# 0.04fF
C2829 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d 6.93fF
C2830 a_338285_n185409# VDD 0.23fF
C2831 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d 13.66fF
C2832 a_223872_n145742# VDD 0.09fF
C2833 dac_8bit_1/amux_2to1_17/SELB q7B 2.36fF
C2834 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp 0.08fF
C2835 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d 0.75fF
C2836 a_242951_n121443# a_243382_n121389# 0.31fF
C2837 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d 1.74fF
C2838 adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp 0.28fF
C2839 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/vom1 5.46fF
C2840 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_241328_n135628# 0.03fF
C2841 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 12.94fF
C2842 sample dac_8bit_1/amux_2to1_3/SELB 2.36fF
C2843 a_236582_n145742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/csinvp 0.08fF
C2844 a_237956_n145742# a_238414_n145742# 0.02fF
C2845 biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail2 biquad_gm_c_filter_0/gm_c_stage_3/vbiasp 0.90fF
C2846 dac_8bit_0/amux_2to1_1/SELB dac_8bit_0/c6m 1.59fF
C2847 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y a_242951_n123369# 0.17fF
C2848 input_amplifier_0/diff_fold_casc_ota_0/M13d input_amplifier_0/diff_fold_casc_ota_0/vcascnm 0.12fF
C2849 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 2.21fF
C2850 a_244783_n121711# a_245649_n121443# 0.11fF
C2851 a_245224_n121599# a_245056_n121345# 0.59fF
C2852 gain_ctrl_0 VDD 0.39fF
C2853 input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc vocm 1.53fF
C2854 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d 1.51fF
C2855 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d 1.84fF
C2856 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y 0.42fF
C2857 vocm_filt biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail1 2.22fF
C2858 a_241919_n120623# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y 0.35fF
C2859 vocm_filt diff_to_se_converter_0/vim 5.88fF
C2860 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout VDD 9.13fF
C2861 input_amplifier_0/vom1 vocm 5.54fF
C2862 a_337592_n185269# VDD 0.45fF
C2863 a_242783_n122433# a_242085_n123337# 0.01fF
C2864 a_242358_n122433# a_242358_n123343# 0.05fF
C2865 a_242951_n122531# VDD 0.45fF
C2866 biquad_gm_c_filter_0/gm_c_stage_2/vbiasp vfiltp 0.10fF
C2867 input_amplifier_0/diff_fold_casc_ota_0/vfoldp input_amplifier_0/vop1 0.28fF
C2868 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout a_238464_n119618# 0.03fF
C2869 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 0.71fF
C2870 input_amplifier_0/ibiasn2 rst_n 0.19fF
C2871 q1B vrefB 0.88fF
C2872 sample dac_8bit_1/amux_2to1_5/B 2.66fF
C2873 a_242867_n120257# VDD 0.02fF
C2874 a_244617_n122249# VDD 0.78fF
C2875 input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc input_amplifier_0/vip2 0.22fF
C2876 diff_to_se_converter_0/vim diff_to_se_converter_0/rst 0.80fF
C2877 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm 16.88fF
C2878 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 vocm 2.22fF
C2879 dac_8bit_0/amux_2to1_8/SELB dac_8bit_0/amux_2to1_9/Y 1.51fF
C2880 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_246080_n122477# 0.37fF
C2881 a_241919_n122799# a_242273_n122799# 0.21fF
C2882 a_236582_n145742# VDD 0.73fF
C2883 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y a_244617_n121161# 0.04fF
C2884 input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc 0.86fF
C2885 a_336955_n185409# adc_clk 0.02fF
C2886 input_amplifier_0/diff_fold_casc_ota_1/vbias2 vampm 5.46fF
C2887 dac_8bit_1/latched_comparator_folded_0/vlatchp dac_8bit_1/latched_comparator_folded_0/vcompp 0.36fF
C2888 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp vpeak 9.44fF
C2889 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d 0.70fF
C2890 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp 0.08fF
C2891 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d 1.26fF
C2892 a_338356_n185269# a_338532_n184877# 0.04fF
C2893 a_338149_n185269# a_338703_n185243# 0.21fF
C2894 biquad_gm_c_filter_0/ibiasn1 rst_n 0.18fF
C2895 low_freq_pll_0/pfd_cp_lpf_0/vRSTN a_242575_n114888# 0.30fF
C2896 a_226954_n122869# a_227412_n122869# 0.02fF
C2897 peak_detector_0/verr peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn 3.39fF
C2898 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 58.37fF
C2899 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm a_230446_n180872# 10.16fF
C2900 q3A q0A 0.10fF
C2901 input_amplifier_0/txgate_5/txb vincm 0.36fF
C2902 q2B vrefB 0.88fF
C2903 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q a_241919_n121711# 0.51fF
C2904 a_245481_n121345# a_245607_n121711# 0.04fF
C2905 a_239883_n115151# VDD 0.37fF
C2906 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 0.97fF
C2907 input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 0.45fF
C2908 a_336116_n185269# a_336359_n184877# 0.05fF
C2909 a_242453_n123343# VDD 0.02fF
C2910 q4B q0B 0.10fF
C2911 a_229244_n119618# vcp 0.03fF
C2912 dac_8bit_0/amux_2to1_6/SELB vcp_sampled 2.07fF
C2913 a_243382_n120301# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_0/A 0.25fF
C2914 biquad_gm_c_filter_0/ibiasn2 biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail1 3.69fF
C2915 diff_to_se_converter_0/ibiasn vpeak_sampled 0.44fF
C2916 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/csinvp a_225730_n140786# 0.08fF
C2917 vocm_filt biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail1 0.32fF
C2918 a_245056_n122433# a_245182_n122799# 0.02fF
C2919 peak_detector_rst q3B 0.12fF
C2920 a_238770_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.03fF
C2921 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d 5.21fF
C2922 a_243138_n114759# VDD 0.60fF
C2923 vrefA dac_8bit_0/amux_2to1_0/B 2.44fF
C2924 vcp a_238770_n132168# 0.03fF
C2925 a_244617_n123337# a_245224_n123369# 0.37fF
C2926 a_338285_n185409# a_338703_n185409# 0.04fF
C2927 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y a_244783_n123337# 0.61fF
C2928 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q low_freq_pll_0/freq_div_0/vout 0.03fF
C2929 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn vfiltm 0.12fF
C2930 input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc input_amplifier_0/vop1 0.96fF
C2931 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d 21.43fF
C2932 a_243382_n120301# a_243382_n121167# 0.04fF
C2933 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp 9.20fF
C2934 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VDD 2.04fF
C2935 a_337864_n185555# a_338156_n185665# 0.44fF
C2936 a_337592_n185460# a_338356_n185510# 0.02fF
C2937 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_227397_n130007# 0.03fF
C2938 sample dac_8bit_1/c3m 2.36fF
C2939 dac_8bit_1/amux_2to1_13/SELB vrefB 2.12fF
C2940 a_222040_n145742# a_222956_n145742# 2.26fF
C2941 a_221582_n145742# a_223414_n145742# 0.65fF
C2942 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror 2.23fF
C2943 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm 4.75fF
C2944 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp a_356329_n113250# 10.36fF
C2945 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 1.13fF
C2946 a_243312_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs 0.03fF
C2947 vampm gain_ctrl_1 0.52fF
C2948 a_242783_n121167# a_243382_n121167# 0.02fF
C2949 low_freq_pll_0/cs_ring_osc_0/vpbias a_228478_n140786# 0.77fF
C2950 a_242951_n121193# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_1/A 0.04fF
C2951 dac_8bit_1/c7m dac_8bit_1/amux_2to1_0/B 2.37fF
C2952 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp 3.66fF
C2953 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror 0.69fF
C2954 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d 7.88fF
C2955 a_243138_n114759# vcomp 0.01fF
C2956 low_freq_pll_0/pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/Q_N low_freq_pll_0/pfd_cp_lpf_0/vQAb 0.08fF
C2957 vpeak_sampled vbiasp 9.07fF
C2958 dac_8bit_0/vcom_buf dac_8bit_0/latched_comparator_folded_0/vlatchm 0.05fF
C2959 biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail1 biquad_gm_c_filter_0/ibiasn4 0.07fF
C2960 dac_8bit_0/amux_2to1_7/SELB sample 2.36fF
C2961 a_335844_n185269# VDD 0.45fF
C2962 vintp biquad_gm_c_filter_0/gm_c_stage_3/vcmcn 0.11fF
C2963 VDD dac_8bit_1/amux_2to1_7/B 4.57fF
C2964 biquad_gm_c_filter_0/ibiasn2 low_freq_pll_0/ibiasn 0.98fF
C2965 biquad_gm_c_filter_0/ibiasn3 biquad_gm_c_filter_0/ibiasn4 0.62fF
C2966 sample_and_hold_1/vholdm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp 1.42fF
C2967 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d vpeak 0.73fF
C2968 q7B vrefB 0.88fF
C2969 vcp_sampled dac_8bit_0/c4m 1.94fF
C2970 a_239251_n114759# a_238793_n115125# 0.12fF
C2971 q7A q6A 11.40fF
C2972 a_242358_n121167# a_242453_n121167# 0.04fF
C2973 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/M13d 1.61fF
C2974 a_241646_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias 0.63fF
C2975 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y a_242951_n121443# 0.17fF
C2976 a_241919_n121711# a_242783_n121345# 0.09fF
C2977 vintm biquad_gm_c_filter_0/gm_c_stage_2/vbiasp 0.34fF
C2978 vlowB dac_8bit_1/amux_2to1_2/B 1.86fF
C2979 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_244783_n122249# 0.03fF
C2980 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp 6.59fF
C2981 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d 5.99fF
C2982 a_336401_n185269# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.19fF
C2983 a_238793_n115125# low_freq_pll_0/pfd_cp_lpf_0/vRSTN 0.33fF
C2984 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/B pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/Q_N 0.13fF
C2985 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin VDD 4.91fF
C2986 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_225412_n135628# 0.03fF
C2987 adc_clk a_336401_n185569# 0.41fF
C2988 a_230412_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.03fF
C2989 dac_8bit_0/ibiasn vlowA 0.54fF
C2990 dac_8bit_0/ibiasp vlowA 17.58fF
C2991 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d 1.26fF
C2992 vocm_filt biquad_gm_c_filter_0/gm_c_stage_1/vcmcn 2.07fF
C2993 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp 0.08fF
C2994 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_10/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/A 0.35fF
C2995 low_freq_pll_0/pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/Q_N low_freq_pll_0/pfd_cp_lpf_0/vQB 0.13fF
C2996 vcp low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/csinvn 0.08fF
C2997 biquad_gm_c_filter_0/gm_c_stage_2/vbiasp biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail2 0.90fF
C2998 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn1 biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail1 0.58fF
C2999 a_244783_n123337# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.03fF
C3000 a_242085_n122799# a_241919_n123337# 0.02fF
C3001 q1A q0A 2.20fF
C3002 a_242783_n122433# a_242909_n122799# 0.04fF
C3003 a_241919_n122799# a_242085_n123337# 0.02fF
C3004 a_245565_n122255# VDD 0.02fF
C3005 dac_8bit_0/c3m dac_8bit_0/c6m 1.31fF
C3006 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_242243_n138121# 0.03fF
C3007 a_227412_n122869# low_freq_pll_0/cs_ring_osc_0/vpbias 0.77fF
C3008 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y 0.29fF
C3009 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d 15.11fF
C3010 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp 7.95fF
C3011 a_242396_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs 0.03fF
C3012 dac_8bit_0/c0m dac_8bit_0/ibiasn 0.19fF
C3013 low_freq_pll_0/cs_ring_osc_0/vosc a_221480_n131500# 0.03fF
C3014 a_227104_n140786# VDD 0.69fF
C3015 dac_8bit_0/c0m dac_8bit_0/ibiasp 9.64fF
C3016 a_236633_n122049# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout 0.03fF
C3017 input_amplifier_0/txgate_7/txb VDD 3.08fF
C3018 peak_detector_rst q1B 0.12fF
C3019 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d 10.82fF
C3020 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d 0.82fF
C3021 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm 1.74fF
C3022 dac_8bit_0/ibiasn sample 0.19fF
C3023 low_freq_pll_0/pfd_cp_lpf_0/VQBb a_240447_n115125# 0.04fF
C3024 biquad_gm_c_filter_0/ibiasn3 input_amplifier_0/ibiasn2 0.20fF
C3025 a_336955_n185409# a_336608_n185510# 0.11fF
C3026 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_2/Q a_336401_n185569# 0.02fF
C3027 sample dac_8bit_0/ibiasp 0.18fF
C3028 peak_detector_0/vpeak peak_detector_rst 0.59fF
C3029 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD 19.81fF
C3030 input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/M13d 3.61fF
C3031 VDD dac_8bit_1/cdumm 2.41fF
C3032 vintp biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail1 2.83fF
C3033 vintm biquad_gm_c_filter_0/gm_c_stage_2/vcmc 0.54fF
C3034 low_freq_pll_0/cs_ring_osc_0/vosc a_223771_n130007# 0.03fF
C3035 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d a_230446_n180872# 0.79fF
C3036 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp 5.37fF
C3037 peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 0.04fF
C3038 q2A q0A 0.10fF
C3039 a_242273_n121167# a_242273_n121711# 0.02fF
C3040 dac_8bit_1/amux_2to1_10/SELB vrefB 2.12fF
C3041 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 8.42fF
C3042 a_242273_n121711# VDD 0.15fF
C3043 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm 4.75fF
C3044 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror 2.23fF
C3045 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 21.43fF
C3046 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn 9.20fF
C3047 q3B q0B 0.10fF
C3048 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/A VDD 0.62fF
C3049 vocm_filt biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail1 2.22fF
C3050 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d 1.51fF
C3051 comparator_0/ibiasn VDD 8.06fF
C3052 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d 1.84fF
C3053 dac_8bit_0/latched_comparator_folded_0/vcompmb dac_8bit_0/latched_comparator_folded_0/vcompm 0.23fF
C3054 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_0/A 0.27fF
C3055 a_338149_n185569# adc_clk 0.66fF
C3056 peak_detector_rst q2B 0.12fF
C3057 dac_8bit_1/latched_comparator_folded_0/vlatchp dac_8bit_1/latched_comparator_folded_0/vcompm 1.33fF
C3058 a_242085_n122249# a_241919_n122799# 0.09fF
C3059 biquad_gm_c_filter_0/ibiasn3 biquad_gm_c_filter_0/ibiasn1 0.35fF
C3060 dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d 5.10fF
C3061 dac_8bit_0/amux_2to1_5/B q2A 1.99fF
C3062 VDD input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc 15.85fF
C3063 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q a_244617_n122799# 0.49fF
C3064 diff_to_se_converter_0/txgate_0/txb VDD 3.10fF
C3065 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_8/A VDD 0.48fF
C3066 a_337592_n185269# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.02fF
C3067 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A a_338149_n185269# 0.02fF
C3068 vpeak_sampled vcp 1.58fF
C3069 dac_8bit_1/amux_2to1_12/SELB vrefB 2.12fF
C3070 a_242783_n122433# a_242867_n122433# 0.05fF
C3071 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VDD 11.66fF
C3072 q4A dac_8bit_0/amux_2to1_3/B 1.99fF
C3073 a_242783_n122255# VDD 0.22fF
C3074 a_226038_n122869# VDD 1.55fF
C3075 dac_8bit_1/amux_2to1_11/SELB dac_8bit_1/amux_2to1_6/B 1.59fF
C3076 dac_8bit_1/vcom_buf dac_8bit_1/latched_comparator_folded_0/vlatchp 3.59fF
C3077 comparator_0/ibiasn vcomp 0.17fF
C3078 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VDD 1.46fF
C3079 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 a_162668_n147576# 8.05fF
C3080 comparator_0/vcompm vfiltp 2.90fF
C3081 a_242951_n120355# VDD 0.45fF
C3082 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 28.69fF
C3083 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn 16.73fF
C3084 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q a_242085_n122799# 0.09fF
C3085 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y a_242783_n121167# 0.14fF
C3086 a_244783_n122249# a_245481_n122255# 0.44fF
C3087 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VDD 2.04fF
C3088 a_245224_n122281# a_245649_n122281# 0.04fF
C3089 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD 6.84fF
C3090 dac_8bit_1/ibiasn dac_8bit_0/c5m 0.20fF
C3091 a_245481_n121167# VDD 0.22fF
C3092 q7A q5A 0.10fF
C3093 a_242526_n121599# a_242273_n121711# 0.04fF
C3094 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn 2.79fF
C3095 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 6.00fF
C3096 vintp biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail1 2.83fF
C3097 a_224330_n127742# VDD 0.06fF
C3098 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin 1.49fF
C3099 a_336537_n185243# VDD 0.23fF
C3100 a_242358_n121167# a_242273_n121167# 0.11fF
C3101 a_242358_n121167# VDD 0.36fF
C3102 vpeak_sampled dac_8bit_1/amux_2to1_0/SELB 2.07fF
C3103 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d 0.73fF
C3104 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm 0.08fF
C3105 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm 20.84fF
C3106 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 1.35fF
C3107 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VDD 12.54fF
C3108 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_236939_n148007# 0.03fF
C3109 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d 0.70fF
C3110 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm 0.51fF
C3111 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d a_356329_n164260# 1.44fF
C3112 peak_detector_rst q7B 16.71fF
C3113 low_freq_pll_0/freq_div_0/vout a_238627_n115125# 0.49fF
C3114 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d 0.12fF
C3115 dac_8bit_1/latched_comparator_folded_0/vlatchm adc_clk 0.68fF
C3116 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d 9.86fF
C3117 vocm input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 2.22fF
C3118 VDD a_246080_n122477# 0.37fF
C3119 a_336401_n185569# a_336608_n185510# 0.63fF
C3120 a_336116_n185555# a_336537_n185409# 0.11fF
C3121 a_245649_n123369# a_245481_n123343# 0.67fF
C3122 vse vfiltm 0.20fF
C3123 low_freq_pll_0/pfd_cp_lpf_0/vswitchh low_freq_pll_0/pfd_cp_lpf_0/vQA 0.18fF
C3124 dac_8bit_1/amux_2to1_17/SELB vrefB 2.12fF
C3125 dac_8bit_1/amux_2to1_6/B vrefB 2.44fF
C3126 a_238414_n127742# a_239330_n127742# 0.79fF
C3127 a_338149_n185269# pulse_generator_0/sky130_fd_sc_hd__inv_1_0/Y 0.51fF
C3128 a_336116_n185269# a_336408_n185665# 0.01fF
C3129 a_338356_n185269# a_338285_n185243# 0.59fF
C3130 a_336408_n184969# a_336401_n185569# 0.02fF
C3131 VDD input_amplifier_0/vim1 0.62fF
C3132 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD 19.81fF
C3133 dac_8bit_1/c3m dac_8bit_1/cdumm 0.07fF
C3134 q1B q0B 2.20fF
C3135 low_freq_pll_0/cs_ring_osc_0/vpbias a_238872_n145742# 0.92fF
C3136 a_221582_n127742# a_223414_n127742# 0.65fF
C3137 a_222040_n127742# a_222956_n127742# 2.26fF
C3138 a_242377_n115125# a_242102_n114873# 0.04fF
C3139 a_242720_n114759# a_242575_n114888# 0.21fF
C3140 a_243138_n114759# a_242419_n114983# 0.23fF
C3141 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn a_356329_n164260# 0.11fF
C3142 vcp a_221480_n150168# 0.03fF
C3143 a_244617_n122249# a_244971_n122255# 0.21fF
C3144 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d VDD 11.46fF
C3145 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d 0.16fF
C3146 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/csinvp VDD 0.48fF
C3147 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn 32.00fF
C3148 vhpf vincm 5.53fF
C3149 vintp biquad_gm_c_filter_0/gm_c_stage_1/vcmcn 1.45fF
C3150 input_amplifier_0/vip1 input_amplifier_0/ibiasn1 0.23fF
C3151 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_242244_n135628# 0.03fF
C3152 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror adc_vcaparrayB 1.41fF
C3153 dac_8bit_1/amux_2to1_9/SELB vrefB 2.12fF
C3154 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD 25.41fF
C3155 sample dac_8bit_1/amux_2to1_5/SELB 2.36fF
C3156 a_237956_n145742# a_239330_n145742# 0.01fF
C3157 a_237498_n145742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/csinvp 0.09fF
C3158 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp 3.66fF
C3159 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d 7.88fF
C3160 a_238414_n145742# a_238872_n145742# 0.01fF
C3161 q7A dac_8bit_1/ibiasn 0.20fF
C3162 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VDD 25.41fF
C3163 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_236582_n145742# 0.90fF
C3164 q2B q0B 0.10fF
C3165 a_245056_n121345# a_245649_n121443# 0.02fF
C3166 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_244971_n121711# 0.02fF
C3167 a_245224_n121599# a_245481_n121345# 0.11fF
C3168 a_245224_n123369# VDD 0.23fF
C3169 vcp a_221480_n132168# 0.03fF
C3170 vcp_sampled dac_8bit_0/amux_2to1_4/SELB 2.07fF
C3171 low_freq_pll_0/ibiasn biquad_gm_c_filter_0/ibiasn4 7.72fF
C3172 biquad_gm_c_filter_0/ibiasn2 vocm_filt 0.15fF
C3173 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_227397_n148007# 0.03fF
C3174 a_338156_n184969# VDD 0.45fF
C3175 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y 0.03fF
C3176 a_242951_n122531# a_242951_n123369# 0.09fF
C3177 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/Q_N a_335844_n185460# 0.02fF
C3178 a_244783_n122799# a_245056_n122433# 0.38fF
C3179 a_337592_n185460# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/D 0.02fF
C3180 a_243382_n122477# VDD 0.37fF
C3181 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout low_freq_pll_0/cs_ring_osc_0/vosc 1.76fF
C3182 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_242273_n121167# 0.02fF
C3183 sample dac_8bit_1/c4m 2.36fF
C3184 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q VDD 0.38fF
C3185 diff_to_se_converter_0/vip diff_to_se_converter_0/txgate_0/txb 0.36fF
C3186 dac_8bit_1/amux_2to1_11/SELB vrefB 2.12fF
C3187 sample_and_hold_1/vholdm VDD 0.76fF
C3188 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y 0.13fF
C3189 pulse_generator_0/sky130_fd_sc_hd__inv_1_1/A pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/B 0.30fF
C3190 a_238627_n115125# a_239883_n115151# 0.12fF
C3191 a_238793_n115125# a_239143_n115125# 0.49fF
C3192 a_242273_n122255# a_242273_n122799# 0.02fF
C3193 comparator_0/vcompp VDD 9.64fF
C3194 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VDD 2.04fF
C3195 dac_8bit_0/c7m dac_8bit_0/c5m 1.37fF
C3196 a_237498_n145742# VDD 0.40fF
C3197 dac_8bit_0/amux_2to1_7/B vcp_sampled 0.38fF
C3198 dac_8bit_0/amux_2to1_9/Y vlowA 1.90fF
C3199 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin VDD 4.83fF
C3200 a_244783_n121711# VDD 0.43fF
C3201 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_2/Q adc_clk 0.07fF
C3202 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d 2.72fF
C3203 a_244617_n122249# a_244783_n122249# 2.23fF
C3204 q7A q4A 0.10fF
C3205 a_245869_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.03fF
C3206 a_244617_n121161# VDD 0.78fF
C3207 dac_8bit_0/amux_2to1_5/B dac_8bit_0/amux_2to1_12/SELB 1.59fF
C3208 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror 5.68fF
C3209 a_226954_n122869# a_228328_n122869# 0.01fF
C3210 a_227412_n122869# a_227870_n122869# 0.01fF
C3211 a_338285_n185243# a_338703_n185243# 0.04fF
C3212 diff_to_se_converter_0/txgate_1/txb VDD 3.26fF
C3213 comparator_0/ibiasn rst_n 0.51fF
C3214 q0B q7B 0.10fF
C3215 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 58.37fF
C3216 comparator_0/vcompm comparator_0/vo1 1.42fF
C3217 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror 17.44fF
C3218 low_freq_pll_0/pfd_cp_lpf_0/vswitchl low_freq_pll_0/ibiasn 0.26fF
C3219 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm 2.41fF
C3220 input_amplifier_0/rst input_amplifier_0/vip1 0.87fF
C3221 dac_8bit_1/ibiasp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d 0.01fF
C3222 a_236582_n145742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs 0.82fF
C3223 a_240447_n115125# VDD 0.29fF
C3224 dac_8bit_0/amux_2to1_14/SELB dac_8bit_0/amux_2to1_3/B 1.59fF
C3225 dac_8bit_0/c0m dac_8bit_0/amux_2to1_9/Y 1.72fF
C3226 diff_to_se_converter_0/txgate_0/txb rst_n 0.18fF
C3227 a_230160_n119618# vcp 0.03fF
C3228 peak_detector_0/ibiasn1 VDD 3.49fF
C3229 dac_8bit_1/amux_2to1_0/SELB dac_8bit_1/c7m 1.59fF
C3230 dac_8bit_0/amux_2to1_9/Y sample 2.66fF
C3231 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/csinvp a_226646_n140786# 0.09fF
C3232 a_226022_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.03fF
C3233 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 12.94fF
C3234 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 3.47fF
C3235 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm 16.88fF
C3236 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_0/vhold 0.86fF
C3237 peak_detector_0/ibiasn2 vse 5.49fF
C3238 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y 0.93fF
C3239 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_224953_n138121# 0.03fF
C3240 input_amplifier_0/ibiasn2 low_freq_pll_0/ibiasn 0.23fF
C3241 a_221481_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin 0.03fF
C3242 VDD dac_8bit_1/amux_2to1_7/SELB 1.15fF
C3243 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y a_245056_n123343# 0.16fF
C3244 a_244617_n123337# a_245649_n123369# 0.11fF
C3245 vrefA q6A 0.88fF
C3246 a_229953_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.03fF
C3247 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VDD 7.64fF
C3248 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn2 vampm 0.10fF
C3249 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_0/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_1/A 0.04fF
C3250 a_338149_n185569# a_338356_n185510# 0.63fF
C3251 a_337864_n185555# a_338285_n185409# 0.11fF
C3252 vse a_162668_n147576# 19.89fF
C3253 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_228313_n130007# 0.03fF
C3254 input_amplifier_0/venm1 input_amplifier_0/vop1 0.78fF
C3255 a_222040_n145742# a_223872_n145742# 0.43fF
C3256 a_221582_n145742# a_224330_n145742# 0.14fF
C3257 a_222498_n145742# a_223414_n145742# 1.92fF
C3258 a_236480_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin 0.03fF
C3259 a_241919_n122249# VDD 0.79fF
C3260 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_0/A 0.35fF
C3261 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_226480_n149500# 0.03fF
C3262 a_243382_n121167# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_1/A 0.25fF
C3263 dac_8bit_0/cdumm vcp_sampled 1.94fF
C3264 biquad_gm_c_filter_0/gm_c_stage_1/vcmc VDD 2.70fF
C3265 vlowA dac_8bit_0/latched_comparator_folded_0/vlatchp 0.16fF
C3266 a_246080_n122255# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/A 0.05fF
C3267 dac_8bit_1/latched_comparator_folded_0/vlatchp VDD 4.86fF
C3268 a_245481_n121167# a_245607_n120789# 0.04fF
C3269 a_338107_n184877# VDD 0.02fF
C3270 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 a_230446_n180872# 8.26fF
C3271 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 44.84fF
C3272 biquad_gm_c_filter_0/ibiasn2 biquad_gm_c_filter_0/ibiasn4 33.88fF
C3273 biquad_gm_c_filter_0/ibiasn1 low_freq_pll_0/ibiasn 3.56fF
C3274 a_239251_n114759# low_freq_pll_0/pfd_cp_lpf_0/vRSTN 0.06fF
C3275 dac_8bit_0/amux_2to1_9/SELB q0A 2.36fF
C3276 a_242562_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias 0.76fF
C3277 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y a_243382_n121389# 0.11fF
C3278 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d VDD 9.36fF
C3279 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp adc_vcaparrayA 28.95fF
C3280 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 3.45fF
C3281 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm 23.84fF
C3282 adc_vcaparrayA dac_8bit_0/c5m 214.58fF
C3283 vlowB dac_8bit_1/amux_2to1_4/B 1.86fF
C3284 VDD input_amplifier_0/txgate_4/txb 3.10fF
C3285 dac_8bit_1/amux_2to1_6/SELB dac_8bit_1/amux_2to1_6/B 1.51fF
C3286 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/vip 0.08fF
C3287 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q low_freq_pll_0/freq_div_0/vin 0.04fF
C3288 dac_8bit_0/c1m dac_8bit_0/c0m 12.39fF
C3289 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_226328_n135628# 0.03fF
C3290 a_231328_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.03fF
C3291 a_244617_n121711# a_245224_n121599# 0.37fF
C3292 rst_n input_amplifier_0/vim1 0.16fF
C3293 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y a_244783_n121711# 0.61fF
C3294 a_241480_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs 0.03fF
C3295 vcp_sampled dac_8bit_1/ibiasp 0.17fF
C3296 dac_8bit_0/c1m sample 2.36fF
C3297 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm 4.75fF
C3298 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 8.42fF
C3299 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_241481_n130007# 0.03fF
C3300 a_241919_n122799# a_242358_n123343# 0.01fF
C3301 a_242358_n122433# a_241919_n123337# 0.01fF
C3302 adc_clk a_336408_n184969# 0.08fF
C3303 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q a_244783_n121711# 0.03fF
C3304 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y VDD 0.91fF
C3305 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d VDD 7.37fF
C3306 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_1/vcom_buf 0.86fF
C3307 dac_8bit_1/adc_run VDD 3.10fF
C3308 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.38fF
C3309 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y a_242085_n122249# 0.61fF
C3310 vcp a_227412_n119618# 0.03fF
C3311 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 5.68fF
C3312 q1B dac_8bit_1/amux_2to1_7/B 1.99fF
C3313 a_228328_n122869# low_freq_pll_0/cs_ring_osc_0/vpbias 0.85fF
C3314 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q a_244617_n121161# 0.51fF
C3315 dac_8bit_0/latched_comparator_folded_0/vcompp adc_clk 0.37fF
C3316 VDD input_amplifier_0/diff_fold_casc_ota_0/vbias1 23.91fF
C3317 a_242085_n122799# a_242358_n122433# 0.38fF
C3318 a_243312_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs 0.03fF
C3319 dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d 9.79fF
C3320 low_freq_pll_0/cs_ring_osc_0/vosc a_222396_n131500# 0.03fF
C3321 a_228020_n140786# VDD 0.09fF
C3322 a_237549_n122049# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout 0.03fF
C3323 biquad_gm_c_filter_0/gm_c_stage_1/vbiasp VDD 3.04fF
C3324 q7A q3A 0.10fF
C3325 biquad_gm_c_filter_0/ibiasn2 input_amplifier_0/ibiasn2 0.19fF
C3326 a_336955_n185409# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/D 0.39fF
C3327 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 28.76fF
C3328 peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 2.30fF
C3329 a_242358_n122255# a_242453_n122255# 0.04fF
C3330 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/Q_N VDD 0.51fF
C3331 a_241188_n140786# VDD 1.55fF
C3332 a_241634_n115151# a_241731_n115151# 0.30fF
C3333 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm adc_vcaparrayA 0.75fF
C3334 vpeak_sampled sample_and_hold_1/vhold 4.86fF
C3335 dac_8bit_0/amux_2to1_2/SELB dac_8bit_0/amux_2to1_2/B 1.51fF
C3336 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_7/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/A 0.35fF
C3337 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 13.36fF
C3338 vcp_sampled VDD 19.27fF
C3339 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/vholdm 5.59fF
C3340 low_freq_pll_0/freq_div_0/vout low_freq_pll_0/ibiasn 0.68fF
C3341 a_338356_n185510# adc_clk 0.11fF
C3342 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/A VDD 0.62fF
C3343 biquad_gm_c_filter_0/ibiasn2 biquad_gm_c_filter_0/ibiasn1 0.48fF
C3344 dac_8bit_0/latched_comparator_folded_0/vcompmb dac_8bit_0/comp_outm 0.03fF
C3345 biquad_gm_c_filter_0/ibiasn3 comparator_0/ibiasn 0.60fF
C3346 vrefA q5A 0.88fF
C3347 a_242085_n122249# a_242273_n122255# 0.26fF
C3348 dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn 14.42fF
C3349 low_freq_pll_0/cs_ring_osc_0/vpbias a_236582_n127742# 0.51fF
C3350 low_freq_pll_0/pfd_cp_lpf_0/vswitchh low_freq_pll_0/pfd_cp_lpf_0/vQAb 1.92fF
C3351 vpeak_sampled dac_8bit_1/amux_2to1_1/B 0.38fF
C3352 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_1/vcom_buf 24.36fF
C3353 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/B pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A 0.43fF
C3354 input_amplifier_0/diff_fold_casc_ota_1/vfoldm VDD 20.43fF
C3355 a_242783_n122433# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q 0.05fF
C3356 dac_8bit_1/c5m dac_8bit_1/c1m 1.12fF
C3357 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_2/A VDD 0.48fF
C3358 dac_8bit_1/c4m dac_8bit_1/cdumm 0.43fF
C3359 dac_8bit_1/c6m dac_8bit_1/c0m 0.85fF
C3360 VDD input_amplifier_0/diff_fold_casc_ota_0/M6d 11.14fF
C3361 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/vbias3 1.29fF
C3362 a_226954_n122869# VDD 0.69fF
C3363 biquad_gm_c_filter_0/gm_c_stage_3/vcmc VDD 2.70fF
C3364 diff_to_se_converter_0/txgate_1/txb rst_n 0.18fF
C3365 dac_8bit_0/c2m dac_8bit_1/ibiasn 2.53fF
C3366 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 16.73fF
C3367 a_243382_n120301# VDD 0.37fF
C3368 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 28.69fF
C3369 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_1/A 0.27fF
C3370 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn1 vfiltp 0.03fF
C3371 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn vocm_filt 2.07fF
C3372 vampp input_amplifier_0/diff_fold_casc_ota_1/vbias3 11.45fF
C3373 a_245056_n122255# a_245481_n122255# 0.03fF
C3374 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/A 1.64fF
C3375 peak_detector_0/ibiasn2 input_amplifier_0/ibiasn1 4.67fF
C3376 vse diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp 21.50fF
C3377 adc_vcaparrayB dac_8bit_1/c7m 854.85fF
C3378 adc_clk a_337497_n185269# 0.13fF
C3379 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_6/A VDD 0.48fF
C3380 vfiltp vfiltm 16.67fF
C3381 vrefA dac_8bit_0/amux_2to1_16/SELB 2.12fF
C3382 a_242358_n121345# a_242453_n121345# 0.04fF
C3383 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 2.79fF
C3384 a_239048_n115125# low_freq_pll_0/freq_div_0/vout 0.01fF
C3385 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y 0.03fF
C3386 peak_detector_0/ibiasn1 rst_n 0.09fF
C3387 a_242783_n121167# VDD 0.22fF
C3388 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn 3.60fF
C3389 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/csinvn low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.09fF
C3390 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_237855_n148007# 0.03fF
C3391 input_amplifier_0/venm2 input_amplifier_0/vim2 1.11fF
C3392 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp 5.37fF
C3393 dac_8bit_1/amux_2to1_9/SELB q0B 2.36fF
C3394 low_freq_pll_0/pfd_cp_lpf_0/VQBb low_freq_pll_0/pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/Q_N 0.08fF
C3395 a_242273_n120623# a_242085_n120623# 0.26fF
C3396 q0A adc_vcaparrayB 1.72fF
C3397 dac_8bit_1/latched_comparator_folded_0/vcompp dac_8bit_1/latched_comparator_folded_0/vcompp_buf 0.02fF
C3398 q7A q1A 0.10fF
C3399 peak_detector_0/ibiasn1 dac_8bit_0/ibiasn 0.01fF
C3400 a_241919_n121161# a_242085_n121161# 2.23fF
C3401 input_amplifier_0/vip2 VDD 3.63fF
C3402 a_336408_n185665# a_336537_n185409# 0.28fF
C3403 a_336401_n185569# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/D 0.59fF
C3404 a_240062_n115125# a_239883_n115151# 0.04fF
C3405 a_239817_n115125# a_239708_n115125# 0.04fF
C3406 a_245649_n123369# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_10/A 0.04fF
C3407 a_245481_n123343# a_246080_n123343# 0.02fF
C3408 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn1 vocm_filt 1.07fF
C3409 input_amplifier_0/diff_fold_casc_ota_1/M13d VDD 1.24fF
C3410 vpeak_sampled dac_8bit_1/c7m 1.94fF
C3411 a_336401_n185269# a_336408_n185665# 0.02fF
C3412 a_336608_n185269# a_336401_n185569# 0.01fF
C3413 a_338285_n185243# pulse_generator_0/sky130_fd_sc_hd__inv_1_0/Y 0.04fF
C3414 sample dac_8bit_1/amux_2to1_6/B 2.66fF
C3415 input_amplifier_0/diff_fold_casc_ota_1/M3d VDD 1.56fF
C3416 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/vcom_buf 15.32fF
C3417 pulse_generator_0/sky130_fd_sc_hd__inv_1_1/A a_335507_n185243# 0.05fF
C3418 a_244783_n121161# a_245056_n121167# 0.38fF
C3419 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn1 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn2 0.17fF
C3420 VDD input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc 5.35fF
C3421 low_freq_pll_0/cs_ring_osc_0/vpbias low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/csinvp 0.31fF
C3422 biquad_gm_c_filter_0/gm_c_stage_3/vbiasp VDD 3.04fF
C3423 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y 0.04fF
C3424 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q a_242085_n121711# 0.03fF
C3425 a_242104_n140786# a_242562_n140786# 0.02fF
C3426 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q a_242085_n122249# 0.08fF
C3427 a_221582_n127742# a_224330_n127742# 0.14fF
C3428 a_222040_n127742# a_223872_n127742# 0.43fF
C3429 a_222498_n127742# a_223414_n127742# 1.92fF
C3430 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm a_356329_n113250# 10.16fF
C3431 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn2 vfiltm 2.12fF
C3432 a_336116_n185269# a_336401_n185269# 0.09fF
C3433 vampp input_amplifier_0/diff_fold_casc_ota_1/vcascnp 7.04fF
C3434 vcp a_222396_n150168# 0.03fF
C3435 q7A q2A 0.10fF
C3436 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/vpeak 1.41fF
C3437 vocm_filt biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail1 0.32fF
C3438 sample_and_hold_1/vhold sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn 2.30fF
C3439 vfiltp biquad_gm_c_filter_0/gm_c_stage_2/vtail_diff 2.64fF
C3440 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 28.76fF
C3441 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp 1.94fF
C3442 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm 23.84fF
C3443 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 3.45fF
C3444 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/vhold 28.95fF
C3445 low_freq_pll_0/pfd_cp_lpf_0/vQA low_freq_pll_0/pfd_cp_lpf_0/vRSTN 1.34fF
C3446 vintp vocm_filt 3.46fF
C3447 a_238414_n145742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/csinvp 0.10fF
C3448 a_238872_n145742# a_239330_n145742# 0.02fF
C3449 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/vim 0.08fF
C3450 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp 6.59fF
C3451 dac_8bit_1/amux_2to1_10/SELB dac_8bit_1/amux_2to1_7/B 1.59fF
C3452 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_237498_n145742# 0.25fF
C3453 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d 0.73fF
C3454 dac_8bit_0/latched_comparator_folded_0/vcompm adc_clk 0.51fF
C3455 biquad_gm_c_filter_0/gm_c_stage_0/vbiasp biquad_gm_c_filter_0/gm_c_stage_0/vcmcn1 0.19fF
C3456 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm 2.00fF
C3457 dac_8bit_0/amux_2to1_7/SELB vcp_sampled 2.07fF
C3458 low_freq_pll_0/cs_ring_osc_0/vpbias VDD 18.73fF
C3459 a_245649_n121443# a_245481_n121345# 0.67fF
C3460 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d 1.51fF
C3461 dac_8bit_1/latched_comparator_folded_0/vcompmb dac_8bit_1/latched_comparator_folded_0/vcompm_buf 0.31fF
C3462 a_245649_n123369# VDD 0.45fF
C3463 vintm biquad_gm_c_filter_0/gm_c_stage_3/vcmcn1 0.12fF
C3464 vcp a_222396_n132168# 0.03fF
C3465 vrefA q4A 0.88fF
C3466 vrefA dac_8bit_0/amux_2to1_1/B 2.44fF
C3467 biquad_gm_c_filter_0/ibiasn1 vocm_filt 0.31fF
C3468 input_amplifier_0/diff_fold_casc_ota_1/vbias3 input_amplifier_0/diff_fold_casc_ota_1/vbias4 36.54fF
C3469 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_228313_n148007# 0.03fF
C3470 a_244783_n121161# low_freq_pll_0/freq_div_0/vout 0.01fF
C3471 a_338356_n185269# VDD 0.36fF
C3472 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm vse 5.69fF
C3473 a_245224_n122687# a_245649_n122531# 0.04fF
C3474 a_244783_n122799# a_245481_n122433# 0.44fF
C3475 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d 3.28fF
C3476 a_239251_n114759# a_239143_n115125# 0.21fF
C3477 low_freq_pll_0/pfd_cp_lpf_0/vQAb vcp 0.08fF
C3478 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 3.02fF
C3479 vintm vfiltm 3.38fF
C3480 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/vcom_buf 22.36fF
C3481 q0B vrefB 0.88fF
C3482 dac_8bit_0/c2m dac_8bit_0/c7m 2.04fF
C3483 input_amplifier_0/ibiasn2 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 3.91fF
C3484 sample dac_8bit_1/c2m 2.36fF
C3485 a_239361_n114883# a_239883_n115151# 0.03fF
C3486 a_238793_n115125# a_239708_n115125# 0.29fF
C3487 low_freq_pll_0/pfd_cp_lpf_0/vRSTN a_239143_n115125# 0.30fF
C3488 a_241919_n122799# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q 0.03fF
C3489 sample vpeak 0.75fF
C3490 dac_8bit_0/amux_2to1_8/SELB dac_8bit_0/c0m 1.59fF
C3491 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD 19.81fF
C3492 adc_compB adc_clk 0.05fF
C3493 a_238414_n145742# VDD 0.14fF
C3494 a_245056_n121345# VDD 0.36fF
C3495 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 21.43fF
C3496 input_amplifier_0/vip1 input_amplifier_0/diff_fold_casc_ota_0/vfoldp 9.23fF
C3497 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y VDD 0.96fF
C3498 dac_8bit_0/amux_2to1_8/SELB sample 2.36fF
C3499 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 33.98fF
C3500 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d VDD 1.27fF
C3501 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_0/vhold 0.75fF
C3502 input_amplifier_0/rst input_amplifier_0/diff_fold_casc_ota_0/vfoldm 0.11fF
C3503 a_242720_n114759# low_freq_pll_0/pfd_cp_lpf_0/vRSTN 0.06fF
C3504 peak_detector_0/ibiasn2 vfiltp 0.18fF
C3505 VDD dac_8bit_1/amux_2to1_9/Y 4.57fF
C3506 a_244617_n122249# a_245056_n122255# 0.63fF
C3507 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y a_245224_n122281# 0.15fF
C3508 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs VDD 4.44fF
C3509 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror 17.44fF
C3510 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/vpeak 0.08fF
C3511 vrefA dac_8bit_0/amux_2to1_15/SELB 2.12fF
C3512 a_246785_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.03fF
C3513 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm 2.41fF
C3514 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn 2.79fF
C3515 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 6.00fF
C3516 dac_8bit_0/amux_2to1_0/B VDD 4.57fF
C3517 a_227870_n122869# a_228328_n122869# 0.02fF
C3518 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d 0.70fF
C3519 vlowB dac_8bit_1/amux_2to1_3/B 1.86fF
C3520 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 1.65fF
C3521 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror 4.50fF
C3522 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm 0.51fF
C3523 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm 0.08fF
C3524 vincm input_amplifier_0/vip1 7.74fF
C3525 a_245481_n123343# a_245607_n122965# 0.04fF
C3526 diff_to_se_converter_0/vim diff_to_se_converter_0/txgate_1/txb 0.36fF
C3527 a_244783_n121711# a_244783_n122249# 0.06fF
C3528 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm 4.75fF
C3529 a_237498_n145742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs 0.22fF
C3530 a_336608_n185269# a_336784_n184877# 0.04fF
C3531 a_336401_n185269# a_336955_n185243# 0.21fF
C3532 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 33.98fF
C3533 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail1 0.58fF
C3534 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/csinvp a_227562_n140786# 0.10fF
C3535 a_226938_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.03fF
C3536 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d 5.21fF
C3537 input_amplifier_0/diff_fold_casc_ota_1/vbias1 vampp 2.53fF
C3538 input_amplifier_0/diff_fold_casc_ota_1/vbias3 a_163060_n102324# 7.49fF
C3539 input_amplifier_0/ibiasn2 biquad_gm_c_filter_0/ibiasn4 0.20fF
C3540 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc input_amplifier_0/diff_fold_casc_ota_0/M3d 0.64fF
C3541 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vbias2 0.63fF
C3542 biquad_gm_c_filter_0/ibiasn3 peak_detector_0/ibiasn1 0.42fF
C3543 input_amplifier_0/diff_fold_casc_ota_1/vbias4 input_amplifier_0/diff_fold_casc_ota_1/vcascnp 17.91fF
C3544 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_225869_n138121# 0.03fF
C3545 diff_to_se_converter_0/ibiasn vfiltm 0.46fF
C3546 a_222397_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin 0.03fF
C3547 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn vintp 1.30fF
C3548 a_230869_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.03fF
C3549 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y a_245481_n123343# 0.14fF
C3550 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 a_356329_n113250# 8.05fF
C3551 a_244783_n123337# a_244783_n122799# 0.06fF
C3552 pulse_generator_0/sky130_fd_sc_hd__inv_1_1/A VDD 0.90fF
C3553 vintm biquad_gm_c_filter_0/gm_c_stage_2/vtail_diff 0.58fF
C3554 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 1.35fF
C3555 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm 20.84fF
C3556 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn biquad_gm_c_filter_0/gm_c_stage_2/vcmcn2 1.28fF
C3557 a_338156_n185665# a_338285_n185409# 0.28fF
C3558 adc_vcaparrayA dac_8bit_0/vcom_buf 15.10fF
C3559 dac_8bit_0/c3m dac_8bit_0/c5m 0.66fF
C3560 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm 16.73fF
C3561 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.38fF
C3562 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VDD 11.66fF
C3563 a_222956_n145742# a_223872_n145742# 1.33fF
C3564 a_237396_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin 0.03fF
C3565 a_222498_n145742# a_224330_n145742# 0.24fF
C3566 dac_8bit_1/ibiasn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp 0.03fF
C3567 input_amplifier_0/txgate_7/txb input_amplifier_0/vom1 0.36fF
C3568 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VDD 6.84fF
C3569 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_227396_n149500# 0.03fF
C3570 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 13.36fF
C3571 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm 5.03fF
C3572 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d 1.26fF
C3573 input_amplifier_0/venp1 VDD 1.25fF
C3574 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc vocm 1.48fF
C3575 low_freq_pll_0/pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/Q_N a_241634_n115151# 0.14fF
C3576 a_245481_n121167# a_245565_n121167# 0.05fF
C3577 input_amplifier_0/rst input_amplifier_0/diff_fold_casc_ota_0/M3d 0.11fF
C3578 a_338703_n185243# VDD 0.15fF
C3579 comparator_0/ibiasn low_freq_pll_0/ibiasn 9.19fF
C3580 biquad_gm_c_filter_0/ibiasn1 biquad_gm_c_filter_0/ibiasn4 27.03fF
C3581 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm peak_detector_0/verr 5.69fF
C3582 VDD dac_8bit_1/c1m 2.47fF
C3583 dac_8bit_0/c2m adc_vcaparrayA 57.70fF
C3584 a_242951_n122281# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q 0.39fF
C3585 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror 14.22fF
C3586 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_1/vholdm 19.15fF
C3587 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d 1.91fF
C3588 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp 1.03fF
C3589 a_243478_n140786# low_freq_pll_0/cs_ring_osc_0/vpbias 0.77fF
C3590 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d 3.60fF
C3591 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/A 0.10fF
C3592 dac_8bit_1/amux_2to1_1/B dac_8bit_1/amux_2to1_16/SELB 1.59fF
C3593 vintp biquad_gm_c_filter_0/gm_c_stage_2/vcmcn1 0.13fF
C3594 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp 13.60fF
C3595 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d 3.07fF
C3596 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp 0.81fF
C3597 input_amplifier_0/diff_fold_casc_ota_0/vbias3 input_amplifier_0/diff_fold_casc_ota_0/vbias4 36.54fF
C3598 a_337864_n185555# a_338156_n184969# 0.01fF
C3599 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_245481_n122255# 0.05fF
C3600 a_236480_n150168# vcp 0.03fF
C3601 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d 3.28fF
C3602 dac_8bit_1/vcom_buf vlowB 1.79fF
C3603 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_227244_n135628# 0.03fF
C3604 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn2 biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail2 0.58fF
C3605 adc_clk pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/D 0.34fF
C3606 a_232244_n135628# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.03fF
C3607 a_225730_n140786# a_226646_n140786# 2.99fF
C3608 adc_compA VDD 2.44fF
C3609 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y a_245056_n121345# 0.16fF
C3610 a_244617_n121711# a_245649_n121443# 0.11fF
C3611 input_amplifier_0/diff_fold_casc_ota_1/M6d vampp 0.31fF
C3612 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/A 0.10fF
C3613 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/vom1 7.09fF
C3614 input_amplifier_0/diff_fold_casc_ota_1/vcascnp a_163060_n102324# 6.65fF
C3615 vrefA q3A 0.88fF
C3616 peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 0.21fF
C3617 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d 7.95fF
C3618 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp a_189446_n180872# 10.36fF
C3619 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 1.13fF
C3620 low_freq_pll_0/freq_div_0/vin low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y 0.05fF
C3621 vcp sample_and_hold_0/vhold 1.71fF
C3622 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_242397_n130007# 0.03fF
C3623 vintm biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail2 0.32fF
C3624 a_245481_n123343# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.05fF
C3625 low_freq_pll_0/pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/Q_N VDD 0.23fF
C3626 a_244617_n122799# a_244783_n122799# 2.23fF
C3627 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin a_236481_n130007# 0.03fF
C3628 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp 21.50fF
C3629 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_5/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/A 0.35fF
C3630 vcp a_228328_n119618# 0.03fF
C3631 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 1.11fF
C3632 dac_8bit_1/cdumm dac_8bit_1/amux_2to1_6/B 1.72fF
C3633 a_335844_n185269# a_336116_n185269# 0.67fF
C3634 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn biquad_gm_c_filter_0/gm_c_stage_3/vcmc 0.05fF
C3635 a_242085_n122799# a_242783_n122433# 0.44fF
C3636 a_242526_n122687# a_242951_n122531# 0.04fF
C3637 dac_8bit_0/latched_comparator_folded_0/vcompm dac_8bit_0/latched_comparator_folded_0/vcompp 1.51fF
C3638 low_freq_pll_0/cs_ring_osc_0/vosc a_223312_n131500# 0.03fF
C3639 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d 1.91fF
C3640 a_238465_n122049# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout 0.03fF
C3641 dac_8bit_0/latched_comparator_folded_0/vlatchm VDD 6.80fF
C3642 peak_detector_0/ibiasn1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 1.43fF
C3643 input_amplifier_0/txgate_0/txb input_amplifier_0/venm1 0.35fF
C3644 biquad_gm_c_filter_0/gm_c_stage_1/vcmc biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail1 0.15fF
C3645 vfiltp biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail2 0.07fF
C3646 peak_detector_rst q0B 0.12fF
C3647 a_245481_n122255# a_245607_n121877# 0.04fF
C3648 biquad_gm_c_filter_0/ibiasn1 biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail1 0.07fF
C3649 biquad_gm_c_filter_0/ibiasn1 input_amplifier_0/ibiasn2 29.04fF
C3650 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_2/Q pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/D 0.06fF
C3651 dac_8bit_1/ibiasn dac_8bit_0/c4m 0.20fF
C3652 vrefA dac_8bit_0/amux_2to1_14/SELB 2.12fF
C3653 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 14.48fF
C3654 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 15.11fF
C3655 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/verr 15.32fF
C3656 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp 0.08fF
C3657 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 3.47fF
C3658 a_242104_n140786# VDD 0.69fF
C3659 a_241731_n115151# a_242102_n114873# 0.62fF
C3660 biquad_gm_c_filter_0/ibiasn1 vintp 0.16fF
C3661 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 13.66fF
C3662 vpeak_sampled dac_8bit_1/amux_2to1_1/SELB 2.07fF
C3663 input_amplifier_0/diff_fold_casc_ota_0/vbias4 input_amplifier_0/diff_fold_casc_ota_0/vcascnp 17.91fF
C3664 input_amplifier_0/diff_fold_casc_ota_0/vbias3 a_217060_n102324# 7.49fF
C3665 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp vse 0.86fF
C3666 gain_ctrl_1 input_amplifier_0/venm2 0.55fF
C3667 adc_compB a_383050_n152139# 0.05fF
C3668 vampm input_amplifier_0/venm2 2.18fF
C3669 dac_8bit_0/vcom_buf a_356329_n113250# 19.89fF
C3670 vampp input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc 4.62fF
C3671 vcp low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin 6.63fF
C3672 input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc vampp 0.60fF
C3673 diff_to_se_converter_0/ibiasn peak_detector_0/ibiasn2 4.18fF
C3674 VDD a_244971_n122799# 0.15fF
C3675 biquad_gm_c_filter_0/ibiasn3 vcp_sampled 0.40fF
C3676 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d 5.03fF
C3677 biquad_gm_c_filter_0/ibiasn2 comparator_0/ibiasn 1.55fF
C3678 a_246080_n122477# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/A 0.05fF
C3679 a_338703_n185409# a_338703_n185243# 0.02fF
C3680 low_freq_pll_0/cs_ring_osc_0/vpbias a_237498_n127742# 0.63fF
C3681 input_amplifier_0/vom1 input_amplifier_0/vim1 1.08fF
C3682 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q a_244783_n123337# 0.06fF
C3683 a_244617_n123337# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y 0.35fF
C3684 dac_8bit_1/amux_2to1_7/B vrefB 2.44fF
C3685 low_freq_pll_0/pfd_cp_lpf_0/vpbias low_freq_pll_0/pfd_cp_lpf_0/vswitchh 0.52fF
C3686 sample_and_hold_0/vholdm VDD 0.76fF
C3687 input_amplifier_0/txgate_5/txb input_amplifier_0/vip1 0.35fF
C3688 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_4/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q 0.07fF
C3689 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin a_244953_n138121# 0.03fF
C3690 a_227870_n122869# VDD 0.09fF
C3691 dac_8bit_0/c5m dac_8bit_0/amux_2to1_2/B 2.37fF
C3692 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn2 biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail2 0.58fF
C3693 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn biquad_gm_c_filter_0/gm_c_stage_3/vbiasp 0.53fF
C3694 dac_8bit_1/c2m dac_8bit_1/cdumm 10.49fF
C3695 dac_8bit_1/c3m dac_8bit_1/c1m 0.07fF
C3696 vlowB q6B 2.75fF
C3697 vfiltm biquad_gm_c_filter_0/gm_c_stage_3/vtail_diff 0.58fF
C3698 biquad_gm_c_filter_0/gm_c_stage_1/vcmc biquad_gm_c_filter_0/gm_c_stage_1/vcmcn 0.05fF
C3699 vrefA q1A 0.88fF
C3700 biquad_gm_c_filter_0/ibiasn3 biquad_gm_c_filter_0/gm_c_stage_3/vcmc 0.11fF
C3701 a_245649_n122281# a_246080_n122255# 0.31fF
C3702 peak_detector_0/ibiasn2 vbiasp 10.06fF
C3703 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/diff_fold_casc_ota_1/vtail_casc 8.06fF
C3704 adc_clk a_337864_n185269# 0.04fF
C3705 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp 19.65fF
C3706 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d 3.28fF
C3707 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 8.42fF
C3708 a_242951_n121193# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q 0.39fF
C3709 a_242783_n121167# a_242909_n120789# 0.04fF
C3710 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_1/A VDD 0.48fF
C3711 input_amplifier_0/diff_fold_casc_ota_0/vcascnp a_217060_n102324# 6.65fF
C3712 a_242526_n122281# a_242951_n122281# 0.04fF
C3713 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 0.56fF
C3714 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 28.76fF
C3715 low_freq_pll_0/pfd_cp_lpf_0/vQAb low_freq_pll_0/pfd_cp_lpf_0/vRSTN 0.29fF
C3716 sample dac_8bit_1/amux_2to1_6/SELB 2.36fF
C3717 a_242909_n120623# a_242783_n120257# 0.04fF
C3718 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin a_238771_n148007# 0.03fF
C3719 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_244617_n122249# 0.03fF
C3720 dac_8bit_0/latched_comparator_folded_0/vcomppb dac_8bit_0/latched_comparator_folded_0/vcompp 0.23fF
C3721 a_242273_n120623# a_242358_n120257# 0.11fF
C3722 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/A VDD 0.62fF
C3723 biquad_gm_c_filter_0/gm_c_stage_0/vbiasp VDD 3.04fF
C3724 dac_8bit_1/amux_2to1_1/SELB dac_8bit_1/amux_2to1_1/B 1.51fF
C3725 a_244783_n121711# a_244971_n121711# 0.26fF
C3726 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 5.47fF
C3727 input_amplifier_0/txgate_1/txb VDD 3.08fF
C3728 a_241919_n121161# a_242358_n121167# 0.63fF
C3729 a_336608_n185510# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/D 0.04fF
C3730 a_242085_n120623# a_242358_n120257# 0.38fF
C3731 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d 3.60fF
C3732 vrefA q2A 0.88fF
C3733 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d 0.75fF
C3734 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp 0.08fF
C3735 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VDD 2.04fF
C3736 a_246080_n123343# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_10/A 0.25fF
C3737 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A VDD 0.48fF
C3738 a_242273_n122799# VDD 0.15fF
C3739 dac_8bit_1/ibiasp vlowB 0.20fF
C3740 a_244617_n123337# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.03fF
C3741 a_241919_n122799# a_241919_n123337# 0.08fF
C3742 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm 0.75fF
C3743 a_336608_n185269# a_336608_n185510# 0.05fF
C3744 a_336408_n184969# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/D 0.02fF
C3745 a_244783_n121161# a_245481_n121167# 0.44fF
C3746 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/M1d 2.72fF
C3747 a_245224_n121193# a_245649_n121193# 0.04fF
C3748 input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/diff_fold_casc_ota_0/vfoldm 10.45fF
C3749 a_241731_n115151# VDD 0.37fF
C3750 a_356329_n113250# dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d 1.44fF
C3751 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 vocm 2.06fF
C3752 dac_8bit_0/c6m dac_8bit_0/c5m 1.39fF
C3753 dac_8bit_0/c7m dac_8bit_0/c4m 1.44fF
C3754 dac_8bit_0/amux_2to1_9/Y vcp_sampled 0.38fF
C3755 a_242867_n121345# a_242783_n121345# 0.05fF
C3756 a_242562_n140786# a_243020_n140786# 0.01fF
C3757 a_242104_n140786# a_243478_n140786# 0.01fF
C3758 a_222498_n127742# a_224330_n127742# 0.24fF
C3759 a_222956_n127742# a_223872_n127742# 1.33fF
C3760 biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail2 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn2 0.58fF
C3761 biquad_gm_c_filter_0/gm_c_stage_1/vbiasp biquad_gm_c_filter_0/gm_c_stage_1/vcmcn 0.53fF
C3762 a_241919_n122799# a_242085_n122799# 2.23fF
C3763 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.07fF
C3764 a_336408_n184969# a_336608_n185269# 0.38fF
C3765 a_336116_n185269# a_336537_n185243# 0.11fF
C3766 biquad_gm_c_filter_0/ibiasn3 biquad_gm_c_filter_0/gm_c_stage_3/vbiasp 0.04fF
C3767 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc input_amplifier_0/diff_fold_casc_ota_1/vtail_casc 23.17fF
C3768 input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_0/vbias3 0.02fF
C3769 input_amplifier_0/diff_fold_casc_ota_1/M13d input_amplifier_0/diff_fold_casc_ota_1/vcascnm 0.12fF
C3770 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/diff_fold_casc_ota_0/vbias4 1.53fF
C3771 vcp a_223312_n150168# 0.03fF
C3772 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vcascnm 0.69fF
C3773 vampm input_amplifier_0/diff_fold_casc_ota_1/vbias3 5.67fF
C3774 peak_detector_0/ibiasn1 low_freq_pll_0/ibiasn 0.47fF
C3775 vrefA dac_8bit_0/amux_2to1_13/SELB 2.12fF
C3776 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror vpeak 22.47fF
C3777 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn VDD 4.05fF
C3778 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 24.81fF
C3779 vbiasn dac_8bit_1/ibiasp 1.52fF
C3780 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp 0.28fF
C3781 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp a_230446_n180872# 10.36fF
C3782 peak_detector_0/verr peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 8.85fF
C3783 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.40fF
C3784 a_239330_n145742# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/csinvp 0.16fF
C3785 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc vocm 0.07fF
C3786 dac_8bit_1/latched_comparator_folded_0/vcompp_buf VDD 0.53fF
C3787 input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 0.10fF
C3788 dac_8bit_0/amux_2to1_4/B vrefA 2.44fF
C3789 a_245481_n121345# a_246080_n121389# 0.02fF
C3790 a_245649_n121443# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_7/A 0.04fF
C3791 dac_8bit_0/comp_outm adc_clk 0.04fF
C3792 a_246080_n123343# VDD 0.37fF
C3793 dac_8bit_1/latched_comparator_folded_0/vcompm dac_8bit_1/latched_comparator_folded_0/vcompm_buf 0.02fF
C3794 vlowB VDD 43.74fF
C3795 vcp a_223312_n132168# 0.03fF
C3796 low_freq_pll_0/cs_ring_osc_0/vosc low_freq_pll_0/cs_ring_osc_0/vpbias 2.76fF
C3797 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d 1.26fF
C3798 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.38fF
C3799 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp 0.08fF
C3800 VDD dac_8bit_1/amux_2to1_8/SELB 1.15fF
C3801 a_242783_n123343# a_242085_n123337# 0.44fF
C3802 pulse_generator_0/sky130_fd_sc_hd__inv_1_0/Y VDD 0.43fF
C3803 a_239251_n114759# a_239708_n115125# 0.01fF
C3804 a_245056_n122433# a_245481_n122433# 0.03fF
C3805 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/M1d 2.72fF
C3806 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/A 1.66fF
C3807 input_amplifier_0/diff_fold_casc_ota_1/M2d input_amplifier_0/diff_fold_casc_ota_1/vfoldm 10.45fF
C3808 low_freq_pll_0/pfd_cp_lpf_0/vpbias vcp 0.08fF
C3809 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 3.28fF
C3810 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp 58.37fF
C3811 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d 8.02fF
C3812 dac_8bit_0/amux_2to1_0/SELB VDD 1.15fF
C3813 input_amplifier_0/diff_fold_casc_ota_0/M2d input_amplifier_0/diff_fold_casc_ota_0/M3d 1.87fF
C3814 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/diff_fold_casc_ota_0/vbias2 11.85fF
C3815 input_amplifier_0/diff_fold_casc_ota_0/M1d input_amplifier_0/diff_fold_casc_ota_0/M6d 5.96fF
C3816 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/diff_fold_casc_ota_0/vfoldp 23.11fF
C3817 low_freq_pll_0/pfd_cp_lpf_0/vRSTN a_239708_n115125# 0.56fF
C3818 gain_ctrl_1 input_amplifier_0/txgate_2/txb 0.48fF
C3819 a_243382_n122477# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/A 0.05fF
C3820 a_239330_n145742# VDD 0.06fF
C3821 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm 3.14fF
C3822 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp 11.53fF
C3823 vampm input_amplifier_0/txgate_2/txb 0.53fF
C3824 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn1 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn2 0.17fF
C3825 vlowB q5B 2.75fF
C3826 dac_8bit_0/c1m vcp_sampled 1.94fF
C3827 a_245481_n121345# VDD 0.22fF
C3828 input_amplifier_0/vom1 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc 1.58fF
C3829 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror 2.23fF
C3830 dac_8bit_0/ibiasp dac_8bit_0/latched_comparator_folded_0/vlatchm 0.04fF
C3831 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q a_241919_n122799# 0.51fF
C3832 vampm input_amplifier_0/diff_fold_casc_ota_1/vcascnp 3.37fF
C3833 diff_to_se_converter_0/rst diff_to_se_converter_0/txgate_0/txb 0.36fF
C3834 a_242137_n115125# low_freq_pll_0/pfd_cp_lpf_0/vRSTN 0.01fF
C3835 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d 0.75fF
C3836 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_241919_n121161# 0.49fF
C3837 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp 0.08fF
C3838 a_244617_n122249# a_245481_n122255# 0.09fF
C3839 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y a_245649_n122281# 0.17fF
C3840 sample vlowA 3.83fF
C3841 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 vpeak 8.16fF
C3842 a_247701_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.03fF
C3843 a_338703_n185409# pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A 0.35fF
C3844 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y a_242273_n121711# 0.38fF
C3845 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin a_244954_n135628# 0.03fF
C3846 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/B a_335844_n185460# 0.37fF
C3847 q6A VDD 3.81fF
C3848 low_freq_pll_0/cs_ring_osc_0/vpbias a_221582_n127742# 0.51fF
C3849 adc_vcaparrayA dac_8bit_0/c4m 111.85fF
C3850 vlowB dac_8bit_1/amux_2to1_5/B 1.86fF
C3851 a_245481_n123343# a_245565_n123343# 0.05fF
C3852 a_245224_n121599# a_245224_n122281# 0.05fF
C3853 a_336537_n185243# a_336955_n185243# 0.04fF
C3854 a_336401_n185269# a_337592_n185269# 0.02fF
C3855 a_242085_n123337# a_242526_n123369# 0.28fF
C3856 VDD a_242085_n123337# 0.43fF
C3857 input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vbias3 11.45fF
C3858 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/csinvp a_228478_n140786# 0.16fF
C3859 a_227854_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.03fF
C3860 vrefA dac_8bit_0/amux_2to1_10/SELB 2.12fF
C3861 dac_8bit_0/c0m sample 2.36fF
C3862 input_amplifier_0/diff_fold_casc_ota_1/M2d input_amplifier_0/diff_fold_casc_ota_1/M13d 0.70fF
C3863 biquad_gm_c_filter_0/ibiasn2 peak_detector_0/ibiasn1 0.40fF
C3864 a_223313_n148007# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin 0.03fF
C3865 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_226785_n138121# 0.03fF
C3866 dac_8bit_0/c3m dac_8bit_0/c2m 0.16fF
C3867 vpeak sample_and_hold_1/vholdm 8.80fF
C3868 input_amplifier_0/diff_fold_casc_ota_1/M1d input_amplifier_0/diff_fold_casc_ota_1/M6d 5.96fF
C3869 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_10/A 0.27fF
C3870 input_amplifier_0/diff_fold_casc_ota_1/M2d input_amplifier_0/diff_fold_casc_ota_1/M3d 1.87fF
C3871 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/vfoldp 23.11fF
C3872 input_amplifier_0/diff_fold_casc_ota_1/vbias1 input_amplifier_0/diff_fold_casc_ota_1/vbias2 11.85fF
C3873 a_231785_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.03fF
C3874 a_245224_n123369# a_245224_n122687# 0.05fF
C3875 a_244783_n121161# a_244783_n121711# 0.05fF
C3876 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp 1.94fF
C3877 input_amplifier_0/diff_fold_casc_ota_0/vbias1 input_amplifier_0/vom1 1.02fF
C3878 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc 0.08fF
C3879 input_amplifier_0/diff_fold_casc_ota_0/M6d input_amplifier_0/diff_fold_casc_ota_0/vbias2 1.00fF
C3880 a_238312_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin 0.03fF
C3881 a_223414_n145742# a_224330_n145742# 0.79fF
C3882 a_244617_n121161# a_244783_n121161# 2.23fF
C3883 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_228312_n149500# 0.03fF
C3884 biquad_gm_c_filter_0/gm_c_stage_3/vcmc biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail1 0.15fF
C3885 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp 6.59fF
C3886 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d 5.99fF
C3887 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp 7.95fF
C3888 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d 15.11fF
C3889 vcp_sampled low_freq_pll_0/ibiasn 0.48fF
C3890 biquad_gm_c_filter_0/ibiasn2 biquad_gm_c_filter_0/gm_c_stage_1/vcmc 0.11fF
C3891 vrefA dac_8bit_0/amux_2to1_12/SELB 2.12fF
C3892 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d 0.16fF
C3893 comparator_0/ibiasn biquad_gm_c_filter_0/ibiasn4 0.91fF
C3894 vse diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm 13.89fF
C3895 input_amplifier_0/diff_fold_casc_ota_1/vfoldm vocm 0.02fF
C3896 low_freq_pll_0/pfd_cp_lpf_0/vQAb low_freq_pll_0/pfd_cp_lpf_0/vQA 3.28fF
C3897 dac_8bit_0/amux_2to1_6/B dac_8bit_0/amux_2to1_11/SELB 1.59fF
C3898 a_243382_n122255# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q 0.37fF
C3899 dac_8bit_1/latched_comparator_folded_0/vtailp dac_8bit_1/latched_comparator_folded_0/vlatchp 2.00fF
C3900 a_222040_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias 0.66fF
C3901 a_243382_n122255# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/A 0.05fF
C3902 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror 19.51fF
C3903 vcp low_freq_pll_0/pfd_cp_lpf_0/vQB 0.07fF
C3904 peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d a_230446_n180872# 1.44fF
C3905 a_338156_n185665# a_338156_n184969# 0.06fF
C3906 a_338149_n185569# a_338149_n185269# 0.08fF
C3907 comparator_0/vcompp comparator_0/vmirror 2.84fF
C3908 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_8/A 0.07fF
C3909 a_237396_n150168# vcp 0.03fF
C3910 dac_8bit_1/amux_2to1_6/SELB dac_8bit_1/cdumm 1.59fF
C3911 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/vip2 9.23fF
C3912 a_242085_n121711# VDD 0.43fF
C3913 a_242085_n122249# VDD 0.43fF
C3914 input_amplifier_0/vop1 input_amplifier_0/diff_fold_casc_ota_0/vcascnp 7.04fF
C3915 low_freq_pll_0/pfd_cp_lpf_0/vndiode VDD 0.32fF
C3916 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp 28.95fF
C3917 a_225730_n140786# a_227562_n140786# 0.65fF
C3918 a_226188_n140786# a_227104_n140786# 2.26fF
C3919 input_amplifier_0/diff_fold_casc_ota_1/vfoldp input_amplifier_0/diff_fold_casc_ota_1/M13d 1.62fF
C3920 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y a_245481_n121345# 0.14fF
C3921 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y VDD 0.93fF
C3922 input_amplifier_0/diff_fold_casc_ota_1/vbias1 vampm 0.93fF
C3923 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc 0.08fF
C3924 input_amplifier_0/diff_fold_casc_ota_1/M6d input_amplifier_0/diff_fold_casc_ota_1/vbias2 1.00fF
C3925 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/A 0.09fF
C3926 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_243313_n130007# 0.03fF
C3927 vhpf input_amplifier_0/vip1 31.09fF
C3928 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_10/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.07fF
C3929 adc_clk pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/D 0.21fF
C3930 vpeak_sampled dac_8bit_1/amux_2to1_2/B 0.38fF
C3931 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin a_237397_n130007# 0.03fF
C3932 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y a_245224_n122687# 0.15fF
C3933 a_244617_n122799# a_245056_n122433# 0.63fF
C3934 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q a_245481_n121345# 0.05fF
C3935 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp 19.65fF
C3936 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d 3.28fF
C3937 adc_vcaparrayA dac_8bit_0/adc_run 0.36fF
C3938 input_amplifier_0/diff_fold_casc_ota_0/vbias2 input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc 2.34fF
C3939 input_amplifier_0/diff_fold_casc_ota_0/M6d input_amplifier_0/vom1 2.11fF
C3940 a_246080_n121167# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/A 0.05fF
C3941 dac_8bit_1/c4m dac_8bit_1/c1m 1.12fF
C3942 dac_8bit_1/c5m dac_8bit_1/c0m 0.43fF
C3943 a_244971_n122255# a_244971_n122799# 0.02fF
C3944 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VDD 1.46fF
C3945 input_amplifier_0/vip2 vocm 0.35fF
C3946 a_337497_n185269# a_337864_n185269# 0.02fF
C3947 vampp biquad_gm_c_filter_0/gm_c_stage_0/vcmc 0.12fF
C3948 a_335844_n185269# a_336401_n185269# 0.11fF
C3949 vlowB q4B 2.75fF
C3950 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/A 1.64fF
C3951 a_242358_n122433# a_242783_n122433# 0.03fF
C3952 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VDD 1.49fF
C3953 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn a_162668_n147576# 0.11fF
C3954 dac_8bit_0/cdumm dac_8bit_1/ibiasn 0.20fF
C3955 input_amplifier_0/diff_fold_casc_ota_0/M13d input_amplifier_0/diff_fold_casc_ota_0/vtail_casc 0.04fF
C3956 dac_8bit_0/comp_outm dac_8bit_0/latched_comparator_folded_0/vcompp 0.08fF
C3957 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror a_230446_n180872# 8.05fF
C3958 a_244617_n121711# VDD 0.78fF
C3959 a_245481_n122255# a_245565_n122255# 0.05fF
C3960 biquad_gm_c_filter_0/ibiasn2 biquad_gm_c_filter_0/gm_c_stage_1/vbiasp 0.04fF
C3961 sample_and_hold_0/vholdm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp 1.42fF
C3962 dac_8bit_0/amux_2to1_5/SELB dac_8bit_0/amux_2to1_5/B 1.51fF
C3963 vse VDD 4.91fF
C3964 comparator_0/ibiasn input_amplifier_0/ibiasn2 0.28fF
C3965 adc_vcaparrayB dac_8bit_1/c6m 427.49fF
C3966 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin VDD 4.26fF
C3967 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d 0.56fF
C3968 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm 0.19fF
C3969 input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc vocm 2.02fF
C3970 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn1 vampp 0.11fF
C3971 a_242102_n114873# a_242380_n114857# 0.29fF
C3972 a_241731_n115151# a_242419_n114983# 0.12fF
C3973 a_243020_n140786# VDD 0.09fF
C3974 input_amplifier_0/diff_fold_casc_ota_0/vfoldm input_amplifier_0/vop1 6.63fF
C3975 q5A VDD 3.81fF
C3976 a_242085_n121711# a_242526_n121599# 0.28fF
C3977 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 9.59fF
C3978 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_2/Q pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/D 0.03fF
C3979 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VDD 6.84fF
C3980 dac_8bit_0/amux_2to1_2/SELB dac_8bit_0/c5m 1.59fF
C3981 input_amplifier_0/vip2 input_amplifier_0/vom1 33.30fF
C3982 vlowB dac_8bit_1/amux_2to1_15/SELB 1.62fF
C3983 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc 0.63fF
C3984 input_amplifier_0/diff_fold_casc_ota_1/M3d input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc 0.64fF
C3985 vrefA dac_8bit_0/amux_2to1_9/SELB 2.12fF
C3986 vocm input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 2.06fF
C3987 dac_8bit_1/ibiasn dac_8bit_1/ibiasp 0.25fF
C3988 biquad_gm_c_filter_0/ibiasn2 vcp_sampled 0.39fF
C3989 diff_to_se_converter_0/rst diff_to_se_converter_0/txgate_1/txb 0.39fF
C3990 input_amplifier_0/diff_fold_casc_ota_1/M6d vampm 2.11fF
C3991 a_245224_n123369# a_244971_n123343# 0.04fF
C3992 input_amplifier_0/diff_fold_casc_ota_1/vbias2 input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc 2.34fF
C3993 biquad_gm_c_filter_0/ibiasn1 comparator_0/ibiasn 10.01fF
C3994 VDD low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.38fF
C3995 low_freq_pll_0/cs_ring_osc_0/vpbias a_238414_n127742# 0.76fF
C3996 low_freq_pll_0/pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/Q_N VDD 0.23fF
C3997 input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc input_amplifier_0/vom1 2.96fF
C3998 vpeak_sampled dac_8bit_1/c6m 1.94fF
C3999 sample dac_8bit_1/amux_2to1_7/B 2.66fF
C4000 dac_8bit_0/amux_2to1_16/SELB VDD 1.15fF
C4001 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/A 0.10fF
C4002 a_236175_n122049# VDD 0.01fF
C4003 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d VDD 11.46fF
C4004 input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 0.37fF
C4005 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q 0.08fF
C4006 dac_8bit_1/latched_comparator_folded_0/vcompm_buf VDD 0.53fF
C4007 input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 0.36fF
C4008 vrefA dac_8bit_0/amux_2to1_11/SELB 2.12fF
C4009 adc_clk a_338149_n185269# 1.31fF
C4010 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VDD 7.64fF
C4011 vbiasn dac_8bit_0/ibiasp 1.23fF
C4012 biquad_gm_c_filter_0/gm_c_stage_2/vbiasp vfiltm 0.10fF
C4013 a_243382_n121167# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q 0.37fF
C4014 input_amplifier_0/diff_fold_casc_ota_0/M3d input_amplifier_0/vop1 1.08fF
C4015 a_242358_n122255# a_242783_n122255# 0.03fF
C4016 vampp biquad_gm_c_filter_0/gm_c_stage_0/vtail_diff 2.73fF
C4017 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d VDD 7.37fF
C4018 a_239143_n115125# a_239708_n115125# 0.01fF
C4019 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d VDD 9.36fF
C4020 a_242867_n121167# VDD 0.02fF
C4021 dac_8bit_1/ibiasn VDD 3.15fF
C4022 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 58.37fF
C4023 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 8.02fF
C4024 dac_8bit_0/amux_2to1_8/SELB vcp_sampled 2.07fF
C4025 a_245056_n121345# a_244971_n121711# 0.11fF
C4026 vampm input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc 7.09fF
C4027 peak_detector_0/ibiasn2 vpeak_sampled 0.46fF
C4028 q7A q0A 0.10fF
C4029 a_241919_n121161# a_242783_n121167# 0.09fF
C4030 input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc vampm 2.96fF
C4031 a_244617_n121711# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y 0.35fF
C4032 a_242526_n120511# a_242951_n120355# 0.04fF
C4033 a_242085_n120623# a_242783_n120257# 0.44fF
C4034 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_244783_n121711# 0.08fF
C4035 vrefA dac_8bit_0/amux_2to1_2/B 2.44fF
C4036 a_242867_n122433# VDD 0.02fF
C4037 a_237040_n127742# VDD 1.55fF
C4038 input_amplifier_0/diff_fold_casc_ota_0/M6d input_amplifier_0/diff_fold_casc_ota_0/M13d 0.56fF
C4039 a_337864_n185555# a_338084_n185421# 0.04fF
C4040 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y 0.13fF
C4041 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q a_244617_n121711# 0.03fF
C4042 dac_8bit_0/c2m dac_8bit_0/c6m 2.04fF
C4043 dac_8bit_0/cdumm dac_8bit_0/c7m 0.86fF
C4044 a_336537_n185243# a_336537_n185409# 0.05fF
C4045 sample dac_8bit_1/cdumm 2.36fF
C4046 vintm biquad_gm_c_filter_0/gm_c_stage_0/vcmc 0.10fF
C4047 a_242783_n123343# a_243382_n123343# 0.02fF
C4048 a_245056_n121167# a_245481_n121167# 0.03fF
C4049 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin a_221480_n149500# 0.03fF
C4050 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/A 1.64fF
C4051 a_242380_n114857# VDD 1.23fF
C4052 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp 7.95fF
C4053 vlowB q3B 2.75fF
C4054 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d 15.11fF
C4055 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q a_242783_n121345# 0.05fF
C4056 a_243020_n140786# a_243478_n140786# 0.02fF
C4057 peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d VDD 1.27fF
C4058 a_223414_n127742# a_224330_n127742# 0.79fF
C4059 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y a_242526_n122687# 0.15fF
C4060 a_241919_n122799# a_242358_n122433# 0.63fF
C4061 dac_8bit_1/c6m dac_8bit_1/amux_2to1_1/B 2.37fF
C4062 a_336401_n185269# a_336537_n185243# 0.37fF
C4063 a_336408_n184969# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/D 0.55fF
C4064 a_242085_n121161# a_242358_n121167# 0.38fF
C4065 vcp low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/csinvn 0.08fF
C4066 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d 5.21fF
C4067 vocm_filt biquad_gm_c_filter_0/gm_c_stage_1/vbiasp 0.10fF
C4068 peak_detector_0/ibiasn1 biquad_gm_c_filter_0/ibiasn4 0.42fF
C4069 vse diff_to_se_converter_0/vip 7.89fF
C4070 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn1 vintm 0.03fF
C4071 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail1 0.58fF
C4072 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q 0.29fF
C4073 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror 28.69fF
C4074 dac_8bit_0/amux_2to1_1/B VDD 4.57fF
C4075 q4A VDD 3.81fF
C4076 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_241481_n148007# 0.03fF
C4077 vcomp a_242380_n114857# 0.04fF
C4078 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/A 1.64fF
C4079 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d 2.72fF
C4080 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 9.20fF
C4081 dac_8bit_1/latched_comparator_folded_0/vcompp_buf dac_8bit_1/latched_comparator_folded_0/vcomppb 0.32fF
C4082 vlowB dac_8bit_1/amux_2to1_14/SELB 1.62fF
C4083 a_246080_n121389# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_7/A 0.25fF
C4084 dac_8bit_0/latched_comparator_folded_0/vlatchp dac_8bit_0/latched_comparator_folded_0/vlatchm 3.86fF
C4085 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm 0.19fF
C4086 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 6.88fF
C4087 VDD input_amplifier_0/ibiasn1 1.56fF
C4088 vcp low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/csinvn 0.08fF
C4089 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y 1.64fF
C4090 a_242783_n123343# a_242358_n123343# 0.03fF
C4091 a_245481_n121167# low_freq_pll_0/freq_div_0/vout 0.04fF
C4092 a_243382_n123343# VDD 0.37fF
C4093 a_245649_n122531# a_246080_n122477# 0.31fF
C4094 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d VDD 9.36fF
C4095 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VDD 12.54fF
C4096 dac_8bit_0/c3m dac_8bit_0/c4m 1.18fF
C4097 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/csinvp low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin 0.10fF
C4098 vintm biquad_gm_c_filter_0/gm_c_stage_2/vcmcn2 2.05fF
C4099 dac_8bit_0/amux_2to1_15/SELB VDD 1.15fF
C4100 peak_detector_0/ibiasn2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 0.60fF
C4101 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d 7.88fF
C4102 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror 0.69fF
C4103 low_freq_pll_0/pfd_cp_lpf_0/vRSTN low_freq_pll_0/pfd_cp_lpf_0/vQB 1.19fF
C4104 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm 5.03fF
C4105 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp 3.66fF
C4106 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 24.81fF
C4107 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_7/A VDD 0.48fF
C4108 dac_8bit_1/c7m dac_8bit_1/c6m 2.04fF
C4109 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp 4.15fF
C4110 vocm_filt biquad_gm_c_filter_0/gm_c_stage_3/vcmc 0.24fF
C4111 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d 0.56fF
C4112 vcp a_230412_n134960# 0.03fF
C4113 peak_detector_0/ibiasn1 input_amplifier_0/ibiasn2 2.69fF
C4114 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y a_246080_n122255# 0.11fF
C4115 dac_8bit_0/amux_2to1_7/B q1A 1.99fF
C4116 VDD dac_8bit_1/c0m 2.48fF
C4117 biquad_gm_c_filter_0/gm_c_stage_2/vcmc biquad_gm_c_filter_0/gm_c_stage_2/vtail_diff 0.03fF
C4118 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn2 biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail2 0.58fF
C4119 dac_8bit_0/cdumm adc_vcaparrayA 11.56fF
C4120 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn a_230446_n180872# 0.11fF
C4121 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/vip 28.95fF
C4122 vintm biquad_gm_c_filter_0/gm_c_stage_0/vtail_diff 2.75fF
C4123 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin a_245870_n135628# 0.03fF
C4124 dac_8bit_0/vcom_buf dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp 23.02fF
C4125 VDD input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc 5.18fF
C4126 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q 0.29fF
C4127 dac_8bit_0/c7m VDD 2.60fF
C4128 low_freq_pll_0/cs_ring_osc_0/vpbias a_222498_n127742# 0.63fF
C4129 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VDD 19.81fF
C4130 a_245056_n121345# a_245056_n122255# 0.05fF
C4131 a_245481_n121345# a_244783_n122249# 0.01fF
C4132 a_244783_n121711# a_245481_n122255# 0.01fF
C4133 vlowB q1B 2.75fF
C4134 dac_8bit_1/amux_2to1_9/SELB dac_8bit_1/amux_2to1_9/Y 1.59fF
C4135 a_242484_n120623# a_242358_n120257# 0.02fF
C4136 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/D a_337497_n185269# 0.46fF
C4137 a_242526_n123369# a_242358_n123343# 0.59fF
C4138 a_242085_n123337# a_242951_n123369# 0.11fF
C4139 VDD a_242358_n123343# 0.36fF
C4140 a_242273_n120623# a_241919_n120623# 0.21fF
C4141 a_228770_n131500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.03fF
C4142 adc_compA dac_8bit_0/latched_comparator_folded_0/vcompp_buf 0.12fF
C4143 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_242085_n121161# 0.08fF
C4144 biquad_gm_c_filter_0/ibiasn1 peak_detector_0/ibiasn1 0.41fF
C4145 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm 3.14fF
C4146 input_amplifier_0/diff_fold_casc_ota_1/vfoldm input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 0.03fF
C4147 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 13.36fF
C4148 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_227701_n138121# 0.03fF
C4149 a_241919_n120623# a_242085_n120623# 2.23fF
C4150 a_232701_n138121# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.03fF
C4151 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VDD 12.54fF
C4152 a_244783_n123337# a_245481_n122433# 0.01fF
C4153 a_245481_n123343# a_244783_n122799# 0.01fF
C4154 a_245056_n123343# a_245056_n122433# 0.05fF
C4155 VDD input_amplifier_0/rst 1.57fF
C4156 a_245224_n121193# a_245224_n121599# 0.03fF
C4157 vintp biquad_gm_c_filter_0/gm_c_stage_1/vcmc 0.10fF
C4158 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VDD 25.41fF
C4159 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d 5.21fF
C4160 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 adc_vcaparrayB 0.08fF
C4161 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm 2.41fF
C4162 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror 17.44fF
C4163 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror a_162668_n147576# 8.05fF
C4164 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 21.43fF
C4165 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 16.73fF
C4166 vlowB q2B 2.75fF
C4167 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y a_245224_n121193# 0.15fF
C4168 a_244617_n121161# a_245056_n121167# 0.63fF
C4169 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d a_356329_n164260# 0.79fF
C4170 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 0.04fF
C4171 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q a_241919_n121711# 0.03fF
C4172 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d 0.82fF
C4173 adc_vcaparrayB dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp 0.28fF
C4174 vocm_filt biquad_gm_c_filter_0/gm_c_stage_3/vbiasp 0.10fF
C4175 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d 1.74fF
C4176 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/csinvp a_240730_n140786# 0.08fF
C4177 vcp_sampled biquad_gm_c_filter_0/ibiasn4 0.41fF
C4178 a_335844_n185460# VDD 0.45fF
C4179 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm a_189446_n180872# 10.16fF
C4180 peak_detector_0/vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 12.64fF
C4181 q3A VDD 3.81fF
C4182 dac_8bit_0/amux_2to1_4/B dac_8bit_0/amux_2to1_4/SELB 1.51fF
C4183 a_222956_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias 0.83fF
C4184 vpeak_sampled dac_8bit_1/amux_2to1_2/SELB 2.07fF
C4185 vampp VDD 8.39fF
C4186 a_245565_n123343# VDD 0.02fF
C4187 a_338356_n185510# a_338149_n185269# 0.01fF
C4188 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y a_242526_n122281# 0.15fF
C4189 a_241919_n122249# a_242358_n122255# 0.63fF
C4190 a_238312_n150168# vcp 0.03fF
C4191 input_amplifier_0/vip2 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 0.07fF
C4192 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q 0.08fF
C4193 a_242358_n121345# VDD 0.36fF
C4194 vlowB dac_8bit_1/amux_2to1_13/SELB 1.62fF
C4195 sample sample_and_hold_1/vholdm 0.82fF
C4196 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 3.60fF
C4197 comparator_0/vcompm vfiltm 0.06fF
C4198 dac_8bit_0/ibiasn dac_8bit_1/ibiasn 6.02fF
C4199 dac_8bit_1/ibiasn dac_8bit_0/ibiasp 0.23fF
C4200 a_226188_n140786# a_228020_n140786# 0.43fF
C4201 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin 0.38fF
C4202 a_225730_n140786# a_228478_n140786# 0.14fF
C4203 a_226646_n140786# a_227562_n140786# 1.92fF
C4204 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_7/A 0.27fF
C4205 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_0/vholdm 4.81fF
C4206 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 a_356329_n164260# 8.26fF
C4207 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 44.84fF
C4208 vfiltp VDD 2.49fF
C4209 adc_vcaparrayA VDD 3.82fF
C4210 a_335749_n185813# a_335844_n185460# 0.31fF
C4211 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn 0.61fF
C4212 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 12.94fF
C4213 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror a_356329_n164260# 8.05fF
C4214 dac_8bit_1/amux_2to1_9/Y vrefB 1.93fF
C4215 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin a_238313_n130007# 0.03fF
C4216 a_244617_n122799# a_245481_n122433# 0.09fF
C4217 vintp biquad_gm_c_filter_0/gm_c_stage_1/vbiasp 0.42fF
C4218 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y a_245649_n122531# 0.17fF
C4219 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_7/A 0.07fF
C4220 vlowB q7B 2.75fF
C4221 dac_8bit_0/amux_2to1_14/SELB VDD 1.15fF
C4222 vpeak_sampled dac_8bit_1/amux_2to1_4/B 0.38fF
C4223 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 3.45fF
C4224 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm 23.84fF
C4225 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp adc_vcaparrayB 28.95fF
C4226 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm 12.61fF
C4227 dac_8bit_1/c3m dac_8bit_1/c0m 0.07fF
C4228 dac_8bit_1/c2m dac_8bit_1/c1m 1.20fF
C4229 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d 1.91fF
C4230 a_336608_n185269# a_336757_n185243# 0.02fF
C4231 a_337592_n185269# a_338156_n184969# 0.11fF
C4232 a_335844_n185269# a_336537_n185243# 0.04fF
C4233 a_242951_n122531# a_243382_n122477# 0.31fF
C4234 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 3.28fF
C4235 vcp_sampled input_amplifier_0/ibiasn2 0.83fF
C4236 a_338107_n185787# VDD 0.02fF
C4237 dac_8bit_0/latched_comparator_folded_0/vcompmb VDD 0.47fF
C4238 a_242526_n122281# a_242273_n122255# 0.04fF
C4239 vse diff_to_se_converter_0/vim 30.71fF
C4240 a_337592_n185460# VDD 0.45fF
C4241 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 5.68fF
C4242 a_221582_n145742# VDD 0.73fF
C4243 a_242102_n114873# a_242575_n114888# 0.01fF
C4244 a_242380_n114857# a_242419_n114983# 1.60fF
C4245 a_241731_n115151# a_242506_n114759# 0.03fF
C4246 a_242526_n121599# a_242358_n121345# 0.59fF
C4247 a_242085_n121711# a_242951_n121443# 0.11fF
C4248 dac_8bit_1/amux_2to1_0/B VDD 4.57fF
C4249 sample dac_8bit_1/amux_2to1_7/SELB 2.36fF
C4250 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 8.90fF
C4251 rst_n input_amplifier_0/ibiasn1 0.19fF
C4252 a_244617_n121711# a_244783_n122249# 0.02fF
C4253 a_244783_n121711# a_244617_n122249# 0.02fF
C4254 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror 19.51fF
C4255 a_236582_n145742# a_237498_n145742# 2.99fF
C4256 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn2 VDD 1.51fF
C4257 biquad_gm_c_filter_0/ibiasn1 vcp_sampled 0.40fF
C4258 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_0/vholdm 0.08fF
C4259 a_245056_n123343# a_245182_n122965# 0.02fF
C4260 dac_8bit_0/c2m dac_8bit_0/amux_2to1_5/B 1.72fF
C4261 dac_8bit_0/amux_2to1_7/B dac_8bit_0/amux_2to1_10/SELB 1.59fF
C4262 q1A VDD 3.81fF
C4263 vintp biquad_gm_c_filter_0/gm_c_stage_3/vcmc 0.51fF
C4264 low_freq_pll_0/cs_ring_osc_0/vpbias a_239330_n127742# 0.77fF
C4265 low_freq_pll_0/pfd_cp_lpf_0/vQA low_freq_pll_0/pfd_cp_lpf_0/vQB 0.15fF
C4266 a_244783_n123337# a_244617_n122799# 0.02fF
C4267 a_244617_n123337# a_244783_n122799# 0.02fF
C4268 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm adc_vcaparrayB 0.75fF
C4269 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout a_236174_n119618# 0.03fF
C4270 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror 4.50fF
C4271 vlowB dac_8bit_1/amux_2to1_10/SELB 1.62fF
C4272 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm 0.08fF
C4273 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 1.65fF
C4274 a_237091_n122049# VDD 0.01fF
C4275 dac_8bit_0/c6m dac_8bit_0/c4m 1.44fF
C4276 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_244783_n122799# 0.03fF
C4277 dac_8bit_1/comp_outm dac_8bit_1/latched_comparator_folded_0/vcompp_buf 0.21fF
C4278 dac_8bit_1/latched_comparator_folded_0/vcompp adc_clk 0.37fF
C4279 vrefA q0A 0.88fF
C4280 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d 2.62fF
C4281 adc_clk a_338285_n185243# 0.06fF
C4282 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm 2.00fF
C4283 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm peak_detector_0/vpeak 6.29fF
C4284 input_amplifier_0/vip2 input_amplifier_0/ibiasn2 0.31fF
C4285 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm a_275374_n180872# 10.16fF
C4286 vintm VDD 2.01fF
C4287 q2A VDD 3.81fF
C4288 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/vim 5.59fF
C4289 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp 4.15fF
C4290 dac_8bit_0/c3m dac_8bit_0/amux_2to1_4/SELB 1.59fF
C4291 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/vhold 1.41fF
C4292 VDD input_amplifier_0/vim2 3.63fF
C4293 a_242951_n122281# a_243382_n122255# 0.31fF
C4294 dac_8bit_0/ibiasn dac_8bit_0/c7m 0.19fF
C4295 dac_8bit_0/ibiasp dac_8bit_0/c7m 0.10fF
C4296 a_225580_n122869# a_226496_n122869# 3.27fF
C4297 a_239883_n115151# a_240447_n115125# 0.30fF
C4298 low_freq_pll_0/pfd_cp_lpf_0/vRSTN a_241634_n115151# 0.10fF
C4299 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp 0.08fF
C4300 vlowB dac_8bit_1/amux_2to1_12/SELB 1.62fF
C4301 a_245151_n121167# VDD 0.02fF
C4302 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 9.59fF
C4303 sample dac_8bit_1/adc_run 0.38fF
C4304 rst_n input_amplifier_0/rst 0.47fF
C4305 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp 0.08fF
C4306 dac_8bit_0/amux_2to1_5/B vrefA 2.44fF
C4307 dac_8bit_1/amux_2to1_1/SELB dac_8bit_1/c6m 1.59fF
C4308 a_242273_n123343# a_242526_n123369# 0.04fF
C4309 a_242273_n123343# VDD 0.15fF
C4310 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 vse 2.45fF
C4311 a_242358_n120257# a_242783_n120257# 0.03fF
C4312 diff_to_se_converter_0/vip vfiltp 31.71fF
C4313 a_245224_n122687# a_244971_n122799# 0.04fF
C4314 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q VDD 0.38fF
C4315 a_237956_n127742# VDD 0.69fF
C4316 a_236480_n149500# low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.03fF
C4317 dac_8bit_0/vcom_buf dac_8bit_0/latched_comparator_folded_0/vtailp 2.62fF
C4318 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 vse 3.16fF
C4319 vcp a_236480_n132168# 0.03fF
C4320 dac_8bit_0/amux_2to1_13/SELB VDD 1.15fF
C4321 dac_8bit_0/amux_2to1_1/SELB VDD 1.15fF
C4322 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/A VDD 0.62fF
C4323 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/D pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/D 0.11fF
C4324 a_243382_n123343# low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_5/A 0.25fF
C4325 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm 0.19fF
C4326 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 6.88fF
C4327 a_337497_n185813# a_337592_n185460# 0.31fF
C4328 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin a_222396_n149500# 0.03fF
C4329 input_amplifier_0/ibiasn2 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 1.79fF
C4330 a_245649_n121193# a_246080_n121167# 0.31fF
C4331 a_242575_n114888# VDD 0.33fF
C4332 comparator_0/vo1 VDD 2.00fF
C4333 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_3/A 0.07fF
C4334 a_241919_n122799# a_242783_n122433# 0.09fF
C4335 dac_8bit_0/c0m vcp_sampled 1.85fF
C4336 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y a_242951_n122531# 0.17fF
C4337 a_336608_n185269# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/D 0.04fF
C4338 peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 0.56fF
C4339 a_242526_n121193# a_242951_n121193# 0.04fF
C4340 a_242085_n121161# a_242783_n121167# 0.44fF
C4341 diff_to_se_converter_0/ibiasn VDD 2.60fF
C4342 low_freq_pll_0/cs_ring_osc_0/vpbias a_226188_n140786# 0.66fF
C4343 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/csinvp VDD 0.48fF
C4344 dac_8bit_0/amux_2to1_4/B VDD 4.57fF
C4345 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 44.84fF
C4346 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 a_275374_n180872# 8.26fF
C4347 dac_8bit_0/latched_comparator_folded_0/vcompm_buf adc_compA 0.20fF
C4348 vcp_sampled sample 14.31fF
C4349 a_245224_n121193# a_244971_n121167# 0.04fF
C4350 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm 0.08fF
C4351 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 1.35fF
C4352 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm 20.84fF
C4353 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn 5.68fF
C4354 vlowB dac_8bit_1/amux_2to1_17/SELB 1.62fF
C4355 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A a_336408_n185665# 0.02fF
C4356 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_242397_n148007# 0.03fF
C4357 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/vhold 0.08fF
C4358 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror 17.44fF
C4359 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm 2.41fF
C4360 peak_detector_0/ibiasn2 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp 0.16fF
C4361 vlowB dac_8bit_1/amux_2to1_6/B 1.86fF
C4362 comparator_0/vo1 vcomp 1.46fF
C4363 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d dac_8bit_1/vcom_buf 15.32fF
C4364 vfiltp rst_n 0.48fF
C4365 vampm biquad_gm_c_filter_0/gm_c_stage_0/vtail_diff 0.33fF
C4366 dac_8bit_1/amux_2to1_7/SELB dac_8bit_1/amux_2to1_7/B 1.51fF
C4367 low_freq_pll_0/pfd_cp_lpf_0/vswitchh VDD 10.21fF
C4368 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A a_336116_n185269# 0.05fF
C4369 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 44.84fF
C4370 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 a_275374_n146348# 8.26fF
C4371 VDD input_amplifier_0/diff_fold_casc_ota_0/M2d 9.25fF
C4372 dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d 5.10fF
C4373 peak_detector_rst pulse_generator_0/sky130_fd_sc_hd__inv_1_1/A 0.27fF
C4374 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp 0.08fF
C4375 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d 1.26fF
C4376 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 13.22fF
C4377 a_336955_n185409# VDD 0.15fF
C4378 VDD vbiasp 49.03fF
C4379 dac_8bit_0/c3m dac_8bit_0/cdumm 0.07fF
C4380 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_6/A low_freq_pll_0/freq_div_0/vout 0.07fF
C4381 dac_8bit_1/latched_comparator_folded_0/vlatchm dac_8bit_1/latched_comparator_folded_0/vcompm 0.54fF
C4382 a_243382_n123343# a_242951_n123369# 0.31fF
C4383 a_239870_n114759# a_239708_n115125# 0.04fF
C4384 adc_vcaparrayA dac_8bit_0/ibiasp 0.18fF
C4385 biquad_gm_c_filter_0/ibiasn3 input_amplifier_0/ibiasn1 0.19fF
C4386 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q a_244617_n123337# 0.41fF
C4387 dac_8bit_1/latched_comparator_folded_0/vtailp vlowB 1.83fF
C4388 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm 16.88fF
C4389 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 3.47fF
C4390 vcomp low_freq_pll_0/pfd_cp_lpf_0/vswitchh 0.10fF
C4391 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 adc_vcaparrayA 0.71fF
C4392 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm 12.94fF
C4393 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 0.61fF
C4394 vlowB dac_8bit_1/amux_2to1_9/SELB 1.62fF
C4395 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VDD 1.46fF
C4396 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_239953_n138121# 0.03fF
C4397 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm 0.08fF
C4398 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d vse 15.32fF
C4399 dac_8bit_1/vcom_buf dac_8bit_1/latched_comparator_folded_0/vlatchm 0.05fF
C4400 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d 5.21fF
C4401 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 8.42fF
C4402 a_238793_n115125# VDD 1.24fF
C4403 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 3.45fF
C4404 dac_8bit_0/amux_2to1_10/SELB VDD 1.15fF
C4405 dac_8bit_1/vcom_buf dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 13.20fF
C4406 a_336336_n185421# a_336116_n185555# 0.04fF
C4407 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d 7.88fF
C4408 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror 0.69fF
C4409 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm 5.03fF
C4410 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 sample_and_hold_1/vholdm 2.37fF
C4411 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q 0.02fF
C4412 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp 3.66fF
C4413 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin a_246786_n135628# 0.03fF
C4414 low_freq_pll_0/cs_ring_osc_0/vpbias a_223414_n127742# 0.76fF
C4415 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_1/vcom_buf 22.36fF
C4416 low_freq_pll_0/cs_ring_osc_0/vosc a_221481_n130007# 0.03fF
C4417 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y 0.03fF
C4418 a_245649_n121443# a_245649_n122281# 0.09fF
C4419 a_338156_n185665# pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A 0.48fF
C4420 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/A 0.03fF
C4421 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror 14.22fF
C4422 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d 1.91fF
C4423 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp 1.03fF
C4424 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_242951_n120355# 0.39fF
C4425 input_amplifier_0/diff_fold_casc_ota_1/M1d VDD 10.42fF
C4426 dac_8bit_0/amux_2to1_3/SELB dac_8bit_0/amux_2to1_3/B 1.51fF
C4427 vlowB dac_8bit_1/amux_2to1_11/SELB 1.62fF
C4428 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/D a_337864_n185269# 0.04fF
C4429 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d 0.82fF
C4430 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d 1.74fF
C4431 VDD input_amplifier_0/diff_fold_casc_ota_0/vfoldp 17.12fF
C4432 a_242358_n123343# a_242951_n123369# 0.02fF
C4433 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q VDD 2.18fF
C4434 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn2 VDD 1.51fF
C4435 a_244617_n121711# a_244971_n121711# 0.21fF
C4436 dac_8bit_1/latched_comparator_folded_0/vcompm adc_clk 0.51fF
C4437 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 5.68fF
C4438 biquad_gm_c_filter_0/gm_c_stage_0/vbiasp vocm_filt 0.10fF
C4439 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn vfiltp 0.42fF
C4440 a_244971_n123343# a_244971_n122799# 0.02fF
C4441 comparator_0/ibiasn peak_detector_0/ibiasn1 0.56fF
C4442 a_241919_n120623# a_242358_n120257# 0.63fF
C4443 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y a_242526_n120511# 0.15fF
C4444 input_amplifier_0/vip2 gain_ctrl_0 0.52fF
C4445 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d a_189446_n180872# 0.79fF
C4446 peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 0.04fF
C4447 a_245649_n123369# a_245649_n122531# 0.09fF
C4448 VDD vincm 2.34fF
C4449 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/A 0.03fF
C4450 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/A low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y 0.03fF
C4451 vpeak_sampled dac_8bit_1/amux_2to1_3/B 0.38fF
C4452 a_245056_n121167# a_245056_n121345# 0.08fF
C4453 dac_8bit_0/amux_2to1_12/SELB VDD 1.15fF
C4454 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_226023_n148007# 0.03fF
C4455 a_244954_n134960# vcp 0.03fF
C4456 vcp_sampled sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d 4.98fF
C4457 a_245224_n122281# VDD 0.23fF
C4458 dac_8bit_1/c4m dac_8bit_1/c0m 0.43fF
C4459 dac_8bit_1/vcom_buf adc_clk 0.24fF
C4460 q0B dac_8bit_1/amux_2to1_9/Y 1.99fF
C4461 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 0.97fF
C4462 a_335844_n185269# pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/Q_N 0.02fF
C4463 a_244617_n121161# a_245481_n121167# 0.09fF
C4464 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y a_245649_n121193# 0.17fF
C4465 a_242526_n122687# a_242273_n122799# 0.04fF
C4466 dac_8bit_0/c1m dac_8bit_1/ibiasn 0.20fF
C4467 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d 3.07fF
C4468 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp 3.66fF
C4469 peak_detector_0/ibiasn1 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm 3.89fF
C4470 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/csinvp a_241646_n140786# 0.09fF
C4471 a_336401_n185569# VDD 0.81fF
C4472 adc_vcaparrayB dac_8bit_1/c5m 214.58fF
C4473 diff_to_se_converter_0/ibiasn diff_to_se_converter_0/vip 0.20fF
C4474 dac_8bit_0/c3m VDD 2.41fF
C4475 vpeak peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 8.94fF
C4476 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp 0.28fF
C4477 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 6.88fF
C4478 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm 0.19fF
C4479 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d 10.82fF
C4480 vlowB vrefB 9.06fF
C4481 low_freq_pll_0/pfd_cp_lpf_0/vQA a_241634_n115151# 0.59fF
C4482 a_223872_n145742# low_freq_pll_0/cs_ring_osc_0/vpbias 0.92fF
C4483 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn vocm_filt 2.07fF
C4484 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp sample_and_hold_1/vholdm 0.86fF
C4485 adc_vcaparrayB dac_8bit_1/vcom_buf 15.10fF
C4486 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d 10.82fF
C4487 a_222040_n127742# VDD 1.55fF
C4488 vpeak_sampled dac_8bit_1/amux_2to1_4/SELB 2.07fF
C4489 vlowA dac_8bit_0/amux_2to1_0/B 1.86fF
C4490 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y a_242951_n122281# 0.17fF
C4491 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VDD 14.23fF
C4492 input_amplifier_0/txgate_2/txb input_amplifier_0/venm2 0.35fF
C4493 a_241919_n122249# a_242783_n122255# 0.09fF
C4494 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 13.66fF
C4495 vcp VDD 5.38fF
C4496 vpeak_sampled sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp 21.50fF
C4497 a_242783_n121345# VDD 0.22fF
C4498 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn biquad_gm_c_filter_0/gm_c_stage_3/vcmcn2 1.28fF
C4499 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc input_amplifier_0/diff_fold_casc_ota_0/vtail_casc 0.01fF
C4500 VDD input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc 8.68fF
C4501 adc_vcaparrayA dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn 2.30fF
C4502 a_226646_n140786# a_228478_n140786# 0.24fF
C4503 a_227104_n140786# a_228020_n140786# 1.33fF
C4504 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 28.76fF
C4505 dac_8bit_1/latched_comparator_folded_0/vcompm_buf dac_8bit_1/comp_outm 0.12fF
C4506 vampp input_amplifier_0/diff_fold_casc_ota_1/vcascnm 11.77fF
C4507 VDD a_244783_n122799# 0.43fF
C4508 a_335844_n185460# a_336116_n185555# 0.67fF
C4509 a_242783_n123343# a_241919_n123337# 0.09fF
C4510 diff_to_se_converter_0/vim vfiltp 4.38fF
C4511 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/csinvp low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin 0.10fF
C4512 a_244783_n123337# a_245056_n123343# 0.38fF
C4513 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y a_246080_n122477# 0.11fF
C4514 a_241919_n121161# a_242085_n121711# 0.09fF
C4515 low_freq_pll_0/pfd_cp_lpf_0/VQBb low_freq_pll_0/pfd_cp_lpf_0/vRSTN 0.20fF
C4516 biquad_gm_c_filter_0/ibiasn3 vfiltp 0.36fF
C4517 vhpf VSS 14.51fF
C4518 m1_326207_n110098# VSS 0.11fF $ **FLOATING
C4519 m1_326207_n59088# VSS 0.11fF $ **FLOATING
C4520 a_338703_n185409# VSS 0.20fF
C4521 a_338505_n185421# VSS 0.01fF
C4522 a_338084_n185421# VSS 0.01fF
C4523 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_2/Q VSS 0.14fF
C4524 a_336955_n185409# VSS 0.20fF
C4525 a_336757_n185421# VSS 0.01fF
C4526 a_336336_n185421# VSS 0.01fF
C4527 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/Q_N VSS 0.40fF
C4528 a_338285_n185409# VSS 0.61fF
C4529 a_338356_n185510# VSS 0.49fF
C4530 a_338156_n185665# VSS 1.18fF
C4531 a_338149_n185569# VSS 1.57fF
C4532 a_337864_n185555# VSS 0.60fF
C4533 a_337592_n185460# VSS 0.28fF
C4534 a_337497_n185813# VSS 0.48fF
C4535 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_3/D VSS 1.22fF
C4536 a_336537_n185409# VSS 0.61fF
C4537 a_336608_n185510# VSS 0.49fF
C4538 a_336408_n185665# VSS 1.17fF
C4539 a_336401_n185569# VSS 1.52fF
C4540 a_336116_n185555# VSS 0.60fF
C4541 a_335844_n185460# VSS 0.28fF
C4542 a_335749_n185813# VSS 0.49fF
C4543 a_338505_n185243# VSS 0.01fF
C4544 a_338084_n185243# VSS 0.01fF
C4545 a_338703_n185243# VSS 0.20fF
C4546 a_336757_n185243# VSS 0.01fF
C4547 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_0/Q_N VSS 0.17fF
C4548 a_336336_n185243# VSS 0.01fF
C4549 pulse_generator_0/sky130_fd_sc_hd__inv_1_0/Y VSS 1.25fF
C4550 a_338285_n185243# VSS 0.61fF
C4551 a_338356_n185269# VSS 0.49fF
C4552 a_338149_n185269# VSS 1.53fF
C4553 a_338156_n184969# VSS 1.18fF
C4554 a_337864_n185269# VSS 0.60fF
C4555 a_337592_n185269# VSS 0.32fF
C4556 a_337497_n185269# VSS 0.31fF
C4557 a_336955_n185243# VSS 0.20fF
C4558 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/Q_N VSS 0.17fF
C4559 pulse_generator_0/sky130_fd_sc_hd__dfxbp_1_1/D VSS 1.43fF
C4560 a_336537_n185243# VSS 0.61fF
C4561 a_336608_n185269# VSS 0.49fF
C4562 a_336401_n185269# VSS 1.52fF
C4563 a_336408_n184969# VSS 1.17fF
C4564 a_336116_n185269# VSS 0.60fF
C4565 a_335844_n185269# VSS 0.32fF
C4566 a_335749_n185269# VSS 0.31fF
C4567 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/A VSS 0.43fF
C4568 pulse_generator_0/sky130_fd_sc_hd__nand2_1_0/B VSS 0.36fF
C4569 pulse_generator_0/sky130_fd_sc_hd__inv_1_1/A VSS 0.31fF
C4570 q0B VSS 0.37fF
C4571 dac_8bit_1/amux_2to1_9/SELB VSS 5.39fF
C4572 q1B VSS 0.37fF
C4573 dac_8bit_1/amux_2to1_10/SELB VSS 5.39fF
C4574 dac_8bit_1/amux_2to1_11/SELB VSS 7.75fF
C4575 q2B VSS 15.35fF
C4576 dac_8bit_1/amux_2to1_12/SELB VSS 5.39fF
C4577 q3B VSS 0.23fF
C4578 dac_8bit_1/amux_2to1_13/SELB VSS 5.39fF
C4579 q4B VSS 0.37fF
C4580 dac_8bit_1/amux_2to1_14/SELB VSS 5.39fF
C4581 q5B VSS 0.36fF
C4582 dac_8bit_1/amux_2to1_15/SELB VSS 5.39fF
C4583 q6B VSS 0.36fF
C4584 dac_8bit_1/amux_2to1_16/SELB VSS 5.39fF
C4585 vrefB VSS 23.40fF
C4586 q7B VSS 0.36fF
C4587 dac_8bit_1/amux_2to1_17/SELB VSS 5.39fF
C4588 dac_8bit_1/amux_2to1_9/Y VSS 10.41fF
C4589 dac_8bit_1/c0m VSS 17.82fF
C4590 dac_8bit_1/amux_2to1_8/SELB VSS 0.26fF
C4591 dac_8bit_1/amux_2to1_7/B VSS 10.41fF
C4592 dac_8bit_1/c1m VSS 18.04fF
C4593 dac_8bit_1/amux_2to1_7/SELB VSS 0.26fF
C4594 dac_8bit_1/amux_2to1_6/B VSS 12.68fF
C4595 dac_8bit_1/cdumm VSS 14.46fF
C4596 dac_8bit_1/amux_2to1_6/SELB VSS 0.17fF
C4597 dac_8bit_1/amux_2to1_5/B VSS 10.41fF
C4598 dac_8bit_1/c2m VSS 32.51fF
C4599 dac_8bit_1/amux_2to1_5/SELB VSS 5.39fF
C4600 dac_8bit_1/amux_2to1_4/B VSS 10.41fF
C4601 dac_8bit_1/c3m VSS 27.21fF
C4602 dac_8bit_1/amux_2to1_4/SELB VSS 0.35fF
C4603 dac_8bit_1/amux_2to1_3/B VSS 10.41fF
C4604 dac_8bit_1/c4m VSS 50.08fF
C4605 dac_8bit_1/amux_2to1_3/SELB VSS 0.35fF
C4606 dac_8bit_1/amux_2to1_2/B VSS 10.41fF
C4607 dac_8bit_1/c5m VSS 81.69fF
C4608 dac_8bit_1/amux_2to1_2/SELB VSS 0.26fF
C4609 dac_8bit_1/amux_2to1_1/B VSS 10.41fF
C4610 dac_8bit_1/c6m VSS 158.36fF
C4611 dac_8bit_1/amux_2to1_1/SELB VSS 0.26fF
C4612 dac_8bit_1/amux_2to1_0/B VSS 10.41fF
C4613 dac_8bit_1/c7m VSS 309.11fF
C4614 dac_8bit_1/amux_2to1_0/SELB VSS 0.26fF
C4615 a_275374_n180872# VSS 36.23fF
C4616 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS 304.65fF
C4617 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS 66.29fF
C4618 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS 132.57fF
C4619 a_230446_n180872# VSS 36.23fF
C4620 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias4 VSS 304.65fF
C4621 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascn VSS 66.29fF
C4622 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias3 VSS 132.57fF
C4623 peak_detector_rst VSS 78.50fF
C4624 a_189446_n180872# VSS 36.23fF
C4625 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS 304.65fF
C4626 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS 66.29fF
C4627 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS 132.57fF
C4628 a_356329_n164260# VSS 36.23fF
C4629 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias4 VSS 304.65fF
C4630 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS 66.29fF
C4631 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias3 VSS 132.57fF
C4632 dac_8bit_1/adc_run VSS 2.54fF
C4633 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M8d VSS 74.42fF
C4634 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS 141.20fF
C4635 sample_and_hold_1/vholdm VSS 75.34fF
C4636 sample_and_hold_1/vhold VSS 111.78fF
C4637 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS 83.16fF
C4638 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS 90.33fF
C4639 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS 48.55fF
C4640 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vmirror VSS 97.87fF
C4641 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS 41.82fF
C4642 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M13d VSS 17.52fF
C4643 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VSS 12.44fF
C4644 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M9d VSS 29.04fF
C4645 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS 138.72fF
C4646 sample_and_hold_1/se_fold_casc_wide_swing_ota_0/M7d VSS 26.00fF
C4647 peak_detector_0/se_fold_casc_wide_swing_ota_1/M16d VSS 11.42fF
C4648 peak_detector_0/se_fold_casc_wide_swing_ota_1/M8d VSS 74.42fF
C4649 peak_detector_0/verr VSS 584.68fF
C4650 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnp VSS 141.20fF
C4651 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascnm VSS 83.16fF
C4652 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias2 VSS 90.33fF
C4653 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpm VSS 48.55fF
C4654 peak_detector_0/se_fold_casc_wide_swing_ota_1/vmirror VSS 97.87fF
C4655 peak_detector_0/se_fold_casc_wide_swing_ota_1/vcascpp VSS 41.82fF
C4656 peak_detector_0/se_fold_casc_wide_swing_ota_1/M13d VSS 17.52fF
C4657 peak_detector_0/se_fold_casc_wide_swing_ota_1/vtail_cascp VSS 12.44fF
C4658 peak_detector_0/se_fold_casc_wide_swing_ota_1/M9d VSS 29.04fF
C4659 peak_detector_0/se_fold_casc_wide_swing_ota_1/vbias1 VSS 138.72fF
C4660 peak_detector_0/se_fold_casc_wide_swing_ota_1/M7d VSS 26.00fF
C4661 peak_detector_0/se_fold_casc_wide_swing_ota_0/M16d VSS 11.42fF
C4662 peak_detector_0/se_fold_casc_wide_swing_ota_0/M8d VSS 74.42fF
C4663 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS 141.20fF
C4664 vpeak VSS 729.19fF
C4665 peak_detector_0/vpeak VSS 570.00fF
C4666 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS 83.14fF
C4667 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS 90.33fF
C4668 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS 48.55fF
C4669 peak_detector_0/se_fold_casc_wide_swing_ota_0/vmirror VSS 97.87fF
C4670 peak_detector_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS 41.82fF
C4671 peak_detector_0/se_fold_casc_wide_swing_ota_0/M13d VSS 17.52fF
C4672 peak_detector_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VSS 12.44fF
C4673 peak_detector_0/se_fold_casc_wide_swing_ota_0/M9d VSS 29.04fF
C4674 peak_detector_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS 138.72fF
C4675 peak_detector_0/se_fold_casc_wide_swing_ota_0/M7d VSS 26.00fF
C4676 dac_8bit_1/latched_comparator_folded_0/vcomppb VSS 0.02fF
C4677 dac_8bit_1/latched_comparator_folded_0/vcompp_buf VSS 0.02fF
C4678 adc_compB VSS 0.14fF
C4679 dac_8bit_1/comp_outm VSS 0.02fF
C4680 dac_8bit_1/latched_comparator_folded_0/vcompm_buf VSS 0.04fF
C4681 dac_8bit_1/latched_comparator_folded_0/vcompmb VSS 0.80fF
C4682 dac_8bit_1/latched_comparator_folded_0/vcompp VSS 6.15fF
C4683 dac_8bit_1/latched_comparator_folded_0/vcompm VSS 5.03fF
C4684 dac_8bit_1/latched_comparator_folded_0/vlatchm VSS 9.90fF
C4685 dac_8bit_1/latched_comparator_folded_0/vlatchp VSS 10.61fF
C4686 vlowB VSS 102.09fF
C4687 dac_8bit_1/latched_comparator_folded_0/vtailp VSS 3.95fF
C4688 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M16d VSS 11.42fF
C4689 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M8d VSS 74.42fF
C4690 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnp VSS 141.20fF
C4691 dac_8bit_1/vcom_buf VSS 619.35fF
C4692 adc_vcaparrayB VSS 428.24fF
C4693 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascnm VSS 83.16fF
C4694 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias2 VSS 90.33fF
C4695 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpm VSS 48.55fF
C4696 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vmirror VSS 97.87fF
C4697 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vcascpp VSS 41.82fF
C4698 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M13d VSS 17.52fF
C4699 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vtail_cascp VSS 12.44fF
C4700 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M9d VSS 29.04fF
C4701 dac_8bit_1/se_fold_casc_wide_swing_ota_0/vbias1 VSS 138.72fF
C4702 dac_8bit_1/se_fold_casc_wide_swing_ota_0/M7d VSS 26.00fF
C4703 a_275374_n146348# VSS 36.23fF
C4704 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS 304.65fF
C4705 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS 67.50fF
C4706 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS 132.57fF
C4707 a_238770_n150168# VSS 0.03fF
C4708 a_238312_n150168# VSS 0.03fF
C4709 a_237854_n150168# VSS 0.03fF
C4710 a_237396_n150168# VSS 0.03fF
C4711 a_236938_n150168# VSS 0.03fF
C4712 a_236480_n150168# VSS 0.03fF
C4713 a_236022_n150168# VSS 0.03fF
C4714 a_243770_n149500# VSS 0.03fF
C4715 a_243312_n149500# VSS 0.03fF
C4716 a_242854_n149500# VSS 0.03fF
C4717 a_242396_n149500# VSS 0.03fF
C4718 a_241938_n149500# VSS 0.03fF
C4719 a_241480_n149500# VSS 0.03fF
C4720 a_241022_n149500# VSS 0.03fF
C4721 a_238770_n149500# VSS 0.03fF
C4722 a_238312_n149500# VSS 0.03fF
C4723 a_237854_n149500# VSS 0.03fF
C4724 a_237396_n149500# VSS 0.03fF
C4725 a_236938_n149500# VSS 0.03fF
C4726 a_236480_n149500# VSS 0.03fF
C4727 a_236022_n149500# VSS 0.03fF
C4728 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/csinvn VSS 0.46fF
C4729 a_223770_n150168# VSS 0.03fF
C4730 a_223312_n150168# VSS 0.03fF
C4731 a_222854_n150168# VSS 0.03fF
C4732 a_222396_n150168# VSS 0.03fF
C4733 a_221938_n150168# VSS 0.03fF
C4734 a_221480_n150168# VSS 0.03fF
C4735 a_228770_n149500# VSS 0.03fF
C4736 a_228312_n149500# VSS 0.03fF
C4737 a_227854_n149500# VSS 0.03fF
C4738 a_227396_n149500# VSS 0.03fF
C4739 a_226938_n149500# VSS 0.03fF
C4740 a_226480_n149500# VSS 0.03fF
C4741 a_226022_n149500# VSS 0.03fF
C4742 a_223770_n149500# VSS 0.03fF
C4743 a_223312_n149500# VSS 0.03fF
C4744 a_222854_n149500# VSS 0.03fF
C4745 a_222396_n149500# VSS 0.03fF
C4746 a_221938_n149500# VSS 0.03fF
C4747 a_221480_n149500# VSS 0.03fF
C4748 a_221022_n149500# VSS 0.03fF
C4749 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/csinvn VSS 0.46fF
C4750 a_243771_n148007# VSS 0.03fF
C4751 a_243313_n148007# VSS 0.03fF
C4752 a_242855_n148007# VSS 0.03fF
C4753 a_242397_n148007# VSS 0.03fF
C4754 a_241939_n148007# VSS 0.03fF
C4755 a_241481_n148007# VSS 0.03fF
C4756 a_241023_n148007# VSS 0.03fF
C4757 a_238771_n148007# VSS 0.03fF
C4758 a_238313_n148007# VSS 0.03fF
C4759 a_237855_n148007# VSS 0.03fF
C4760 a_237397_n148007# VSS 0.03fF
C4761 a_236939_n148007# VSS 0.03fF
C4762 a_236481_n148007# VSS 0.03fF
C4763 a_236023_n148007# VSS 0.03fF
C4764 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/voutcs VSS 20.26fF
C4765 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/csinvp VSS 2.10fF
C4766 a_239330_n145742# VSS 0.62fF
C4767 a_238872_n145742# VSS 1.00fF
C4768 a_238414_n145742# VSS 1.48fF
C4769 a_237956_n145742# VSS 1.86fF
C4770 a_237498_n145742# VSS 2.33fF
C4771 a_237040_n145742# VSS 2.71fF
C4772 a_236582_n145742# VSS 3.19fF
C4773 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_3/vin VSS 43.02fF
C4774 a_228771_n148007# VSS 0.03fF
C4775 a_228313_n148007# VSS 0.03fF
C4776 a_227855_n148007# VSS 0.03fF
C4777 a_227397_n148007# VSS 0.03fF
C4778 a_226939_n148007# VSS 0.03fF
C4779 a_226481_n148007# VSS 0.03fF
C4780 a_226023_n148007# VSS 0.03fF
C4781 a_223771_n148007# VSS 0.03fF
C4782 a_223313_n148007# VSS 0.03fF
C4783 a_222855_n148007# VSS 0.03fF
C4784 a_222397_n148007# VSS 0.03fF
C4785 a_221939_n148007# VSS 0.03fF
C4786 a_221481_n148007# VSS 0.03fF
C4787 a_221023_n148007# VSS 0.03fF
C4788 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/voutcs VSS 20.26fF
C4789 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/csinvp VSS 2.10fF
C4790 a_224330_n145742# VSS 0.62fF
C4791 a_223872_n145742# VSS 1.00fF
C4792 a_223414_n145742# VSS 1.48fF
C4793 a_222956_n145742# VSS 1.86fF
C4794 a_222498_n145742# VSS 2.33fF
C4795 a_222040_n145742# VSS 2.71fF
C4796 a_221582_n145742# VSS 3.19fF
C4797 a_243478_n140786# VSS 0.62fF
C4798 a_243020_n140786# VSS 1.00fF
C4799 a_242562_n140786# VSS 1.48fF
C4800 a_242104_n140786# VSS 1.86fF
C4801 a_241646_n140786# VSS 2.33fF
C4802 a_241188_n140786# VSS 2.71fF
C4803 a_240730_n140786# VSS 3.19fF
C4804 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/csinvp VSS 2.10fF
C4805 a_247701_n138121# VSS 0.03fF
C4806 a_247243_n138121# VSS 0.03fF
C4807 a_246785_n138121# VSS 0.03fF
C4808 a_246327_n138121# VSS 0.03fF
C4809 a_245869_n138121# VSS 0.03fF
C4810 a_245411_n138121# VSS 0.03fF
C4811 a_244953_n138121# VSS 0.03fF
C4812 a_242701_n138121# VSS 0.03fF
C4813 a_242243_n138121# VSS 0.03fF
C4814 a_241785_n138121# VSS 0.03fF
C4815 a_241327_n138121# VSS 0.03fF
C4816 a_240869_n138121# VSS 0.03fF
C4817 a_240411_n138121# VSS 0.03fF
C4818 a_239953_n138121# VSS 0.03fF
C4819 a_228478_n140786# VSS 0.62fF
C4820 a_228020_n140786# VSS 1.00fF
C4821 a_227562_n140786# VSS 1.48fF
C4822 a_227104_n140786# VSS 1.86fF
C4823 a_226646_n140786# VSS 2.33fF
C4824 a_226188_n140786# VSS 2.71fF
C4825 a_225730_n140786# VSS 3.19fF
C4826 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/csinvp VSS 2.10fF
C4827 a_232701_n138121# VSS 0.03fF
C4828 a_232243_n138121# VSS 0.03fF
C4829 a_231785_n138121# VSS 0.03fF
C4830 a_231327_n138121# VSS 0.03fF
C4831 a_230869_n138121# VSS 0.03fF
C4832 a_230411_n138121# VSS 0.03fF
C4833 a_229953_n138121# VSS 0.03fF
C4834 a_227701_n138121# VSS 0.03fF
C4835 a_227243_n138121# VSS 0.03fF
C4836 a_226785_n138121# VSS 0.03fF
C4837 a_226327_n138121# VSS 0.03fF
C4838 a_225869_n138121# VSS 0.03fF
C4839 a_225411_n138121# VSS 0.03fF
C4840 a_224953_n138121# VSS 0.03fF
C4841 q0A VSS 0.50fF
C4842 dac_8bit_0/amux_2to1_9/SELB VSS 0.26fF
C4843 q1A VSS 0.50fF
C4844 dac_8bit_0/amux_2to1_10/SELB VSS 0.26fF
C4845 dac_8bit_0/amux_2to1_11/SELB VSS 0.17fF
C4846 q2A VSS 0.43fF
C4847 dac_8bit_0/amux_2to1_12/SELB VSS 5.39fF
C4848 q3A VSS 0.25fF
C4849 dac_8bit_0/amux_2to1_13/SELB VSS 0.35fF
C4850 q4A VSS 0.50fF
C4851 dac_8bit_0/amux_2to1_14/SELB VSS 0.35fF
C4852 q5A VSS 0.49fF
C4853 dac_8bit_0/amux_2to1_15/SELB VSS 0.26fF
C4854 q6A VSS 0.48fF
C4855 dac_8bit_0/amux_2to1_16/SELB VSS 0.26fF
C4856 vrefA VSS 23.46fF
C4857 q7A VSS 0.51fF
C4858 dac_8bit_0/amux_2to1_17/SELB VSS 0.26fF
C4859 dac_8bit_0/amux_2to1_9/Y VSS 10.41fF
C4860 dac_8bit_0/c0m VSS 14.69fF
C4861 dac_8bit_0/amux_2to1_8/SELB VSS 0.26fF
C4862 dac_8bit_0/amux_2to1_7/B VSS 10.41fF
C4863 dac_8bit_0/c1m VSS 17.78fF
C4864 dac_8bit_0/amux_2to1_7/SELB VSS 0.26fF
C4865 dac_8bit_0/amux_2to1_6/B VSS 12.68fF
C4866 dac_8bit_0/cdumm VSS 14.11fF
C4867 dac_8bit_0/amux_2to1_6/SELB VSS 0.17fF
C4868 dac_8bit_0/amux_2to1_5/B VSS 10.41fF
C4869 dac_8bit_0/c2m VSS 31.13fF
C4870 dac_8bit_0/amux_2to1_5/SELB VSS 5.39fF
C4871 dac_8bit_0/amux_2to1_4/B VSS 10.41fF
C4872 dac_8bit_0/c3m VSS 26.95fF
C4873 dac_8bit_0/amux_2to1_4/SELB VSS 0.36fF
C4874 dac_8bit_0/amux_2to1_3/B VSS 10.41fF
C4875 dac_8bit_0/c4m VSS 49.83fF
C4876 dac_8bit_0/amux_2to1_3/SELB VSS 0.36fF
C4877 dac_8bit_0/amux_2to1_2/B VSS 10.41fF
C4878 dac_8bit_0/c5m VSS 81.43fF
C4879 dac_8bit_0/amux_2to1_2/SELB VSS 0.26fF
C4880 dac_8bit_0/amux_2to1_1/B VSS 10.41fF
C4881 dac_8bit_0/c6m VSS 158.09fF
C4882 dac_8bit_0/amux_2to1_1/SELB VSS 0.26fF
C4883 dac_8bit_0/amux_2to1_0/B VSS 10.41fF
C4884 dac_8bit_0/c7m VSS 308.90fF
C4885 dac_8bit_0/amux_2to1_0/SELB VSS 0.26fF
C4886 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M8d VSS 74.42fF
C4887 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS 141.20fF
C4888 sample_and_hold_0/vholdm VSS 75.34fF
C4889 sample_and_hold_0/vhold VSS 111.78fF
C4890 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS 83.16fF
C4891 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS 90.33fF
C4892 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS 48.55fF
C4893 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vmirror VSS 97.87fF
C4894 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS 41.82fF
C4895 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M13d VSS 17.52fF
C4896 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VSS 12.44fF
C4897 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M9d VSS 29.04fF
C4898 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS 138.72fF
C4899 sample_and_hold_0/se_fold_casc_wide_swing_ota_0/M7d VSS 26.00fF
C4900 a_247702_n135628# VSS 0.03fF
C4901 a_247244_n135628# VSS 0.03fF
C4902 a_246786_n135628# VSS 0.03fF
C4903 a_246328_n135628# VSS 0.03fF
C4904 a_245870_n135628# VSS 0.03fF
C4905 a_245412_n135628# VSS 0.03fF
C4906 a_244954_n135628# VSS 0.03fF
C4907 a_242702_n135628# VSS 0.03fF
C4908 a_242244_n135628# VSS 0.03fF
C4909 a_241786_n135628# VSS 0.03fF
C4910 a_241328_n135628# VSS 0.03fF
C4911 a_240870_n135628# VSS 0.03fF
C4912 a_240412_n135628# VSS 0.03fF
C4913 a_239954_n135628# VSS 0.03fF
C4914 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/vin VSS 48.60fF
C4915 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/voutcs VSS 20.26fF
C4916 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_4/csinvn VSS 0.46fF
C4917 a_247702_n134960# VSS 0.03fF
C4918 a_247244_n134960# VSS 0.03fF
C4919 a_246786_n134960# VSS 0.03fF
C4920 a_246328_n134960# VSS 0.03fF
C4921 a_245870_n134960# VSS 0.03fF
C4922 a_245412_n134960# VSS 0.03fF
C4923 a_244954_n134960# VSS 0.03fF
C4924 a_232702_n135628# VSS 0.03fF
C4925 a_232244_n135628# VSS 0.03fF
C4926 a_231786_n135628# VSS 0.03fF
C4927 a_231328_n135628# VSS 0.03fF
C4928 a_230870_n135628# VSS 0.03fF
C4929 a_230412_n135628# VSS 0.03fF
C4930 a_229954_n135628# VSS 0.03fF
C4931 a_227702_n135628# VSS 0.03fF
C4932 a_227244_n135628# VSS 0.03fF
C4933 a_226786_n135628# VSS 0.03fF
C4934 a_226328_n135628# VSS 0.03fF
C4935 a_225870_n135628# VSS 0.03fF
C4936 a_225412_n135628# VSS 0.03fF
C4937 a_224954_n135628# VSS 0.03fF
C4938 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS 48.61fF
C4939 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/voutcs VSS 20.26fF
C4940 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/csinvn VSS 0.46fF
C4941 a_232702_n134960# VSS 0.03fF
C4942 a_232244_n134960# VSS 0.03fF
C4943 a_231786_n134960# VSS 0.03fF
C4944 a_231328_n134960# VSS 0.03fF
C4945 a_230870_n134960# VSS 0.03fF
C4946 a_230412_n134960# VSS 0.03fF
C4947 a_229954_n134960# VSS 0.03fF
C4948 a_162668_n147576# VSS 36.23fF
C4949 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS 66.29fF
C4950 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS 304.65fF
C4951 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS 132.57fF
C4952 diff_to_se_converter_0/txgate_0/txb VSS 2.49fF
C4953 diff_to_se_converter_0/txgate_1/txb VSS 2.50fF
C4954 diff_to_se_converter_0/rst VSS 11.25fF
C4955 a_238770_n132168# VSS 0.03fF
C4956 a_238312_n132168# VSS 0.03fF
C4957 a_237854_n132168# VSS 0.03fF
C4958 a_237396_n132168# VSS 0.03fF
C4959 a_236938_n132168# VSS 0.03fF
C4960 a_236480_n132168# VSS 0.03fF
C4961 a_236022_n132168# VSS 0.03fF
C4962 a_243770_n131500# VSS 0.03fF
C4963 a_243312_n131500# VSS 0.03fF
C4964 a_242854_n131500# VSS 0.03fF
C4965 a_242396_n131500# VSS 0.03fF
C4966 a_241938_n131500# VSS 0.03fF
C4967 a_241480_n131500# VSS 0.03fF
C4968 a_241022_n131500# VSS 0.03fF
C4969 a_238770_n131500# VSS 0.03fF
C4970 a_238312_n131500# VSS 0.03fF
C4971 a_237854_n131500# VSS 0.03fF
C4972 a_237396_n131500# VSS 0.03fF
C4973 a_236938_n131500# VSS 0.03fF
C4974 a_236480_n131500# VSS 0.03fF
C4975 a_236022_n131500# VSS 0.03fF
C4976 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/csinvn VSS 0.46fF
C4977 a_223770_n132168# VSS 0.03fF
C4978 a_223312_n132168# VSS 0.03fF
C4979 a_222854_n132168# VSS 0.03fF
C4980 a_222396_n132168# VSS 0.03fF
C4981 a_221938_n132168# VSS 0.03fF
C4982 a_221480_n132168# VSS 0.03fF
C4983 a_228770_n131500# VSS 0.03fF
C4984 a_228312_n131500# VSS 0.03fF
C4985 a_227854_n131500# VSS 0.03fF
C4986 a_227396_n131500# VSS 0.03fF
C4987 a_226938_n131500# VSS 0.03fF
C4988 a_226480_n131500# VSS 0.03fF
C4989 a_226022_n131500# VSS 0.03fF
C4990 a_223770_n131500# VSS 0.03fF
C4991 a_223312_n131500# VSS 0.03fF
C4992 a_222854_n131500# VSS 0.03fF
C4993 a_222396_n131500# VSS 0.03fF
C4994 a_221938_n131500# VSS 0.03fF
C4995 a_221480_n131500# VSS 0.03fF
C4996 a_221022_n131500# VSS 0.03fF
C4997 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/csinvn VSS 0.46fF
C4998 a_243771_n130007# VSS 0.03fF
C4999 a_243313_n130007# VSS 0.03fF
C5000 a_242855_n130007# VSS 0.03fF
C5001 a_242397_n130007# VSS 0.03fF
C5002 a_241939_n130007# VSS 0.03fF
C5003 a_241481_n130007# VSS 0.03fF
C5004 a_241023_n130007# VSS 0.03fF
C5005 a_238771_n130007# VSS 0.03fF
C5006 a_238313_n130007# VSS 0.03fF
C5007 a_237855_n130007# VSS 0.03fF
C5008 a_237397_n130007# VSS 0.03fF
C5009 a_236939_n130007# VSS 0.03fF
C5010 a_236481_n130007# VSS 0.03fF
C5011 a_236023_n130007# VSS 0.03fF
C5012 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/voutcs VSS 20.26fF
C5013 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS 46.10fF
C5014 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/csinvp VSS 2.10fF
C5015 a_239330_n127742# VSS 0.62fF
C5016 a_238872_n127742# VSS 1.00fF
C5017 a_238414_n127742# VSS 1.48fF
C5018 a_237956_n127742# VSS 1.86fF
C5019 a_237498_n127742# VSS 2.33fF
C5020 a_237040_n127742# VSS 2.71fF
C5021 a_236582_n127742# VSS 3.19fF
C5022 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_1/vin VSS 47.79fF
C5023 a_228771_n130007# VSS 0.03fF
C5024 a_228313_n130007# VSS 0.03fF
C5025 a_227855_n130007# VSS 0.03fF
C5026 a_227397_n130007# VSS 0.03fF
C5027 a_226939_n130007# VSS 0.03fF
C5028 a_226481_n130007# VSS 0.03fF
C5029 a_226023_n130007# VSS 0.03fF
C5030 a_223771_n130007# VSS 0.03fF
C5031 a_223313_n130007# VSS 0.03fF
C5032 a_222855_n130007# VSS 0.03fF
C5033 a_222397_n130007# VSS 0.03fF
C5034 a_221939_n130007# VSS 0.03fF
C5035 a_221481_n130007# VSS 0.03fF
C5036 a_221023_n130007# VSS 0.03fF
C5037 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/voutcs VSS 20.26fF
C5038 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_0/csinvp VSS 2.10fF
C5039 a_224330_n127742# VSS 0.62fF
C5040 a_223872_n127742# VSS 1.00fF
C5041 a_223414_n127742# VSS 1.48fF
C5042 a_222956_n127742# VSS 1.86fF
C5043 a_222498_n127742# VSS 2.33fF
C5044 a_222040_n127742# VSS 2.71fF
C5045 a_221582_n127742# VSS 3.19fF
C5046 a_245607_n122965# VSS 0.01fF
C5047 a_245182_n122965# VSS 0.01fF
C5048 a_244971_n123343# VSS 0.20fF
C5049 a_242909_n122965# VSS 0.01fF
C5050 a_242484_n122965# VSS 0.01fF
C5051 a_242273_n123343# VSS 0.20fF
C5052 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/A VSS 0.77fF
C5053 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_10/A VSS 0.41fF
C5054 a_246080_n123343# VSS 0.31fF
C5055 a_245481_n123343# VSS 0.60fF
C5056 a_245649_n123369# VSS 1.13fF
C5057 a_245056_n123343# VSS 0.49fF
C5058 a_245224_n123369# VSS 0.61fF
C5059 a_244783_n123337# VSS 0.16fF
C5060 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_10/Y VSS 0.25fF
C5061 a_244617_n123337# VSS 0.34fF
C5062 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q VSS 0.74fF
C5063 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/A VSS 0.52fF
C5064 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_5/A VSS 0.41fF
C5065 a_243382_n123343# VSS 0.31fF
C5066 a_242783_n123343# VSS 0.60fF
C5067 a_242951_n123369# VSS 1.13fF
C5068 a_242358_n123343# VSS 0.49fF
C5069 a_242526_n123369# VSS 0.61fF
C5070 a_242085_n123337# VSS 0.16fF
C5071 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_5/Y VSS 0.25fF
C5072 a_241919_n123337# VSS 0.34fF
C5073 a_245607_n122799# VSS 0.01fF
C5074 a_245182_n122799# VSS 0.01fF
C5075 a_242909_n122799# VSS 0.01fF
C5076 a_244971_n122799# VSS 0.20fF
C5077 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/A VSS 0.04fF
C5078 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_9/A VSS 0.04fF
C5079 a_246080_n122477# VSS 0.24fF
C5080 a_245481_n122433# VSS 0.60fF
C5081 a_245649_n122531# VSS 1.13fF
C5082 a_245056_n122433# VSS 0.49fF
C5083 a_245224_n122687# VSS 0.61fF
C5084 a_244783_n122799# VSS 0.03fF
C5085 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_9/Y VSS 0.20fF
C5086 a_244617_n122799# VSS 0.02fF
C5087 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q VSS 0.26fF
C5088 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q VSS 0.40fF
C5089 a_242484_n122799# VSS 0.01fF
C5090 a_242273_n122799# VSS 0.20fF
C5091 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/A VSS 0.04fF
C5092 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_4/A VSS 0.04fF
C5093 a_243382_n122477# VSS 0.24fF
C5094 a_242783_n122433# VSS 0.60fF
C5095 a_242951_n122531# VSS 1.13fF
C5096 a_242358_n122433# VSS 0.49fF
C5097 a_242526_n122687# VSS 0.61fF
C5098 a_242085_n122799# VSS 1.17fF
C5099 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_4/Y VSS 0.19fF
C5100 a_241919_n122799# VSS 1.52fF
C5101 a_245607_n121877# VSS 0.01fF
C5102 a_245182_n121877# VSS 0.01fF
C5103 a_244971_n122255# VSS 0.20fF
C5104 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q VSS 0.43fF
C5105 a_242909_n121877# VSS 0.01fF
C5106 a_242484_n121877# VSS 0.01fF
C5107 a_242273_n122255# VSS 0.20fF
C5108 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/A VSS 0.77fF
C5109 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_8/A VSS 0.41fF
C5110 a_246080_n122255# VSS 0.31fF
C5111 a_245481_n122255# VSS 0.60fF
C5112 a_245649_n122281# VSS 1.13fF
C5113 a_245056_n122255# VSS 0.49fF
C5114 a_245224_n122281# VSS 0.61fF
C5115 a_244783_n122249# VSS 0.16fF
C5116 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_8/Y VSS 0.25fF
C5117 a_244617_n122249# VSS 0.34fF
C5118 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q VSS 0.30fF
C5119 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/A VSS 0.52fF
C5120 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_2/A VSS 0.41fF
C5121 a_243382_n122255# VSS 0.31fF
C5122 a_242783_n122255# VSS 0.60fF
C5123 a_242951_n122281# VSS 1.13fF
C5124 a_242358_n122255# VSS 0.49fF
C5125 a_242526_n122281# VSS 0.61fF
C5126 a_242085_n122249# VSS 0.16fF
C5127 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_2/Y VSS 0.25fF
C5128 a_241919_n122249# VSS 0.34fF
C5129 a_245607_n121711# VSS 0.01fF
C5130 a_245182_n121711# VSS 0.01fF
C5131 a_242909_n121711# VSS 0.01fF
C5132 a_244971_n121711# VSS 0.20fF
C5133 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/A VSS 0.67fF
C5134 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_7/A VSS 0.36fF
C5135 a_246080_n121389# VSS 0.49fF
C5136 a_245481_n121345# VSS 0.60fF
C5137 a_245649_n121443# VSS 1.13fF
C5138 a_245056_n121345# VSS 0.49fF
C5139 a_245224_n121599# VSS 0.61fF
C5140 a_244783_n121711# VSS 0.14fF
C5141 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_7/Y VSS 0.24fF
C5142 a_244617_n121711# VSS 0.25fF
C5143 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q VSS 0.27fF
C5144 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q VSS 0.30fF
C5145 a_242484_n121711# VSS 0.01fF
C5146 a_242273_n121711# VSS 0.20fF
C5147 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/A VSS 0.47fF
C5148 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_3/A VSS 0.36fF
C5149 a_243382_n121389# VSS 0.49fF
C5150 a_242783_n121345# VSS 0.60fF
C5151 a_242951_n121443# VSS 1.13fF
C5152 a_242358_n121345# VSS 0.49fF
C5153 a_242526_n121599# VSS 0.61fF
C5154 a_242085_n121711# VSS 0.08fF
C5155 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_3/Y VSS 1.30fF
C5156 a_241919_n121711# VSS 0.19fF
C5157 a_245607_n120789# VSS 0.01fF
C5158 a_245182_n120789# VSS 0.01fF
C5159 a_244971_n121167# VSS 0.20fF
C5160 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q VSS 0.21fF
C5161 a_242909_n120789# VSS 0.01fF
C5162 a_242484_n120789# VSS 0.01fF
C5163 a_242273_n121167# VSS 0.20fF
C5164 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/A VSS 0.77fF
C5165 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_6/A VSS 0.41fF
C5166 a_246080_n121167# VSS 0.31fF
C5167 a_245481_n121167# VSS 0.60fF
C5168 a_245649_n121193# VSS 1.13fF
C5169 a_245056_n121167# VSS 0.49fF
C5170 a_245224_n121193# VSS 0.61fF
C5171 a_244783_n121161# VSS 0.16fF
C5172 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_6/Y VSS 0.25fF
C5173 a_244617_n121161# VSS 0.34fF
C5174 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q VSS 0.39fF
C5175 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/A VSS 0.52fF
C5176 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_1/A VSS 0.41fF
C5177 a_243382_n121167# VSS 0.31fF
C5178 a_242783_n121167# VSS 0.60fF
C5179 a_242951_n121193# VSS 1.13fF
C5180 a_242358_n121167# VSS 0.49fF
C5181 a_242526_n121193# VSS 0.61fF
C5182 a_242085_n121161# VSS 0.16fF
C5183 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_1/Y VSS 0.25fF
C5184 a_241919_n121161# VSS 0.34fF
C5185 a_242909_n120623# VSS 0.01fF
C5186 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q VSS 0.30fF
C5187 a_242484_n120623# VSS 0.01fF
C5188 a_238923_n122049# VSS 0.03fF
C5189 a_238465_n122049# VSS 0.03fF
C5190 a_238007_n122049# VSS 0.03fF
C5191 a_237549_n122049# VSS 0.03fF
C5192 a_237091_n122049# VSS 0.03fF
C5193 a_236633_n122049# VSS 0.03fF
C5194 a_236175_n122049# VSS 0.03fF
C5195 a_228328_n122869# VSS 0.62fF
C5196 a_227870_n122869# VSS 1.00fF
C5197 a_227412_n122869# VSS 1.48fF
C5198 a_226954_n122869# VSS 1.86fF
C5199 a_226496_n122869# VSS 2.33fF
C5200 a_226038_n122869# VSS 2.70fF
C5201 a_225580_n122869# VSS 3.19fF
C5202 a_242273_n120623# VSS 0.20fF
C5203 low_freq_pll_0/cs_ring_osc_0/vosc2 VSS 0.87fF
C5204 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/A VSS 0.52fF
C5205 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_1_0/A VSS 0.41fF
C5206 a_243382_n120301# VSS 0.31fF
C5207 a_242783_n120257# VSS 0.60fF
C5208 a_242951_n120355# VSS 1.13fF
C5209 a_242358_n120257# VSS 0.49fF
C5210 a_242526_n120511# VSS 0.61fF
C5211 a_242085_n120623# VSS 0.16fF
C5212 low_freq_pll_0/freq_div_0/sky130_fd_sc_hd__inv_4_0/Y VSS 0.25fF
C5213 a_241919_n120623# VSS 0.34fF
C5214 low_freq_pll_0/freq_div_0/vin VSS 0.24fF
C5215 low_freq_pll_0/cs_ring_osc_0/vosc VSS 32.85fF
C5216 a_238922_n119618# VSS 0.03fF
C5217 a_238464_n119618# VSS 0.03fF
C5218 a_238006_n119618# VSS 0.03fF
C5219 a_237548_n119618# VSS 0.03fF
C5220 a_237090_n119618# VSS 0.03fF
C5221 a_236632_n119618# VSS 0.03fF
C5222 a_236174_n119618# VSS 0.03fF
C5223 low_freq_pll_0/cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS 48.36fF
C5224 a_230160_n119618# VSS 0.03fF
C5225 a_229702_n119618# VSS 0.03fF
C5226 a_229244_n119618# VSS 0.03fF
C5227 a_228786_n119618# VSS 0.03fF
C5228 a_228328_n119618# VSS 0.03fF
C5229 a_227870_n119618# VSS 0.03fF
C5230 a_227412_n119618# VSS 0.03fF
C5231 low_freq_pll_0/cs_ring_osc_0/vpbias VSS 128.39fF
C5232 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M16d VSS 11.42fF
C5233 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS 83.16fF
C5234 diff_to_se_converter_0/vip VSS 68.00fF
C5235 diff_to_se_converter_0/vim VSS 77.24fF
C5236 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS 141.20fF
C5237 vse VSS 658.66fF
C5238 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M8d VSS 74.42fF
C5239 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS 90.33fF
C5240 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS 48.55fF
C5241 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vmirror VSS 97.87fF
C5242 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS 41.82fF
C5243 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M13d VSS 17.52fF
C5244 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VSS 12.44fF
C5245 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M7d VSS 26.00fF
C5246 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS 138.72fF
C5247 diff_to_se_converter_0/se_fold_casc_wide_swing_ota_0/M9d VSS 29.04fF
C5248 a_356329_n113250# VSS 36.23fF
C5249 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias4 VSS 304.65fF
C5250 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascn VSS 66.29fF
C5251 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias3 VSS 132.57fF
C5252 sample VSS 294.58fF
C5253 dac_8bit_0/adc_run VSS 2.54fF
C5254 a_242885_n115125# VSS -0.03fF
C5255 a_242377_n115125# VSS -0.01fF
C5256 a_243138_n114759# VSS 0.08fF
C5257 a_242720_n114759# VSS -0.03fF
C5258 a_240062_n115125# VSS -0.01fF
C5259 a_239817_n115125# VSS -0.01fF
C5260 low_freq_pll_0/pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/Q_N VSS 0.16fF
C5261 low_freq_pll_0/pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/Q_N VSS 0.16fF
C5262 low_freq_pll_0/pfd_cp_lpf_0/VQBb VSS 4.27fF
C5263 low_freq_pll_0/pfd_cp_lpf_0/vswitchl VSS 0.15fF
C5264 a_239251_n114759# VSS 0.09fF
C5265 a_239048_n115125# VSS 0.08fF
C5266 a_242506_n114759# VSS -0.38fF
C5267 a_242575_n114888# VSS -0.26fF
C5268 a_242419_n114983# VSS -0.90fF
C5269 a_242380_n114857# VSS -0.63fF
C5270 a_242102_n114873# VSS 0.47fF
C5271 a_241731_n115151# VSS 1.03fF
C5272 a_241634_n115151# VSS 0.30fF
C5273 low_freq_pll_0/pfd_cp_lpf_0/vQB VSS 0.29fF
C5274 a_240447_n115125# VSS 0.30fF
C5275 a_239708_n115125# VSS -0.40fF
C5276 a_239883_n115151# VSS -0.42fF
C5277 a_239143_n115125# VSS 0.46fF
C5278 low_freq_pll_0/pfd_cp_lpf_0/vRSTN VSS 0.15fF
C5279 a_239361_n114883# VSS 0.40fF
C5280 a_238793_n115125# VSS 0.98fF
C5281 a_238627_n115125# VSS 1.19fF
C5282 low_freq_pll_0/freq_div_0/vout VSS 0.45fF
C5283 low_freq_pll_0/pfd_cp_lpf_0/vndiode VSS 1.36fF
C5284 low_freq_pll_0/pfd_cp_lpf_0/vpdiode VSS 0.90fF
C5285 low_freq_pll_0/pfd_cp_lpf_0/vQA VSS 2.66fF
C5286 vcp VSS 0.74fF
C5287 low_freq_pll_0/pfd_cp_lpf_0/vQAb VSS 2.62fF
C5288 comparator_0/vtail VSS 12.57fF
C5289 low_freq_pll_0/pfd_cp_lpf_0/vswitchh VSS 7.07fF
C5290 low_freq_pll_0/pfd_cp_lpf_0/vpbias VSS 24.46fF
C5291 vcomp VSS 0.81fF
C5292 comparator_0/vo1 VSS 7.36fF
C5293 comparator_0/vmirror VSS 5.68fF
C5294 comparator_0/vcompm VSS 10.90fF
C5295 comparator_0/vcompp VSS 11.89fF
C5296 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn2 VSS 3.23fF
C5297 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn1 VSS 0.09fF
C5298 biquad_gm_c_filter_0/gm_c_stage_3/vcmcn VSS 10.01fF
C5299 biquad_gm_c_filter_0/gm_c_stage_3/vbiasp VSS 5.02fF
C5300 biquad_gm_c_filter_0/gm_c_stage_3/vtail_diff VSS 3.39fF
C5301 biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail2 VSS 0.10fF
C5302 biquad_gm_c_filter_0/gm_c_stage_3/vcmn_tail1 VSS 10.52fF
C5303 biquad_gm_c_filter_0/gm_c_stage_3/vcmc VSS 6.85fF
C5304 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn2 VSS 3.23fF
C5305 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn1 VSS 0.15fF
C5306 biquad_gm_c_filter_0/gm_c_stage_1/vcmcn VSS 10.01fF
C5307 biquad_gm_c_filter_0/gm_c_stage_1/vbiasp VSS 5.02fF
C5308 biquad_gm_c_filter_0/gm_c_stage_1/vtail_diff VSS 3.39fF
C5309 biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail2 VSS 0.65fF
C5310 biquad_gm_c_filter_0/gm_c_stage_1/vcmn_tail1 VSS 0.69fF
C5311 biquad_gm_c_filter_0/gm_c_stage_1/vcmc VSS 6.85fF
C5312 biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail2 VSS 0.10fF
C5313 biquad_gm_c_filter_0/gm_c_stage_2/vtail_diff VSS 3.39fF
C5314 biquad_gm_c_filter_0/gm_c_stage_2/vcmn_tail1 VSS 10.52fF
C5315 vfiltm VSS 64.38fF
C5316 vfiltp VSS 63.22fF
C5317 biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail2 VSS 0.10fF
C5318 biquad_gm_c_filter_0/gm_c_stage_0/vtail_diff VSS 3.39fF
C5319 biquad_gm_c_filter_0/gm_c_stage_0/vcmn_tail1 VSS 0.10fF
C5320 vocm_filt VSS 0.87fF
C5321 dac_8bit_1/ibiasp VSS 80.87fF
C5322 vbiasn VSS 9.59fF
C5323 biquad_gm_c_filter_0/gm_c_stage_2/vcmc VSS 6.85fF
C5324 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn2 VSS 3.23fF
C5325 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn1 VSS 0.44fF
C5326 biquad_gm_c_filter_0/gm_c_stage_2/vcmcn VSS 10.01fF
C5327 biquad_gm_c_filter_0/gm_c_stage_2/vbiasp VSS 5.02fF
C5328 biquad_gm_c_filter_0/gm_c_stage_0/vcmc VSS 6.85fF
C5329 vintm VSS 37.79fF
C5330 vintp VSS 36.94fF
C5331 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn2 VSS 3.23fF
C5332 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn1 VSS 0.15fF
C5333 biquad_gm_c_filter_0/gm_c_stage_0/vcmcn VSS 10.01fF
C5334 biquad_gm_c_filter_0/gm_c_stage_0/vbiasp VSS 5.02fF
C5335 dac_8bit_0/latched_comparator_folded_0/vcomppb VSS 0.43fF
C5336 dac_8bit_0/latched_comparator_folded_0/vcompp_buf VSS 0.44fF
C5337 adc_compA VSS 0.45fF
C5338 dac_8bit_0/comp_outm VSS 0.30fF
C5339 dac_8bit_0/latched_comparator_folded_0/vcompm_buf VSS 0.44fF
C5340 dac_8bit_0/latched_comparator_folded_0/vcompmb VSS 0.28fF
C5341 adc_clk VSS 90.49fF
C5342 dac_8bit_0/latched_comparator_folded_0/vcompp VSS 6.15fF
C5343 dac_8bit_0/latched_comparator_folded_0/vcompm VSS 5.03fF
C5344 dac_8bit_0/latched_comparator_folded_0/vlatchm VSS 9.90fF
C5345 dac_8bit_0/latched_comparator_folded_0/vlatchp VSS 10.61fF
C5346 vlowA VSS 102.43fF
C5347 dac_8bit_0/ibiasp VSS 75.23fF
C5348 dac_8bit_0/latched_comparator_folded_0/vtailp VSS 3.95fF
C5349 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M16d VSS 11.42fF
C5350 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M8d VSS 74.42fF
C5351 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnp VSS 141.20fF
C5352 dac_8bit_0/vcom_buf VSS 619.37fF
C5353 adc_vcaparrayA VSS 436.43fF
C5354 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascnm VSS 83.16fF
C5355 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias2 VSS 90.33fF
C5356 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpm VSS 48.55fF
C5357 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vmirror VSS 97.87fF
C5358 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vcascpp VSS 41.82fF
C5359 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M13d VSS 17.52fF
C5360 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vtail_cascp VSS 12.44fF
C5361 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M9d VSS 29.04fF
C5362 dac_8bit_0/se_fold_casc_wide_swing_ota_0/vbias1 VSS 138.72fF
C5363 dac_8bit_0/se_fold_casc_wide_swing_ota_0/M7d VSS 26.00fF
C5364 dac_8bit_1/ibiasn VSS 77.26fF
C5365 vpeak_sampled VSS 723.79fF
C5366 dac_8bit_0/ibiasn VSS 61.12fF
C5367 vcp_sampled VSS 713.74fF
C5368 peak_detector_0/ibiasn2 VSS 96.88fF
C5369 peak_detector_0/ibiasn1 VSS 74.75fF
C5370 diff_to_se_converter_0/ibiasn VSS 77.04fF
C5371 comparator_0/ibiasn VSS 47.65fF
C5372 biquad_gm_c_filter_0/ibiasn1 VSS 64.24fF
C5373 biquad_gm_c_filter_0/ibiasn2 VSS 69.86fF
C5374 biquad_gm_c_filter_0/ibiasn3 VSS 60.28fF
C5375 biquad_gm_c_filter_0/ibiasn4 VSS 56.07fF
C5376 low_freq_pll_0/ibiasn VSS 43.21fF
C5377 vbiasp VSS 73.17fF
C5378 input_amplifier_0/ibiasn1 VSS 55.37fF
C5379 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail1 VSS 9.65fF
C5380 input_amplifier_0/diff_fold_casc_ota_0/vcmn_casc_tail2 VSS 14.09fF
C5381 a_217060_n102324# VSS 35.46fF
C5382 input_amplifier_0/diff_fold_casc_ota_0/vcascnp VSS 40.40fF
C5383 input_amplifier_0/diff_fold_casc_ota_0/vcascnm VSS 45.20fF
C5384 input_amplifier_0/diff_fold_casc_ota_0/vtail_casc VSS 47.41fF
C5385 input_amplifier_0/diff_fold_casc_ota_0/vbias4 VSS 214.47fF
C5386 input_amplifier_0/diff_fold_casc_ota_0/vbias3 VSS 140.70fF
C5387 input_amplifier_0/txgate_6/txb VSS 0.42fF
C5388 input_amplifier_0/venp1 VSS 7.64fF
C5389 input_amplifier_0/txgate_1/txb VSS 2.60fF
C5390 input_amplifier_0/venm1 VSS 7.64fF
C5391 input_amplifier_0/txgate_0/txb VSS 0.42fF
C5392 gain_ctrl_0 VSS 10.39fF
C5393 input_amplifier_0/txgate_7/txb VSS 0.18fF
C5394 input_amplifier_0/ibiasn2 VSS 78.84fF
C5395 input_amplifier_0/vip2 VSS 69.56fF
C5396 input_amplifier_0/vim2 VSS 68.82fF
C5397 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail1 VSS 0.44fF
C5398 input_amplifier_0/diff_fold_casc_ota_1/vcmn_casc_tail2 VSS 0.09fF
C5399 vocm VSS 0.78fF
C5400 a_163060_n102324# VSS 35.46fF
C5401 input_amplifier_0/diff_fold_casc_ota_1/vcascnp VSS 40.40fF
C5402 input_amplifier_0/diff_fold_casc_ota_1/vcascnm VSS 45.20fF
C5403 input_amplifier_0/diff_fold_casc_ota_1/vtail_casc VSS 47.41fF
C5404 input_amplifier_0/diff_fold_casc_ota_1/vbias4 VSS 214.47fF
C5405 input_amplifier_0/diff_fold_casc_ota_1/vbias3 VSS 140.70fF
C5406 input_amplifier_0/vim1 VSS 47.97fF
C5407 input_amplifier_0/txgate_4/txb VSS 0.42fF
C5408 input_amplifier_0/vip1 VSS 45.92fF
C5409 vincm VSS 26.77fF
C5410 input_amplifier_0/txgate_5/txb VSS 0.42fF
C5411 input_amplifier_0/rst VSS 0.24fF
C5412 rst_n VSS 49.54fF
C5413 input_amplifier_0/diff_fold_casc_ota_0/vcmcn_casc VSS 20.10fF
C5414 input_amplifier_0/diff_fold_casc_ota_0/vcmc_casc VSS 116.91fF
C5415 input_amplifier_0/diff_fold_casc_ota_0/M13d VSS 11.37fF
C5416 input_amplifier_0/vop1 VSS 252.20fF
C5417 input_amplifier_0/vom1 VSS 253.53fF
C5418 input_amplifier_0/diff_fold_casc_ota_0/vcmcn2_casc VSS 17.40fF
C5419 input_amplifier_0/diff_fold_casc_ota_0/vcmcn1_casc VSS 14.98fF
C5420 input_amplifier_0/diff_fold_casc_ota_0/M3d VSS 121.32fF
C5421 input_amplifier_0/diff_fold_casc_ota_0/vbias2 VSS 77.67fF
C5422 input_amplifier_0/diff_fold_casc_ota_0/M6d VSS 16.33fF
C5423 input_amplifier_0/diff_fold_casc_ota_0/vfoldp VSS 34.92fF
C5424 input_amplifier_0/diff_fold_casc_ota_0/vfoldm VSS 35.62fF
C5425 input_amplifier_0/diff_fold_casc_ota_0/M1d VSS 25.43fF
C5426 input_amplifier_0/diff_fold_casc_ota_0/vbias1 VSS 144.76fF
C5427 input_amplifier_0/diff_fold_casc_ota_0/M2d VSS 24.87fF
C5428 input_amplifier_0/venm2 VSS 10.22fF
C5429 input_amplifier_0/txgate_2/txb VSS 0.43fF
C5430 input_amplifier_0/venp2 VSS 11.42fF
C5431 input_amplifier_0/txgate_3/txb VSS 0.14fF
C5432 gain_ctrl_1 VSS 0.63fF
C5433 input_amplifier_0/diff_fold_casc_ota_1/vcmcn_casc VSS 20.10fF
C5434 input_amplifier_0/diff_fold_casc_ota_1/vcmc_casc VSS 116.91fF
C5435 input_amplifier_0/diff_fold_casc_ota_1/M13d VSS 11.37fF
C5436 vampp VSS 221.12fF
C5437 vampm VSS 216.07fF
C5438 input_amplifier_0/diff_fold_casc_ota_1/vcmcn2_casc VSS 17.40fF
C5439 input_amplifier_0/diff_fold_casc_ota_1/vcmcn1_casc VSS 14.98fF
C5440 input_amplifier_0/diff_fold_casc_ota_1/M3d VSS 121.32fF
C5441 input_amplifier_0/diff_fold_casc_ota_1/vbias2 VSS 77.67fF
C5442 input_amplifier_0/diff_fold_casc_ota_1/M6d VSS 16.33fF
C5443 input_amplifier_0/diff_fold_casc_ota_1/vfoldp VSS 34.92fF
C5444 input_amplifier_0/diff_fold_casc_ota_1/vfoldm VSS 35.62fF
C5445 input_amplifier_0/diff_fold_casc_ota_1/M1d VSS 25.43fF
C5446 input_amplifier_0/diff_fold_casc_ota_1/vbias1 VSS 144.76fF
C5447 input_amplifier_0/diff_fold_casc_ota_1/M2d VSS 24.87fF
C5448 VDD VSS 16228.00fF
.ends

