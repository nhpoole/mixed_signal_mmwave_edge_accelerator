* NGSPICE file created from deconv_kernel_estimator_top_level.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A VPB VNB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_2 A Y VPB VNB VPWR VGND
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__ha_2 VNB VPB VGND VPWR A COUT SUM B
X0 VPWR A a_342_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_766_47# B a_342_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND B a_389_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 COUT a_342_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND A a_766_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_342_199# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 a_468_369# B a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 a_389_47# a_342_199# a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_79_21# a_342_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 COUT a_342_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_389_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_342_199# COUT VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND a_79_21# SUM VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR a_79_21# SUM VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND a_342_199# COUT VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 SUM a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A a_468_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 SUM a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 X A VNB VPB VGND VPWR
X0 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__sdlclkp_4 SCE CLK GCLK GATE VGND VPWR VPB VNB
X0 a_257_147# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_109_369# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_465_315# a_287_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_1045_47# GCLK VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_287_413# a_257_147# a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5 VPWR a_257_147# a_257_243# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 GCLK a_1045_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_257_147# a_257_243# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR a_1045_47# GCLK VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND a_1045_47# GCLK VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_465_315# a_383_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_1127_47# a_465_315# a_1045_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_27_47# GATE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 GCLK a_1045_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_287_413# a_257_243# a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_383_413# a_257_147# a_287_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VGND CLK a_1127_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_257_147# CLK VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 GCLK a_1045_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 GCLK a_1045_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_27_47# GATE a_109_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 VPWR CLK a_1045_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1045_47# a_465_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_395_47# a_257_243# a_287_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 VGND a_1045_47# GCLK VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VGND a_465_315# a_395_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND SCE a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_465_315# a_287_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_1 B Y A VPB VNB VGND VPWR
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_1 Y A VPB VNB VGND VPWR w_84_21#
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22oi_1 B1 A1 B2 A2 Y VPWR VGND VPB VNB
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_381_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_12 A X VGND VPWR VPB VNB
X0 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND X A VPB VNB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xnor2_1 VGND VPWR B Y A VPB VNB
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_4 A Y VNB VPB VPWR VGND w_82_21#
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_16 Y A VPB VNB VGND VPWR
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR A2 A1 B1 Y VPB VNB
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21oi_1 A1 B1 Y A2 VPWR VGND VPB VNB
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xor2_1 B X A VNB VPB VPWR VGND
X0 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 VPB VNB Q CLK D VPWR VGND
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a32o_1 X A3 B2 B1 A1 A2 VGND VPWR VPB VNB
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 X A VGND VPWR VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2_0 VNB VPB VPWR VGND X B A
X0 VPWR B a_40_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_40_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VGND B a_123_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_40_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_123_47# A a_40_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_40_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2_0 A X B VNB VPB VGND VPWR
X0 VGND A a_68_355# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_150_355# B a_68_355# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_68_355# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_68_355# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR A a_150_355# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_68_355# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a211o_1 VNB VPB VGND VPWR X A2 B1 A1 C1
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21a_1 X A1 B1 A2 VPB VNB VGND VPWR
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_2 VGND VPWR A1 A0 S X VPB VNB
X0 VPWR S a_591_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_591_369# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_79_21# A1 a_306_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND S a_578_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_306_369# a_257_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 a_79_21# A0 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_288_47# a_257_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_257_199# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_578_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_257_199# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__fa_2 COUT SUM A B CIN VGND VPWR VPB VNB
X0 VGND CIN a_829_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VGND a_1086_47# SUM VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 COUT a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_829_369# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 VPWR CIN a_829_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_473_371# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X6 a_294_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR A a_473_371# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X8 a_829_369# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 a_829_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_829_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_473_371# CIN a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X12 a_473_47# CIN a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VPWR a_1086_47# SUM VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_473_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VGND a_80_21# COUT VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 COUT a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 SUM a_1086_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_80_21# B a_289_371# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X19 a_80_21# B a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 SUM a_1086_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND A a_473_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR a_80_21# COUT VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_289_371# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X24 a_1194_47# CIN a_1086_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_1086_47# a_80_21# a_829_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND A a_1266_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_1266_371# B a_1171_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X28 VPWR A a_1266_371# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X29 a_1266_47# B a_1194_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 a_1086_47# a_80_21# a_829_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X31 a_1171_369# CIN a_1086_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3_1 Y A C B VPB VNB VGND VPWR
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__sdlclkp_1 SCE CLK GCLK GATE VGND VPWR VPB VNB
X0 a_464_315# a_286_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_1094_47# a_464_315# a_1012_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_464_315# a_286_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR CLK a_1012_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_1012_47# a_464_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_109_369# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 VPWR a_464_315# a_382_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_382_413# a_256_147# a_286_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_286_413# a_256_243# a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_27_47# GATE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_256_147# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 VGND a_256_147# a_256_243# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 GCLK a_1012_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_27_47# GATE a_109_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 a_256_147# CLK VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 GCLK a_1012_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR a_256_147# a_256_243# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 a_286_413# a_256_147# a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18 VGND CLK a_1094_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_394_47# a_256_243# a_286_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20 VGND a_464_315# a_394_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND SCE a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21bai_1 A1 Y B1_N A2 VPB VNB VPWR VGND
X0 a_105_352# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_297_47# a_105_352# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A1 a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR B1_N a_105_352# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y a_105_352# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_388_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__maj3_1 C X B A VPB VNB VGND VPWR
X0 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_109_341# C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_27_47# B a_265_341# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_265_341# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A a_109_341# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_421_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_265_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND C a_421_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR C a_421_341# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_27_47# B a_265_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_421_341# B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_109_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22ai_1 A2 B1 Y A1 B2 VPB VNB VGND VPWR
X0 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR A1 a_307_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_307_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_1 Y B A VPB VNB VGND VPWR
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2b_1 B_N Y A VPB VNB VGND VPWR
X0 Y a_74_47# a_265_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR B_N a_74_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_265_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND B_N a_74_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND a_74_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o31ai_1 Y A2 A1 A3 B1 VPB VNB VPWR VGND
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y A3 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_297# A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A VPB VNB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3_1 A X B C VPWR VGND VPB VNB
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3_1 C Y A B VPB VNB VGND VPWR
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_6 VPWR VGND X A VPB VNB
X0 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR VPB VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=5.36e+06u area=4.347e+11p
.ends

.subckt sky130_fd_sc_hd__a21boi_1 Y A1 B1_N A2 VPWR VGND VPB VNB
X0 a_300_297# a_27_413# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Y a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A1 a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_384_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_300_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 Y C1 B1 VPB VNB VGND VPWR
X0 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_326_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y C1 a_326_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2bb2ai_1 Y A1_N A2_N B2 B1 VPB VNB VGND VPWR
X0 Y a_112_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND B2 a_394_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_112_297# A2_N a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_112_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_112_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR B1 a_478_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_394_47# a_112_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_394_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_478_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A2_N a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_8 X A VPB VNB VGND VPWR
X0 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3_2 A Y B C VNB VPB VGND VPWR
X0 VGND C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_277_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_277_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_8 Y A VNB VPB VGND VPWR w_189_21#
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21o_2 X B1 A1 A2 VNB VPB VGND VPWR
X0 X a_80_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_80_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_386_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_80_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_80_199# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_386_297# B1 a_80_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_458_47# A1 a_80_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A1 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A2 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR a_80_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 Y VPWR VGND VPB VNB
X0 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_467_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_467_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A1 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_109_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A2 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22o_1 A1 A2 X B2 B1 VPWR VGND VPB VNB
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21oi_2 B1 A2 A1 Y VNB VPB VGND VPWR
X0 VGND A2 a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A1 a_114_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_114_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_285_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_8 A X VGND VPWR VPB VNB
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_12 A Y VNB VPB VGND VPWR
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_8 A Y VNB VPB VGND VPWR
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__bufbuf_8 A X VNB VPB VGND VPWR
X0 VPWR a_206_47# a_318_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_318_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_318_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_318_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_318_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_206_47# a_318_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR a_318_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_318_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_318_47# a_206_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_318_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_206_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_318_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_206_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR a_318_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND a_206_47# a_318_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND a_318_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND a_318_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND a_318_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 X a_318_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND a_318_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VPWR a_206_47# a_318_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 X a_318_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_318_47# a_206_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VPWR a_318_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__bufinv_8 A Y VNB VPB VGND VPWR
X0 VPWR a_215_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_109_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND a_109_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND a_215_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_215_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_215_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND a_215_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND a_215_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR a_109_47# a_215_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_215_47# a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR a_215_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_215_47# a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR a_109_47# a_215_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR a_215_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 Y a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o32ai_1 A2 Y A1 A3 B2 B1 VPB VNB VGND VPWR
X0 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_333_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A1 a_461_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_461_297# A2 a_333_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand4_1 C B Y D A VPB VNB VPWR VGND
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_193_47# C a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y A a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_277_47# B a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

* Black-box entry subcircuit for sky130_sram_2kbyte_1rw1r_32x512_8 abstract view
.subckt sky130_sram_2kbyte_1rw1r_32x512_8 din0[0] din0[1] din0[2] din0[3] din0[4]
+ din0[5] din0[6] din0[7] din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14]
+ din0[15] din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22] din0[23]
+ din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[30] din0[31] addr0[0]
+ addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] addr0[8] addr1[0]
+ addr1[1] addr1[2] addr1[3] addr1[4] addr1[5] addr1[6] addr1[7] addr1[8] csb0 csb1
+ web0 clk0 clk1 wmask0[0] wmask0[1] wmask0[2] wmask0[3] dout0[0] dout0[1] dout0[2]
+ dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9] dout0[10] dout0[11]
+ dout0[12] dout0[13] dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19]
+ dout0[20] dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27]
+ dout0[28] dout0[29] dout0[30] dout0[31] dout1[0] dout1[1] dout1[2] dout1[3] dout1[4]
+ dout1[5] dout1[6] dout1[7] dout1[8] dout1[9] dout1[10] dout1[11] dout1[12] dout1[13]
+ dout1[14] dout1[15] dout1[16] dout1[17] dout1[18] dout1[19] dout1[20] dout1[21]
+ dout1[22] dout1[23] dout1[24] dout1[25] dout1[26] dout1[27] dout1[28] dout1[29]
+ dout1[30] dout1[31] vccd1 vssd1
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND X B A VPB VNB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_2 Y A B VPB VNB VGND VPWR
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_2 Y A VNB VPB VPWR VGND w_94_21#
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_4 Y A VPB VNB VPWR VGND
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2b_2 B_N A Y VPB VNB VGND VPWR
X0 Y a_251_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y a_251_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND a_251_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR B_N a_251_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND B_N a_251_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_27_297# a_251_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3_2 C Y A B VPB VNB VGND VPWR
X0 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_281_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2111ai_1 D1 C1 A2 A1 B1 Y VPB VNB VGND VPWR
X0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_235_47# C1 a_163_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_343_47# B1 a_235_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_454_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A1 a_454_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_163_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND A2 a_343_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_343_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2_1 A X B VPB VNB VGND VPWR
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__sdlclkp_2 SCE CLK GCLK GATE VGND VPWR VPB VNB
X0 GCLK a_1020_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_109_369# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_465_315# a_287_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_257_147# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_1102_47# a_465_315# a_1020_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND a_1020_47# GCLK VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_287_413# a_257_147# a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X7 VGND a_257_147# a_257_243# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND CLK a_1102_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR a_465_315# a_383_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_27_47# GATE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR CLK a_1020_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 GCLK a_1020_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_287_413# a_257_243# a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_383_413# a_257_147# a_287_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_257_147# CLK VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_27_47# GATE a_109_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 VPWR a_257_147# a_257_243# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X18 a_1020_47# a_465_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 a_395_47# a_257_243# a_287_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20 VGND a_465_315# a_395_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR a_1020_47# GCLK VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND SCE a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_465_315# a_287_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2b_1 Y A_N B VPB VNB VGND VPWR
X0 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Y a_27_93# a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_206_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_8 Y A B VPB VNB VGND VPWR
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_4 Y A B VPB VNB VGND VPWR
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21boi_0 B1_N Y A1 A2 VNB VPB VPWR VGND
X0 a_300_369# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_400_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND A2 a_400_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND B1_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR B1_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_300_369# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 VPWR A1 a_300_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hd__bufbuf_16 A X VNB VPB VGND VPWR
X0 VPWR a_215_47# a_549_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_109_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_109_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_215_47# a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_549_47# a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_215_47# a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_549_47# a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_549_47# a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_549_47# a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR a_215_47# a_549_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_549_47# a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VGND a_215_47# a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 VPWR a_109_47# a_215_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 a_215_47# a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X38 a_215_47# a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 VPWR a_109_47# a_215_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X41 VPWR a_215_47# a_549_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X43 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X44 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X45 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X46 a_549_47# a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X47 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X48 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X49 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X50 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X51 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3b_1 B C A_N Y VPB VNB VGND VPWR
X0 Y a_53_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_232_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A_N a_53_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND A_N a_53_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_316_47# B a_232_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y a_53_93# a_316_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22o_4 B1 B2 X A2 A1 VNB VPB VGND VPWR
X0 a_484_297# B2 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND B2 a_566_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_96_21# B1 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_484_297# B1 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_484_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_96_21# B2 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_96_21# B1 a_566_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A2 a_918_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_484_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A1 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_96_21# A1 a_918_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR A2 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_566_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_918_47# A1 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_566_47# B1 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_918_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__conb_1 LO HI VPB VNB VGND VPWR
R0 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
.ends

.subckt sky130_fd_sc_hd__a22o_2 A1 A2 X B2 B1 VPWR VGND VPB VNB
X0 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_381_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor4_1 D C Y A B VPB VNB VGND VPWR
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2_4 X B A VNB VPB VGND VPWR
X0 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND B a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_110_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a222oi_1 VNB VPB VPWR VGND C2 C1 B1 A2 A1 Y B2
X0 Y B1 a_393_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 VGND A2 a_561_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VGND C2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 Y C2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A1 a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_311_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_311_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_297# B2 a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_109_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_393_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_109_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 a_561_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a211oi_1 A1 C1 B1 Y A2 VPWR VGND VPB VNB
X0 a_56_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A2 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_139_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_311_297# B1 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y C1 a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A1 a_139_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_2 B Y A VPB VNB VGND VPWR
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2_2 VPWR VGND A X B VPB VNB
X0 X a_61_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_61_75# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B a_61_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND B a_147_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_61_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND a_61_75# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_61_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_147_75# A a_61_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4_1 C A X B D VPWR VGND VPB VNB
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a221oi_1 Y C1 A1 A2 B2 B1 VGND VPWR VPB VNB
X0 a_465_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_204_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y B1 a_204_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_109_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31oi_1 VGND VPWR Y B1 A2 A1 A3 VPB VNB
X0 a_181_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A1 a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_2 B1 Y A2 A1 VGND VPWR VPB VNB
X0 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__edfxtp_1 VPWR VGND CLK DE D Q VPB VNB
X0 a_381_369# D a_299_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 VGND a_1591_413# a_791_264# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 VPWR DE a_423_343# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_1591_413# a_193_47# a_1514_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5 a_1101_47# a_193_47# a_986_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X6 Q a_1591_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_986_413# a_193_47# a_299_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_1500_413# a_1150_159# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_1514_47# a_1150_159# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND DE a_423_343# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_1675_413# a_193_47# a_1591_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_1591_413# a_27_47# a_1500_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_729_47# a_423_343# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_729_369# DE VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X16 a_1077_413# a_27_47# a_986_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_791_264# a_1675_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 Q a_1591_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_299_47# a_791_264# a_729_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR a_1591_413# a_791_264# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 VGND a_791_264# a_1717_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 a_1717_47# a_27_47# a_1591_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 VPWR a_1150_159# a_1077_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_1150_159# a_986_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X26 a_986_413# a_27_47# a_299_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X27 a_299_47# a_791_264# a_729_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X28 a_381_47# D a_299_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 VGND a_1150_159# a_1101_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VPWR a_423_343# a_381_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X31 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VGND DE a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 a_1150_159# a_986_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3_4 Y A B C VNB VPB VGND VPWR
X0 a_27_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_445_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_445_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_445_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_445_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_27_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22a_1 A2 X B1 A1 B2 VPB VNB VGND VPWR
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3b_2 Y C A_N B VNB VPB VGND VPWR
X0 a_408_47# B a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_408_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y a_27_47# a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND C a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_218_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_218_47# B a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a221o_1 X B1 A1 B2 A2 VGND VPWR C1 VPB VNB
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o221ai_1 A2 Y B1 C1 A1 B2 VPB VNB VGND VPWR
X0 a_109_47# B1 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B2 a_295_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_213_123# B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_295_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_493_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A2 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_213_123# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__bufinv_16 A Y VNB VPB VGND VPWR
X0 a_361_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR a_27_47# a_361_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_361_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_361_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR a_27_47# a_361_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_361_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 VGND a_27_47# a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 VPWR a_27_47# a_361_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 VGND a_27_47# a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 VGND a_27_47# a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X38 a_361_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X41 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X43 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X44 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X45 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X46 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X47 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X48 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X49 a_361_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt deconv_kernel_estimator_top_level clk rst_n load_en debug_en serial_in sram_select[1]
+ sram_select[0] frequency_adc_done amplitude_adc_done sig_frequency[7] sig_frequency[6]
+ sig_frequency[5] sig_frequency[4] sig_frequency[3] sig_frequency[2] sig_frequency[1]
+ sig_frequency[0] sig_amplitude[7] sig_amplitude[6] sig_amplitude[5] sig_amplitude[4]
+ sig_amplitude[3] sig_amplitude[2] sig_amplitude[1] sig_amplitude[0] adc_bypass_en
+ serial_out serial_out_valid freq_eval_done VSS VDD
Xsky130_fd_sc_hd__clkbuf_1_508 VSS VDD sky130_fd_sc_hd__buf_8_218/A sky130_fd_sc_hd__buf_2_161/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_519 VSS VDD sky130_fd_sc_hd__clkbuf_1_519/X sky130_fd_sc_hd__nand3_1_37/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__inv_2_90 sky130_fd_sc_hd__inv_2_90/A sky130_fd_sc_hd__inv_2_90/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__ha_2_109 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_112/B sky130_fd_sc_hd__maj3_1_81/C
+ sky130_fd_sc_hd__ha_2_109/SUM sky130_fd_sc_hd__ha_2_109/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_11 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_11/A sky130_fd_sc_hd__ha_2_10/B
+ sky130_fd_sc_hd__ha_2_11/SUM sky130_fd_sc_hd__ha_2_11/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_22 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_22/A sky130_fd_sc_hd__ha_2_21/B
+ sky130_fd_sc_hd__ha_2_22/SUM sky130_fd_sc_hd__ha_2_22/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_33 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_33/A sky130_fd_sc_hd__ha_2_32/B
+ sky130_fd_sc_hd__ha_2_33/SUM sky130_fd_sc_hd__ha_2_33/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_44 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_44/A sky130_fd_sc_hd__ha_2_43/B
+ sky130_fd_sc_hd__ha_2_44/SUM sky130_fd_sc_hd__ha_2_44/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_55 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_55/A sky130_fd_sc_hd__ha_2_54/B
+ sky130_fd_sc_hd__ha_2_55/SUM sky130_fd_sc_hd__ha_2_55/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_66 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_66/A sky130_fd_sc_hd__ha_2_65/B
+ sky130_fd_sc_hd__ha_2_66/SUM sky130_fd_sc_hd__ha_2_66/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_77 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_77/A sky130_fd_sc_hd__ha_2_76/B
+ sky130_fd_sc_hd__ha_2_77/SUM sky130_fd_sc_hd__ha_2_77/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_88 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_88/A sky130_fd_sc_hd__ha_2_87/B
+ sky130_fd_sc_hd__ha_2_88/SUM sky130_fd_sc_hd__ha_2_88/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_99 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_99/A sky130_fd_sc_hd__maj3_1_55/C
+ sky130_fd_sc_hd__ha_2_99/SUM sky130_fd_sc_hd__ha_2_99/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_16_11 sky130_fd_sc_hd__clkbuf_4_210/A sky130_fd_sc_hd__buf_2_146/X
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__clkbuf_1_7 VSS VDD sky130_fd_sc_hd__buf_4_6/A sky130_fd_sc_hd__clkbuf_1_7/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__sdlclkp_4_40 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_72/A
+ sky130_fd_sc_hd__dfxtp_1_380/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_51 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_53/A
+ sky130_fd_sc_hd__dfxtp_1_473/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_62 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__clkinv_8_61/Y
+ sky130_fd_sc_hd__dfxtp_1_591/CLK sky130_fd_sc_hd__nand2b_1_5/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_73 sky130_fd_sc_hd__conb_1_23/LO sky130_fd_sc_hd__clkinv_8_53/A
+ sky130_fd_sc_hd__dfxtp_1_606/CLK sky130_fd_sc_hd__or2_0_6/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_84 sky130_fd_sc_hd__conb_1_26/LO sky130_fd_sc_hd__clkinv_8_68/Y
+ sky130_fd_sc_hd__dfxtp_1_1026/CLK sky130_fd_sc_hd__or2_0_10/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_120 sky130_fd_sc_hd__nor2_1_120/B sky130_fd_sc_hd__o21a_1_15/A1
+ sky130_fd_sc_hd__nor2_1_120/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_131 sky130_fd_sc_hd__nor2_1_131/B sky130_fd_sc_hd__nor2_1_131/Y
+ sky130_fd_sc_hd__nor2_1_131/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_142 sky130_fd_sc_hd__nor2_1_176/A sky130_fd_sc_hd__o21a_1_17/A1
+ sky130_fd_sc_hd__o21a_1_18/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_153 sky130_fd_sc_hd__nor2_1_153/B sky130_fd_sc_hd__o21a_1_26/A1
+ sky130_fd_sc_hd__o21a_1_27/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_1_7 sky130_fd_sc_hd__nor3_2_1/A sky130_fd_sc_hd__o21ai_1_0/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_7/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22oi_1_40 sky130_fd_sc_hd__a22oi_1_81/B1 sky130_fd_sc_hd__clkbuf_1_99/X
+ sky130_fd_sc_hd__clkbuf_1_47/X sky130_fd_sc_hd__clkbuf_4_22/X sky130_fd_sc_hd__nand4_1_3/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_164 sky130_fd_sc_hd__nor2_1_164/B sky130_fd_sc_hd__nor2_1_164/Y
+ sky130_fd_sc_hd__nor2_1_182/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_51 sky130_fd_sc_hd__nor2_2_2/Y sky130_fd_sc_hd__a22oi_1_82/A1
+ sky130_fd_sc_hd__clkbuf_1_64/X sky130_fd_sc_hd__a22oi_1_51/A2 sky130_fd_sc_hd__nand4_1_6/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_175 sky130_fd_sc_hd__nor2_1_175/B sky130_fd_sc_hd__nor2_1_175/Y
+ sky130_fd_sc_hd__nor2_1_183/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_186 sky130_fd_sc_hd__nor2_1_186/B sky130_fd_sc_hd__o21a_1_32/A1
+ sky130_fd_sc_hd__o21a_1_33/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_62 sky130_fd_sc_hd__a22oi_1_81/B1 sky130_fd_sc_hd__clkbuf_1_99/X
+ sky130_fd_sc_hd__clkbuf_1_40/X sky130_fd_sc_hd__clkbuf_4_15/X sky130_fd_sc_hd__nand4_1_10/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_197 sky130_fd_sc_hd__nor2_1_197/B sky130_fd_sc_hd__nor2_1_197/Y
+ sky130_fd_sc_hd__o21a_1_41/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_73 sky130_fd_sc_hd__a22oi_1_81/B1 sky130_fd_sc_hd__clkbuf_1_99/X
+ sky130_fd_sc_hd__clkbuf_1_37/X sky130_fd_sc_hd__clkbuf_4_12/X sky130_fd_sc_hd__nand4_1_13/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_84 sky130_fd_sc_hd__a22oi_1_96/B1 sky130_fd_sc_hd__a22oi_1_96/A1
+ sky130_fd_sc_hd__a22oi_1_84/B2 sky130_fd_sc_hd__a22oi_1_84/A2 sky130_fd_sc_hd__nand4_1_16/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_95 sky130_fd_sc_hd__clkbuf_4_72/X sky130_fd_sc_hd__clkbuf_4_73/X
+ sky130_fd_sc_hd__a22oi_1_95/B2 sky130_fd_sc_hd__buf_2_95/X sky130_fd_sc_hd__buf_2_110/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_360 sky130_fd_sc_hd__buf_12_360/A sky130_fd_sc_hd__buf_8_179/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_371 sky130_fd_sc_hd__buf_12_371/A sky130_fd_sc_hd__buf_12_371/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_230 sky130_fd_sc_hd__nor3_1_21/Y sky130_fd_sc_hd__nor2_4_8/Y
+ sky130_fd_sc_hd__clkbuf_1_422/X sky130_fd_sc_hd__buf_2_231/X sky130_fd_sc_hd__nand4_1_54/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_382 sky130_fd_sc_hd__inv_2_120/Y sky130_fd_sc_hd__buf_12_488/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_241 sky130_fd_sc_hd__a22oi_2_25/B1 sky130_fd_sc_hd__a22oi_2_25/A1
+ sky130_fd_sc_hd__clkbuf_1_386/X sky130_fd_sc_hd__a22oi_1_241/A2 sky130_fd_sc_hd__a22oi_1_241/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_393 sky130_fd_sc_hd__inv_2_129/Y sky130_fd_sc_hd__buf_12_393/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_252 sky130_fd_sc_hd__nor2_4_7/Y sky130_fd_sc_hd__buf_2_165/X
+ sky130_fd_sc_hd__clkbuf_1_492/X sky130_fd_sc_hd__clkbuf_1_440/X sky130_fd_sc_hd__nand4_1_62/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_263 sky130_fd_sc_hd__nor2_2_4/Y sky130_fd_sc_hd__clkbuf_1_377/X
+ sky130_fd_sc_hd__a22oi_1_263/B2 sky130_fd_sc_hd__clkbuf_4_191/X sky130_fd_sc_hd__nand4_1_65/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_274 sky130_fd_sc_hd__clkbuf_1_378/X sky130_fd_sc_hd__clkbuf_1_379/X
+ sky130_fd_sc_hd__clkbuf_4_172/X sky130_fd_sc_hd__buf_2_198/X sky130_fd_sc_hd__nand4_1_68/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_285 sky130_fd_sc_hd__clkbuf_4_165/X sky130_fd_sc_hd__clkinv_2_23/Y
+ sky130_fd_sc_hd__clkbuf_1_406/X sky130_fd_sc_hd__a22oi_1_285/A2 sky130_fd_sc_hd__a22oi_1_285/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_4_103 VDD VSS sky130_fd_sc_hd__buf_4_103/X sky130_fd_sc_hd__buf_4_103/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__a22oi_1_296 sky130_fd_sc_hd__clkbuf_1_376/X sky130_fd_sc_hd__nor2_2_5/Y
+ sky130_fd_sc_hd__buf_2_208/X sky130_fd_sc_hd__clkbuf_1_464/X sky130_fd_sc_hd__nand4_1_73/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_4_114 VDD VSS sky130_fd_sc_hd__buf_4_114/X sky130_fd_sc_hd__buf_8_201/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__xnor2_1_101 VSS VDD sky130_fd_sc_hd__o21a_1_62/B1 sky130_fd_sc_hd__xnor2_1_101/Y
+ sky130_fd_sc_hd__fa_2_1310/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_560 sky130_fd_sc_hd__nor2_1_70/B sky130_fd_sc_hd__fa_2_976/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_560/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_571 sky130_fd_sc_hd__nand2_1_275/A sky130_fd_sc_hd__a211oi_1_5/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_571/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_582 sky130_fd_sc_hd__o21ai_1_153/A2 sky130_fd_sc_hd__fa_2_1005/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_582/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_593 sky130_fd_sc_hd__nor2_1_90/B sky130_fd_sc_hd__nor2_4_9/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_593/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_4_40 sky130_fd_sc_hd__clkinv_4_40/A sky130_fd_sc_hd__buf_6_56/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_40/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_51 sky130_fd_sc_hd__clkinv_4_51/A sky130_fd_sc_hd__clkinv_8_63/A
+ VSS VDD VDD VSS VSS sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_62 sky130_fd_sc_hd__clkinv_4_0/A sky130_fd_sc_hd__clkinv_4_63/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_62/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_73 sky130_fd_sc_hd__clkinv_4_73/A sky130_fd_sc_hd__clkinv_4_73/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_73/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__o21ai_1_507 VSS VDD sky130_fd_sc_hd__nand2_1_568/A sky130_fd_sc_hd__o21ai_1_507/A1
+ sky130_fd_sc_hd__nand2_1_568/Y sky130_fd_sc_hd__and2_0_352/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a21oi_1_490 sky130_fd_sc_hd__or2_0_13/B sky130_fd_sc_hd__or2_0_0/B
+ sky130_fd_sc_hd__nand2_1_558/A sky130_fd_sc_hd__nor2_1_317/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__xor2_1_301 sky130_fd_sc_hd__nor2_4_20/Y sky130_fd_sc_hd__fa_2_1309/B
+ sky130_fd_sc_hd__xor2_1_301/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_312 sky130_fd_sc_hd__nor2_4_20/Y sky130_fd_sc_hd__fa_2_1298/B
+ sky130_fd_sc_hd__xor2_1_312/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_707 VDD VSS sky130_fd_sc_hd__mux2_2_19/A1 sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__o21ai_1_47/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_718 VDD VSS sky130_fd_sc_hd__mux2_2_28/A1 sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__nor2_1_41/B VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_729 VDD VSS sky130_fd_sc_hd__mux2_2_14/A1 sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__o21ai_1_66/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_305 VSS VDD sky130_fd_sc_hd__nand4_1_40/D sky130_fd_sc_hd__a22oi_1_179/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_316 VSS VDD sky130_fd_sc_hd__buf_2_126/A sky130_fd_sc_hd__buf_8_140/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_327 VSS VDD sky130_fd_sc_hd__buf_12_275/A sky130_fd_sc_hd__buf_8_124/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_338 VSS VDD sky130_fd_sc_hd__buf_8_149/A sky130_fd_sc_hd__buf_4_68/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_349 VSS VDD sky130_fd_sc_hd__buf_8_163/A sky130_fd_sc_hd__buf_8_158/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a32o_1_0 sky130_fd_sc_hd__a32o_1_0/X sky130_fd_sc_hd__a32o_1_0/A3
+ sky130_fd_sc_hd__nor2_1_71/Y sky130_fd_sc_hd__nor2_2_7/A sky130_fd_sc_hd__nor2_4_10/B
+ sky130_fd_sc_hd__nor2_2_9/A VSS VDD VDD VSS sky130_fd_sc_hd__a32o_1
Xsky130_fd_sc_hd__dfxtp_1_20 VDD VSS sky130_fd_sc_hd__ha_2_114/A sky130_fd_sc_hd__dfxtp_1_29/CLK
+ sky130_fd_sc_hd__nand4_1_38/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_31 VDD VSS sky130_fd_sc_hd__ha_2_168/B sky130_fd_sc_hd__clkinv_4_80/Y
+ sky130_fd_sc_hd__dfxtp_1_63/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_42 VDD VSS sky130_fd_sc_hd__fa_2_913/CIN sky130_fd_sc_hd__clkinv_4_80/Y
+ sky130_fd_sc_hd__buf_2_286/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_53 VDD VSS sky130_fd_sc_hd__fa_2_535/A sky130_fd_sc_hd__dfxtp_1_60/CLK
+ sky130_fd_sc_hd__nand4_1_39/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_64 VDD VSS sky130_fd_sc_hd__ha_2_99/B sky130_fd_sc_hd__dfxtp_1_77/CLK
+ sky130_fd_sc_hd__nand4_1_34/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_75 VDD VSS sky130_fd_sc_hd__buf_2_259/A sky130_fd_sc_hd__dfxtp_1_77/CLK
+ sky130_fd_sc_hd__dfxtp_1_75/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_86 VDD VSS sky130_fd_sc_hd__a22o_1_2/B2 sky130_fd_sc_hd__dfxtp_1_93/CLK
+ sky130_fd_sc_hd__buf_6_56/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_97 VDD VSS sky130_fd_sc_hd__ha_2_7/A sky130_fd_sc_hd__dfxtp_1_99/CLK
+ sky130_fd_sc_hd__and2_0_12/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_4_110 sky130_fd_sc_hd__clkbuf_4_110/X sky130_fd_sc_hd__nand3_4_1/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_121 sky130_fd_sc_hd__clkbuf_4_121/X sky130_fd_sc_hd__clkbuf_4_121/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_132 sky130_fd_sc_hd__clkbuf_4_132/X sky130_fd_sc_hd__clkbuf_4_132/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_303 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_303/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_303/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_143 sky130_fd_sc_hd__nand4_1_42/B sky130_fd_sc_hd__a22oi_1_189/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_314 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_314/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_314/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_154 sky130_fd_sc_hd__buf_8_127/A sky130_fd_sc_hd__buf_8_140/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_325 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_325/X sky130_fd_sc_hd__mux2_2_171/S
+ sky130_fd_sc_hd__and2_0_325/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_165 sky130_fd_sc_hd__clkbuf_4_165/X sky130_fd_sc_hd__nor3_2_10/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_336 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_336/X sky130_fd_sc_hd__inv_2_140/Y
+ sky130_fd_sc_hd__and2_0_336/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_176 sky130_fd_sc_hd__clkbuf_4_176/X sky130_fd_sc_hd__clkbuf_4_176/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_347 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_347/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_347/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_187 sky130_fd_sc_hd__clkbuf_4_187/X sky130_fd_sc_hd__clkbuf_4_187/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_198 sky130_fd_sc_hd__nand4_1_71/D sky130_fd_sc_hd__a22oi_1_285/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__inv_2_103 sky130_fd_sc_hd__inv_2_103/A sky130_fd_sc_hd__inv_2_103/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_114 sky130_fd_sc_hd__inv_4_0/Y sky130_fd_sc_hd__inv_2_114/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__or2_0_5 sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__or2_0_5/X sky130_fd_sc_hd__or2_0_5/B
+ VSS VDD VSS VDD sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__inv_2_125 sky130_fd_sc_hd__inv_2_125/A sky130_fd_sc_hd__inv_2_125/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_136 sky130_fd_sc_hd__inv_2_136/A sky130_fd_sc_hd__inv_2_136/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_12_190 sky130_fd_sc_hd__bufinv_8_1/Y sky130_fd_sc_hd__buf_12_190/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_390 sky130_fd_sc_hd__fa_2_882/B sky130_fd_sc_hd__nand2_1_35/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_390/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a211o_1_4 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_51/A sky130_fd_sc_hd__a211o_1_4/A2
+ sky130_fd_sc_hd__nor2_1_73/Y sky130_fd_sc_hd__a211o_1_6/A1 sky130_fd_sc_hd__o22ai_1_92/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o21ai_1_304 VSS VDD sky130_fd_sc_hd__o21ai_1_304/A2 sky130_fd_sc_hd__o22ai_1_265/A2
+ sky130_fd_sc_hd__a22oi_1_376/Y sky130_fd_sc_hd__o21ai_1_304/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_20 sky130_fd_sc_hd__o21a_1_20/X sky130_fd_sc_hd__o21a_1_20/A1
+ sky130_fd_sc_hd__o21a_1_20/B1 sky130_fd_sc_hd__fa_2_1132/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21ai_1_315 VSS VDD sky130_fd_sc_hd__a21oi_1_290/Y sky130_fd_sc_hd__nor2_1_172/A
+ sky130_fd_sc_hd__o21ai_1_317/B1 sky130_fd_sc_hd__o21ai_1_315/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_31 sky130_fd_sc_hd__o21a_1_31/X sky130_fd_sc_hd__o21a_1_31/A1
+ sky130_fd_sc_hd__o21a_1_31/B1 sky130_fd_sc_hd__fa_2_1187/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21ai_1_326 VSS VDD sky130_fd_sc_hd__o22ai_1_261/A2 sky130_fd_sc_hd__o21a_1_29/A2
+ sky130_fd_sc_hd__a21oi_1_295/Y sky130_fd_sc_hd__o21ai_1_326/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_337 VSS VDD sky130_fd_sc_hd__o22ai_1_292/A1 sky130_fd_sc_hd__nor2_1_204/Y
+ sky130_fd_sc_hd__or3_1_3/X sky130_fd_sc_hd__o21ai_1_337/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_42 sky130_fd_sc_hd__o21a_1_42/X sky130_fd_sc_hd__o21a_1_42/A1
+ sky130_fd_sc_hd__o21a_1_42/B1 sky130_fd_sc_hd__o21a_1_42/A2 VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21ai_1_348 VSS VDD sky130_fd_sc_hd__o22ai_1_304/A1 sky130_fd_sc_hd__o21a_1_42/A1
+ sky130_fd_sc_hd__a21oi_1_326/Y sky130_fd_sc_hd__o21ai_1_348/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_53 sky130_fd_sc_hd__o21a_1_53/X sky130_fd_sc_hd__o21a_1_53/A1
+ sky130_fd_sc_hd__o21a_1_53/B1 sky130_fd_sc_hd__fa_2_1250/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21ai_1_359 VSS VDD sky130_fd_sc_hd__o22ai_1_309/B1 sky130_fd_sc_hd__o21a_1_42/A1
+ sky130_fd_sc_hd__a21oi_1_337/Y sky130_fd_sc_hd__o21ai_1_359/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_64 sky130_fd_sc_hd__o21a_1_64/X sky130_fd_sc_hd__o21a_1_64/A1
+ sky130_fd_sc_hd__o21a_1_64/B1 sky130_fd_sc_hd__fa_2_1305/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__mux2_2_17 VSS VDD sky130_fd_sc_hd__mux2_2_17/A1 sky130_fd_sc_hd__mux2_2_17/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_17/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_28 VSS VDD sky130_fd_sc_hd__mux2_2_28/A1 sky130_fd_sc_hd__xor2_1_84/X
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_28/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_39 VSS VDD sky130_fd_sc_hd__mux2_2_39/A1 sky130_fd_sc_hd__mux2_2_39/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_39/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__xor2_1_120 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1086/B
+ sky130_fd_sc_hd__xor2_1_120/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_131 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1075/B
+ sky130_fd_sc_hd__xor2_1_131/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_142 sky130_fd_sc_hd__xor2_1_143/X sky130_fd_sc_hd__xor2_1_142/X
+ sky130_fd_sc_hd__xor2_1_164/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_153 sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__fa_2_1130/B
+ sky130_fd_sc_hd__xor2_1_153/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_504 VDD VSS sky130_fd_sc_hd__o21ai_1_35/A1 sky130_fd_sc_hd__edfxtp_1_0/CLK
+ sky130_fd_sc_hd__nor2b_1_80/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_164 sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__xor2_1_164/X
+ sky130_fd_sc_hd__xor2_1_164/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_515 VDD VSS sky130_fd_sc_hd__nor4_1_9/A sky130_fd_sc_hd__dfxtp_1_595/CLK
+ sky130_fd_sc_hd__a22o_1_56/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_175 sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__fa_2_1147/B
+ sky130_fd_sc_hd__xor2_1_175/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_186 sky130_fd_sc_hd__xor2_1_186/B sky130_fd_sc_hd__xor2_1_186/X
+ sky130_fd_sc_hd__xor2_1_187/X VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_526 VDD VSS sky130_fd_sc_hd__fa_2_965/A sky130_fd_sc_hd__dfxtp_1_526/CLK
+ sky130_fd_sc_hd__and2_0_265/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_537 VDD VSS sky130_fd_sc_hd__fa_2_954/A sky130_fd_sc_hd__dfxtp_1_538/CLK
+ sky130_fd_sc_hd__a22o_1_48/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_197 sky130_fd_sc_hd__fa_2_1173/A sky130_fd_sc_hd__fa_2_1182/B
+ sky130_fd_sc_hd__xor2_1_197/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_548 VDD VSS sky130_fd_sc_hd__xor2_1_31/A sky130_fd_sc_hd__dfxtp_1_548/CLK
+ sky130_fd_sc_hd__a22o_1_37/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_559 VDD VSS sky130_fd_sc_hd__and2_0_220/A sky130_fd_sc_hd__dfxtp_1_571/CLK
+ sky130_fd_sc_hd__dfxtp_1_560/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_102 VSS VDD sky130_fd_sc_hd__buf_8_9/A sky130_fd_sc_hd__ha_2_11/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_113 VSS VDD sky130_fd_sc_hd__clkbuf_1_98/A sky130_fd_sc_hd__clkinv_1_54/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_124 VSS VDD sky130_fd_sc_hd__clkbuf_1_124/X sky130_fd_sc_hd__buf_8_44/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_135 VSS VDD sky130_fd_sc_hd__a22oi_1_97/B1 sky130_fd_sc_hd__nor3_1_11/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_146 VSS VDD sky130_fd_sc_hd__clkbuf_1_146/X sky130_fd_sc_hd__buf_2_122/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_157 VSS VDD sky130_fd_sc_hd__clkbuf_1_157/X sky130_fd_sc_hd__clkbuf_1_157/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_4 VDD VSS sky130_fd_sc_hd__dfxtp_1_4/Q sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__a22o_1_1/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_168 VSS VDD sky130_fd_sc_hd__clkbuf_1_168/X sky130_fd_sc_hd__buf_2_123/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_179 VSS VDD sky130_fd_sc_hd__nand4_1_27/B sky130_fd_sc_hd__a22oi_2_12/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_409 sky130_fd_sc_hd__fa_2_411/CIN sky130_fd_sc_hd__fa_2_406/A
+ sky130_fd_sc_hd__fa_2_409/A sky130_fd_sc_hd__fa_2_409/B sky130_fd_sc_hd__fa_2_409/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nand3_1_13 sky130_fd_sc_hd__nand3_1_13/Y sky130_fd_sc_hd__a22oi_2_1/Y
+ sky130_fd_sc_hd__nand3_1_13/C sky130_fd_sc_hd__nand3_1_13/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_24 sky130_fd_sc_hd__buf_2_25/A sky130_fd_sc_hd__ha_2_20/A
+ sky130_fd_sc_hd__nand3_2_0/C sky130_fd_sc_hd__nor2_4_3/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_35 sky130_fd_sc_hd__buf_2_124/A sky130_fd_sc_hd__nand3_4_1/A
+ sky130_fd_sc_hd__nand3_1_35/C sky130_fd_sc_hd__nand3_4_1/C VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_46 sky130_fd_sc_hd__nand3_1_46/Y sky130_fd_sc_hd__or4_1_2/D
+ sky130_fd_sc_hd__nor3_1_32/Y sky130_fd_sc_hd__or4_1_2/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__dfxtp_1_1400 VDD VSS sky130_fd_sc_hd__mux2_2_243/A0 sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__o22ai_1_389/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1411 VDD VSS sky130_fd_sc_hd__mux2_2_267/A0 sky130_fd_sc_hd__clkinv_8_102/Y
+ sky130_fd_sc_hd__dfxtp_1_426/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1422 VDD VSS sky130_fd_sc_hd__mux2_2_244/A0 sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__dfxtp_1_437/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1433 VDD VSS sky130_fd_sc_hd__mux2_2_237/A0 sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__o22ai_1_400/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1444 VDD VSS serial_out_valid sky130_fd_sc_hd__clkinv_8_124/Y
+ sky130_fd_sc_hd__inv_2_141/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1455 VDD VSS sky130_fd_sc_hd__buf_6_84/A sky130_fd_sc_hd__dfxtp_1_1458/CLK
+ sky130_fd_sc_hd__and2_0_349/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1466 VDD VSS sky130_fd_sc_hd__nor2_1_320/A sky130_fd_sc_hd__clkinv_2_41/Y
+ sky130_fd_sc_hd__nor2b_1_139/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_100 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_100/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__fa_2_582/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_111 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_111/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__fa_2_864/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_122 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_122/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_891/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_30 sky130_fd_sc_hd__inv_2_19/A sky130_fd_sc_hd__inv_2_8/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_30/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_133 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_133/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_855/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_41 sky130_fd_sc_hd__inv_2_30/A sky130_fd_sc_hd__ha_2_12/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_41/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_144 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_144/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_843/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_52 sky130_fd_sc_hd__inv_2_41/A sky130_fd_sc_hd__inv_2_24/Y
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_155 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_155/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_926/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_63 sky130_fd_sc_hd__nor3_2_4/C sky130_fd_sc_hd__nor3_1_9/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_63/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_166 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_166/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_166/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_74 sky130_fd_sc_hd__inv_2_48/A sky130_fd_sc_hd__dfxtp_1_258/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_74/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_177 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_177/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_177/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_85 sky130_fd_sc_hd__buf_8_69/A sky130_fd_sc_hd__clkinv_1_86/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_85/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_188 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_188/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_927/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_96 sky130_fd_sc_hd__inv_2_60/A sky130_fd_sc_hd__ha_2_39/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_96/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_199 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_199/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__ha_2_165/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__fa_2_910 sky130_fd_sc_hd__fa_2_892/A sky130_fd_sc_hd__fa_2_893/B
+ sky130_fd_sc_hd__fa_2_910/A sky130_fd_sc_hd__fa_2_910/B sky130_fd_sc_hd__fa_2_910/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_921 sky130_fd_sc_hd__fa_2_920/CIN sky130_fd_sc_hd__fa_2_921/SUM
+ sky130_fd_sc_hd__fa_2_921/A sky130_fd_sc_hd__fa_2_921/B sky130_fd_sc_hd__fa_2_921/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_932 sky130_fd_sc_hd__fa_2_926/A sky130_fd_sc_hd__fa_2_927/B
+ sky130_fd_sc_hd__fa_2_932/A sky130_fd_sc_hd__fa_2_932/B sky130_fd_sc_hd__ha_2_121/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_943 sky130_fd_sc_hd__xnor2_1_25/A sky130_fd_sc_hd__fa_2_916/B
+ sky130_fd_sc_hd__fa_2_943/A sky130_fd_sc_hd__fa_2_943/B sky130_fd_sc_hd__ha_2_125/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_954 sky130_fd_sc_hd__fa_2_953/CIN sky130_fd_sc_hd__fa_2_954/SUM
+ sky130_fd_sc_hd__fa_2_954/A sky130_fd_sc_hd__fa_2_954/B sky130_fd_sc_hd__fa_2_954/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_965 sky130_fd_sc_hd__fa_2_964/CIN sky130_fd_sc_hd__fa_2_965/SUM
+ sky130_fd_sc_hd__fa_2_965/A sky130_fd_sc_hd__fa_2_965/B sky130_fd_sc_hd__fa_2_965/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_976 sky130_fd_sc_hd__fa_2_977/CIN sky130_fd_sc_hd__mux2_2_37/A1
+ sky130_fd_sc_hd__fa_2_976/A sky130_fd_sc_hd__fa_2_976/B sky130_fd_sc_hd__fa_2_976/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_987 sky130_fd_sc_hd__fa_2_988/CIN sky130_fd_sc_hd__mux2_2_13/A0
+ sky130_fd_sc_hd__fa_2_987/A sky130_fd_sc_hd__fa_2_987/B sky130_fd_sc_hd__fa_2_987/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_998 sky130_fd_sc_hd__fa_2_999/CIN sky130_fd_sc_hd__fa_2_998/SUM
+ sky130_fd_sc_hd__fa_2_998/A sky130_fd_sc_hd__fa_2_998/B sky130_fd_sc_hd__fa_2_998/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_1_5 sky130_fd_sc_hd__conb_1_27/LO sky130_fd_sc_hd__clkinv_4_60/A
+ sky130_fd_sc_hd__clkinv_2_36/A sky130_fd_sc_hd__or2_0_11/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_1
Xsky130_fd_sc_hd__mux2_2_210 VSS VDD sky130_fd_sc_hd__mux2_2_210/A1 sky130_fd_sc_hd__mux2_2_210/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_210/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_221 VSS VDD sky130_fd_sc_hd__mux2_2_221/A1 sky130_fd_sc_hd__xor2_1_276/X
+ sky130_fd_sc_hd__nor2_8_2/A sky130_fd_sc_hd__mux2_2_221/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_232 VSS VDD sky130_fd_sc_hd__mux2_2_232/A1 sky130_fd_sc_hd__mux2_2_232/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_232/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_243 VSS VDD sky130_fd_sc_hd__mux2_2_243/A1 sky130_fd_sc_hd__mux2_2_243/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_243/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_254 VSS VDD sky130_fd_sc_hd__mux2_2_254/A1 sky130_fd_sc_hd__mux2_2_254/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_254/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_265 VSS VDD sky130_fd_sc_hd__mux2_2_265/A1 sky130_fd_sc_hd__mux2_2_265/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_265/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__o21ai_1_101 VSS VDD sky130_fd_sc_hd__nor2_1_82/Y sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__a21oi_1_87/Y sky130_fd_sc_hd__xor2_1_70/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_112 VSS VDD sky130_fd_sc_hd__o21a_1_8/A2 sky130_fd_sc_hd__o21ai_1_112/A1
+ sky130_fd_sc_hd__a22oi_1_327/Y sky130_fd_sc_hd__o21ai_1_112/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_123 VSS VDD sky130_fd_sc_hd__a222oi_1_1/Y sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__nand2_1_273/Y sky130_fd_sc_hd__xor2_1_36/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_134 VSS VDD sky130_fd_sc_hd__a21oi_1_119/Y sky130_fd_sc_hd__nor2_1_76/A
+ sky130_fd_sc_hd__nand2b_1_13/Y sky130_fd_sc_hd__o21ai_1_134/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_145 VSS VDD sky130_fd_sc_hd__nor2_1_77/A sky130_fd_sc_hd__a21oi_1_134/Y
+ sky130_fd_sc_hd__a21oi_1_121/Y sky130_fd_sc_hd__xor2_1_53/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_156 VSS VDD sky130_fd_sc_hd__o21ai_1_156/A2 sky130_fd_sc_hd__o21ai_1_92/A1
+ sky130_fd_sc_hd__a22oi_1_345/Y sky130_fd_sc_hd__o21ai_1_156/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_167 VSS VDD sky130_fd_sc_hd__o21ai_1_171/A2 sky130_fd_sc_hd__xnor2_1_81/Y
+ sky130_fd_sc_hd__a21oi_1_144/Y sky130_fd_sc_hd__o21ai_1_167/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_178 VSS VDD sky130_fd_sc_hd__nand2_2_5/Y sky130_fd_sc_hd__xnor2_1_69/Y
+ sky130_fd_sc_hd__a21oi_1_153/Y sky130_fd_sc_hd__o21ai_1_178/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_189 VSS VDD sky130_fd_sc_hd__o21ai_1_189/A2 sky130_fd_sc_hd__nand2_1_284/Y
+ sky130_fd_sc_hd__a21oi_1_164/Y sky130_fd_sc_hd__o21ai_1_189/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21bai_1_2 sky130_fd_sc_hd__buf_2_263/A sky130_fd_sc_hd__o21bai_1_2/Y
+ sky130_fd_sc_hd__buf_2_262/X sky130_fd_sc_hd__o21bai_1_2/A2 VDD VSS VDD VSS sky130_fd_sc_hd__o21bai_1
Xsky130_fd_sc_hd__maj3_1_40 sky130_fd_sc_hd__maj3_1_41/X sky130_fd_sc_hd__maj3_1_40/X
+ sky130_fd_sc_hd__maj3_1_40/B sky130_fd_sc_hd__maj3_1_40/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_51 sky130_fd_sc_hd__maj3_1_52/X sky130_fd_sc_hd__maj3_1_51/X
+ sky130_fd_sc_hd__maj3_1_51/B sky130_fd_sc_hd__maj3_1_51/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_430 sky130_fd_sc_hd__o22ai_1_432/A2 sky130_fd_sc_hd__o22ai_1_430/B1
+ sky130_fd_sc_hd__o22ai_1_430/Y sky130_fd_sc_hd__nor2_1_277/B sky130_fd_sc_hd__o32ai_1_11/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_62 sky130_fd_sc_hd__maj3_1_63/X sky130_fd_sc_hd__maj3_1_62/X
+ sky130_fd_sc_hd__maj3_1_62/B sky130_fd_sc_hd__maj3_1_62/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_505 sky130_fd_sc_hd__o21a_1_62/B1 sky130_fd_sc_hd__fa_2_1309/A
+ sky130_fd_sc_hd__o21a_1_62/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_73 sky130_fd_sc_hd__maj3_1_74/X sky130_fd_sc_hd__maj3_1_73/X
+ sky130_fd_sc_hd__maj3_1_73/B sky130_fd_sc_hd__maj3_1_73/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_516 sky130_fd_sc_hd__nand2_1_516/Y sky130_fd_sc_hd__nor2_1_290/B
+ sky130_fd_sc_hd__nor2_1_287/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_84 sky130_fd_sc_hd__maj3_1_85/X sky130_fd_sc_hd__maj3_1_84/X
+ sky130_fd_sc_hd__maj3_1_84/B sky130_fd_sc_hd__maj3_1_84/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_527 sky130_fd_sc_hd__nor2_1_296/B sky130_fd_sc_hd__nand2_1_527/B
+ sky130_fd_sc_hd__nor2_1_297/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_95 sky130_fd_sc_hd__maj3_1_96/X sky130_fd_sc_hd__maj3_1_95/X
+ sky130_fd_sc_hd__maj3_1_95/B sky130_fd_sc_hd__maj3_1_95/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_538 sky130_fd_sc_hd__nand2_1_538/Y sky130_fd_sc_hd__xor2_1_298/A
+ sky130_fd_sc_hd__nor2_1_309/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_549 sky130_fd_sc_hd__a31oi_1_3/A3 sky130_fd_sc_hd__nand3_1_4/Y
+ sky130_fd_sc_hd__nor2_1_312/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_7 sky130_fd_sc_hd__ha_2_26/SUM sky130_fd_sc_hd__nor2b_1_7/Y
+ sky130_fd_sc_hd__or2_0_1/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1107 sky130_fd_sc_hd__nor2_1_280/B sky130_fd_sc_hd__fa_2_1302/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1107/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1118 sky130_fd_sc_hd__o21ai_1_507/A1 serial_in VDD VSS
+ VSS VDD sky130_fd_sc_hd__clkinv_1_1118/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1129 sky130_fd_sc_hd__clkinv_4_38/A sky130_fd_sc_hd__buf_4_121/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1129/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_90 sky130_fd_sc_hd__nand2_1_90/Y sky130_fd_sc_hd__nand2_1_91/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_301 VDD VSS sky130_fd_sc_hd__a22o_1_48/A1 sky130_fd_sc_hd__dfxtp_1_304/CLK
+ sky130_fd_sc_hd__and2_0_97/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_312 VDD VSS sky130_fd_sc_hd__a22o_1_37/A1 sky130_fd_sc_hd__dfxtp_1_477/CLK
+ sky130_fd_sc_hd__and2_0_86/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_323 VDD VSS sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__dfxtp_1_325/CLK
+ sky130_fd_sc_hd__and2_0_160/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_334 VDD VSS sky130_fd_sc_hd__a22o_2_10/B2 sky130_fd_sc_hd__clkinv_4_27/Y
+ sky130_fd_sc_hd__o21ai_1_26/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_345 VDD VSS sky130_fd_sc_hd__ha_2_155/A sky130_fd_sc_hd__dfxtp_1_347/CLK
+ sky130_fd_sc_hd__o2bb2ai_1_6/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_356 VDD VSS sky130_fd_sc_hd__a22o_2_4/B2 sky130_fd_sc_hd__dfxtp_1_360/CLK
+ sky130_fd_sc_hd__ha_2_149/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_367 VDD VSS sky130_fd_sc_hd__fa_2_1111/A sky130_fd_sc_hd__dfxtp_1_393/CLK
+ sky130_fd_sc_hd__and2_0_154/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_378 VDD VSS sky130_fd_sc_hd__ha_2_201/B sky130_fd_sc_hd__dfxtp_1_380/CLK
+ sky130_fd_sc_hd__and2_0_185/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_389 VDD VSS sky130_fd_sc_hd__fa_2_1117/B sky130_fd_sc_hd__dfxtp_1_391/CLK
+ sky130_fd_sc_hd__and2_0_120/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_9 sky130_fd_sc_hd__nand3_1_9/C sky130_fd_sc_hd__nand2_1_9/B
+ sky130_fd_sc_hd__nand2_1_9/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o31ai_1_12 sky130_fd_sc_hd__o31ai_1_12/Y sky130_fd_sc_hd__o31ai_1_12/A2
+ sky130_fd_sc_hd__nor2_1_287/A sky130_fd_sc_hd__o31ai_1_12/A3 sky130_fd_sc_hd__o31ai_1_12/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__o31ai_1
Xsky130_fd_sc_hd__fa_2_206 sky130_fd_sc_hd__fa_2_211/B sky130_fd_sc_hd__fa_2_206/SUM
+ sky130_fd_sc_hd__fa_2_206/A sky130_fd_sc_hd__fa_2_206/B sky130_fd_sc_hd__fa_2_206/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_217 sky130_fd_sc_hd__fa_2_214/A sky130_fd_sc_hd__fa_2_217/SUM
+ sky130_fd_sc_hd__fa_2_242/B sky130_fd_sc_hd__fa_2_247/A sky130_fd_sc_hd__fa_2_209/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_228 sky130_fd_sc_hd__fa_2_230/CIN sky130_fd_sc_hd__fa_2_221/B
+ sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__fa_2_280/A sky130_fd_sc_hd__fa_2_265/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_239 sky130_fd_sc_hd__fa_2_241/CIN sky130_fd_sc_hd__fa_2_236/A
+ sky130_fd_sc_hd__fa_2_239/A sky130_fd_sc_hd__fa_2_239/B sky130_fd_sc_hd__fa_2_247/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_20 sky130_fd_sc_hd__fa_2_16/B sky130_fd_sc_hd__fa_2_19/B sky130_fd_sc_hd__fa_2_20/A
+ sky130_fd_sc_hd__fa_2_20/B sky130_fd_sc_hd__fa_2_20/CIN VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_31 sky130_fd_sc_hd__maj3_1_28/B sky130_fd_sc_hd__maj3_1_29/A
+ sky130_fd_sc_hd__fa_2_31/A sky130_fd_sc_hd__ha_2_99/B sky130_fd_sc_hd__fa_2_67/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_42 sky130_fd_sc_hd__fa_2_44/B sky130_fd_sc_hd__fa_2_42/SUM
+ sky130_fd_sc_hd__ha_2_96/B sky130_fd_sc_hd__fa_2_96/A sky130_fd_sc_hd__fa_2_42/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_53 sky130_fd_sc_hd__fa_2_52/CIN sky130_fd_sc_hd__fa_2_53/SUM
+ sky130_fd_sc_hd__fa_2_82/A sky130_fd_sc_hd__ha_2_91/A sky130_fd_sc_hd__fa_2_96/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_64 sky130_fd_sc_hd__fa_2_69/B sky130_fd_sc_hd__fa_2_64/SUM
+ sky130_fd_sc_hd__fa_2_64/A sky130_fd_sc_hd__fa_2_64/B sky130_fd_sc_hd__fa_2_64/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_75 sky130_fd_sc_hd__fa_2_72/A sky130_fd_sc_hd__fa_2_75/SUM
+ sky130_fd_sc_hd__ha_2_96/B sky130_fd_sc_hd__ha_2_97/A sky130_fd_sc_hd__fa_2_67/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_86 sky130_fd_sc_hd__fa_2_88/CIN sky130_fd_sc_hd__fa_2_79/B
+ sky130_fd_sc_hd__fa_2_86/A sky130_fd_sc_hd__fa_2_91/A sky130_fd_sc_hd__fa_2_76/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_97 sky130_fd_sc_hd__fa_2_99/CIN sky130_fd_sc_hd__fa_2_94/A
+ sky130_fd_sc_hd__fa_2_97/A sky130_fd_sc_hd__fa_2_97/B sky130_fd_sc_hd__fa_2_97/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_201 VDD VSS sky130_fd_sc_hd__buf_2_201/X sky130_fd_sc_hd__buf_2_201/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_212 VDD VSS sky130_fd_sc_hd__buf_2_212/X sky130_fd_sc_hd__buf_2_212/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_223 VDD VSS sky130_fd_sc_hd__buf_2_223/X sky130_fd_sc_hd__buf_2_223/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_234 VDD VSS sky130_fd_sc_hd__buf_2_234/X sky130_fd_sc_hd__buf_2_234/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_245 VDD VSS sky130_fd_sc_hd__buf_2_245/X sky130_fd_sc_hd__inv_2_112/Y
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_256 VDD VSS sky130_fd_sc_hd__buf_2_256/X sky130_fd_sc_hd__inv_4_1/Y
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_267 VDD VSS sky130_fd_sc_hd__buf_2_267/X sky130_fd_sc_hd__buf_2_267/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_278 VDD VSS sky130_fd_sc_hd__buf_2_278/X amplitude_adc_done
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_289 VDD VSS sky130_fd_sc_hd__buf_2_289/X sky130_fd_sc_hd__buf_2_289/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1230 VDD VSS sky130_fd_sc_hd__xor2_1_254/A sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__mux2_2_173/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1241 VDD VSS sky130_fd_sc_hd__fa_2_1270/A sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__mux2_2_199/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1252 VDD VSS sky130_fd_sc_hd__nor2_4_18/A sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__nor2b_1_122/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1263 VDD VSS sky130_fd_sc_hd__mux2_2_185/A0 sky130_fd_sc_hd__clkinv_8_75/Y
+ sky130_fd_sc_hd__o22ai_1_328/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1274 VDD VSS sky130_fd_sc_hd__mux2_2_215/A0 sky130_fd_sc_hd__clkinv_8_63/Y
+ sky130_fd_sc_hd__dfxtp_1_430/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1285 VDD VSS sky130_fd_sc_hd__mux2_2_209/A0 sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__a21oi_1_379/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1296 VDD VSS sky130_fd_sc_hd__mux2_2_180/A1 sky130_fd_sc_hd__clkinv_8_116/Y
+ sky130_fd_sc_hd__o22ai_1_339/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_890 VDD VSS sky130_fd_sc_hd__fa_2_852/A sky130_fd_sc_hd__clkinv_4_22/Y
+ sky130_fd_sc_hd__o21a_1_24/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__or3_1_0 sky130_fd_sc_hd__or3_1_0/A sky130_fd_sc_hd__or3_1_0/X sky130_fd_sc_hd__or3_1_0/B
+ sky130_fd_sc_hd__or3_1_0/C VDD VSS VDD VSS sky130_fd_sc_hd__or3_1
Xsky130_fd_sc_hd__a21oi_1_14 sky130_fd_sc_hd__xor2_1_21/X sky130_fd_sc_hd__a21oi_1_14/B1
+ sky130_fd_sc_hd__a21oi_1_14/Y sky130_fd_sc_hd__nor2_1_13/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_25 sky130_fd_sc_hd__nand2b_1_8/Y sky130_fd_sc_hd__o21ai_1_39/Y
+ sky130_fd_sc_hd__a21oi_1_25/Y sky130_fd_sc_hd__or3_1_1/X VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_36 sky130_fd_sc_hd__nor2_1_41/Y sky130_fd_sc_hd__o22ai_1_69/Y
+ sky130_fd_sc_hd__a21oi_1_36/Y sky130_fd_sc_hd__fa_2_1039/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_47 sky130_fd_sc_hd__nor2_2_6/Y sky130_fd_sc_hd__o22ai_1_79/Y
+ sky130_fd_sc_hd__a21oi_1_47/Y sky130_fd_sc_hd__fa_2_1035/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_58 sky130_fd_sc_hd__nor2_2_6/Y sky130_fd_sc_hd__o22ai_1_89/Y
+ sky130_fd_sc_hd__a21oi_1_58/Y sky130_fd_sc_hd__nor2_1_91/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__fa_2_740 sky130_fd_sc_hd__fa_2_742/B sky130_fd_sc_hd__fa_2_738/A
+ sky130_fd_sc_hd__fa_2_832/A sky130_fd_sc_hd__fa_2_823/B sky130_fd_sc_hd__fa_2_826/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a21oi_1_69 sky130_fd_sc_hd__nand2_1_247/Y sky130_fd_sc_hd__nor2_1_52/Y
+ sky130_fd_sc_hd__xnor2_1_47/A sky130_fd_sc_hd__xnor2_1_45/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__fa_2_751 sky130_fd_sc_hd__fa_2_750/CIN sky130_fd_sc_hd__fa_2_751/SUM
+ sky130_fd_sc_hd__fa_2_835/B sky130_fd_sc_hd__fa_2_801/B sky130_fd_sc_hd__fa_2_812/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_762 sky130_fd_sc_hd__fa_2_761/A sky130_fd_sc_hd__fa_2_757/A
+ sky130_fd_sc_hd__fa_2_832/A sky130_fd_sc_hd__ha_2_140/A sky130_fd_sc_hd__fa_2_817/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_773 sky130_fd_sc_hd__fa_2_775/B sky130_fd_sc_hd__fa_2_773/SUM
+ sky130_fd_sc_hd__fa_2_773/A sky130_fd_sc_hd__fa_2_773/B sky130_fd_sc_hd__fa_2_777/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_784 sky130_fd_sc_hd__fa_2_786/B sky130_fd_sc_hd__fa_2_784/SUM
+ sky130_fd_sc_hd__fa_2_784/A sky130_fd_sc_hd__fa_2_784/B sky130_fd_sc_hd__fa_2_788/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_795 sky130_fd_sc_hd__fa_2_715/A sky130_fd_sc_hd__fa_2_716/B
+ sky130_fd_sc_hd__fa_2_795/A sky130_fd_sc_hd__fa_2_795/B sky130_fd_sc_hd__fa_2_800/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor3_1_6 sky130_fd_sc_hd__nor3_2_2/C sky130_fd_sc_hd__nor3_1_6/Y
+ sky130_fd_sc_hd__nor3_2_2/B sky130_fd_sc_hd__nor3_1_8/C VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__buf_6_10 VDD VSS sky130_fd_sc_hd__buf_8_56/A sky130_fd_sc_hd__inv_2_3/Y
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_21 VDD VSS sky130_fd_sc_hd__buf_6_21/X sky130_fd_sc_hd__inv_2_59/Y
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_32 VDD VSS sky130_fd_sc_hd__buf_6_40/A sky130_fd_sc_hd__inv_2_98/Y
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_43 VDD VSS sky130_fd_sc_hd__buf_6_43/X sky130_fd_sc_hd__buf_6_43/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_54 VDD VSS sky130_fd_sc_hd__buf_6_54/X sky130_fd_sc_hd__buf_6_54/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_65 VDD VSS sky130_fd_sc_hd__buf_6_65/X sky130_fd_sc_hd__buf_6_65/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_76 VDD VSS sky130_fd_sc_hd__buf_6_76/X sky130_fd_sc_hd__buf_6_77/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_12 sky130_fd_sc_hd__clkbuf_1_247/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__buf_6_87 VDD VSS sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__buf_6_87/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_23 sky130_fd_sc_hd__buf_2_59/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_308 sky130_fd_sc_hd__nor2_1_191/A sky130_fd_sc_hd__nor2_1_191/Y
+ sky130_fd_sc_hd__a21oi_1_308/Y sky130_fd_sc_hd__nor2_1_191/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_34 sky130_fd_sc_hd__nand4_1_23/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_319 sky130_fd_sc_hd__or3_1_3/C sky130_fd_sc_hd__o21ai_1_338/Y
+ sky130_fd_sc_hd__a21oi_1_319/Y sky130_fd_sc_hd__nor2_1_205/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_45 sky130_fd_sc_hd__buf_2_80/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_56 sky130_fd_sc_hd__buf_2_101/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_67 sky130_fd_sc_hd__buf_2_81/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_78 sky130_fd_sc_hd__buf_8_63/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_89 sky130_fd_sc_hd__clkbuf_1_535/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__nand2_1_302 sky130_fd_sc_hd__nand2_1_302/Y sky130_fd_sc_hd__nor2_1_104/B
+ sky130_fd_sc_hd__fa_2_1109/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_901 sky130_fd_sc_hd__clkinv_1_901/Y sky130_fd_sc_hd__nand2_1_428/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_901/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_313 sky130_fd_sc_hd__o21a_1_14/B1 sky130_fd_sc_hd__fa_2_1055/A
+ sky130_fd_sc_hd__o21a_1_14/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_912 sky130_fd_sc_hd__nor2_1_188/B sky130_fd_sc_hd__fa_2_1180/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_912/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_260 sky130_fd_sc_hd__o32ai_1_2/A3 sky130_fd_sc_hd__o22ai_1_265/B1
+ sky130_fd_sc_hd__o22ai_1_260/Y sky130_fd_sc_hd__nor2_1_151/B sky130_fd_sc_hd__o21a_1_29/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_324 sky130_fd_sc_hd__nand3_1_50/C sky130_fd_sc_hd__fa_2_1062/A
+ sky130_fd_sc_hd__nor2_4_12/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_271 sky130_fd_sc_hd__nand2_1_410/Y sky130_fd_sc_hd__nand2_1_409/Y
+ sky130_fd_sc_hd__o22ai_1_271/Y sky130_fd_sc_hd__nand2_1_421/B sky130_fd_sc_hd__o21ai_1_333/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_923 sky130_fd_sc_hd__nor2_1_220/A sky130_fd_sc_hd__xor2_1_208/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_923/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_335 sky130_fd_sc_hd__nand2_1_335/Y sky130_fd_sc_hd__fa_2_1091/A
+ sky130_fd_sc_hd__nor2_4_12/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_934 sky130_fd_sc_hd__o21ai_1_382/A1 sky130_fd_sc_hd__fa_2_1205/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_934/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_282 sky130_fd_sc_hd__nand2_1_412/Y sky130_fd_sc_hd__nand2_1_411/Y
+ sky130_fd_sc_hd__o22ai_1_282/Y sky130_fd_sc_hd__nand2_1_420/B sky130_fd_sc_hd__o21ai_1_332/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_346 sky130_fd_sc_hd__o21a_1_21/B1 sky130_fd_sc_hd__fa_2_1130/A
+ sky130_fd_sc_hd__o21a_1_21/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_293 sky130_fd_sc_hd__nor2_1_225/A sky130_fd_sc_hd__nor2_1_222/A
+ sky130_fd_sc_hd__o22ai_1_293/Y sky130_fd_sc_hd__a21boi_1_4/Y sky130_fd_sc_hd__nor2_1_206/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_945 sky130_fd_sc_hd__nor2_1_226/B sky130_fd_sc_hd__nor2_8_1/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_945/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_357 sky130_fd_sc_hd__nand2_1_357/Y sky130_fd_sc_hd__xnor2_1_93/Y
+ sky130_fd_sc_hd__xor2_1_140/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_956 sky130_fd_sc_hd__nor2_1_231/A sky130_fd_sc_hd__nor2_1_232/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_956/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_368 sky130_fd_sc_hd__a21o_2_6/A2 sky130_fd_sc_hd__nand2_1_368/B
+ sky130_fd_sc_hd__a21o_2_7/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_967 sky130_fd_sc_hd__o22ai_1_342/A1 sky130_fd_sc_hd__nor2_1_253/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_967/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_379 sky130_fd_sc_hd__nand2_1_379/Y sky130_fd_sc_hd__nor2b_1_104/Y
+ sky130_fd_sc_hd__o21ai_1_301/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_978 sky130_fd_sc_hd__nor2_1_248/B sky130_fd_sc_hd__xor2_1_275/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_978/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_989 sky130_fd_sc_hd__nor2_1_258/A sky130_fd_sc_hd__xor2_1_254/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_989/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_120 VDD VSS sky130_fd_sc_hd__inv_2_3/A sky130_fd_sc_hd__dfxtp_1_129/CLK
+ sky130_fd_sc_hd__and2_0_17/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_131 VDD VSS sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__clkinv_2_2/Y
+ sky130_fd_sc_hd__and2_0_21/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_142 VDD VSS sky130_fd_sc_hd__ha_2_20/A sky130_fd_sc_hd__dfxtp_1_143/CLK
+ sky130_fd_sc_hd__nor2b_1_11/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_153 VDD VSS sky130_fd_sc_hd__ha_2_34/A sky130_fd_sc_hd__dfxtp_1_155/CLK
+ sky130_fd_sc_hd__and2_0_27/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_164 VDD VSS sky130_fd_sc_hd__ha_2_45/A sky130_fd_sc_hd__clkinv_8_14/Y
+ sky130_fd_sc_hd__nor2b_1_21/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_175 VDD VSS sky130_fd_sc_hd__ha_2_59/A sky130_fd_sc_hd__dfxtp_1_185/CLK
+ sky130_fd_sc_hd__and2_0_56/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_186 VDD VSS sky130_fd_sc_hd__ha_2_69/B sky130_fd_sc_hd__dfxtp_1_195/CLK
+ sky130_fd_sc_hd__nor2b_1_26/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_197 VDD VSS sky130_fd_sc_hd__xor2_1_6/B sky130_fd_sc_hd__dfxtp_1_197/CLK
+ sky130_fd_sc_hd__nor2b_1_25/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a21boi_1_7 sky130_fd_sc_hd__a21boi_1_7/Y sky130_fd_sc_hd__nor2_2_18/Y
+ sky130_fd_sc_hd__a21oi_1_448/Y sky130_fd_sc_hd__fa_2_1288/A VDD VSS VDD VSS sky130_fd_sc_hd__a21boi_1
Xsky130_fd_sc_hd__fa_2_1230 sky130_fd_sc_hd__fa_2_1231/CIN sky130_fd_sc_hd__mux2_2_201/A1
+ sky130_fd_sc_hd__fa_2_1230/A sky130_fd_sc_hd__fa_2_1230/B sky130_fd_sc_hd__fa_2_1230/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o211ai_1_17 sky130_fd_sc_hd__nor2_1_126/A sky130_fd_sc_hd__nor2_1_129/Y
+ sky130_fd_sc_hd__xor2_1_134/A sky130_fd_sc_hd__nand2_1_326/Y sky130_fd_sc_hd__a22oi_1_353/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_28 sky130_fd_sc_hd__a21oi_1_275/Y sky130_fd_sc_hd__nor2_1_182/A
+ sky130_fd_sc_hd__xor2_1_175/A sky130_fd_sc_hd__a211oi_1_11/Y sky130_fd_sc_hd__nand2_1_379/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__fa_2_1241 sky130_fd_sc_hd__xor2_1_231/B sky130_fd_sc_hd__mux2_2_175/A0
+ sky130_fd_sc_hd__fa_2_1241/A sky130_fd_sc_hd__fa_2_1241/B sky130_fd_sc_hd__fa_2_1241/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o211ai_1_39 sky130_fd_sc_hd__nor2_1_214/A sky130_fd_sc_hd__a222oi_1_16/Y
+ sky130_fd_sc_hd__xor2_1_219/A sky130_fd_sc_hd__nand2_1_430/Y sky130_fd_sc_hd__a21oi_1_327/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__fa_2_1252 sky130_fd_sc_hd__fa_2_1253/CIN sky130_fd_sc_hd__mux2_2_189/A1
+ sky130_fd_sc_hd__fa_2_1252/A sky130_fd_sc_hd__fa_2_1252/B sky130_fd_sc_hd__fa_2_1252/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1263 sky130_fd_sc_hd__fa_2_1264/CIN sky130_fd_sc_hd__mux2_2_216/A1
+ sky130_fd_sc_hd__fa_2_1263/A sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1263/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1274 sky130_fd_sc_hd__xor2_1_273/B sky130_fd_sc_hd__nand2_1_469/A
+ sky130_fd_sc_hd__fa_2_1274/A sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1274/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1285 sky130_fd_sc_hd__fa_2_1286/CIN sky130_fd_sc_hd__mux2_2_238/A1
+ sky130_fd_sc_hd__fa_2_1285/A sky130_fd_sc_hd__fa_2_1285/B sky130_fd_sc_hd__fa_2_1285/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1296 sky130_fd_sc_hd__fa_2_1297/CIN sky130_fd_sc_hd__mux2_2_257/A1
+ sky130_fd_sc_hd__fa_2_1296/A sky130_fd_sc_hd__fa_2_1296/B sky130_fd_sc_hd__fa_2_1296/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1060 VDD VSS sky130_fd_sc_hd__fa_2_1199/A sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__mux2_2_146/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1071 VDD VSS sky130_fd_sc_hd__fa_2_1173/B sky130_fd_sc_hd__clkinv_4_23/Y
+ sky130_fd_sc_hd__and2_0_324/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_80 VSS VDD sky130_fd_sc_hd__xnor2_1_36/A sky130_fd_sc_hd__o21ai_1_80/A1
+ sky130_fd_sc_hd__o21ai_1_80/B1 sky130_fd_sc_hd__xnor2_1_38/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1082 VDD VSS sky130_fd_sc_hd__fa_2_1184/A sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__mux2_2_139/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_91 VSS VDD sky130_fd_sc_hd__o21ai_1_91/A2 sky130_fd_sc_hd__o21ai_1_92/A1
+ sky130_fd_sc_hd__o21ai_1_91/B1 sky130_fd_sc_hd__o21ai_1_91/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1093 VDD VSS sky130_fd_sc_hd__fa_2_1212/A sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__mux2_2_168/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o2bb2ai_1_11 sky130_fd_sc_hd__dfxtp_1_339/D sky130_fd_sc_hd__o21ai_1_28/A1
+ sky130_fd_sc_hd__nor2_1_18/Y sky130_fd_sc_hd__o21ai_1_31/A1 sky130_fd_sc_hd__o21ai_1_28/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__o2bb2ai_1_22 sky130_fd_sc_hd__dfxtp_1_564/D sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__dfxtp_1_564/Q sky130_fd_sc_hd__nand2_1_210/Y sky130_fd_sc_hd__nand3_1_46/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__o2bb2ai_1_33 sky130_fd_sc_hd__o2bb2ai_1_33/Y sky130_fd_sc_hd__nor4_1_13/B
+ sky130_fd_sc_hd__nor2_1_311/Y sky130_fd_sc_hd__nor2_1_311/Y sky130_fd_sc_hd__nor4_1_13/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_570 sky130_fd_sc_hd__fa_2_569/CIN sky130_fd_sc_hd__and2_0_88/A
+ sky130_fd_sc_hd__fa_2_570/A sky130_fd_sc_hd__fa_2_570/B sky130_fd_sc_hd__fa_2_570/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_581 sky130_fd_sc_hd__fa_2_580/CIN sky130_fd_sc_hd__and2_0_99/A
+ sky130_fd_sc_hd__fa_2_581/A sky130_fd_sc_hd__fa_2_581/B sky130_fd_sc_hd__fa_2_581/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_592 sky130_fd_sc_hd__maj3_1_126/B sky130_fd_sc_hd__maj3_1_127/A
+ sky130_fd_sc_hd__fa_2_592/A sky130_fd_sc_hd__fa_2_592/B sky130_fd_sc_hd__fa_2_593/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_1_208 sky130_fd_sc_hd__clkinv_1_208/Y sky130_fd_sc_hd__clkinv_2_22/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_208/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_219 sky130_fd_sc_hd__buf_4_106/A sky130_fd_sc_hd__clkinv_1_219/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_219/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_105 sky130_fd_sc_hd__a21o_2_3/A2 sky130_fd_sc_hd__o22ai_1_118/Y
+ sky130_fd_sc_hd__a21oi_1_105/Y sky130_fd_sc_hd__fa_2_972/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_116 sky130_fd_sc_hd__a211o_1_3/A1 sky130_fd_sc_hd__o22ai_1_124/Y
+ sky130_fd_sc_hd__a21oi_1_116/Y sky130_fd_sc_hd__nand2_1_275/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_127 sky130_fd_sc_hd__a21o_2_3/A2 sky130_fd_sc_hd__o21ai_1_151/Y
+ sky130_fd_sc_hd__a21oi_1_127/Y sky130_fd_sc_hd__fa_2_1008/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_138 sky130_fd_sc_hd__nor2_2_10/Y sky130_fd_sc_hd__o22ai_1_138/Y
+ sky130_fd_sc_hd__a21oi_1_138/Y sky130_fd_sc_hd__fa_2_1110/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nor2_1_302 sky130_fd_sc_hd__nor2_1_302/B sky130_fd_sc_hd__nor2_1_302/Y
+ sky130_fd_sc_hd__nor2_1_310/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a21oi_1_149 sky130_fd_sc_hd__clkinv_1_626/Y sky130_fd_sc_hd__a22o_1_72/X
+ sky130_fd_sc_hd__a21oi_1_149/Y sky130_fd_sc_hd__o21ai_1_199/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nor2_1_313 sky130_fd_sc_hd__nor2_1_315/A sky130_fd_sc_hd__nor2_1_313/Y
+ sky130_fd_sc_hd__nor2_1_314/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_401 sky130_fd_sc_hd__nor2_1_307/Y sky130_fd_sc_hd__nor2_1_309/Y
+ sky130_fd_sc_hd__fa_2_1302/A sky130_fd_sc_hd__fa_2_1298/A sky130_fd_sc_hd__a22oi_1_401/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkbuf_8_1 sky130_fd_sc_hd__buf_2_144/A sky130_fd_sc_hd__buf_2_143/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkbuf_8
Xsky130_fd_sc_hd__nand2_1_110 sky130_fd_sc_hd__nand2_1_110/Y sky130_fd_sc_hd__nand2_1_111/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_121 sky130_fd_sc_hd__nand2_1_121/Y sky130_fd_sc_hd__nand2_1_122/Y
+ sky130_fd_sc_hd__buf_2_264/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_720 sky130_fd_sc_hd__o22ai_1_193/A1 sky130_fd_sc_hd__fa_2_1055/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_720/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_132 sky130_fd_sc_hd__nand2_1_132/Y sky130_fd_sc_hd__fa_2_709/SUM
+ sky130_fd_sc_hd__and2_0_235/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_731 sky130_fd_sc_hd__clkinv_1_731/Y sky130_fd_sc_hd__nor2_1_123/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_731/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_143 sky130_fd_sc_hd__nand2_1_143/Y sky130_fd_sc_hd__nand2_1_144/Y
+ sky130_fd_sc_hd__buf_2_264/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_742 sky130_fd_sc_hd__o22ai_1_206/B2 sky130_fd_sc_hd__fa_2_1085/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_742/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_154 sky130_fd_sc_hd__fa_2_120/B sky130_fd_sc_hd__fa_2_91/A
+ sky130_fd_sc_hd__fa_2_2/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_753 sky130_fd_sc_hd__ha_2_197/B sky130_fd_sc_hd__fa_2_1110/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_753/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_165 sky130_fd_sc_hd__fa_2_276/A sky130_fd_sc_hd__fa_2_265/B
+ sky130_fd_sc_hd__fa_2_2/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_764 sky130_fd_sc_hd__ha_2_196/B sky130_fd_sc_hd__fa_2_1111/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_764/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_176 sky130_fd_sc_hd__fa_2_458/B sky130_fd_sc_hd__fa_2_559/B
+ sky130_fd_sc_hd__ha_2_125/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_775 sky130_fd_sc_hd__o22ai_1_204/B1 sky130_fd_sc_hd__nor2_4_12/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_775/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_187 sky130_fd_sc_hd__fa_2_625/B sky130_fd_sc_hd__ha_2_126/A
+ sky130_fd_sc_hd__ha_2_131/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_786 sky130_fd_sc_hd__nor2_1_180/A sky130_fd_sc_hd__nor2b_1_104/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_786/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_198 sky130_fd_sc_hd__fa_2_798/B sky130_fd_sc_hd__fa_2_834/B
+ sky130_fd_sc_hd__ha_2_140/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_797 sky130_fd_sc_hd__nor2_1_161/B sky130_fd_sc_hd__xor2_1_140/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_797/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor2_1_3 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__xor2_1_3/X
+ sky130_fd_sc_hd__xor2_1_3/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand3_2_4 sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__nand3_2_4/Y
+ sky130_fd_sc_hd__nand3_2_4/B sky130_fd_sc_hd__nand3_2_4/C VSS VDD VSS VDD sky130_fd_sc_hd__nand3_2
Xsky130_fd_sc_hd__clkinv_8_1 sky130_fd_sc_hd__clkinv_8_1/Y sky130_fd_sc_hd__clkinv_8_1/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_1/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__xor2_1_18 sky130_fd_sc_hd__xor2_1_18/B sky130_fd_sc_hd__nor4_1_3/C
+ sky130_fd_sc_hd__ha_2_153/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_29 sky130_fd_sc_hd__xor2_1_29/B sky130_fd_sc_hd__xor2_1_29/X
+ sky130_fd_sc_hd__or4_1_2/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nor3_1_20 sky130_fd_sc_hd__nor3_1_21/C sky130_fd_sc_hd__nor3_1_20/Y
+ sky130_fd_sc_hd__nor3_2_8/A sky130_fd_sc_hd__nor3_2_8/C VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_31 sky130_fd_sc_hd__nor3_1_31/C sky130_fd_sc_hd__nor3_1_31/Y
+ sky130_fd_sc_hd__or4_1_2/D sky130_fd_sc_hd__nor3_1_31/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__a21o_2_8 sky130_fd_sc_hd__a21o_2_8/X sky130_fd_sc_hd__a21o_2_8/B1
+ sky130_fd_sc_hd__a21o_2_8/A1 sky130_fd_sc_hd__a21o_2_8/A2 VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__fa_2_1060 sky130_fd_sc_hd__fa_2_1061/CIN sky130_fd_sc_hd__mux2_2_57/A0
+ sky130_fd_sc_hd__fa_2_1060/A sky130_fd_sc_hd__xor2_1_97/X sky130_fd_sc_hd__fa_2_1060/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1071 sky130_fd_sc_hd__fa_2_1072/CIN sky130_fd_sc_hd__and2_0_308/A
+ sky130_fd_sc_hd__fa_2_1071/A sky130_fd_sc_hd__fa_2_1071/B sky130_fd_sc_hd__fa_2_1071/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1082 sky130_fd_sc_hd__fa_2_1083/CIN sky130_fd_sc_hd__mux2_2_58/A0
+ sky130_fd_sc_hd__fa_2_1082/A sky130_fd_sc_hd__fa_2_1082/B sky130_fd_sc_hd__fa_2_1082/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1093 sky130_fd_sc_hd__fa_2_1094/CIN sky130_fd_sc_hd__and2_0_295/A
+ sky130_fd_sc_hd__fa_2_1093/A sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1093/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_509 VSS VDD sky130_fd_sc_hd__buf_12_397/A sky130_fd_sc_hd__buf_2_161/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__inv_2_80 sky130_fd_sc_hd__inv_2_80/A sky130_fd_sc_hd__inv_2_80/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_91 sky130_fd_sc_hd__inv_2_91/A sky130_fd_sc_hd__inv_2_91/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__ha_2_12 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_12/A sky130_fd_sc_hd__ha_2_11/B
+ sky130_fd_sc_hd__ha_2_12/SUM sky130_fd_sc_hd__ha_2_12/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_23 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_23/A sky130_fd_sc_hd__ha_2_22/B
+ sky130_fd_sc_hd__ha_2_23/SUM sky130_fd_sc_hd__ha_2_23/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_34 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_34/A sky130_fd_sc_hd__ha_2_33/B
+ sky130_fd_sc_hd__ha_2_34/SUM sky130_fd_sc_hd__ha_2_34/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_45 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_45/A sky130_fd_sc_hd__ha_2_44/B
+ sky130_fd_sc_hd__ha_2_45/SUM sky130_fd_sc_hd__ha_2_45/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_56 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_56/A sky130_fd_sc_hd__ha_2_55/B
+ sky130_fd_sc_hd__ha_2_56/SUM sky130_fd_sc_hd__ha_2_56/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_67 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_67/A sky130_fd_sc_hd__ha_2_66/B
+ sky130_fd_sc_hd__ha_2_67/SUM sky130_fd_sc_hd__ha_2_67/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_78 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_78/A sky130_fd_sc_hd__ha_2_77/B
+ sky130_fd_sc_hd__ha_2_78/SUM sky130_fd_sc_hd__ha_2_78/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_89 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_89/A sky130_fd_sc_hd__ha_2_88/B
+ sky130_fd_sc_hd__ha_2_89/SUM sky130_fd_sc_hd__ha_2_89/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__a22oi_2_0 sky130_fd_sc_hd__nor3_2_0/A sky130_fd_sc_hd__a22o_1_3/A1
+ sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__dfxtp_1_66/D sky130_fd_sc_hd__a22oi_2_0/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__sdlclkp_4_30 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_53/A
+ sky130_fd_sc_hd__dfxtp_1_277/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__clkbuf_1_8 VSS VDD sky130_fd_sc_hd__buf_6_5/A sky130_fd_sc_hd__clkbuf_1_8/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_16_12 sky130_fd_sc_hd__buf_12_508/A sky130_fd_sc_hd__clkinv_1_238/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__sdlclkp_4_41 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_72/A
+ sky130_fd_sc_hd__dfxtp_1_393/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_52 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_96/A
+ sky130_fd_sc_hd__dfxtp_1_462/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_63 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__clkinv_8_61/Y
+ sky130_fd_sc_hd__dfxtp_1_594/CLK sky130_fd_sc_hd__nand2b_1_5/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_74 sky130_fd_sc_hd__conb_1_24/LO sky130_fd_sc_hd__clkinv_8_58/A
+ sky130_fd_sc_hd__dfxtp_1_764/CLK sky130_fd_sc_hd__or2_0_8/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_85 sky130_fd_sc_hd__conb_1_27/LO sky130_fd_sc_hd__clkinv_2_35/Y
+ sky130_fd_sc_hd__dfxtp_1_1179/CLK sky130_fd_sc_hd__or2_0_11/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_110 sky130_fd_sc_hd__nor2_1_110/B sky130_fd_sc_hd__nor2_1_110/Y
+ sky130_fd_sc_hd__fa_2_1116/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_121 sky130_fd_sc_hd__nor2_1_121/B sky130_fd_sc_hd__a32o_1_1/B2
+ sky130_fd_sc_hd__nor2_4_12/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_132 sky130_fd_sc_hd__nor2_1_132/B sky130_fd_sc_hd__nor2_1_132/Y
+ sky130_fd_sc_hd__nor2_1_132/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_143 sky130_fd_sc_hd__nor2_1_143/B sky130_fd_sc_hd__o21a_1_18/A1
+ sky130_fd_sc_hd__o21a_1_19/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_30 sky130_fd_sc_hd__nor2_2_2/Y sky130_fd_sc_hd__a22oi_1_82/A1
+ sky130_fd_sc_hd__clkbuf_1_70/X sky130_fd_sc_hd__a22oi_1_30/A2 sky130_fd_sc_hd__nand4_1_0/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_154 sky130_fd_sc_hd__nor2_1_154/B sky130_fd_sc_hd__o21a_1_27/A1
+ sky130_fd_sc_hd__nor2_1_154/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_1_8 sky130_fd_sc_hd__and2_0_2/A sky130_fd_sc_hd__ha_2_9/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_8/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_165 sky130_fd_sc_hd__nor2_1_165/B sky130_fd_sc_hd__nor2_1_165/Y
+ sky130_fd_sc_hd__nor2_1_182/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_41 sky130_fd_sc_hd__nor2_2_2/Y sky130_fd_sc_hd__a22oi_1_82/A1
+ sky130_fd_sc_hd__clkbuf_1_67/X sky130_fd_sc_hd__a22oi_1_41/A2 sky130_fd_sc_hd__nand4_1_3/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_52 sky130_fd_sc_hd__clkbuf_4_8/X sky130_fd_sc_hd__clkbuf_4_9/X
+ sky130_fd_sc_hd__clkbuf_1_27/X sky130_fd_sc_hd__a22oi_1_52/A2 sky130_fd_sc_hd__a22oi_1_52/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_176 sky130_fd_sc_hd__o21a_1_29/A1 sky130_fd_sc_hd__nor2_1_176/Y
+ sky130_fd_sc_hd__nor2_1_176/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_187 sky130_fd_sc_hd__nor2_1_187/B sky130_fd_sc_hd__o21a_1_33/A1
+ sky130_fd_sc_hd__o21a_1_34/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_63 sky130_fd_sc_hd__nor2_2_2/Y sky130_fd_sc_hd__a22oi_1_82/A1
+ sky130_fd_sc_hd__clkbuf_1_60/X sky130_fd_sc_hd__a22oi_1_63/A2 sky130_fd_sc_hd__nand4_1_10/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_198 sky130_fd_sc_hd__nor2_1_198/B sky130_fd_sc_hd__o21a_1_41/A1
+ sky130_fd_sc_hd__nor2_1_198/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_74 sky130_fd_sc_hd__nor2_2_2/Y sky130_fd_sc_hd__a22oi_1_82/A1
+ sky130_fd_sc_hd__clkbuf_1_57/X sky130_fd_sc_hd__clkbuf_1_53/X sky130_fd_sc_hd__nand4_1_13/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_85 sky130_fd_sc_hd__nor3_1_11/Y sky130_fd_sc_hd__nor3_1_12/Y
+ sky130_fd_sc_hd__buf_2_65/X sky130_fd_sc_hd__clkbuf_4_89/X sky130_fd_sc_hd__nand4_1_16/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_96 sky130_fd_sc_hd__a22oi_1_96/B1 sky130_fd_sc_hd__a22oi_1_96/A1
+ sky130_fd_sc_hd__a22oi_1_96/B2 sky130_fd_sc_hd__a22oi_1_96/A2 sky130_fd_sc_hd__nand4_1_19/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_350 sky130_fd_sc_hd__buf_6_44/X sky130_fd_sc_hd__buf_12_350/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_361 sky130_fd_sc_hd__buf_12_361/A sky130_fd_sc_hd__buf_12_361/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_220 sky130_fd_sc_hd__buf_2_164/X sky130_fd_sc_hd__nor2_4_8/Y
+ sky130_fd_sc_hd__clkbuf_1_423/X sky130_fd_sc_hd__buf_2_232/X sky130_fd_sc_hd__nand4_1_51/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_372 sky130_fd_sc_hd__buf_12_372/A sky130_fd_sc_hd__buf_12_374/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_231 sky130_fd_sc_hd__nor3_2_8/Y sky130_fd_sc_hd__nor3_2_7/Y
+ sky130_fd_sc_hd__clkbuf_1_390/X sky130_fd_sc_hd__a22oi_1_231/A2 sky130_fd_sc_hd__a22oi_1_231/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_383 sky130_fd_sc_hd__inv_2_118/Y sky130_fd_sc_hd__buf_12_475/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_242 sky130_fd_sc_hd__buf_2_166/X sky130_fd_sc_hd__buf_2_167/X
+ sky130_fd_sc_hd__clkbuf_1_430/X sky130_fd_sc_hd__buf_2_172/X sky130_fd_sc_hd__nand4_1_59/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_394 sky130_fd_sc_hd__buf_6_58/X sky130_fd_sc_hd__buf_12_491/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_253 sky130_fd_sc_hd__buf_2_164/X sky130_fd_sc_hd__nor2_4_8/Y
+ sky130_fd_sc_hd__buf_2_184/X sky130_fd_sc_hd__clkbuf_1_455/X sky130_fd_sc_hd__nand4_1_62/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_264 sky130_fd_sc_hd__clkbuf_1_376/X sky130_fd_sc_hd__nor2_2_5/Y
+ sky130_fd_sc_hd__buf_2_216/X sky130_fd_sc_hd__clkbuf_1_472/X sky130_fd_sc_hd__nand4_1_65/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_275 sky130_fd_sc_hd__nor2_2_4/Y sky130_fd_sc_hd__clkbuf_1_377/X
+ sky130_fd_sc_hd__a22oi_1_275/B2 sky130_fd_sc_hd__clkbuf_4_188/X sky130_fd_sc_hd__nand4_1_68/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_286 sky130_fd_sc_hd__clkbuf_1_378/X sky130_fd_sc_hd__clkbuf_1_379/X
+ sky130_fd_sc_hd__buf_2_221/X sky130_fd_sc_hd__buf_2_195/X sky130_fd_sc_hd__nand4_1_71/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_4_104 VDD VSS sky130_fd_sc_hd__buf_4_104/X sky130_fd_sc_hd__buf_4_104/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__a22oi_1_297 sky130_fd_sc_hd__clkbuf_4_165/X sky130_fd_sc_hd__clkinv_2_23/Y
+ sky130_fd_sc_hd__clkbuf_1_403/X sky130_fd_sc_hd__a22oi_1_297/A2 sky130_fd_sc_hd__a22oi_1_297/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_4_115 VDD VSS sky130_fd_sc_hd__buf_4_115/X sky130_fd_sc_hd__buf_8_200/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__xnor2_1_102 VSS VDD sky130_fd_sc_hd__xor2_1_275/A sky130_fd_sc_hd__nor2_1_286/A
+ sky130_fd_sc_hd__xnor2_1_99/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_550 sky130_fd_sc_hd__a21oi_1_96/A1 sky130_fd_sc_hd__nor2_1_84/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_550/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_561 sky130_fd_sc_hd__o22ai_1_121/B2 sky130_fd_sc_hd__fa_2_974/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_561/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_572 sky130_fd_sc_hd__o21a_1_8/A1 sky130_fd_sc_hd__fa_2_1015/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_572/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_583 sky130_fd_sc_hd__o21ai_1_155/A1 sky130_fd_sc_hd__fa_2_1007/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_583/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_594 sky130_fd_sc_hd__ha_2_181/B sky130_fd_sc_hd__fa_2_1034/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_594/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_4_30 sky130_fd_sc_hd__clkinv_4_30/A sky130_fd_sc_hd__clkinv_4_31/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_30/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_41 sky130_fd_sc_hd__clkinv_4_41/A sky130_fd_sc_hd__buf_6_57/A
+ VSS VDD VDD VSS VSS sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_52 sky130_fd_sc_hd__clkinv_8_99/A sky130_fd_sc_hd__clkinv_4_53/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_52/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_63 sky130_fd_sc_hd__clkinv_4_63/A sky130_fd_sc_hd__clkinv_4_63/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_63/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_74 sky130_fd_sc_hd__clkinv_4_74/A sky130_fd_sc_hd__clkinv_4_9/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_74/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__inv_16_4 sky130_fd_sc_hd__inv_16_4/Y sky130_fd_sc_hd__inv_16_4/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__o21ai_1_508 VSS VDD sky130_fd_sc_hd__nor2_1_322/B sky130_fd_sc_hd__nor2_1_321/Y
+ sky130_fd_sc_hd__nand2_1_569/Y sky130_fd_sc_hd__o21ai_1_508/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a21oi_1_480 sky130_fd_sc_hd__or2_0_12/B sky130_fd_sc_hd__nor3_1_41/C
+ sky130_fd_sc_hd__o21bai_1_5/A2 sky130_fd_sc_hd__nor3_1_41/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_491 sky130_fd_sc_hd__or2_0_13/A sky130_fd_sc_hd__or2_0_0/B
+ sky130_fd_sc_hd__nand2_1_559/A sky130_fd_sc_hd__nor2_1_317/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__xor2_1_302 sky130_fd_sc_hd__nor2_4_20/Y sky130_fd_sc_hd__fa_2_1308/B
+ sky130_fd_sc_hd__xor2_1_302/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_313 sky130_fd_sc_hd__nor2_4_20/Y sky130_fd_sc_hd__fa_2_1297/B
+ sky130_fd_sc_hd__xor2_1_313/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_708 VDD VSS sky130_fd_sc_hd__mux2_2_17/A1 sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__o21ai_1_48/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_719 VDD VSS sky130_fd_sc_hd__mux2_2_36/A0 sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__a22o_1_68/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_306 VSS VDD sky130_fd_sc_hd__nand4_1_39/D sky130_fd_sc_hd__a22oi_1_175/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_317 VSS VDD sky130_fd_sc_hd__clkinv_1_169/A sky130_fd_sc_hd__clkbuf_1_366/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_328 VSS VDD sky130_fd_sc_hd__buf_4_67/A sky130_fd_sc_hd__nand2_1_568/B
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_339 VSS VDD sky130_fd_sc_hd__buf_6_34/A sky130_fd_sc_hd__inv_2_84/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a32o_1_1 sky130_fd_sc_hd__a32o_1_1/X sky130_fd_sc_hd__a32o_1_1/A3
+ sky130_fd_sc_hd__a32o_1_1/B2 sky130_fd_sc_hd__nor2_4_13/A sky130_fd_sc_hd__nor2_4_12/B
+ sky130_fd_sc_hd__nor2_2_13/A VSS VDD VDD VSS sky130_fd_sc_hd__a32o_1
Xsky130_fd_sc_hd__dfxtp_1_10 VDD VSS sky130_fd_sc_hd__dfxtp_1_10/Q sky130_fd_sc_hd__dfxtp_1_8/CLK
+ sky130_fd_sc_hd__a22o_1_7/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_21 VDD VSS sky130_fd_sc_hd__fa_2_393/A sky130_fd_sc_hd__dfxtp_1_29/CLK
+ sky130_fd_sc_hd__nand4_1_39/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_32 VDD VSS sky130_fd_sc_hd__fa_2_903/CIN sky130_fd_sc_hd__dfxtp_1_39/CLK
+ sky130_fd_sc_hd__nand4_1_34/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_43 VDD VSS sky130_fd_sc_hd__fa_2_914/CIN sky130_fd_sc_hd__clkinv_4_80/Y
+ sky130_fd_sc_hd__dfxtp_1_75/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_54 VDD VSS sky130_fd_sc_hd__ha_2_123/B sky130_fd_sc_hd__dfxtp_1_60/CLK
+ sky130_fd_sc_hd__buf_2_290/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_65 VDD VSS sky130_fd_sc_hd__ha_2_99/A sky130_fd_sc_hd__dfxtp_1_73/CLK
+ sky130_fd_sc_hd__nand4_1_35/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_76 VDD VSS sky130_fd_sc_hd__fa_2_247/A sky130_fd_sc_hd__dfxtp_1_77/CLK
+ sky130_fd_sc_hd__nand4_1_46/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_87 VDD VSS sky130_fd_sc_hd__a22o_1_3/B2 sky130_fd_sc_hd__dfxtp_1_93/CLK
+ sky130_fd_sc_hd__dfxtp_1_87/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_98 VDD VSS sky130_fd_sc_hd__ha_2_6/A sky130_fd_sc_hd__dfxtp_1_99/CLK
+ sky130_fd_sc_hd__and2_0_11/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_4_100 sky130_fd_sc_hd__buf_4_34/A sky130_fd_sc_hd__dfxtp_1_250/Q
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_111 sky130_fd_sc_hd__clkbuf_4_111/X sky130_fd_sc_hd__nor2_1_5/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_122 sky130_fd_sc_hd__clkbuf_4_122/X sky130_fd_sc_hd__clkbuf_4_122/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_133 sky130_fd_sc_hd__clkbuf_4_133/X sky130_fd_sc_hd__clkbuf_4_133/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_304 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_304/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_304/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_144 sky130_fd_sc_hd__nand4_1_41/B sky130_fd_sc_hd__a22oi_1_185/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_315 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_315/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_315/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_155 sky130_fd_sc_hd__clkbuf_4_155/X sky130_fd_sc_hd__clkbuf_4_155/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_326 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_326/X sky130_fd_sc_hd__mux2_2_171/S
+ sky130_fd_sc_hd__and2_0_326/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_166 sky130_fd_sc_hd__clkbuf_4_166/X sky130_fd_sc_hd__clkbuf_4_166/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_337 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_337/X sky130_fd_sc_hd__inv_2_140/Y
+ sky130_fd_sc_hd__and2_0_337/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_177 sky130_fd_sc_hd__clkbuf_4_177/X sky130_fd_sc_hd__clkbuf_4_177/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_348 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_348/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_348/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_188 sky130_fd_sc_hd__clkbuf_4_188/X sky130_fd_sc_hd__clkbuf_4_188/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_199 sky130_fd_sc_hd__nand4_1_69/D sky130_fd_sc_hd__a22oi_1_277/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__inv_2_104 sky130_fd_sc_hd__buf_6_38/A sky130_fd_sc_hd__inv_2_104/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_115 sky130_fd_sc_hd__inv_4_0/Y sky130_fd_sc_hd__inv_2_115/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__or2_0_6 sky130_fd_sc_hd__or2_0_6/A sky130_fd_sc_hd__or2_0_6/X sky130_fd_sc_hd__or2_0_6/B
+ VSS VDD VSS VDD sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__inv_2_126 sky130_fd_sc_hd__inv_2_126/A sky130_fd_sc_hd__buf_6_58/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_137 sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_37/S
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_12_180 sky130_fd_sc_hd__buf_8_95/X sky130_fd_sc_hd__buf_12_211/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_191 sky130_fd_sc_hd__bufinv_8_2/Y sky130_fd_sc_hd__buf_12_191/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_380 sky130_fd_sc_hd__fa_2_868/B sky130_fd_sc_hd__dfxtp_1_268/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_380/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_391 sky130_fd_sc_hd__fa_2_881/B sky130_fd_sc_hd__nor2_1_22/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_391/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a211o_1_5 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_79/A sky130_fd_sc_hd__a211o_1_5/A2
+ sky130_fd_sc_hd__nor2_1_74/Y sky130_fd_sc_hd__a211o_1_6/A1 sky130_fd_sc_hd__o22ai_1_93/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o21a_1_10 sky130_fd_sc_hd__o21a_1_10/X sky130_fd_sc_hd__o21a_1_10/A1
+ sky130_fd_sc_hd__o21a_1_10/B1 sky130_fd_sc_hd__fa_2_1064/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21ai_1_305 VSS VDD sky130_fd_sc_hd__o22ai_1_252/B1 sky130_fd_sc_hd__o21a_1_29/A1
+ sky130_fd_sc_hd__a21oi_1_277/Y sky130_fd_sc_hd__o21ai_1_305/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_316 VSS VDD sky130_fd_sc_hd__o22ai_1_258/B1 sky130_fd_sc_hd__o21a_1_29/A1
+ sky130_fd_sc_hd__a21oi_1_283/Y sky130_fd_sc_hd__o21ai_1_316/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_21 sky130_fd_sc_hd__o21a_1_21/X sky130_fd_sc_hd__o21a_1_21/A1
+ sky130_fd_sc_hd__o21a_1_21/B1 sky130_fd_sc_hd__fa_2_1130/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_32 sky130_fd_sc_hd__o21a_1_32/X sky130_fd_sc_hd__o21a_1_32/A1
+ sky130_fd_sc_hd__o21a_1_32/B1 sky130_fd_sc_hd__fa_2_1185/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21ai_1_327 VSS VDD sky130_fd_sc_hd__nor2_1_172/A sky130_fd_sc_hd__o21a_1_29/X
+ sky130_fd_sc_hd__a211oi_1_17/Y sky130_fd_sc_hd__xor2_1_160/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_43 sky130_fd_sc_hd__o21a_1_43/X sky130_fd_sc_hd__o21a_1_43/A1
+ sky130_fd_sc_hd__xnor2_1_97/B sky130_fd_sc_hd__fa_2_1240/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21ai_1_338 VSS VDD sky130_fd_sc_hd__nor2_1_205/Y sky130_fd_sc_hd__or3_1_3/C
+ sky130_fd_sc_hd__o31ai_1_8/A1 sky130_fd_sc_hd__o21ai_1_338/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_54 sky130_fd_sc_hd__o21a_1_54/X sky130_fd_sc_hd__o21a_1_54/A1
+ sky130_fd_sc_hd__o21a_1_54/B1 sky130_fd_sc_hd__fa_2_1247/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21ai_1_349 VSS VDD sky130_fd_sc_hd__nor2_1_224/A sky130_fd_sc_hd__a21oi_1_338/Y
+ sky130_fd_sc_hd__a21oi_1_329/Y sky130_fd_sc_hd__xor2_1_221/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_65 sky130_fd_sc_hd__o21a_1_65/X sky130_fd_sc_hd__o21a_1_65/A1
+ sky130_fd_sc_hd__o21a_1_65/B1 sky130_fd_sc_hd__fa_2_1303/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__mux2_2_18 VSS VDD sky130_fd_sc_hd__mux2_2_18/A1 sky130_fd_sc_hd__mux2_2_18/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_18/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_29 VSS VDD sky130_fd_sc_hd__mux2_2_29/A1 sky130_fd_sc_hd__mux2_2_29/A0
+ sky130_fd_sc_hd__mux2_2_37/S sky130_fd_sc_hd__mux2_2_29/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__xor2_1_110 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1047/B
+ sky130_fd_sc_hd__xor2_1_110/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_121 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1085/B
+ sky130_fd_sc_hd__xor2_1_121/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_132 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1074/B
+ sky130_fd_sc_hd__xor2_1_132/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_143 sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__xor2_1_143/X
+ sky130_fd_sc_hd__xor2_1_163/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_154 sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__fa_2_1129/B
+ sky130_fd_sc_hd__xor2_1_154/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_505 VDD VSS sky130_fd_sc_hd__xnor2_1_32/A sky130_fd_sc_hd__edfxtp_1_0/CLK
+ sky130_fd_sc_hd__nor2b_1_73/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_165 sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__fa_2_1157/B
+ sky130_fd_sc_hd__xor2_1_165/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_516 VDD VSS sky130_fd_sc_hd__nor4_1_10/B sky130_fd_sc_hd__dfxtp_1_520/CLK
+ sky130_fd_sc_hd__a22o_1_55/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_176 sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__fa_2_1146/B
+ sky130_fd_sc_hd__xor2_1_176/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_187 sky130_fd_sc_hd__xor2_1_188/X sky130_fd_sc_hd__xor2_1_187/X
+ sky130_fd_sc_hd__xor2_1_209/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_527 VDD VSS sky130_fd_sc_hd__fa_2_964/A sky130_fd_sc_hd__dfxtp_1_533/CLK
+ sky130_fd_sc_hd__and2_0_263/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_198 sky130_fd_sc_hd__fa_2_1173/A sky130_fd_sc_hd__fa_2_1181/B
+ sky130_fd_sc_hd__xor2_1_198/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_538 VDD VSS sky130_fd_sc_hd__fa_2_953/A sky130_fd_sc_hd__dfxtp_1_538/CLK
+ sky130_fd_sc_hd__a22o_1_47/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_549 VDD VSS sky130_fd_sc_hd__and2_0_225/A sky130_fd_sc_hd__dfxtp_1_577/CLK
+ sky130_fd_sc_hd__a22o_1_33/B1 VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_103 VSS VDD sky130_fd_sc_hd__buf_12_15/A sky130_fd_sc_hd__clkbuf_1_119/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_114 VSS VDD sky130_fd_sc_hd__bufinv_16_0/A sky130_fd_sc_hd__inv_2_43/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_125 VSS VDD sky130_fd_sc_hd__clkbuf_1_27/A sky130_fd_sc_hd__clkbuf_1_125/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_136 VSS VDD sky130_fd_sc_hd__a22oi_1_97/A1 sky130_fd_sc_hd__nor3_1_12/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_147 VSS VDD sky130_fd_sc_hd__clkbuf_1_147/X sky130_fd_sc_hd__clkbuf_1_147/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_158 VSS VDD sky130_fd_sc_hd__clkbuf_1_158/X sky130_fd_sc_hd__clkbuf_1_158/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_5 VDD VSS sky130_fd_sc_hd__dfxtp_1_5/Q sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__a22o_1_2/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_169 VSS VDD sky130_fd_sc_hd__a22oi_1_98/A2 sky130_fd_sc_hd__clkbuf_1_169/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__nand3_1_14 sky130_fd_sc_hd__nand3_1_14/Y sky130_fd_sc_hd__a22oi_2_2/Y
+ sky130_fd_sc_hd__nand3_1_14/C sky130_fd_sc_hd__nand3_1_14/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_25 sky130_fd_sc_hd__buf_2_22/A sky130_fd_sc_hd__nand3_2_2/A
+ sky130_fd_sc_hd__nand3_1_25/C sky130_fd_sc_hd__nand3_1_25/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_36 sky130_fd_sc_hd__nand3_1_36/Y sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__a22o_2_6/B1 sky130_fd_sc_hd__nor2_4_0/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_47 sky130_fd_sc_hd__nor4_1_5/B sky130_fd_sc_hd__nor4_1_8/Y
+ sky130_fd_sc_hd__nor4_1_6/Y sky130_fd_sc_hd__nor4_1_7/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__dfxtp_1_1401 VDD VSS sky130_fd_sc_hd__mux2_2_240/A0 sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__o22ai_1_388/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1412 VDD VSS sky130_fd_sc_hd__mux2_2_266/A0 sky130_fd_sc_hd__clkinv_8_102/Y
+ sky130_fd_sc_hd__dfxtp_1_427/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1423 VDD VSS sky130_fd_sc_hd__mux2_2_241/A0 sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__dfxtp_1_438/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1434 VDD VSS sky130_fd_sc_hd__mux2_2_234/A0 sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__o22ai_1_399/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1445 VDD VSS sky130_fd_sc_hd__o22ai_1_437/A1 sky130_fd_sc_hd__clkinv_8_116/Y
+ sky130_fd_sc_hd__nor2b_1_136/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1456 VDD VSS sky130_fd_sc_hd__dfxtp_1_1456/Q sky130_fd_sc_hd__dfxtp_1_1458/CLK
+ sky130_fd_sc_hd__and2_0_350/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1467 VDD VSS sky130_fd_sc_hd__nor2_1_318/A sky130_fd_sc_hd__clkinv_2_41/Y
+ sky130_fd_sc_hd__nor2b_1_140/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_101 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_101/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__xor2_1_25/X sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_112 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_112/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_889/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_20 sky130_fd_sc_hd__inv_2_9/A sky130_fd_sc_hd__ha_2_25/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_20/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_123 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_123/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_839/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_31 sky130_fd_sc_hd__inv_2_20/A sky130_fd_sc_hd__buf_8_23/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_31/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_134 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_134/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_841/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_42 sky130_fd_sc_hd__inv_2_31/A sky130_fd_sc_hd__buf_2_32/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_42/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_145 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_145/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_924/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_53 sky130_fd_sc_hd__inv_2_42/A sky130_fd_sc_hd__buf_2_12/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_53/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_156 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_156/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__fa_2_873/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_64 sky130_fd_sc_hd__nor3_1_13/C sky130_fd_sc_hd__nor3_2_4/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_64/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_167 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_167/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_167/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_75 sky130_fd_sc_hd__clkinv_1_76/A sky130_fd_sc_hd__dfxtp_1_259/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_75/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_178 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_178/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__ha_2_147/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_86 sky130_fd_sc_hd__buf_2_47/A sky130_fd_sc_hd__clkinv_1_86/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_86/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_189 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_189/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__edfxtp_1_0/Q sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_97 sky130_fd_sc_hd__inv_2_61/A sky130_fd_sc_hd__buf_2_45/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_97/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_900 sky130_fd_sc_hd__fa_2_899/CIN sky130_fd_sc_hd__fa_2_900/SUM
+ sky130_fd_sc_hd__fa_2_900/A sky130_fd_sc_hd__fa_2_900/B sky130_fd_sc_hd__fa_2_900/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_911 sky130_fd_sc_hd__fa_2_891/A sky130_fd_sc_hd__fa_2_892/B
+ sky130_fd_sc_hd__fa_2_911/A sky130_fd_sc_hd__fa_2_911/B sky130_fd_sc_hd__fa_2_911/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_922 sky130_fd_sc_hd__fa_2_921/CIN sky130_fd_sc_hd__fa_2_922/SUM
+ sky130_fd_sc_hd__fa_2_922/A sky130_fd_sc_hd__fa_2_922/B sky130_fd_sc_hd__fa_2_922/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_933 sky130_fd_sc_hd__fa_2_925/A sky130_fd_sc_hd__fa_2_926/B
+ sky130_fd_sc_hd__fa_2_933/A sky130_fd_sc_hd__fa_2_933/B sky130_fd_sc_hd__fa_2_502/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_944 sky130_fd_sc_hd__xor2_1_31/B sky130_fd_sc_hd__fa_2_944/SUM
+ sky130_fd_sc_hd__fa_2_944/A sky130_fd_sc_hd__fa_2_944/B sky130_fd_sc_hd__fa_2_944/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_955 sky130_fd_sc_hd__fa_2_954/CIN sky130_fd_sc_hd__fa_2_955/SUM
+ sky130_fd_sc_hd__fa_2_955/A sky130_fd_sc_hd__fa_2_955/B sky130_fd_sc_hd__fa_2_955/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_966 sky130_fd_sc_hd__fa_2_965/CIN sky130_fd_sc_hd__fa_2_966/SUM
+ sky130_fd_sc_hd__fa_2_966/A sky130_fd_sc_hd__fa_2_966/B sky130_fd_sc_hd__fa_2_966/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_977 sky130_fd_sc_hd__fa_2_978/CIN sky130_fd_sc_hd__mux2_2_35/A1
+ sky130_fd_sc_hd__fa_2_977/A sky130_fd_sc_hd__fa_2_977/B sky130_fd_sc_hd__fa_2_977/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_988 sky130_fd_sc_hd__fa_2_989/CIN sky130_fd_sc_hd__mux2_2_11/A0
+ sky130_fd_sc_hd__fa_2_988/A sky130_fd_sc_hd__fa_2_988/B sky130_fd_sc_hd__fa_2_988/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_999 sky130_fd_sc_hd__fa_2_999/COUT sky130_fd_sc_hd__mux2_2_36/A1
+ sky130_fd_sc_hd__fa_2_999/A sky130_fd_sc_hd__fa_2_999/B sky130_fd_sc_hd__fa_2_999/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_1_6 sky130_fd_sc_hd__conb_1_29/LO sky130_fd_sc_hd__clkinv_4_33/Y
+ sky130_fd_sc_hd__sdlclkp_1_6/GCLK sky130_fd_sc_hd__nand2b_1_18/Y VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_1
Xsky130_fd_sc_hd__mux2_2_200 VSS VDD sky130_fd_sc_hd__mux2_2_200/A1 sky130_fd_sc_hd__mux2_2_200/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_200/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_211 VSS VDD sky130_fd_sc_hd__mux2_2_211/A1 sky130_fd_sc_hd__mux2_2_211/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_211/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_222 VSS VDD sky130_fd_sc_hd__mux2_2_222/A1 sky130_fd_sc_hd__mux2_2_222/A0
+ sky130_fd_sc_hd__nor2_8_2/A sky130_fd_sc_hd__mux2_2_222/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_233 VSS VDD sky130_fd_sc_hd__mux2_2_233/A1 sky130_fd_sc_hd__mux2_2_233/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_233/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_244 VSS VDD sky130_fd_sc_hd__mux2_2_244/A1 sky130_fd_sc_hd__mux2_2_244/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_244/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_255 VSS VDD sky130_fd_sc_hd__mux2_2_255/A1 sky130_fd_sc_hd__mux2_2_255/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_255/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_266 VSS VDD sky130_fd_sc_hd__mux2_2_266/A1 sky130_fd_sc_hd__mux2_2_266/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_266/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__a22o_1_0 sky130_fd_sc_hd__buf_2_280/X sky130_fd_sc_hd__nor2_1_1/Y
+ sky130_fd_sc_hd__a22o_1_0/X sky130_fd_sc_hd__a22o_1_0/B2 sky130_fd_sc_hd__nor2_1_0/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__o21ai_1_102 VSS VDD sky130_fd_sc_hd__a21oi_1_95/Y sky130_fd_sc_hd__nor2_1_77/A
+ sky130_fd_sc_hd__nand2_1_264/Y sky130_fd_sc_hd__o21ai_1_102/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_113 VSS VDD sky130_fd_sc_hd__o22ai_1_119/A1 sky130_fd_sc_hd__o21a_1_8/A2
+ sky130_fd_sc_hd__a21oi_1_98/Y sky130_fd_sc_hd__a211o_1_8/A1 VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_124 VSS VDD sky130_fd_sc_hd__o21a_1_8/X sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__nand2_1_273/Y sky130_fd_sc_hd__xor2_1_37/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_135 VSS VDD sky130_fd_sc_hd__nor2_1_74/A sky130_fd_sc_hd__o21ai_1_135/A1
+ sky130_fd_sc_hd__a21oi_1_112/Y sky130_fd_sc_hd__xor2_1_47/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_146 VSS VDD sky130_fd_sc_hd__a21oi_1_124/Y sky130_fd_sc_hd__nor2_1_77/A
+ sky130_fd_sc_hd__a21oi_1_122/Y sky130_fd_sc_hd__xor2_1_54/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_157 VSS VDD sky130_fd_sc_hd__o22ai_1_123/A2 sky130_fd_sc_hd__o21ai_1_92/A1
+ sky130_fd_sc_hd__a22oi_1_346/Y sky130_fd_sc_hd__o21ai_1_157/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_168 VSS VDD sky130_fd_sc_hd__o21ai_1_171/A2 sky130_fd_sc_hd__xnor2_1_83/Y
+ sky130_fd_sc_hd__a21oi_1_145/Y sky130_fd_sc_hd__o21ai_1_168/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_179 VSS VDD sky130_fd_sc_hd__nand2_2_5/Y sky130_fd_sc_hd__xnor2_1_71/Y
+ sky130_fd_sc_hd__a21oi_1_154/Y sky130_fd_sc_hd__o21ai_1_179/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21bai_1_3 sky130_fd_sc_hd__buf_2_263/X sky130_fd_sc_hd__o21bai_1_3/Y
+ sky130_fd_sc_hd__buf_2_262/X sky130_fd_sc_hd__o21bai_1_3/A2 VDD VSS VDD VSS sky130_fd_sc_hd__o21bai_1
Xsky130_fd_sc_hd__maj3_1_30 sky130_fd_sc_hd__maj3_1_31/X sky130_fd_sc_hd__maj3_1_30/X
+ sky130_fd_sc_hd__maj3_1_30/B sky130_fd_sc_hd__maj3_1_30/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_41 sky130_fd_sc_hd__maj3_1_42/X sky130_fd_sc_hd__maj3_1_41/X
+ sky130_fd_sc_hd__maj3_1_41/B sky130_fd_sc_hd__maj3_1_41/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_420 sky130_fd_sc_hd__nor2_1_276/B sky130_fd_sc_hd__nor2_1_309/A
+ sky130_fd_sc_hd__o22ai_1_420/Y sky130_fd_sc_hd__o22ai_1_433/A1 sky130_fd_sc_hd__a222oi_1_39/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_52 sky130_fd_sc_hd__maj3_1_53/X sky130_fd_sc_hd__maj3_1_52/X
+ sky130_fd_sc_hd__maj3_1_52/B sky130_fd_sc_hd__maj3_1_52/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_431 sky130_fd_sc_hd__o32ai_1_11/A3 sky130_fd_sc_hd__o22ai_1_436/B1
+ sky130_fd_sc_hd__o22ai_1_431/Y sky130_fd_sc_hd__nor2_1_278/B sky130_fd_sc_hd__o21a_1_68/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_63 sky130_fd_sc_hd__maj3_1_64/X sky130_fd_sc_hd__maj3_1_63/X
+ sky130_fd_sc_hd__maj3_1_63/B sky130_fd_sc_hd__maj3_1_63/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_506 sky130_fd_sc_hd__o21a_1_63/B1 sky130_fd_sc_hd__fa_2_1307/A
+ sky130_fd_sc_hd__o21a_1_63/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_74 sky130_fd_sc_hd__maj3_1_75/X sky130_fd_sc_hd__maj3_1_74/X
+ sky130_fd_sc_hd__maj3_1_74/B sky130_fd_sc_hd__maj3_1_74/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_517 sky130_fd_sc_hd__nand2_1_517/Y sky130_fd_sc_hd__nand2_1_520/Y
+ sky130_fd_sc_hd__nand2_1_518/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_85 sky130_fd_sc_hd__maj3_1_86/X sky130_fd_sc_hd__maj3_1_85/X
+ sky130_fd_sc_hd__maj3_1_85/B sky130_fd_sc_hd__maj3_1_85/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_528 sky130_fd_sc_hd__nor2_1_297/B sky130_fd_sc_hd__nand2_1_528/B
+ sky130_fd_sc_hd__nor2_1_298/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_96 sky130_fd_sc_hd__maj3_1_97/X sky130_fd_sc_hd__maj3_1_96/X
+ sky130_fd_sc_hd__maj3_1_96/B sky130_fd_sc_hd__maj3_1_96/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_539 sky130_fd_sc_hd__nand2_1_539/Y sky130_fd_sc_hd__nand2_1_543/B
+ sky130_fd_sc_hd__o21ai_1_490/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_8 sky130_fd_sc_hd__ha_2_22/SUM sky130_fd_sc_hd__nor2b_1_8/Y
+ sky130_fd_sc_hd__or2_0_1/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1108 sky130_fd_sc_hd__o21a_1_68/A2 sky130_fd_sc_hd__fa_2_1304/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1108/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1119 sky130_fd_sc_hd__nand2_1_569/A sky130_fd_sc_hd__nor2_1_321/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1119/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_80 sky130_fd_sc_hd__nand2_1_80/Y sky130_fd_sc_hd__nand2_1_81/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_91 sky130_fd_sc_hd__nand2_1_91/Y sky130_fd_sc_hd__nand2_1_91/B
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_302 VDD VSS sky130_fd_sc_hd__a22o_1_47/A1 sky130_fd_sc_hd__dfxtp_1_304/CLK
+ sky130_fd_sc_hd__and2_0_96/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_313 VDD VSS sky130_fd_sc_hd__xor2_1_27/B sky130_fd_sc_hd__dfxtp_1_313/CLK
+ sky130_fd_sc_hd__and2_0_85/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_324 VDD VSS sky130_fd_sc_hd__or4_1_0/A sky130_fd_sc_hd__dfxtp_1_457/CLK
+ sky130_fd_sc_hd__and2_0_158/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_335 VDD VSS sky130_fd_sc_hd__a22o_4_0/B2 sky130_fd_sc_hd__clkinv_4_27/Y
+ sky130_fd_sc_hd__o21ai_1_27/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_346 VDD VSS sky130_fd_sc_hd__a22o_1_25/B2 sky130_fd_sc_hd__dfxtp_1_354/CLK
+ sky130_fd_sc_hd__ha_2_154/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_357 VDD VSS sky130_fd_sc_hd__ha_2_149/A sky130_fd_sc_hd__dfxtp_1_361/CLK
+ sky130_fd_sc_hd__o2bb2ai_1_3/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_368 VDD VSS sky130_fd_sc_hd__fa_2_1112/A sky130_fd_sc_hd__dfxtp_1_393/CLK
+ sky130_fd_sc_hd__and2_0_149/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_379 VDD VSS sky130_fd_sc_hd__fa_2_1107/B sky130_fd_sc_hd__dfxtp_1_380/CLK
+ sky130_fd_sc_hd__and2_0_186/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_207 sky130_fd_sc_hd__fa_2_204/B sky130_fd_sc_hd__fa_2_207/SUM
+ sky130_fd_sc_hd__fa_2_5/B sky130_fd_sc_hd__fa_2_247/A sky130_fd_sc_hd__fa_2_283/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_218 sky130_fd_sc_hd__fa_2_219/CIN sky130_fd_sc_hd__fa_2_212/A
+ sky130_fd_sc_hd__fa_2_265/B sky130_fd_sc_hd__fa_2_258/A sky130_fd_sc_hd__fa_2_277/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_229 sky130_fd_sc_hd__fa_2_230/B sky130_fd_sc_hd__fa_2_221/A
+ sky130_fd_sc_hd__fa_2_242/A sky130_fd_sc_hd__fa_2_273/A sky130_fd_sc_hd__fa_2_238/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_10 sky130_fd_sc_hd__fa_2_1/A sky130_fd_sc_hd__fa_2_8/B sky130_fd_sc_hd__fa_2_91/A
+ sky130_fd_sc_hd__fa_2_10/B sky130_fd_sc_hd__fa_2_13/SUM VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_21 sky130_fd_sc_hd__fa_2_18/B sky130_fd_sc_hd__fa_2_20/B sky130_fd_sc_hd__ha_2_97/B
+ sky130_fd_sc_hd__ha_2_94/B sky130_fd_sc_hd__fa_2_139/B VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_32 sky130_fd_sc_hd__fa_2_33/CIN sky130_fd_sc_hd__maj3_1_28/A
+ sky130_fd_sc_hd__fa_2_32/A sky130_fd_sc_hd__ha_2_99/A sky130_fd_sc_hd__fa_2_31/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_43 sky130_fd_sc_hd__fa_2_45/CIN sky130_fd_sc_hd__fa_2_41/A
+ sky130_fd_sc_hd__ha_2_97/B sky130_fd_sc_hd__ha_2_95/B sky130_fd_sc_hd__fa_2_87/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_54 sky130_fd_sc_hd__maj3_1_18/B sky130_fd_sc_hd__maj3_1_19/A
+ sky130_fd_sc_hd__fa_2_54/A sky130_fd_sc_hd__fa_2_54/B sky130_fd_sc_hd__fa_2_55/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_65 sky130_fd_sc_hd__fa_2_62/B sky130_fd_sc_hd__fa_2_65/SUM
+ sky130_fd_sc_hd__fa_2_82/A sky130_fd_sc_hd__ha_2_97/A sky130_fd_sc_hd__fa_2_49/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_76 sky130_fd_sc_hd__fa_2_77/CIN sky130_fd_sc_hd__fa_2_70/A
+ sky130_fd_sc_hd__fa_2_76/A sky130_fd_sc_hd__fa_2_76/B sky130_fd_sc_hd__fa_2_86/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_87 sky130_fd_sc_hd__fa_2_88/B sky130_fd_sc_hd__fa_2_79/A sky130_fd_sc_hd__fa_2_87/A
+ sky130_fd_sc_hd__fa_2_87/B sky130_fd_sc_hd__fa_2_9/A VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_98 sky130_fd_sc_hd__maj3_1_9/B sky130_fd_sc_hd__maj3_1_10/A
+ sky130_fd_sc_hd__fa_2_98/A sky130_fd_sc_hd__fa_2_98/B sky130_fd_sc_hd__fa_2_99/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_202 VDD VSS sky130_fd_sc_hd__buf_2_202/X sky130_fd_sc_hd__buf_2_202/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_213 VDD VSS sky130_fd_sc_hd__buf_2_213/X sky130_fd_sc_hd__buf_2_213/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_224 VDD VSS sky130_fd_sc_hd__buf_2_224/X sky130_fd_sc_hd__buf_2_224/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_235 VDD VSS sky130_fd_sc_hd__buf_2_235/X sky130_fd_sc_hd__buf_2_235/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_246 VDD VSS sky130_fd_sc_hd__buf_2_246/X sky130_fd_sc_hd__buf_2_246/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_257 VDD VSS sky130_fd_sc_hd__buf_2_257/X sky130_fd_sc_hd__inv_4_1/Y
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_268 VDD VSS sky130_fd_sc_hd__buf_2_268/X sky130_fd_sc_hd__buf_2_268/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_279 VDD VSS sky130_fd_sc_hd__buf_2_279/X sig_frequency[2]
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1220 VDD VSS sky130_fd_sc_hd__fa_2_1232/A sky130_fd_sc_hd__clkinv_8_78/Y
+ sky130_fd_sc_hd__mux2_2_195/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1231 VDD VSS sky130_fd_sc_hd__fa_2_1260/B sky130_fd_sc_hd__clkinv_8_63/Y
+ sky130_fd_sc_hd__mux2_2_219/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1242 VDD VSS sky130_fd_sc_hd__fa_2_1271/A sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__mux2_2_196/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1253 VDD VSS sky130_fd_sc_hd__mux2_2_213/A0 sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__nor2_1_245/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1264 VDD VSS sky130_fd_sc_hd__mux2_2_183/A1 sky130_fd_sc_hd__clkinv_8_116/Y
+ sky130_fd_sc_hd__o22ai_1_327/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1275 VDD VSS sky130_fd_sc_hd__mux2_2_214/A0 sky130_fd_sc_hd__clkinv_8_63/Y
+ sky130_fd_sc_hd__dfxtp_1_431/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1286 VDD VSS sky130_fd_sc_hd__mux2_2_206/A0 sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__o22ai_1_349/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1297 VDD VSS sky130_fd_sc_hd__mux2_2_178/A1 sky130_fd_sc_hd__clkinv_8_116/Y
+ sky130_fd_sc_hd__o22ai_1_338/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_880 VDD VSS sky130_fd_sc_hd__fa_2_862/A sky130_fd_sc_hd__dfxtp_1_902/CLK
+ sky130_fd_sc_hd__dfxtp_1_880/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_891 VDD VSS sky130_fd_sc_hd__fa_2_851/A sky130_fd_sc_hd__clkinv_4_22/Y
+ sky130_fd_sc_hd__dfxtp_1_891/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__or3_1_1 sky130_fd_sc_hd__or3_1_1/A sky130_fd_sc_hd__or3_1_1/X sky130_fd_sc_hd__or3_1_1/B
+ sky130_fd_sc_hd__or3_1_1/C VDD VSS VDD VSS sky130_fd_sc_hd__or3_1
Xsky130_fd_sc_hd__a21oi_1_15 sky130_fd_sc_hd__nor3_1_27/A sky130_fd_sc_hd__or2_0_0/B
+ sky130_fd_sc_hd__a21oi_1_15/Y sky130_fd_sc_hd__nor3_1_26/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_26 sky130_fd_sc_hd__nor2_1_37/B sky130_fd_sc_hd__nor3_1_36/Y
+ sky130_fd_sc_hd__a21oi_1_26/Y sky130_fd_sc_hd__nor2_1_37/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_37 sky130_fd_sc_hd__nor2_1_41/Y sky130_fd_sc_hd__o22ai_1_70/Y
+ sky130_fd_sc_hd__a21oi_1_37/Y sky130_fd_sc_hd__fa_2_1040/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_48 sky130_fd_sc_hd__nor2_2_6/Y sky130_fd_sc_hd__o22ai_1_80/Y
+ sky130_fd_sc_hd__a21oi_1_48/Y sky130_fd_sc_hd__fa_2_1036/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__fa_2_730 sky130_fd_sc_hd__fa_2_732/B sky130_fd_sc_hd__fa_2_730/SUM
+ sky130_fd_sc_hd__fa_2_826/A sky130_fd_sc_hd__fa_2_730/B sky130_fd_sc_hd__fa_2_730/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a21oi_1_59 sky130_fd_sc_hd__a21oi_1_59/A1 sky130_fd_sc_hd__nor2_1_48/B
+ sky130_fd_sc_hd__xnor2_1_60/A sky130_fd_sc_hd__xnor2_1_58/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__fa_2_741 sky130_fd_sc_hd__maj3_1_148/B sky130_fd_sc_hd__maj3_1_149/A
+ sky130_fd_sc_hd__fa_2_741/A sky130_fd_sc_hd__fa_2_741/B sky130_fd_sc_hd__fa_2_742/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_752 sky130_fd_sc_hd__maj3_1_145/B sky130_fd_sc_hd__maj3_1_146/A
+ sky130_fd_sc_hd__fa_2_752/A sky130_fd_sc_hd__fa_2_752/B sky130_fd_sc_hd__fa_2_753/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_763 sky130_fd_sc_hd__fa_2_764/A sky130_fd_sc_hd__fa_2_760/A
+ sky130_fd_sc_hd__fa_2_829/A sky130_fd_sc_hd__fa_2_823/B sky130_fd_sc_hd__fa_2_817/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_774 sky130_fd_sc_hd__fa_2_773/A sky130_fd_sc_hd__fa_2_774/SUM
+ sky130_fd_sc_hd__fa_2_820/B sky130_fd_sc_hd__ha_2_144/A sky130_fd_sc_hd__ha_2_140/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_785 sky130_fd_sc_hd__fa_2_784/A sky130_fd_sc_hd__fa_2_785/SUM
+ sky130_fd_sc_hd__ha_2_145/B sky130_fd_sc_hd__fa_2_793/A sky130_fd_sc_hd__ha_2_140/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_796 sky130_fd_sc_hd__fa_2_795/B sky130_fd_sc_hd__fa_2_796/SUM
+ sky130_fd_sc_hd__fa_2_796/A sky130_fd_sc_hd__fa_2_796/B sky130_fd_sc_hd__fa_2_796/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor3_1_7 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__nor3_1_7/Y
+ sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__nor3_2_2/C VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__buf_6_11 VDD VSS sky130_fd_sc_hd__buf_8_34/A sky130_fd_sc_hd__buf_6_11/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_22 VDD VSS sky130_fd_sc_hd__buf_6_22/X sky130_fd_sc_hd__buf_6_22/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_33 VDD VSS sky130_fd_sc_hd__buf_6_33/X sky130_fd_sc_hd__buf_6_33/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_44 VDD VSS sky130_fd_sc_hd__buf_6_44/X sky130_fd_sc_hd__inv_16_5/Y
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_55 VDD VSS sky130_fd_sc_hd__buf_6_55/X sky130_fd_sc_hd__buf_6_55/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_66 VDD VSS sky130_fd_sc_hd__buf_6_67/A sky130_fd_sc_hd__buf_6_66/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_77 VDD VSS sky130_fd_sc_hd__buf_6_77/X sky130_fd_sc_hd__buf_6_77/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_88 VDD VSS sky130_fd_sc_hd__buf_6_88/X sky130_fd_sc_hd__buf_6_88/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_13 sky130_fd_sc_hd__buf_2_123/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_24 sky130_fd_sc_hd__buf_4_34/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_309 sky130_fd_sc_hd__o21a_1_37/B1 sky130_fd_sc_hd__o21a_1_36/A1
+ sky130_fd_sc_hd__a21oi_1_309/Y sky130_fd_sc_hd__nor2_1_192/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_35 sky130_fd_sc_hd__buf_2_108/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_46 sky130_fd_sc_hd__buf_2_79/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_57 sky130_fd_sc_hd__buf_2_101/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_68 sky130_fd_sc_hd__clkbuf_4_88/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_79 sky130_fd_sc_hd__inv_12_0/Y VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__nand2_1_303 sky130_fd_sc_hd__nand2_1_303/Y sky130_fd_sc_hd__nor2_1_103/B
+ sky130_fd_sc_hd__fa_2_1111/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_902 sky130_fd_sc_hd__clkinv_1_902/Y sky130_fd_sc_hd__a21boi_1_3/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_902/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_250 sky130_fd_sc_hd__o22ai_1_265/A2 sky130_fd_sc_hd__o22ai_1_250/B1
+ sky130_fd_sc_hd__o22ai_1_250/Y sky130_fd_sc_hd__nor2_1_143/B sky130_fd_sc_hd__o32ai_1_2/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_314 sky130_fd_sc_hd__o21a_1_15/B1 sky130_fd_sc_hd__fa_2_1053/A
+ sky130_fd_sc_hd__o21a_1_15/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_913 sky130_fd_sc_hd__o22ai_1_308/A1 sky130_fd_sc_hd__fa_2_1181/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_913/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_261 sky130_fd_sc_hd__o22ai_1_261/A2 sky130_fd_sc_hd__nor2_1_153/B
+ sky130_fd_sc_hd__o22ai_1_261/Y sky130_fd_sc_hd__nor2_1_154/B sky130_fd_sc_hd__o32ai_1_2/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_325 sky130_fd_sc_hd__nand3_1_50/A sky130_fd_sc_hd__fa_2_1064/A
+ sky130_fd_sc_hd__a21o_2_5/A2 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_924 sky130_fd_sc_hd__o22ai_1_315/B1 sky130_fd_sc_hd__fa_2_1201/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_924/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_272 sky130_fd_sc_hd__nand2_1_410/Y sky130_fd_sc_hd__nand2_1_409/Y
+ sky130_fd_sc_hd__o22ai_1_272/Y sky130_fd_sc_hd__o22ai_1_285/A1 sky130_fd_sc_hd__a21o_2_14/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_336 sky130_fd_sc_hd__nor2_1_126/A sky130_fd_sc_hd__nand2_1_339/B
+ sky130_fd_sc_hd__nand2_2_6/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_935 sky130_fd_sc_hd__nor2_1_196/B sky130_fd_sc_hd__fa_2_1198/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_935/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_283 sky130_fd_sc_hd__nand2_1_412/Y sky130_fd_sc_hd__nand2_1_411/Y
+ sky130_fd_sc_hd__o22ai_1_283/Y sky130_fd_sc_hd__o22ai_1_283/A1 sky130_fd_sc_hd__a21o_2_13/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_347 sky130_fd_sc_hd__o21a_1_22/B1 sky130_fd_sc_hd__fa_2_1127/A
+ sky130_fd_sc_hd__o21a_1_22/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_294 sky130_fd_sc_hd__o32ai_1_4/B2 sky130_fd_sc_hd__nor2_1_224/A
+ sky130_fd_sc_hd__o22ai_1_294/Y sky130_fd_sc_hd__o22ai_1_319/A1 sky130_fd_sc_hd__a222oi_1_14/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_946 sky130_fd_sc_hd__clkinv_1_946/Y sky130_fd_sc_hd__o21a_1_55/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_946/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_358 sky130_fd_sc_hd__nand2_1_358/Y sky130_fd_sc_hd__nor2_1_161/B
+ sky130_fd_sc_hd__xnor2_1_93/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_957 sky130_fd_sc_hd__nor2_1_233/A sky130_fd_sc_hd__nor2_1_234/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_957/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_369 sky130_fd_sc_hd__a21o_2_7/A2 sky130_fd_sc_hd__nand2_1_369/B
+ sky130_fd_sc_hd__a21o_2_8/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_968 sky130_fd_sc_hd__o22ai_1_344/A1 sky130_fd_sc_hd__nor2_1_254/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_968/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_979 sky130_fd_sc_hd__o31ai_1_9/A3 sky130_fd_sc_hd__xnor2_1_1/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_979/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_110 VDD VSS sky130_fd_sc_hd__nand2_1_36/A sky130_fd_sc_hd__dfxtp_1_111/CLK
+ sky130_fd_sc_hd__ha_2_6/SUM VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_121 VDD VSS sky130_fd_sc_hd__ha_2_19/A sky130_fd_sc_hd__dfxtp_1_129/CLK
+ sky130_fd_sc_hd__and2_0_19/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_132 VDD VSS sky130_fd_sc_hd__ha_2_29/B sky130_fd_sc_hd__dfxtp_1_140/CLK
+ sky130_fd_sc_hd__nor2b_1_3/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_143 VDD VSS sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__dfxtp_1_143/CLK
+ sky130_fd_sc_hd__nor2b_1_2/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_154 VDD VSS sky130_fd_sc_hd__ha_2_33/A sky130_fd_sc_hd__dfxtp_1_158/CLK
+ sky130_fd_sc_hd__and2_0_35/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_165 VDD VSS sky130_fd_sc_hd__ha_2_44/A sky130_fd_sc_hd__clkinv_8_14/Y
+ sky130_fd_sc_hd__nor2b_2_0/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_176 VDD VSS sky130_fd_sc_hd__ha_2_58/A sky130_fd_sc_hd__dfxtp_1_185/CLK
+ sky130_fd_sc_hd__and2_0_52/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_187 VDD VSS sky130_fd_sc_hd__ha_2_69/A sky130_fd_sc_hd__dfxtp_1_195/CLK
+ sky130_fd_sc_hd__nor2b_1_35/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_198 VDD VSS sky130_fd_sc_hd__nor3_2_5/A sky130_fd_sc_hd__clkinv_2_17/Y
+ sky130_fd_sc_hd__a22o_1_17/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a21boi_1_8 sky130_fd_sc_hd__a21boi_1_8/Y sky130_fd_sc_hd__nor2_2_18/Y
+ sky130_fd_sc_hd__a21oi_1_465/Y sky130_fd_sc_hd__fa_2_1306/A VDD VSS VDD VSS sky130_fd_sc_hd__a21boi_1
Xsky130_fd_sc_hd__fa_2_1220 sky130_fd_sc_hd__fa_2_1221/CIN sky130_fd_sc_hd__mux2_2_148/A1
+ sky130_fd_sc_hd__fa_2_1220/A sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__fa_2_1220/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o211ai_1_18 sky130_fd_sc_hd__nor2_1_131/Y sky130_fd_sc_hd__nor2_1_126/A
+ sky130_fd_sc_hd__xor2_1_135/A sky130_fd_sc_hd__a22oi_1_355/Y sky130_fd_sc_hd__nand2_1_327/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__fa_2_1231 sky130_fd_sc_hd__fa_2_1232/CIN sky130_fd_sc_hd__mux2_2_198/A1
+ sky130_fd_sc_hd__fa_2_1231/A sky130_fd_sc_hd__fa_2_1231/B sky130_fd_sc_hd__fa_2_1231/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o211ai_1_29 sky130_fd_sc_hd__a21oi_1_275/Y sky130_fd_sc_hd__nor2_1_180/A
+ sky130_fd_sc_hd__xor2_1_179/A sky130_fd_sc_hd__a21oi_1_272/Y sky130_fd_sc_hd__nand2_1_381/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__fa_2_1242 sky130_fd_sc_hd__fa_2_1243/CIN sky130_fd_sc_hd__and2_0_330/A
+ sky130_fd_sc_hd__fa_2_1242/A sky130_fd_sc_hd__fa_2_1242/B sky130_fd_sc_hd__xor2_1_272/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1253 sky130_fd_sc_hd__fa_2_1254/CIN sky130_fd_sc_hd__mux2_2_186/A1
+ sky130_fd_sc_hd__fa_2_1253/A sky130_fd_sc_hd__fa_2_1253/B sky130_fd_sc_hd__fa_2_1253/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1264 sky130_fd_sc_hd__fa_2_1265/CIN sky130_fd_sc_hd__mux2_2_215/A1
+ sky130_fd_sc_hd__fa_2_1264/A sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1264/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1275 sky130_fd_sc_hd__fa_2_1276/CIN sky130_fd_sc_hd__and2_0_334/A
+ sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1275/B sky130_fd_sc_hd__xor2_1_296/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1286 sky130_fd_sc_hd__fa_2_1287/CIN sky130_fd_sc_hd__mux2_2_235/A1
+ sky130_fd_sc_hd__fa_2_1286/A sky130_fd_sc_hd__fa_2_1286/B sky130_fd_sc_hd__fa_2_1286/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1297 sky130_fd_sc_hd__fa_2_1298/CIN sky130_fd_sc_hd__mux2_2_254/A1
+ sky130_fd_sc_hd__fa_2_1297/A sky130_fd_sc_hd__fa_2_1297/B sky130_fd_sc_hd__fa_2_1297/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1050 VDD VSS sky130_fd_sc_hd__xor2_1_23/A sky130_fd_sc_hd__dfxtp_1_1050/CLK
+ sky130_fd_sc_hd__xnor2_1_94/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1061 VDD VSS sky130_fd_sc_hd__fa_2_1200/A sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__mux2_2_143/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_70 VSS VDD sky130_fd_sc_hd__nand2_2_3/Y sky130_fd_sc_hd__xnor2_1_60/Y
+ sky130_fd_sc_hd__a21oi_1_56/Y sky130_fd_sc_hd__o21ai_1_70/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1072 VDD VSS sky130_fd_sc_hd__fa_2_1174/A sky130_fd_sc_hd__clkinv_4_23/Y
+ sky130_fd_sc_hd__and2_0_327/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_81 VSS VDD sky130_fd_sc_hd__xnor2_1_59/A sky130_fd_sc_hd__nor2_1_62/Y
+ sky130_fd_sc_hd__o21ai_1_81/B1 sky130_fd_sc_hd__o21ai_1_81/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1083 VDD VSS sky130_fd_sc_hd__fa_2_1185/A sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__mux2_2_137/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_92 VSS VDD sky130_fd_sc_hd__o21ai_1_92/A2 sky130_fd_sc_hd__o21ai_1_92/A1
+ sky130_fd_sc_hd__o21ai_1_92/B1 sky130_fd_sc_hd__o21ai_1_92/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1094 VDD VSS sky130_fd_sc_hd__fa_2_1213/A sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__mux2_2_167/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o2bb2ai_1_12 sky130_fd_sc_hd__xnor2_1_12/B sky130_fd_sc_hd__nand2_1_202/B
+ sky130_fd_sc_hd__nor2_1_22/Y sky130_fd_sc_hd__nor2_1_22/Y sky130_fd_sc_hd__nand2_1_202/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__o2bb2ai_1_23 sky130_fd_sc_hd__dfxtp_1_552/D sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__dfxtp_1_552/Q sky130_fd_sc_hd__nand2_1_210/Y sky130_fd_sc_hd__nand2b_1_4/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_560 sky130_fd_sc_hd__fa_2_464/A sky130_fd_sc_hd__maj3_1_82/A
+ sky130_fd_sc_hd__fa_2_560/A sky130_fd_sc_hd__fa_2_560/B sky130_fd_sc_hd__fa_2_562/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_571 sky130_fd_sc_hd__fa_2_570/CIN sky130_fd_sc_hd__and2_0_89/A
+ sky130_fd_sc_hd__fa_2_571/A sky130_fd_sc_hd__fa_2_571/B sky130_fd_sc_hd__fa_2_571/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_582 sky130_fd_sc_hd__fa_2_581/CIN sky130_fd_sc_hd__fa_2_582/SUM
+ sky130_fd_sc_hd__fa_2_582/A sky130_fd_sc_hd__fa_2_582/B sky130_fd_sc_hd__maj3_1_108/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_593 sky130_fd_sc_hd__fa_2_595/B sky130_fd_sc_hd__fa_2_593/SUM
+ sky130_fd_sc_hd__ha_2_132/A sky130_fd_sc_hd__fa_2_624/B sky130_fd_sc_hd__fa_2_602/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_1_209 sky130_fd_sc_hd__clkinv_2_23/A sky130_fd_sc_hd__nor3_1_18/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_209/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_106 sky130_fd_sc_hd__fa_2_978/A sky130_fd_sc_hd__o22ai_1_119/Y
+ sky130_fd_sc_hd__a21oi_1_106/Y sky130_fd_sc_hd__nor2_4_10/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_117 sky130_fd_sc_hd__nand2_1_276/A sky130_fd_sc_hd__o22ai_1_125/Y
+ sky130_fd_sc_hd__a21oi_1_117/Y sky130_fd_sc_hd__a211o_1_3/A1 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_128 sky130_fd_sc_hd__a21o_2_3/A2 sky130_fd_sc_hd__o21ai_1_152/Y
+ sky130_fd_sc_hd__a21oi_1_128/Y sky130_fd_sc_hd__fa_2_1000/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_139 sky130_fd_sc_hd__nor2_2_10/Y sky130_fd_sc_hd__o22ai_1_139/Y
+ sky130_fd_sc_hd__a21oi_1_139/Y sky130_fd_sc_hd__fa_2_1111/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nor2_1_303 sky130_fd_sc_hd__o21a_1_68/A1 sky130_fd_sc_hd__nor2_1_303/Y
+ sky130_fd_sc_hd__nor2_1_303/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_314 sky130_fd_sc_hd__nor2_1_314/B sky130_fd_sc_hd__nor2_1_314/Y
+ sky130_fd_sc_hd__nor2_1_314/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_510 sky130_fd_sc_hd__buf_12_510/A sky130_fd_sc_hd__buf_12_510/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_402 sky130_fd_sc_hd__nor2_1_307/Y sky130_fd_sc_hd__nor2_1_309/Y
+ sky130_fd_sc_hd__fa_2_1301/A sky130_fd_sc_hd__fa_2_1297/A sky130_fd_sc_hd__a22oi_1_402/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkbuf_8_2 sky130_fd_sc_hd__buf_2_147/A sky130_fd_sc_hd__dfxtp_1_93/D
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkbuf_8
Xsky130_fd_sc_hd__nand2_1_100 sky130_fd_sc_hd__nand2_1_100/Y sky130_fd_sc_hd__nand2_1_101/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_111 sky130_fd_sc_hd__nand2_1_111/Y sky130_fd_sc_hd__nand2_1_111/B
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_710 sky130_fd_sc_hd__nor2_1_119/B sky130_fd_sc_hd__fa_2_1054/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_710/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_122 sky130_fd_sc_hd__nand2_1_122/Y sky130_fd_sc_hd__fa_2_704/SUM
+ sky130_fd_sc_hd__and2_0_235/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_721 sky130_fd_sc_hd__nor2_1_118/B sky130_fd_sc_hd__fa_2_1056/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_721/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_133 sky130_fd_sc_hd__nand2_1_133/Y sky130_fd_sc_hd__nand2_1_134/Y
+ sky130_fd_sc_hd__buf_2_264/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_732 sky130_fd_sc_hd__o21ai_1_253/A1 sky130_fd_sc_hd__a211o_1_9/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_732/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_144 sky130_fd_sc_hd__nand2_1_144/Y sky130_fd_sc_hd__fa_2_715/SUM
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_743 sky130_fd_sc_hd__o21ai_1_270/A2 sky130_fd_sc_hd__fa_2_1077/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_743/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_155 sky130_fd_sc_hd__fa_2_124/CIN sky130_fd_sc_hd__fa_2_9/A
+ sky130_fd_sc_hd__fa_2_5/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_754 sky130_fd_sc_hd__ha_2_186/B sky130_fd_sc_hd__a22o_1_72/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_754/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_166 sky130_fd_sc_hd__fa_2_279/B sky130_fd_sc_hd__fa_2_266/B
+ sky130_fd_sc_hd__ha_2_97/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_765 sky130_fd_sc_hd__ha_2_198/B sky130_fd_sc_hd__fa_2_1109/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_765/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_177 sky130_fd_sc_hd__fa_2_469/B sky130_fd_sc_hd__fa_2_543/A
+ sky130_fd_sc_hd__fa_2_537/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_776 sky130_fd_sc_hd__mux2_2_75/S sky130_fd_sc_hd__or2_0_7/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_776/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_188 sky130_fd_sc_hd__fa_2_642/A sky130_fd_sc_hd__fa_2_683/B
+ sky130_fd_sc_hd__ha_2_128/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_787 sky130_fd_sc_hd__o32ai_1_0/A3 sky130_fd_sc_hd__fa_2_1123/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_787/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_199 sky130_fd_sc_hd__fa_2_817/CIN sky130_fd_sc_hd__ha_2_141/A
+ sky130_fd_sc_hd__ha_2_142/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_798 sky130_fd_sc_hd__o22ai_1_224/A1 sky130_fd_sc_hd__a21o_2_6/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_798/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor2_1_4 sky130_fd_sc_hd__xor2_1_4/B sky130_fd_sc_hd__xor2_1_4/X
+ sky130_fd_sc_hd__xor2_1_4/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand3_2_5 sky130_fd_sc_hd__or2_1_2/A sky130_fd_sc_hd__nand3_2_5/Y
+ sky130_fd_sc_hd__nor2_1_7/A sky130_fd_sc_hd__nor2_1_7/B VSS VDD VSS VDD sky130_fd_sc_hd__nand3_2
Xsky130_fd_sc_hd__clkinv_8_2 sky130_fd_sc_hd__clkinv_8_3/A sky130_fd_sc_hd__clkinv_8_2/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_2/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__xor2_1_19 sky130_fd_sc_hd__xor2_1_19/B sky130_fd_sc_hd__nor4_1_3/B
+ sky130_fd_sc_hd__ha_2_152/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nor3_1_10 sky130_fd_sc_hd__nor2_4_6/A sky130_fd_sc_hd__nor3_1_10/Y
+ sky130_fd_sc_hd__nor3_1_9/B sky130_fd_sc_hd__nor3_2_4/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_21 sky130_fd_sc_hd__nor3_1_21/C sky130_fd_sc_hd__nor3_1_21/Y
+ sky130_fd_sc_hd__nor3_2_9/A sky130_fd_sc_hd__nor3_2_8/A VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_32 sky130_fd_sc_hd__nor3_1_32/C sky130_fd_sc_hd__nor3_1_32/Y
+ sky130_fd_sc_hd__or4_1_2/A sky130_fd_sc_hd__nor4_1_5/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__a21o_2_9 sky130_fd_sc_hd__a21o_2_9/X sky130_fd_sc_hd__a21o_2_9/B1
+ sky130_fd_sc_hd__a21o_2_9/A1 sky130_fd_sc_hd__a21o_2_9/A2 VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__fa_2_1050 sky130_fd_sc_hd__fa_2_1051/CIN sky130_fd_sc_hd__and2_0_313/A
+ sky130_fd_sc_hd__fa_2_1050/A sky130_fd_sc_hd__fa_2_1050/B sky130_fd_sc_hd__fa_2_1050/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1061 sky130_fd_sc_hd__fa_2_1062/CIN sky130_fd_sc_hd__mux2_2_55/A0
+ sky130_fd_sc_hd__fa_2_1061/A sky130_fd_sc_hd__xor2_1_96/X sky130_fd_sc_hd__fa_2_1061/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1072 sky130_fd_sc_hd__fa_2_1073/CIN sky130_fd_sc_hd__and2_0_311/A
+ sky130_fd_sc_hd__fa_2_1072/A sky130_fd_sc_hd__fa_2_1072/B sky130_fd_sc_hd__fa_2_1072/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1083 sky130_fd_sc_hd__fa_2_1084/CIN sky130_fd_sc_hd__mux2_2_56/A0
+ sky130_fd_sc_hd__fa_2_1083/A sky130_fd_sc_hd__fa_2_1083/B sky130_fd_sc_hd__fa_2_1083/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1094 sky130_fd_sc_hd__fa_2_1095/CIN sky130_fd_sc_hd__and2_0_296/A
+ sky130_fd_sc_hd__fa_2_1094/A sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1094/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_70 sky130_fd_sc_hd__inv_2_70/A sky130_fd_sc_hd__inv_2_70/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_81 sky130_fd_sc_hd__inv_2_81/A sky130_fd_sc_hd__inv_2_81/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_92 sky130_fd_sc_hd__inv_2_92/A sky130_fd_sc_hd__inv_2_92/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__ha_2_13 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_13/A sky130_fd_sc_hd__ha_2_12/B
+ sky130_fd_sc_hd__ha_2_13/SUM sky130_fd_sc_hd__ha_2_13/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_24 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_24/A sky130_fd_sc_hd__ha_2_23/B
+ sky130_fd_sc_hd__ha_2_24/SUM sky130_fd_sc_hd__ha_2_24/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_35 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_35/A sky130_fd_sc_hd__ha_2_34/B
+ sky130_fd_sc_hd__ha_2_35/SUM sky130_fd_sc_hd__ha_2_35/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_46 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_46/A sky130_fd_sc_hd__ha_2_45/B
+ sky130_fd_sc_hd__ha_2_46/SUM sky130_fd_sc_hd__ha_2_46/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_57 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_57/A sky130_fd_sc_hd__ha_2_56/B
+ sky130_fd_sc_hd__ha_2_57/SUM sky130_fd_sc_hd__ha_2_57/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_68 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_68/A sky130_fd_sc_hd__ha_2_67/B
+ sky130_fd_sc_hd__ha_2_68/SUM sky130_fd_sc_hd__ha_2_68/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_79 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_79/A sky130_fd_sc_hd__ha_2_78/B
+ sky130_fd_sc_hd__ha_2_79/SUM sky130_fd_sc_hd__ha_2_79/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__sdlclkp_4_20 sky130_fd_sc_hd__conb_1_12/LO sky130_fd_sc_hd__clkinv_2_7/Y
+ sky130_fd_sc_hd__dfxtp_1_185/CLK sky130_fd_sc_hd__nand3b_1_0/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_390 sky130_fd_sc_hd__fa_2_392/CIN sky130_fd_sc_hd__fa_2_387/A
+ sky130_fd_sc_hd__fa_2_390/A sky130_fd_sc_hd__fa_2_390/B sky130_fd_sc_hd__fa_2_398/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22oi_2_1 sky130_fd_sc_hd__nor3_2_0/A sky130_fd_sc_hd__buf_2_279/X
+ sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__nand4_1_34/Y sky130_fd_sc_hd__a22oi_2_1/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__sdlclkp_4_31 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_96/A
+ sky130_fd_sc_hd__dfxtp_1_472/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__clkbuf_16_13 sky130_fd_sc_hd__buf_12_510/A sky130_fd_sc_hd__clkinv_1_248/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__clkbuf_1_9 VSS VDD sky130_fd_sc_hd__buf_6_7/A sky130_fd_sc_hd__clkbuf_1_9/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__sdlclkp_4_42 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_72/A
+ sky130_fd_sc_hd__dfxtp_1_391/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_53 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_53/A
+ sky130_fd_sc_hd__dfxtp_1_266/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_64 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__clkinv_8_61/Y
+ sky130_fd_sc_hd__dfxtp_1_576/CLK sky130_fd_sc_hd__nand2b_1_5/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_75 sky130_fd_sc_hd__conb_1_24/LO sky130_fd_sc_hd__clkinv_8_53/A
+ sky130_fd_sc_hd__dfxtp_1_755/CLK sky130_fd_sc_hd__or2_0_8/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_86 sky130_fd_sc_hd__conb_1_27/LO sky130_fd_sc_hd__clkinv_8_118/Y
+ sky130_fd_sc_hd__dfxtp_1_1180/CLK sky130_fd_sc_hd__or2_0_11/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_100 sky130_fd_sc_hd__nor2_1_100/B sky130_fd_sc_hd__nor2_1_97/A
+ sky130_fd_sc_hd__fa_2_1117/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_111 sky130_fd_sc_hd__nor2_1_111/B sky130_fd_sc_hd__nor2_1_111/Y
+ sky130_fd_sc_hd__fa_2_1118/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_122 sky130_fd_sc_hd__nor2_1_123/B sky130_fd_sc_hd__nor2_1_122/Y
+ sky130_fd_sc_hd__nor2_2_13/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_133 sky130_fd_sc_hd__nor2_1_133/B sky130_fd_sc_hd__nor2_1_133/Y
+ sky130_fd_sc_hd__nor2_1_133/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_20 sky130_fd_sc_hd__nor2_2_0/Y sky130_fd_sc_hd__clkinv_1_4/Y
+ sky130_fd_sc_hd__nand4_1_21/Y sky130_fd_sc_hd__nand4_1_5/Y sky130_fd_sc_hd__a22oi_1_20/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_144 sky130_fd_sc_hd__nor2_1_144/B sky130_fd_sc_hd__o21a_1_19/A1
+ sky130_fd_sc_hd__o21a_1_20/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_31 sky130_fd_sc_hd__clkbuf_4_8/X sky130_fd_sc_hd__clkbuf_4_9/X
+ sky130_fd_sc_hd__clkbuf_1_33/X sky130_fd_sc_hd__a22oi_1_31/A2 sky130_fd_sc_hd__a22oi_1_31/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_155 sky130_fd_sc_hd__nor2_1_155/B sky130_fd_sc_hd__nor2_1_155/Y
+ sky130_fd_sc_hd__o21a_1_28/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_1_9 sky130_fd_sc_hd__and2_0_17/A sky130_fd_sc_hd__inv_2_3/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_9/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22oi_1_42 sky130_fd_sc_hd__a22oi_2_9/B1 sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__clkbuf_4_38/X sky130_fd_sc_hd__a22oi_1_42/A2 sky130_fd_sc_hd__a22oi_1_42/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_166 sky130_fd_sc_hd__a21o_2_6/A2 sky130_fd_sc_hd__a21o_2_6/B1
+ sky130_fd_sc_hd__a21o_2_6/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_53 sky130_fd_sc_hd__a22oi_1_81/B1 sky130_fd_sc_hd__clkbuf_1_99/X
+ sky130_fd_sc_hd__clkbuf_1_43/X sky130_fd_sc_hd__clkbuf_4_18/X sky130_fd_sc_hd__nand4_1_7/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_177 sky130_fd_sc_hd__nor2_1_183/A sky130_fd_sc_hd__nor2_1_177/Y
+ sky130_fd_sc_hd__nor2_1_178/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_188 sky130_fd_sc_hd__nor2_1_188/B sky130_fd_sc_hd__o21a_1_34/A1
+ sky130_fd_sc_hd__nor2_1_188/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_64 sky130_fd_sc_hd__clkbuf_4_8/X sky130_fd_sc_hd__clkbuf_4_9/X
+ sky130_fd_sc_hd__clkbuf_1_23/X sky130_fd_sc_hd__a22oi_1_64/A2 sky130_fd_sc_hd__a22oi_1_64/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_199 sky130_fd_sc_hd__nor2_1_199/B sky130_fd_sc_hd__nor2_1_199/Y
+ sky130_fd_sc_hd__nor2_1_199/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_75 sky130_fd_sc_hd__a22oi_2_9/B1 sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__clkbuf_4_28/X sky130_fd_sc_hd__a22oi_1_75/A2 sky130_fd_sc_hd__a22oi_1_75/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_86 sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__a22oi_2_12/A1
+ sky130_fd_sc_hd__buf_2_81/X sky130_fd_sc_hd__a22oi_1_86/A2 sky130_fd_sc_hd__a22oi_1_86/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_97 sky130_fd_sc_hd__a22oi_1_97/B1 sky130_fd_sc_hd__a22oi_1_97/A1
+ sky130_fd_sc_hd__buf_2_62/X sky130_fd_sc_hd__clkbuf_4_86/X sky130_fd_sc_hd__nand4_1_19/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_340 sky130_fd_sc_hd__buf_8_168/X sky130_fd_sc_hd__buf_12_340/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_351 sky130_fd_sc_hd__buf_6_45/X sky130_fd_sc_hd__buf_12_351/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_210 sky130_fd_sc_hd__clkbuf_1_264/X sky130_fd_sc_hd__nor2_2_3/Y
+ sky130_fd_sc_hd__a22oi_1_210/B2 sky130_fd_sc_hd__clkbuf_4_122/X sky130_fd_sc_hd__nand4_1_47/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_362 sky130_fd_sc_hd__buf_12_362/A sky130_fd_sc_hd__buf_8_174/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_221 sky130_fd_sc_hd__buf_2_166/X sky130_fd_sc_hd__buf_2_167/X
+ sky130_fd_sc_hd__clkbuf_1_521/X sky130_fd_sc_hd__buf_2_179/X sky130_fd_sc_hd__nand4_1_52/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_373 sky130_fd_sc_hd__buf_12_373/A sky130_fd_sc_hd__buf_12_375/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_232 sky130_fd_sc_hd__buf_2_166/X sky130_fd_sc_hd__buf_2_167/X
+ sky130_fd_sc_hd__clkbuf_1_433/X sky130_fd_sc_hd__buf_2_176/X sky130_fd_sc_hd__nand4_1_55/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_384 sky130_fd_sc_hd__inv_2_114/Y sky130_fd_sc_hd__buf_12_498/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_243 sky130_fd_sc_hd__buf_2_164/X sky130_fd_sc_hd__nor2_4_8/Y
+ sky130_fd_sc_hd__clkbuf_1_417/X sky130_fd_sc_hd__buf_2_226/X sky130_fd_sc_hd__nand4_1_59/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_395 sky130_fd_sc_hd__buf_12_395/A sky130_fd_sc_hd__buf_12_511/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_254 sky130_fd_sc_hd__a22oi_2_25/B1 sky130_fd_sc_hd__a22oi_2_25/A1
+ sky130_fd_sc_hd__clkbuf_1_382/X sky130_fd_sc_hd__a22oi_1_254/A2 sky130_fd_sc_hd__a22oi_1_254/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_265 sky130_fd_sc_hd__clkbuf_4_165/X sky130_fd_sc_hd__clkinv_2_23/Y
+ sky130_fd_sc_hd__clkbuf_1_411/X sky130_fd_sc_hd__a22oi_1_265/A2 sky130_fd_sc_hd__a22oi_1_265/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_276 sky130_fd_sc_hd__clkbuf_1_376/X sky130_fd_sc_hd__nor2_2_5/Y
+ sky130_fd_sc_hd__buf_2_213/X sky130_fd_sc_hd__clkbuf_1_469/X sky130_fd_sc_hd__nand4_1_68/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_287 sky130_fd_sc_hd__nor2_2_4/Y sky130_fd_sc_hd__clkbuf_1_377/X
+ sky130_fd_sc_hd__a22oi_1_287/B2 sky130_fd_sc_hd__clkbuf_4_185/X sky130_fd_sc_hd__nand4_1_71/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_4_105 VDD VSS sky130_fd_sc_hd__buf_4_105/X sky130_fd_sc_hd__buf_4_105/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__a22oi_1_298 sky130_fd_sc_hd__clkbuf_1_378/X sky130_fd_sc_hd__clkbuf_1_379/X
+ sky130_fd_sc_hd__clkbuf_4_168/X sky130_fd_sc_hd__buf_2_192/X sky130_fd_sc_hd__nand4_1_74/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_4_116 VDD VSS sky130_fd_sc_hd__buf_4_116/X sky130_fd_sc_hd__buf_4_116/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__clkinv_1_540 sky130_fd_sc_hd__nor2_1_63/B sky130_fd_sc_hd__fa_2_989/A
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_551 sky130_fd_sc_hd__nor2_1_65/B sky130_fd_sc_hd__fa_2_985/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_551/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_562 sky130_fd_sc_hd__nor2_1_70/A sky130_fd_sc_hd__fa_2_975/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_562/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_573 sky130_fd_sc_hd__nand2_1_276/A sky130_fd_sc_hd__a211oi_1_6/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_573/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_584 sky130_fd_sc_hd__nand2_2_4/B sky130_fd_sc_hd__nand2_1_282/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_584/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_595 sky130_fd_sc_hd__ha_2_170/B sky130_fd_sc_hd__a22o_1_67/A2
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_4_20 sky130_fd_sc_hd__clkinv_8_38/A sky130_fd_sc_hd__clkinv_4_20/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_20/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_31 sky130_fd_sc_hd__clkinv_4_31/A sky130_fd_sc_hd__clkinv_4_31/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_31/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_42 sky130_fd_sc_hd__clkinv_8_80/Y sky130_fd_sc_hd__clkinv_8_81/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_42/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_53 sky130_fd_sc_hd__clkinv_4_53/A sky130_fd_sc_hd__clkinv_4_53/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_53/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_64 sky130_fd_sc_hd__clkinv_4_64/A sky130_fd_sc_hd__clkinv_4_64/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_64/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_75 sky130_fd_sc_hd__clkinv_8_18/A sky130_fd_sc_hd__clkinv_4_75/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_75/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__inv_16_5 sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_5/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__a21oi_1_470 sky130_fd_sc_hd__fa_2_1310/A sky130_fd_sc_hd__nor2_1_305/Y
+ sky130_fd_sc_hd__a21oi_1_470/Y sky130_fd_sc_hd__nor3_1_41/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_481 sky130_fd_sc_hd__nor2_1_311/A sky130_fd_sc_hd__nor2_1_311/Y
+ sky130_fd_sc_hd__a21oi_1_481/Y sky130_fd_sc_hd__nor4_1_13/D VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_492 sky130_fd_sc_hd__nor2_1_319/Y sky130_fd_sc_hd__or2_0_0/B
+ sky130_fd_sc_hd__nand2_1_560/A sky130_fd_sc_hd__nor2_1_317/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__xor2_1_303 sky130_fd_sc_hd__nor2_4_20/Y sky130_fd_sc_hd__fa_2_1307/B
+ sky130_fd_sc_hd__xor2_1_303/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_314 sky130_fd_sc_hd__nor2_4_20/Y sky130_fd_sc_hd__fa_2_1296/B
+ sky130_fd_sc_hd__xor2_1_314/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_709 VDD VSS sky130_fd_sc_hd__mux2_2_15/A1 sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__o21ai_1_49/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_307 VSS VDD sky130_fd_sc_hd__nand4_1_38/D sky130_fd_sc_hd__a22oi_1_171/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_318 VSS VDD sky130_fd_sc_hd__buf_8_133/A sky130_fd_sc_hd__and2_0_36/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_329 VSS VDD sky130_fd_sc_hd__buf_4_57/A sky130_fd_sc_hd__dfxtp_1_1463/Q
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_11 VDD VSS sky130_fd_sc_hd__dfxtp_1_11/Q sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__a22o_1_8/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_22 VDD VSS sky130_fd_sc_hd__ha_2_114/B sky130_fd_sc_hd__dfxtp_1_26/CLK
+ sky130_fd_sc_hd__buf_2_290/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_33 VDD VSS sky130_fd_sc_hd__fa_2_904/CIN sky130_fd_sc_hd__dfxtp_1_39/CLK
+ sky130_fd_sc_hd__nand4_1_35/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_44 VDD VSS sky130_fd_sc_hd__fa_2_915/CIN sky130_fd_sc_hd__clkinv_4_80/Y
+ sky130_fd_sc_hd__dfxtp_1_60/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_55 VDD VSS sky130_fd_sc_hd__ha_2_119/B sky130_fd_sc_hd__dfxtp_1_60/CLK
+ sky130_fd_sc_hd__buf_2_289/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_66 VDD VSS sky130_fd_sc_hd__fa_2_67/B sky130_fd_sc_hd__dfxtp_1_73/CLK
+ sky130_fd_sc_hd__dfxtp_1_66/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_77 VDD VSS sky130_fd_sc_hd__fa_2_5/A sky130_fd_sc_hd__dfxtp_1_77/CLK
+ sky130_fd_sc_hd__dfxtp_1_77/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_88 VDD VSS sky130_fd_sc_hd__a22o_1_4/B2 sky130_fd_sc_hd__dfxtp_1_93/CLK
+ sky130_fd_sc_hd__buf_6_55/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_99 VDD VSS sky130_fd_sc_hd__ha_2_5/A sky130_fd_sc_hd__dfxtp_1_99/CLK
+ sky130_fd_sc_hd__and2_0_10/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_4_101 sky130_fd_sc_hd__clkbuf_4_101/X sky130_fd_sc_hd__buf_8_103/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_112 sky130_fd_sc_hd__clkbuf_4_112/X sky130_fd_sc_hd__nor3_1_16/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_123 sky130_fd_sc_hd__clkbuf_4_123/X sky130_fd_sc_hd__clkbuf_4_123/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_134 sky130_fd_sc_hd__clkbuf_4_134/X sky130_fd_sc_hd__clkbuf_4_134/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_305 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_305/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_305/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_145 sky130_fd_sc_hd__nand4_1_40/B sky130_fd_sc_hd__a22oi_1_181/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_316 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_316/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_316/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_156 sky130_fd_sc_hd__inv_2_79/A sky130_fd_sc_hd__a22o_1_13/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_327 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_327/X sky130_fd_sc_hd__mux2_2_171/S
+ sky130_fd_sc_hd__and2_0_327/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_167 sky130_fd_sc_hd__clkbuf_4_167/X sky130_fd_sc_hd__clkbuf_4_167/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_338 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_338/X sky130_fd_sc_hd__buf_2_263/X
+ sky130_fd_sc_hd__nor3_1_41/C sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_178 sky130_fd_sc_hd__clkbuf_4_178/X sky130_fd_sc_hd__clkbuf_4_178/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_349 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_349/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_349/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_189 sky130_fd_sc_hd__clkbuf_4_189/X sky130_fd_sc_hd__clkbuf_4_189/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__inv_2_105 sky130_fd_sc_hd__inv_2_105/A sky130_fd_sc_hd__inv_2_105/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_116 sky130_fd_sc_hd__inv_2_116/A sky130_fd_sc_hd__inv_2_117/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__or2_0_7 sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__or2_0_7/X sky130_fd_sc_hd__or2_0_7/B
+ VSS VDD VSS VDD sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__inv_2_127 sky130_fd_sc_hd__inv_2_127/A sky130_fd_sc_hd__inv_2_127/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_138 sky130_fd_sc_hd__nor2_4_15/A sky130_fd_sc_hd__mux2_2_99/S
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_12_170 sky130_fd_sc_hd__buf_8_107/X sky130_fd_sc_hd__buf_6_29/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_181 sky130_fd_sc_hd__buf_8_106/X sky130_fd_sc_hd__buf_12_181/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_192 sky130_fd_sc_hd__buf_4_44/X sky130_fd_sc_hd__buf_12_192/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_370 sky130_fd_sc_hd__fa_2_758/B sky130_fd_sc_hd__fa_2_801/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_370/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_381 sky130_fd_sc_hd__fa_2_867/B sky130_fd_sc_hd__dfxtp_1_267/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_381/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_392 sky130_fd_sc_hd__fa_2_880/B sky130_fd_sc_hd__nand2_1_34/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_392/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_2_0 sky130_fd_sc_hd__nor3_1_28/B sky130_fd_sc_hd__a21oi_2_0/A2
+ sky130_fd_sc_hd__maj3_1_0/X sky130_fd_sc_hd__a21oi_2_0/Y VSS VDD VSS VDD sky130_fd_sc_hd__a21oi_2
Xsky130_fd_sc_hd__a211o_1_6 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_78/A sky130_fd_sc_hd__a211o_1_6/A2
+ sky130_fd_sc_hd__nor2_1_75/Y sky130_fd_sc_hd__a211o_1_6/A1 sky130_fd_sc_hd__o22ai_1_94/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o21a_1_11 sky130_fd_sc_hd__o21a_1_11/X sky130_fd_sc_hd__o21a_1_11/A1
+ sky130_fd_sc_hd__o21a_1_11/B1 sky130_fd_sc_hd__fa_2_1062/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21ai_1_306 VSS VDD sky130_fd_sc_hd__nor2_1_172/A sky130_fd_sc_hd__o21ai_1_306/A1
+ sky130_fd_sc_hd__a211oi_1_13/Y sky130_fd_sc_hd__xor2_1_181/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_317 VSS VDD sky130_fd_sc_hd__o22ai_1_262/A1 sky130_fd_sc_hd__nor2_1_153/B
+ sky130_fd_sc_hd__o21ai_1_317/B1 sky130_fd_sc_hd__o21ai_1_317/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_22 sky130_fd_sc_hd__o21a_1_22/X sky130_fd_sc_hd__o21a_1_22/A1
+ sky130_fd_sc_hd__o21a_1_22/B1 sky130_fd_sc_hd__fa_2_1127/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_33 sky130_fd_sc_hd__o21a_1_33/X sky130_fd_sc_hd__o21a_1_33/A1
+ sky130_fd_sc_hd__o21a_1_33/B1 sky130_fd_sc_hd__fa_2_1183/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21ai_1_328 VSS VDD sky130_fd_sc_hd__o22ai_1_261/A2 sky130_fd_sc_hd__o21ai_1_328/A1
+ sky130_fd_sc_hd__a21oi_1_297/Y sky130_fd_sc_hd__o21ai_1_328/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_339 VSS VDD sky130_fd_sc_hd__nor2_1_198/B sky130_fd_sc_hd__o22ai_1_322/A2
+ sky130_fd_sc_hd__a22oi_1_379/Y sky130_fd_sc_hd__o21ai_1_339/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_44 sky130_fd_sc_hd__o21a_1_44/X sky130_fd_sc_hd__o21a_1_44/A1
+ sky130_fd_sc_hd__o21a_1_44/B1 sky130_fd_sc_hd__fa_2_1238/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_55 sky130_fd_sc_hd__o21a_1_55/X sky130_fd_sc_hd__o21a_1_55/A1
+ sky130_fd_sc_hd__o21a_1_55/B1 sky130_fd_sc_hd__o21a_1_55/A2 VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_66 sky130_fd_sc_hd__o21a_1_66/X sky130_fd_sc_hd__o21a_1_66/A1
+ sky130_fd_sc_hd__o21a_1_66/B1 sky130_fd_sc_hd__fa_2_1301/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__mux2_2_19 VSS VDD sky130_fd_sc_hd__mux2_2_19/A1 sky130_fd_sc_hd__mux2_2_19/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_19/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__xor2_1_100 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1057/B
+ sky130_fd_sc_hd__xor2_1_100/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_111 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__xor2_1_111/X
+ sky130_fd_sc_hd__xor2_1_111/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_122 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1084/B
+ sky130_fd_sc_hd__xor2_1_122/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_133 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1073/B
+ sky130_fd_sc_hd__xor2_1_133/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_144 sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__fa_2_1139/B
+ sky130_fd_sc_hd__xor2_1_144/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_155 sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__fa_2_1128/B
+ sky130_fd_sc_hd__xor2_1_155/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_506 VDD VSS sky130_fd_sc_hd__nor4_1_12/B sky130_fd_sc_hd__edfxtp_1_0/CLK
+ sky130_fd_sc_hd__a22o_1_65/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_166 sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__fa_2_1156/B
+ sky130_fd_sc_hd__xor2_1_166/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_517 VDD VSS sky130_fd_sc_hd__nor4_1_10/A sky130_fd_sc_hd__dfxtp_1_520/CLK
+ sky130_fd_sc_hd__a22o_1_54/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_177 sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__fa_2_1145/B
+ sky130_fd_sc_hd__xor2_1_177/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_188 sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__xor2_1_188/X
+ sky130_fd_sc_hd__xor2_1_208/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_528 VDD VSS sky130_fd_sc_hd__fa_2_963/A sky130_fd_sc_hd__dfxtp_1_533/CLK
+ sky130_fd_sc_hd__and2_0_262/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_539 VDD VSS sky130_fd_sc_hd__fa_2_952/A sky130_fd_sc_hd__dfxtp_1_544/CLK
+ sky130_fd_sc_hd__a22o_1_46/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_199 sky130_fd_sc_hd__fa_2_1173/A sky130_fd_sc_hd__fa_2_1180/B
+ sky130_fd_sc_hd__xor2_1_199/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_104 VSS VDD sky130_fd_sc_hd__buf_12_10/A sky130_fd_sc_hd__ha_2_16/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_115 VSS VDD sky130_fd_sc_hd__buf_4_13/A sky130_fd_sc_hd__buf_12_82/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_126 VSS VDD sky130_fd_sc_hd__clkbuf_1_126/X sky130_fd_sc_hd__nand3_1_22/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_137 VSS VDD sky130_fd_sc_hd__a22oi_1_96/B1 sky130_fd_sc_hd__nor3_1_10/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_148 VSS VDD sky130_fd_sc_hd__clkbuf_1_148/X sky130_fd_sc_hd__clkbuf_1_148/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_159 VSS VDD sky130_fd_sc_hd__clkbuf_1_159/X sky130_fd_sc_hd__clkbuf_1_159/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_6 VDD VSS sky130_fd_sc_hd__dfxtp_1_6/Q sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__a22o_1_3/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand3_1_15 sky130_fd_sc_hd__nand3_1_15/Y sky130_fd_sc_hd__nand3_1_15/A
+ sky130_fd_sc_hd__nand3_1_15/C sky130_fd_sc_hd__a22oi_2_3/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_26 sky130_fd_sc_hd__nand3_1_26/Y sky130_fd_sc_hd__nand2_2_0/B
+ sky130_fd_sc_hd__xor2_1_4/B sky130_fd_sc_hd__ha_2_40/A VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_37 sky130_fd_sc_hd__nand3_1_37/Y sky130_fd_sc_hd__nor2_1_7/B
+ sky130_fd_sc_hd__or2_1_2/X sky130_fd_sc_hd__nor2_1_7/A VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_48 sky130_fd_sc_hd__nand3_1_48/Y sky130_fd_sc_hd__nand3_1_48/A
+ sky130_fd_sc_hd__nand3_1_48/C sky130_fd_sc_hd__nand3_1_48/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__dfxtp_1_1402 VDD VSS sky130_fd_sc_hd__mux2_2_238/A0 sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__o22ai_1_387/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1413 VDD VSS sky130_fd_sc_hd__mux2_2_265/A0 sky130_fd_sc_hd__clkinv_8_102/Y
+ sky130_fd_sc_hd__dfxtp_1_428/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1424 VDD VSS sky130_fd_sc_hd__nand2_1_520/B sky130_fd_sc_hd__clkinv_8_75/Y
+ sky130_fd_sc_hd__xnor2_1_99/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1435 VDD VSS sky130_fd_sc_hd__mux2_2_232/A0 sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__o22ai_1_398/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1446 VDD VSS sky130_fd_sc_hd__nand3_1_52/B sky130_fd_sc_hd__clkinv_8_116/Y
+ sky130_fd_sc_hd__nor2b_1_134/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1457 VDD VSS sky130_fd_sc_hd__buf_6_89/A sky130_fd_sc_hd__dfxtp_1_1464/CLK
+ sky130_fd_sc_hd__and2_0_351/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1468 VDD VSS sky130_fd_sc_hd__nor2_1_323/A sky130_fd_sc_hd__clkinv_2_41/Y
+ sky130_fd_sc_hd__nor2b_1_142/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_102 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_102/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__xor2_1_23/X sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_10 sky130_fd_sc_hd__nor2b_1_3/B_N sky130_fd_sc_hd__ha_2_29/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_10/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_113 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_113/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_851/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_21 sky130_fd_sc_hd__inv_2_10/A sky130_fd_sc_hd__clkinv_1_21/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_21/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_124 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_124/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_853/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_32 sky130_fd_sc_hd__inv_2_21/A sky130_fd_sc_hd__buf_8_43/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_32/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_135 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_135/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_922/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_43 sky130_fd_sc_hd__inv_2_32/A sky130_fd_sc_hd__ha_2_11/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_43/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_146 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_146/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__fa_2_871/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_54 sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__clkinv_1_54/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_54/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_157 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_157/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__xor2_1_13/X sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_65 sky130_fd_sc_hd__nand3_1_30/C sky130_fd_sc_hd__xor2_1_3/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_65/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_168 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_168/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_168/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_76 sky130_fd_sc_hd__clkinv_1_76/Y sky130_fd_sc_hd__clkinv_1_76/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_76/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_179 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_179/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_179/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_87 sky130_fd_sc_hd__clkinv_1_88/A sky130_fd_sc_hd__ha_2_42/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_87/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_98 sky130_fd_sc_hd__inv_2_62/A sky130_fd_sc_hd__ha_2_38/A
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_901 sky130_fd_sc_hd__fa_2_900/CIN sky130_fd_sc_hd__fa_2_901/SUM
+ sky130_fd_sc_hd__fa_2_901/A sky130_fd_sc_hd__fa_2_901/B sky130_fd_sc_hd__fa_2_901/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_912 sky130_fd_sc_hd__fa_2_890/A sky130_fd_sc_hd__fa_2_891/B
+ sky130_fd_sc_hd__fa_2_912/A sky130_fd_sc_hd__fa_2_912/B sky130_fd_sc_hd__fa_2_912/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_923 sky130_fd_sc_hd__fa_2_922/CIN sky130_fd_sc_hd__fa_2_923/SUM
+ sky130_fd_sc_hd__fa_2_923/A sky130_fd_sc_hd__fa_2_923/B sky130_fd_sc_hd__fa_2_923/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_934 sky130_fd_sc_hd__fa_2_924/A sky130_fd_sc_hd__fa_2_925/B
+ sky130_fd_sc_hd__fa_2_934/A sky130_fd_sc_hd__fa_2_934/B sky130_fd_sc_hd__ha_2_122/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_945 sky130_fd_sc_hd__fa_2_944/CIN sky130_fd_sc_hd__fa_2_945/SUM
+ sky130_fd_sc_hd__fa_2_945/A sky130_fd_sc_hd__fa_2_945/B sky130_fd_sc_hd__fa_2_945/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_956 sky130_fd_sc_hd__fa_2_955/CIN sky130_fd_sc_hd__fa_2_956/SUM
+ sky130_fd_sc_hd__fa_2_956/A sky130_fd_sc_hd__fa_2_956/B sky130_fd_sc_hd__fa_2_956/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_967 sky130_fd_sc_hd__fa_2_966/CIN sky130_fd_sc_hd__fa_2_967/SUM
+ sky130_fd_sc_hd__fa_2_967/A sky130_fd_sc_hd__fa_2_967/B sky130_fd_sc_hd__fa_2_967/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_978 sky130_fd_sc_hd__fa_2_979/CIN sky130_fd_sc_hd__mux2_2_33/A1
+ sky130_fd_sc_hd__fa_2_978/A sky130_fd_sc_hd__fa_2_978/B sky130_fd_sc_hd__fa_2_978/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_989 sky130_fd_sc_hd__fa_2_990/CIN sky130_fd_sc_hd__mux2_2_9/A0
+ sky130_fd_sc_hd__fa_2_989/A sky130_fd_sc_hd__fa_2_989/B sky130_fd_sc_hd__fa_2_989/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__mux2_2_201 VSS VDD sky130_fd_sc_hd__mux2_2_201/A1 sky130_fd_sc_hd__mux2_2_201/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_201/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_212 VSS VDD sky130_fd_sc_hd__mux2_2_212/A1 sky130_fd_sc_hd__mux2_2_212/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_212/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_223 VSS VDD sky130_fd_sc_hd__mux2_2_223/A1 sky130_fd_sc_hd__mux2_2_223/A0
+ sky130_fd_sc_hd__nor2_8_2/A sky130_fd_sc_hd__mux2_2_223/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_234 VSS VDD sky130_fd_sc_hd__mux2_2_234/A1 sky130_fd_sc_hd__mux2_2_234/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_234/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_245 VSS VDD sky130_fd_sc_hd__mux2_2_245/A1 sky130_fd_sc_hd__mux2_2_245/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_245/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_256 VSS VDD sky130_fd_sc_hd__mux2_2_256/A1 sky130_fd_sc_hd__mux2_2_256/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_256/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_267 VSS VDD sky130_fd_sc_hd__mux2_2_267/A1 sky130_fd_sc_hd__mux2_2_267/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_267/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__a22o_1_1 sky130_fd_sc_hd__buf_2_279/X sky130_fd_sc_hd__nor2_1_1/Y
+ sky130_fd_sc_hd__a22o_1_1/X sky130_fd_sc_hd__a22o_1_1/B2 sky130_fd_sc_hd__nor2_1_0/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__o21ai_1_103 VSS VDD sky130_fd_sc_hd__nor2_1_84/Y sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__a21oi_1_88/Y sky130_fd_sc_hd__xor2_1_71/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_114 VSS VDD sky130_fd_sc_hd__o21a_1_8/A2 sky130_fd_sc_hd__nor2_1_64/B
+ sky130_fd_sc_hd__a22oi_1_330/Y sky130_fd_sc_hd__o21ai_1_114/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_125 VSS VDD sky130_fd_sc_hd__a21oi_1_119/Y sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__nand2_1_273/Y sky130_fd_sc_hd__xor2_1_38/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_136 VSS VDD sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_1_90/B
+ sky130_fd_sc_hd__nand2_1_278/Y sky130_fd_sc_hd__o21ai_1_136/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_147 VSS VDD sky130_fd_sc_hd__o21ai_1_147/A2 sky130_fd_sc_hd__o21ai_1_92/A1
+ sky130_fd_sc_hd__a22oi_1_338/Y sky130_fd_sc_hd__o21ai_1_147/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_158 VSS VDD sky130_fd_sc_hd__o21ai_1_171/A2 sky130_fd_sc_hd__xnor2_1_63/Y
+ sky130_fd_sc_hd__a21oi_1_135/Y sky130_fd_sc_hd__o21ai_1_158/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_169 VSS VDD sky130_fd_sc_hd__o21ai_1_171/A2 sky130_fd_sc_hd__xnor2_1_85/Y
+ sky130_fd_sc_hd__a21oi_1_146/Y sky130_fd_sc_hd__o21ai_1_169/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21bai_1_4 sky130_fd_sc_hd__buf_2_263/X sky130_fd_sc_hd__o21bai_1_4/Y
+ sky130_fd_sc_hd__buf_2_262/A sky130_fd_sc_hd__o21bai_1_4/A2 VDD VSS VDD VSS sky130_fd_sc_hd__o21bai_1
Xsky130_fd_sc_hd__maj3_1_20 sky130_fd_sc_hd__maj3_1_21/X sky130_fd_sc_hd__maj3_1_20/X
+ sky130_fd_sc_hd__maj3_1_20/B sky130_fd_sc_hd__maj3_1_20/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_31 sky130_fd_sc_hd__maj3_1_32/X sky130_fd_sc_hd__maj3_1_31/X
+ sky130_fd_sc_hd__maj3_1_31/B sky130_fd_sc_hd__maj3_1_31/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_410 sky130_fd_sc_hd__nor2_1_310/A sky130_fd_sc_hd__nor2_1_307/A
+ sky130_fd_sc_hd__o22ai_1_410/Y sky130_fd_sc_hd__a21boi_1_7/Y sky130_fd_sc_hd__nor2_1_292/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_42 sky130_fd_sc_hd__maj3_1_43/X sky130_fd_sc_hd__maj3_1_42/X
+ sky130_fd_sc_hd__maj3_1_42/B sky130_fd_sc_hd__maj3_1_42/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_421 sky130_fd_sc_hd__o22ai_1_436/A2 sky130_fd_sc_hd__o22ai_1_421/B1
+ sky130_fd_sc_hd__o22ai_1_421/Y sky130_fd_sc_hd__nor2_1_270/B sky130_fd_sc_hd__o32ai_1_11/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_53 sky130_fd_sc_hd__maj3_1_54/X sky130_fd_sc_hd__maj3_1_53/X
+ sky130_fd_sc_hd__maj3_1_53/B sky130_fd_sc_hd__maj3_1_53/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_432 sky130_fd_sc_hd__o22ai_1_432/A2 sky130_fd_sc_hd__nor2_1_280/B
+ sky130_fd_sc_hd__o22ai_1_432/Y sky130_fd_sc_hd__nor2_1_281/B sky130_fd_sc_hd__o32ai_1_11/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_64 sky130_fd_sc_hd__maj3_1_65/X sky130_fd_sc_hd__maj3_1_64/X
+ sky130_fd_sc_hd__maj3_1_64/B sky130_fd_sc_hd__maj3_1_64/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_507 sky130_fd_sc_hd__o21a_1_64/B1 sky130_fd_sc_hd__fa_2_1305/A
+ sky130_fd_sc_hd__o21a_1_64/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_75 sky130_fd_sc_hd__maj3_1_76/X sky130_fd_sc_hd__maj3_1_75/X
+ sky130_fd_sc_hd__maj3_1_75/B sky130_fd_sc_hd__maj3_1_75/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_518 sky130_fd_sc_hd__nand2_1_518/Y sky130_fd_sc_hd__inv_2_140/Y
+ sky130_fd_sc_hd__nand2_1_518/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_86 sky130_fd_sc_hd__maj3_1_87/X sky130_fd_sc_hd__maj3_1_86/X
+ sky130_fd_sc_hd__maj3_1_86/B sky130_fd_sc_hd__maj3_1_86/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_97 sky130_fd_sc_hd__maj3_1_98/X sky130_fd_sc_hd__maj3_1_97/X
+ sky130_fd_sc_hd__maj3_1_97/B sky130_fd_sc_hd__maj3_1_97/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_529 sky130_fd_sc_hd__nand2_1_529/Y sky130_fd_sc_hd__xor2_1_299/A
+ sky130_fd_sc_hd__nor2_1_309/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_9 sky130_fd_sc_hd__ha_2_21/SUM sky130_fd_sc_hd__nor2b_1_9/Y
+ sky130_fd_sc_hd__or2_0_1/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1109 sky130_fd_sc_hd__nor2_1_285/B sky130_fd_sc_hd__o21bai_1_5/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1109/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_70 sky130_fd_sc_hd__nand2_1_70/Y sky130_fd_sc_hd__nand2_1_71/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_81 sky130_fd_sc_hd__nand2_1_81/Y sky130_fd_sc_hd__nand4_1_64/Y
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_92 sky130_fd_sc_hd__nand2_1_92/Y sky130_fd_sc_hd__nand2_1_93/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_303 VDD VSS sky130_fd_sc_hd__a22o_1_46/A1 sky130_fd_sc_hd__dfxtp_1_304/CLK
+ sky130_fd_sc_hd__and2_0_95/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_314 VDD VSS sky130_fd_sc_hd__ha_2_167/B sky130_fd_sc_hd__dfxtp_1_347/CLK
+ sky130_fd_sc_hd__nor2_1_15/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_325 VDD VSS sky130_fd_sc_hd__or4_1_1/A sky130_fd_sc_hd__dfxtp_1_325/CLK
+ sky130_fd_sc_hd__and2_0_157/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_336 VDD VSS sky130_fd_sc_hd__a22o_2_11/B2 sky130_fd_sc_hd__dfxtp_1_360/CLK
+ sky130_fd_sc_hd__o21ai_1_28/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_347 VDD VSS sky130_fd_sc_hd__ha_2_154/A sky130_fd_sc_hd__dfxtp_1_347/CLK
+ sky130_fd_sc_hd__o2bb2ai_1_4/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_358 VDD VSS sky130_fd_sc_hd__a22o_2_6/B2 sky130_fd_sc_hd__dfxtp_1_360/CLK
+ sky130_fd_sc_hd__ha_2_148/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_369 VDD VSS sky130_fd_sc_hd__fa_2_1113/A sky130_fd_sc_hd__clkinv_4_32/Y
+ sky130_fd_sc_hd__and2_0_143/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_208 sky130_fd_sc_hd__fa_2_206/B sky130_fd_sc_hd__fa_2_202/B
+ sky130_fd_sc_hd__fa_2_258/A sky130_fd_sc_hd__fa_2_250/A sky130_fd_sc_hd__ha_2_102/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_219 sky130_fd_sc_hd__fa_2_221/CIN sky130_fd_sc_hd__fa_2_215/A
+ sky130_fd_sc_hd__fa_2_219/A sky130_fd_sc_hd__fa_2_219/B sky130_fd_sc_hd__fa_2_219/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_11 sky130_fd_sc_hd__fa_2_6/A sky130_fd_sc_hd__fa_2_0/B sky130_fd_sc_hd__fa_2_91/A
+ sky130_fd_sc_hd__fa_2_11/B sky130_fd_sc_hd__fa_2_99/B VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_22 sky130_fd_sc_hd__fa_2_19/CIN sky130_fd_sc_hd__fa_2_22/SUM
+ sky130_fd_sc_hd__fa_2_22/A sky130_fd_sc_hd__fa_2_22/B sky130_fd_sc_hd__fa_2_22/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_33 sky130_fd_sc_hd__maj3_1_26/B sky130_fd_sc_hd__maj3_1_27/A
+ sky130_fd_sc_hd__fa_2_67/B sky130_fd_sc_hd__fa_2_76/A sky130_fd_sc_hd__fa_2_33/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_44 sky130_fd_sc_hd__maj3_1_21/B sky130_fd_sc_hd__maj3_1_22/A
+ sky130_fd_sc_hd__fa_2_44/A sky130_fd_sc_hd__fa_2_44/B sky130_fd_sc_hd__fa_2_45/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_55 sky130_fd_sc_hd__fa_2_59/B sky130_fd_sc_hd__fa_2_55/SUM
+ sky130_fd_sc_hd__fa_2_55/A sky130_fd_sc_hd__fa_2_55/B sky130_fd_sc_hd__fa_2_55/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_66 sky130_fd_sc_hd__fa_2_64/B sky130_fd_sc_hd__fa_2_60/B sky130_fd_sc_hd__fa_2_76/B
+ sky130_fd_sc_hd__fa_2_66/B sky130_fd_sc_hd__ha_2_93/SUM VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_77 sky130_fd_sc_hd__fa_2_79/CIN sky130_fd_sc_hd__fa_2_73/A
+ sky130_fd_sc_hd__fa_2_77/A sky130_fd_sc_hd__fa_2_77/B sky130_fd_sc_hd__fa_2_77/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_88 sky130_fd_sc_hd__fa_2_90/CIN sky130_fd_sc_hd__fa_2_84/A
+ sky130_fd_sc_hd__fa_2_88/A sky130_fd_sc_hd__fa_2_88/B sky130_fd_sc_hd__fa_2_88/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_99 sky130_fd_sc_hd__fa_2_103/B sky130_fd_sc_hd__fa_2_99/SUM
+ sky130_fd_sc_hd__fa_2_99/A sky130_fd_sc_hd__fa_2_99/B sky130_fd_sc_hd__fa_2_99/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_203 VDD VSS sky130_fd_sc_hd__buf_2_203/X sky130_fd_sc_hd__buf_2_203/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_214 VDD VSS sky130_fd_sc_hd__buf_2_214/X sky130_fd_sc_hd__buf_2_214/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_225 VDD VSS sky130_fd_sc_hd__buf_2_225/X sky130_fd_sc_hd__buf_2_225/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_236 VDD VSS sky130_fd_sc_hd__buf_2_236/X sky130_fd_sc_hd__buf_2_236/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_247 VDD VSS sky130_fd_sc_hd__buf_2_247/X sky130_fd_sc_hd__buf_2_247/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_258 VDD VSS sky130_fd_sc_hd__ha_2_97/A sky130_fd_sc_hd__fa_2_247/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_269 VDD VSS sky130_fd_sc_hd__buf_2_269/X sky130_fd_sc_hd__buf_2_269/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1210 VDD VSS sky130_fd_sc_hd__fa_2_1259/A sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__mux2_2_174/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1221 VDD VSS sky130_fd_sc_hd__fa_2_1233/A sky130_fd_sc_hd__clkinv_8_78/Y
+ sky130_fd_sc_hd__mux2_2_192/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1232 VDD VSS sky130_fd_sc_hd__fa_2_1261/A sky130_fd_sc_hd__clkinv_8_63/Y
+ sky130_fd_sc_hd__mux2_2_218/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1243 VDD VSS sky130_fd_sc_hd__fa_2_1272/A sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__mux2_2_193/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1254 VDD VSS sky130_fd_sc_hd__mux2_2_210/A0 sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__a21oi_1_378/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1265 VDD VSS sky130_fd_sc_hd__mux2_2_181/A1 sky130_fd_sc_hd__clkinv_8_116/Y
+ sky130_fd_sc_hd__o22ai_1_326/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1276 VDD VSS sky130_fd_sc_hd__mux2_2_211/A0 sky130_fd_sc_hd__clkinv_8_63/Y
+ sky130_fd_sc_hd__dfxtp_1_432/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1287 VDD VSS sky130_fd_sc_hd__mux2_2_203/A0 sky130_fd_sc_hd__clkinv_8_116/Y
+ sky130_fd_sc_hd__o22ai_1_348/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1298 VDD VSS sky130_fd_sc_hd__mux2_2_176/A1 sky130_fd_sc_hd__clkinv_8_116/Y
+ sky130_fd_sc_hd__o22ai_1_337/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_870 VDD VSS sky130_fd_sc_hd__mux2_2_52/A1 sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__o21ai_1_184/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_881 VDD VSS sky130_fd_sc_hd__fa_2_861/A sky130_fd_sc_hd__dfxtp_1_902/CLK
+ sky130_fd_sc_hd__o21a_1_28/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_892 VDD VSS sky130_fd_sc_hd__fa_2_850/A sky130_fd_sc_hd__clkinv_4_22/Y
+ sky130_fd_sc_hd__o21a_1_23/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__or3_1_2 sky130_fd_sc_hd__or3_1_2/A sky130_fd_sc_hd__or3_1_2/X sky130_fd_sc_hd__or3_1_2/B
+ sky130_fd_sc_hd__or3_1_2/C VDD VSS VDD VSS sky130_fd_sc_hd__or3_1
Xsky130_fd_sc_hd__clkbuf_1_490 VSS VDD sky130_fd_sc_hd__a22oi_2_30/B2 sky130_fd_sc_hd__clkbuf_1_490/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a21oi_1_16 sky130_fd_sc_hd__inv_4_1/A sky130_fd_sc_hd__or2_0_0/B
+ sky130_fd_sc_hd__a21oi_1_16/Y sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_27 sky130_fd_sc_hd__fa_2_968/A sky130_fd_sc_hd__nor3_1_37/C
+ sky130_fd_sc_hd__a221o_1_0/B1 sky130_fd_sc_hd__nor3_1_37/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_38 sky130_fd_sc_hd__nor2_1_41/Y sky130_fd_sc_hd__o22ai_1_71/Y
+ sky130_fd_sc_hd__a21oi_1_38/Y sky130_fd_sc_hd__fa_2_1041/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__fa_2_720 sky130_fd_sc_hd__maj3_1_156/B sky130_fd_sc_hd__maj3_1_157/A
+ sky130_fd_sc_hd__fa_2_758/B sky130_fd_sc_hd__fa_2_720/B sky130_fd_sc_hd__fa_2_721/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a21oi_1_49 sky130_fd_sc_hd__nor2_2_6/Y sky130_fd_sc_hd__o22ai_1_81/Y
+ sky130_fd_sc_hd__a21oi_1_49/Y sky130_fd_sc_hd__fa_2_1037/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__fa_2_731 sky130_fd_sc_hd__fa_2_733/CIN sky130_fd_sc_hd__fa_2_729/A
+ sky130_fd_sc_hd__ha_2_138/A sky130_fd_sc_hd__ha_2_136/A sky130_fd_sc_hd__fa_2_817/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_742 sky130_fd_sc_hd__fa_2_744/B sky130_fd_sc_hd__fa_2_742/SUM
+ sky130_fd_sc_hd__fa_2_742/A sky130_fd_sc_hd__fa_2_742/B sky130_fd_sc_hd__fa_2_746/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_753 sky130_fd_sc_hd__fa_2_756/B sky130_fd_sc_hd__fa_2_753/SUM
+ sky130_fd_sc_hd__fa_2_753/A sky130_fd_sc_hd__fa_2_753/B sky130_fd_sc_hd__o22ai_1_51/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_764 sky130_fd_sc_hd__maj3_1_142/B sky130_fd_sc_hd__maj3_1_143/A
+ sky130_fd_sc_hd__fa_2_764/A sky130_fd_sc_hd__fa_2_764/B sky130_fd_sc_hd__fa_2_764/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_775 sky130_fd_sc_hd__maj3_1_139/B sky130_fd_sc_hd__maj3_1_140/A
+ sky130_fd_sc_hd__fa_2_775/A sky130_fd_sc_hd__fa_2_775/B sky130_fd_sc_hd__fa_2_776/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_786 sky130_fd_sc_hd__maj3_1_136/B sky130_fd_sc_hd__maj3_1_137/A
+ sky130_fd_sc_hd__fa_2_786/A sky130_fd_sc_hd__fa_2_786/B sky130_fd_sc_hd__fa_2_787/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_797 sky130_fd_sc_hd__fa_2_798/CIN sky130_fd_sc_hd__fa_2_791/B
+ sky130_fd_sc_hd__fa_2_834/A sky130_fd_sc_hd__fa_2_823/B sky130_fd_sc_hd__fa_2_817/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor3_1_8 sky130_fd_sc_hd__nor3_1_8/C sky130_fd_sc_hd__nor3_1_8/Y
+ sky130_fd_sc_hd__nor3_2_3/A sky130_fd_sc_hd__nor3_2_2/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__buf_6_12 VDD VSS sky130_fd_sc_hd__buf_6_12/X sky130_fd_sc_hd__buf_8_18/X
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_23 VDD VSS sky130_fd_sc_hd__buf_6_23/X sky130_fd_sc_hd__buf_8_65/X
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_34 VDD VSS sky130_fd_sc_hd__buf_6_34/X sky130_fd_sc_hd__buf_6_34/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_45 VDD VSS sky130_fd_sc_hd__buf_6_45/X sky130_fd_sc_hd__buf_6_45/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_56 VDD VSS sky130_fd_sc_hd__buf_6_56/X sky130_fd_sc_hd__buf_6_56/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_67 VDD VSS sky130_fd_sc_hd__buf_6_67/X sky130_fd_sc_hd__buf_6_67/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_78 VDD VSS sky130_fd_sc_hd__buf_6_78/X sky130_fd_sc_hd__buf_6_78/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_89 VDD VSS sky130_fd_sc_hd__buf_6_89/X sky130_fd_sc_hd__buf_6_89/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_14 sky130_fd_sc_hd__buf_2_123/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_25 sky130_fd_sc_hd__clkinv_1_76/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_36 sky130_fd_sc_hd__buf_2_108/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_47 sky130_fd_sc_hd__buf_2_79/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_58 sky130_fd_sc_hd__nand4_1_25/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_69 sky130_fd_sc_hd__clkbuf_4_88/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__o22ai_1_240 sky130_fd_sc_hd__o32ai_1_0/B2 sky130_fd_sc_hd__nor2_1_182/A
+ sky130_fd_sc_hd__o22ai_1_240/Y sky130_fd_sc_hd__o22ai_1_262/A1 sky130_fd_sc_hd__a222oi_1_5/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_304 sky130_fd_sc_hd__nand2_1_304/Y sky130_fd_sc_hd__nor2_1_102/B
+ sky130_fd_sc_hd__fa_2_1113/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_903 sky130_fd_sc_hd__o22ai_1_301/A1 sky130_fd_sc_hd__o21ai_1_352/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_903/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_251 sky130_fd_sc_hd__o32ai_1_2/A3 sky130_fd_sc_hd__nor2_1_146/B
+ sky130_fd_sc_hd__o22ai_1_251/Y sky130_fd_sc_hd__o22ai_1_251/A1 sky130_fd_sc_hd__o21a_1_29/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_315 sky130_fd_sc_hd__nand2_1_315/Y sky130_fd_sc_hd__nand2_1_339/B
+ sky130_fd_sc_hd__o21ai_1_208/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_914 sky130_fd_sc_hd__nor2_1_189/B sky130_fd_sc_hd__fa_2_1179/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_914/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_262 sky130_fd_sc_hd__nor2_1_157/B sky130_fd_sc_hd__nor2_1_182/A
+ sky130_fd_sc_hd__o22ai_1_262/Y sky130_fd_sc_hd__o22ai_1_262/A1 sky130_fd_sc_hd__a222oi_1_13/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_326 sky130_fd_sc_hd__nand2_1_326/Y sky130_fd_sc_hd__nand2_1_331/B
+ sky130_fd_sc_hd__o21ai_1_231/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_273 sky130_fd_sc_hd__nand2_1_410/Y sky130_fd_sc_hd__nand2_1_409/Y
+ sky130_fd_sc_hd__o22ai_1_273/Y sky130_fd_sc_hd__nand2_1_422/B sky130_fd_sc_hd__o21ai_1_334/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_925 sky130_fd_sc_hd__o22ai_1_316/B1 sky130_fd_sc_hd__fa_2_1208/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_925/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_337 sky130_fd_sc_hd__o21a_1_16/A2 sky130_fd_sc_hd__nor2_4_13/B
+ sky130_fd_sc_hd__nor2_4_13/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_936 sky130_fd_sc_hd__o22ai_1_321/A1 sky130_fd_sc_hd__fa_2_1199/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_936/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_284 sky130_fd_sc_hd__nand2_1_412/Y sky130_fd_sc_hd__nand2_1_411/Y
+ sky130_fd_sc_hd__o22ai_1_284/Y sky130_fd_sc_hd__nand2_1_421/B sky130_fd_sc_hd__o21ai_1_333/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_348 sky130_fd_sc_hd__nor2_1_149/A sky130_fd_sc_hd__fa_2_1124/A
+ sky130_fd_sc_hd__fa_2_1123/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_295 sky130_fd_sc_hd__nor2_1_214/A sky130_fd_sc_hd__nor2_1_225/A
+ sky130_fd_sc_hd__o22ai_1_295/Y sky130_fd_sc_hd__a21boi_1_4/Y sky130_fd_sc_hd__a222oi_1_20/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_947 sky130_fd_sc_hd__o22ai_1_375/A2 sky130_fd_sc_hd__nor2_2_17/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_947/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_359 sky130_fd_sc_hd__nand2_1_359/Y sky130_fd_sc_hd__xor2_1_185/B
+ sky130_fd_sc_hd__o31ai_1_6/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_958 sky130_fd_sc_hd__o32ai_1_7/A3 sky130_fd_sc_hd__fa_2_1243/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_958/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_969 sky130_fd_sc_hd__o22ai_1_346/A1 sky130_fd_sc_hd__nor2_1_255/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_969/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_100 VDD VSS sky130_fd_sc_hd__ha_2_4/A sky130_fd_sc_hd__dfxtp_1_99/CLK
+ sky130_fd_sc_hd__and2_0_9/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_111 VDD VSS sky130_fd_sc_hd__nor2_1_23/A sky130_fd_sc_hd__dfxtp_1_111/CLK
+ sky130_fd_sc_hd__ha_2_5/SUM VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_122 VDD VSS sky130_fd_sc_hd__ha_2_18/A sky130_fd_sc_hd__dfxtp_1_129/CLK
+ sky130_fd_sc_hd__and2_0_20/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_133 VDD VSS sky130_fd_sc_hd__ha_2_29/A sky130_fd_sc_hd__dfxtp_1_138/CLK
+ sky130_fd_sc_hd__nor2b_1_5/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_144 VDD VSS sky130_fd_sc_hd__nor3_2_3/A sky130_fd_sc_hd__clkinv_4_2/Y
+ sky130_fd_sc_hd__ha_2_29/B VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_155 VDD VSS sky130_fd_sc_hd__ha_2_32/A sky130_fd_sc_hd__dfxtp_1_155/CLK
+ sky130_fd_sc_hd__and2_0_24/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_166 VDD VSS sky130_fd_sc_hd__ha_2_43/A sky130_fd_sc_hd__dfxtp_1_166/CLK
+ sky130_fd_sc_hd__nor2b_2_1/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_177 VDD VSS sky130_fd_sc_hd__ha_2_57/A sky130_fd_sc_hd__dfxtp_1_185/CLK
+ sky130_fd_sc_hd__and2_0_50/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_188 VDD VSS sky130_fd_sc_hd__ha_2_68/A sky130_fd_sc_hd__dfxtp_1_197/CLK
+ sky130_fd_sc_hd__nor2b_1_32/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_199 VDD VSS sky130_fd_sc_hd__nor3_2_6/B sky130_fd_sc_hd__clkinv_2_17/Y
+ sky130_fd_sc_hd__nand3_4_0/B VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_1210 sky130_fd_sc_hd__fa_2_1211/CIN sky130_fd_sc_hd__mux2_2_170/A1
+ sky130_fd_sc_hd__fa_2_1210/A sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__fa_2_1210/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1221 sky130_fd_sc_hd__fa_2_1222/CIN sky130_fd_sc_hd__mux2_2_145/A1
+ sky130_fd_sc_hd__fa_2_1221/A sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__fa_2_1221/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o211ai_1_19 sky130_fd_sc_hd__nor2_1_133/Y sky130_fd_sc_hd__nor2_1_127/A
+ sky130_fd_sc_hd__xor2_1_136/A sky130_fd_sc_hd__a22oi_1_356/Y sky130_fd_sc_hd__nand2_1_328/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__fa_2_1232 sky130_fd_sc_hd__fa_2_1233/CIN sky130_fd_sc_hd__mux2_2_195/A1
+ sky130_fd_sc_hd__fa_2_1232/A sky130_fd_sc_hd__fa_2_1232/B sky130_fd_sc_hd__fa_2_1232/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1243 sky130_fd_sc_hd__fa_2_1244/CIN sky130_fd_sc_hd__and2_0_332/A
+ sky130_fd_sc_hd__fa_2_1243/A sky130_fd_sc_hd__fa_2_1243/B sky130_fd_sc_hd__fa_2_1243/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1254 sky130_fd_sc_hd__fa_2_1255/CIN sky130_fd_sc_hd__mux2_2_184/A1
+ sky130_fd_sc_hd__fa_2_1254/A sky130_fd_sc_hd__fa_2_1254/B sky130_fd_sc_hd__fa_2_1254/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1265 sky130_fd_sc_hd__fa_2_1266/CIN sky130_fd_sc_hd__mux2_2_214/A1
+ sky130_fd_sc_hd__fa_2_1265/A sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1265/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1276 sky130_fd_sc_hd__fa_2_1277/CIN sky130_fd_sc_hd__and2_0_337/A
+ sky130_fd_sc_hd__fa_2_1276/A sky130_fd_sc_hd__fa_2_1276/B sky130_fd_sc_hd__fa_2_1276/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1287 sky130_fd_sc_hd__fa_2_1288/CIN sky130_fd_sc_hd__mux2_2_233/A1
+ sky130_fd_sc_hd__fa_2_1287/A sky130_fd_sc_hd__fa_2_1287/B sky130_fd_sc_hd__fa_2_1287/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1040 VDD VSS sky130_fd_sc_hd__fa_2_906/B sky130_fd_sc_hd__dfxtp_1_1047/CLK
+ sky130_fd_sc_hd__a21oi_1_305/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_1298 sky130_fd_sc_hd__fa_2_1299/CIN sky130_fd_sc_hd__mux2_2_251/A1
+ sky130_fd_sc_hd__fa_2_1298/A sky130_fd_sc_hd__fa_2_1298/B sky130_fd_sc_hd__fa_2_1298/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1051 VDD VSS sky130_fd_sc_hd__or2_0_10/A sky130_fd_sc_hd__clkinv_8_78/Y
+ sky130_fd_sc_hd__nor2b_1_113/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_60 VSS VDD sky130_fd_sc_hd__nand2_2_3/Y sky130_fd_sc_hd__xnor2_1_40/Y
+ sky130_fd_sc_hd__a21oi_1_46/Y sky130_fd_sc_hd__o21ai_1_60/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1062 VDD VSS sky130_fd_sc_hd__fa_2_1201/A sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__mux2_2_141/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_71 VSS VDD sky130_fd_sc_hd__o21ai_1_71/A2 sky130_fd_sc_hd__o22ai_1_88/B1
+ sky130_fd_sc_hd__a21oi_1_57/Y sky130_fd_sc_hd__o21ai_1_71/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1073 VDD VSS sky130_fd_sc_hd__fa_2_1175/A sky130_fd_sc_hd__clkinv_4_23/Y
+ sky130_fd_sc_hd__mux2_2_165/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_82 VSS VDD sky130_fd_sc_hd__xnor2_1_55/A sky130_fd_sc_hd__nor2_1_61/Y
+ sky130_fd_sc_hd__o21ai_1_82/B1 sky130_fd_sc_hd__xnor2_1_57/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1084 VDD VSS sky130_fd_sc_hd__fa_2_1186/A sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__mux2_2_135/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_93 VSS VDD sky130_fd_sc_hd__a21oi_1_93/Y sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__o21ai_1_96/B1 sky130_fd_sc_hd__xor2_1_61/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1095 VDD VSS sky130_fd_sc_hd__fa_2_1214/A sky130_fd_sc_hd__clkinv_8_64/Y
+ sky130_fd_sc_hd__mux2_2_166/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o2bb2ai_1_13 sky130_fd_sc_hd__maj3_1_1/A sky130_fd_sc_hd__nand2_1_201/B
+ sky130_fd_sc_hd__nor2_1_21/Y sky130_fd_sc_hd__nor2_1_21/Y sky130_fd_sc_hd__nand2_1_201/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__o2bb2ai_1_24 sky130_fd_sc_hd__and2_0_250/A sky130_fd_sc_hd__nand2_1_213/B
+ sky130_fd_sc_hd__nor2_1_31/Y sky130_fd_sc_hd__nor2_1_31/Y sky130_fd_sc_hd__nand2_1_213/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_550 sky130_fd_sc_hd__fa_2_551/CIN sky130_fd_sc_hd__fa_2_545/B
+ sky130_fd_sc_hd__ha_2_124/A sky130_fd_sc_hd__fa_2_559/B sky130_fd_sc_hd__fa_2_537/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_561 sky130_fd_sc_hd__fa_2_460/A sky130_fd_sc_hd__fa_2_464/B
+ sky130_fd_sc_hd__fa_2_561/A sky130_fd_sc_hd__fa_2_561/B sky130_fd_sc_hd__fa_2_565/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_572 sky130_fd_sc_hd__fa_2_571/CIN sky130_fd_sc_hd__and2_0_90/A
+ sky130_fd_sc_hd__fa_2_572/A sky130_fd_sc_hd__fa_2_572/B sky130_fd_sc_hd__fa_2_572/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_583 sky130_fd_sc_hd__maj3_1_132/B sky130_fd_sc_hd__maj3_1_133/A
+ sky130_fd_sc_hd__ha_2_133/A sky130_fd_sc_hd__ha_2_131/B sky130_fd_sc_hd__fa_2_624/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_594 sky130_fd_sc_hd__fa_2_596/CIN sky130_fd_sc_hd__fa_2_592/A
+ sky130_fd_sc_hd__ha_2_135/B sky130_fd_sc_hd__ha_2_132/B sky130_fd_sc_hd__ha_2_129/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a21oi_1_107 sky130_fd_sc_hd__clkinv_1_566/Y sky130_fd_sc_hd__clkinv_1_563/Y
+ sky130_fd_sc_hd__a21oi_1_107/Y sky130_fd_sc_hd__a211o_1_8/A2 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_118 sky130_fd_sc_hd__a21o_2_3/X sky130_fd_sc_hd__o22ai_1_126/Y
+ sky130_fd_sc_hd__a21oi_1_118/Y sky130_fd_sc_hd__a211o_1_6/A1 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_129 sky130_fd_sc_hd__a21o_2_3/A2 sky130_fd_sc_hd__o21ai_1_153/Y
+ sky130_fd_sc_hd__a21oi_1_129/Y sky130_fd_sc_hd__fa_2_1004/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nor2_1_304 sky130_fd_sc_hd__nor2_1_310/A sky130_fd_sc_hd__nor2_1_304/Y
+ sky130_fd_sc_hd__nor2_1_305/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_315 sky130_fd_sc_hd__nor2_1_315/B sky130_fd_sc_hd__nor2_1_315/Y
+ sky130_fd_sc_hd__nor2_1_315/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_500 sky130_fd_sc_hd__buf_12_500/A sky130_fd_sc_hd__buf_12_500/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_511 sky130_fd_sc_hd__buf_12_511/A sky130_fd_sc_hd__buf_6_83/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_403 sky130_fd_sc_hd__nor2_1_315/Y sky130_fd_sc_hd__nor2_1_313/Y
+ sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__nand3_1_3/Y sky130_fd_sc_hd__nand3_1_51/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkbuf_8_3 sky130_fd_sc_hd__clkbuf_8_3/X sky130_fd_sc_hd__dfxtp_1_92/D
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkbuf_8
Xsky130_fd_sc_hd__nand2_1_101 sky130_fd_sc_hd__nand2_1_101/Y sky130_fd_sc_hd__nand2_1_101/B
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_700 sky130_fd_sc_hd__clkinv_1_700/Y sky130_fd_sc_hd__nor2_1_131/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_700/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_112 sky130_fd_sc_hd__nand2_1_112/Y sky130_fd_sc_hd__nand2_1_113/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_711 sky130_fd_sc_hd__clkinv_1_711/Y sky130_fd_sc_hd__nor2_1_134/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_711/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_123 sky130_fd_sc_hd__nand2_1_123/Y sky130_fd_sc_hd__nand2_1_124/Y
+ sky130_fd_sc_hd__buf_2_264/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_722 sky130_fd_sc_hd__o22ai_1_194/B1 sky130_fd_sc_hd__fa_2_1053/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_722/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_134 sky130_fd_sc_hd__nand2_1_134/Y sky130_fd_sc_hd__fa_2_710/SUM
+ sky130_fd_sc_hd__and2_0_235/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_733 sky130_fd_sc_hd__nand2_1_332/A sky130_fd_sc_hd__a211oi_1_8/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_733/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_145 sky130_fd_sc_hd__nand2_1_145/Y sky130_fd_sc_hd__nand2_1_146/Y
+ sky130_fd_sc_hd__buf_2_264/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_744 sky130_fd_sc_hd__o21ai_1_271/A2 sky130_fd_sc_hd__fa_2_1081/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_744/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_156 sky130_fd_sc_hd__fa_2_134/A sky130_fd_sc_hd__fa_2_76/A
+ sky130_fd_sc_hd__fa_2_2/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_755 sky130_fd_sc_hd__ha_2_187/B sky130_fd_sc_hd__fa_2_1120/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_755/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_167 sky130_fd_sc_hd__fa_2_316/B sky130_fd_sc_hd__fa_2_417/B
+ sky130_fd_sc_hd__ha_2_116/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_766 sky130_fd_sc_hd__ha_2_199/B sky130_fd_sc_hd__fa_2_1108/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_766/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_178 sky130_fd_sc_hd__fa_2_474/CIN sky130_fd_sc_hd__fa_2_555/A
+ sky130_fd_sc_hd__fa_2_551/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_777 sky130_fd_sc_hd__nor2_2_11/B sky130_fd_sc_hd__nor2_2_10/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_777/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_189 sky130_fd_sc_hd__fa_2_653/A sky130_fd_sc_hd__fa_2_692/A
+ sky130_fd_sc_hd__fa_2_689/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_788 sky130_fd_sc_hd__o32ai_1_0/A2 sky130_fd_sc_hd__fa_2_1122/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_788/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_799 sky130_fd_sc_hd__o22ai_1_226/A1 sky130_fd_sc_hd__a21o_2_7/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_799/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor2_1_5 sky130_fd_sc_hd__xor2_1_5/B sky130_fd_sc_hd__xor2_1_5/X
+ sky130_fd_sc_hd__xor2_1_5/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand3_2_6 sky130_fd_sc_hd__nor2_1_7/A sky130_fd_sc_hd__nand3_2_6/Y
+ sky130_fd_sc_hd__nor2_1_6/B sky130_fd_sc_hd__or2_1_2/X VSS VDD VSS VDD sky130_fd_sc_hd__nand3_2
Xsky130_fd_sc_hd__clkinv_8_3 sky130_fd_sc_hd__clkinv_8_5/A sky130_fd_sc_hd__clkinv_8_3/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_3/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__nor3_1_11 sky130_fd_sc_hd__nor2_4_6/A sky130_fd_sc_hd__nor3_1_11/Y
+ sky130_fd_sc_hd__nor3_2_4/B sky130_fd_sc_hd__nor3_2_4/C VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_22 sky130_fd_sc_hd__nor2_2_4/A sky130_fd_sc_hd__nor3_1_22/Y
+ sky130_fd_sc_hd__nor3_2_10/B sky130_fd_sc_hd__nor3_1_24/C VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_33 sky130_fd_sc_hd__or4_1_2/D sky130_fd_sc_hd__xor2_1_29/B
+ sky130_fd_sc_hd__or4_1_2/B sky130_fd_sc_hd__or4_1_2/C VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__fa_2_1040 sky130_fd_sc_hd__fa_2_1041/CIN sky130_fd_sc_hd__fa_2_1040/SUM
+ sky130_fd_sc_hd__nor2_1_60/A sky130_fd_sc_hd__fa_2_1040/B sky130_fd_sc_hd__fa_2_1040/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1051 sky130_fd_sc_hd__fa_2_1052/CIN sky130_fd_sc_hd__and2_0_314/A
+ sky130_fd_sc_hd__fa_2_1051/A sky130_fd_sc_hd__fa_2_1051/B sky130_fd_sc_hd__fa_2_1051/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1062 sky130_fd_sc_hd__fa_2_1063/CIN sky130_fd_sc_hd__mux2_2_53/A0
+ sky130_fd_sc_hd__fa_2_1062/A sky130_fd_sc_hd__xor2_1_95/X sky130_fd_sc_hd__fa_2_1062/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1073 sky130_fd_sc_hd__fa_2_1074/CIN sky130_fd_sc_hd__and2_0_312/A
+ sky130_fd_sc_hd__fa_2_1073/A sky130_fd_sc_hd__fa_2_1073/B sky130_fd_sc_hd__fa_2_1073/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1084 sky130_fd_sc_hd__fa_2_1085/CIN sky130_fd_sc_hd__mux2_2_54/A0
+ sky130_fd_sc_hd__fa_2_1084/A sky130_fd_sc_hd__fa_2_1084/B sky130_fd_sc_hd__fa_2_1084/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1095 sky130_fd_sc_hd__fa_2_1096/CIN sky130_fd_sc_hd__and2_0_297/A
+ sky130_fd_sc_hd__fa_2_1095/A sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1095/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_60 sky130_fd_sc_hd__inv_2_60/A sky130_fd_sc_hd__inv_2_60/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_71 sky130_fd_sc_hd__inv_2_71/A sky130_fd_sc_hd__inv_2_71/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_82 sky130_fd_sc_hd__inv_2_82/A sky130_fd_sc_hd__inv_2_82/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_93 sky130_fd_sc_hd__inv_2_93/A sky130_fd_sc_hd__inv_2_93/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__ha_2_14 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_14/A sky130_fd_sc_hd__ha_2_13/B
+ sky130_fd_sc_hd__and2_1_0/A sky130_fd_sc_hd__ha_2_14/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_25 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_25/A sky130_fd_sc_hd__ha_2_24/B
+ sky130_fd_sc_hd__ha_2_25/SUM sky130_fd_sc_hd__ha_2_25/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_36 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_36/A sky130_fd_sc_hd__ha_2_35/B
+ sky130_fd_sc_hd__ha_2_36/SUM sky130_fd_sc_hd__ha_2_36/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_47 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_47/A sky130_fd_sc_hd__ha_2_46/B
+ sky130_fd_sc_hd__ha_2_47/SUM sky130_fd_sc_hd__ha_2_47/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_58 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_58/A sky130_fd_sc_hd__ha_2_57/B
+ sky130_fd_sc_hd__ha_2_58/SUM sky130_fd_sc_hd__ha_2_58/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_69 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_69/A sky130_fd_sc_hd__ha_2_68/B
+ sky130_fd_sc_hd__ha_2_69/SUM sky130_fd_sc_hd__ha_2_69/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__sdlclkp_4_10 sky130_fd_sc_hd__conb_1_5/LO sky130_fd_sc_hd__clkinv_8_112/A
+ sky130_fd_sc_hd__dfxtp_1_93/CLK sky130_fd_sc_hd__nor3_1_0/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_380 sky130_fd_sc_hd__fa_2_381/B sky130_fd_sc_hd__fa_2_372/A
+ sky130_fd_sc_hd__fa_2_393/A sky130_fd_sc_hd__fa_2_425/A sky130_fd_sc_hd__fa_2_389/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_21 sky130_fd_sc_hd__conb_1_13/LO sky130_fd_sc_hd__clkinv_8_112/A
+ sky130_fd_sc_hd__dfxtp_1_195/CLK sky130_fd_sc_hd__or2_0_2/X VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_391 sky130_fd_sc_hd__maj3_1_61/B sky130_fd_sc_hd__maj3_1_62/A
+ sky130_fd_sc_hd__fa_2_391/A sky130_fd_sc_hd__fa_2_391/B sky130_fd_sc_hd__fa_2_392/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22oi_2_2 sky130_fd_sc_hd__nor3_2_0/A sky130_fd_sc_hd__buf_2_280/X
+ sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__dfxtp_1_63/D sky130_fd_sc_hd__a22oi_2_2/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__sdlclkp_4_32 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_62/Y
+ sky130_fd_sc_hd__dfxtp_1_477/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__clkbuf_16_14 sky130_fd_sc_hd__buf_12_509/A sky130_fd_sc_hd__buf_6_69/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__sdlclkp_4_43 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_68/Y
+ sky130_fd_sc_hd__dfxtp_1_419/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_54 sky130_fd_sc_hd__conb_1_20/LO sky130_fd_sc_hd__clkinv_8_62/Y
+ sky130_fd_sc_hd__dfxtp_1_544/CLK sky130_fd_sc_hd__o21ai_1_32/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__diode_2_230 adc_bypass_en VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__sdlclkp_4_65 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__clkinv_8_62/Y
+ sky130_fd_sc_hd__dfxtp_1_483/CLK sky130_fd_sc_hd__nand2b_1_5/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_76 sky130_fd_sc_hd__conb_1_24/LO sky130_fd_sc_hd__clkinv_8_58/A
+ sky130_fd_sc_hd__dfxtp_1_768/CLK sky130_fd_sc_hd__or2_0_8/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_87 sky130_fd_sc_hd__conb_1_27/LO sky130_fd_sc_hd__clkinv_8_118/Y
+ sky130_fd_sc_hd__dfxtp_1_1184/CLK sky130_fd_sc_hd__or2_0_11/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_101 sky130_fd_sc_hd__nor2_1_101/B sky130_fd_sc_hd__nor2_1_96/A
+ sky130_fd_sc_hd__fa_2_1115/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_112 sky130_fd_sc_hd__nor2_1_112/B sky130_fd_sc_hd__nor2_1_112/Y
+ sky130_fd_sc_hd__fa_2_1120/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_123 sky130_fd_sc_hd__nor2_1_123/B sky130_fd_sc_hd__nor2_1_123/Y
+ sky130_fd_sc_hd__nor2_1_126/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_10 sky130_fd_sc_hd__nor2_2_0/Y sky130_fd_sc_hd__clkinv_1_4/Y
+ sky130_fd_sc_hd__nand4_1_26/Y sky130_fd_sc_hd__nand4_1_10/Y sky130_fd_sc_hd__a22oi_1_10/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_134 sky130_fd_sc_hd__nor2_1_134/B sky130_fd_sc_hd__nor2_1_134/Y
+ sky130_fd_sc_hd__nor2_1_134/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_21 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__nor3_2_0/A
+ sky130_fd_sc_hd__nand4_1_37/Y sig_frequency[5] sky130_fd_sc_hd__a22oi_1_21/Y VDD
+ VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_145 sky130_fd_sc_hd__nor2_1_145/B sky130_fd_sc_hd__o21a_1_20/A1
+ sky130_fd_sc_hd__o21a_1_21/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_156 sky130_fd_sc_hd__nor2_1_156/B sky130_fd_sc_hd__o21a_1_28/A1
+ sky130_fd_sc_hd__nor2_1_156/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_32 sky130_fd_sc_hd__a22oi_1_81/B1 sky130_fd_sc_hd__clkbuf_1_99/X
+ sky130_fd_sc_hd__clkbuf_1_49/X sky130_fd_sc_hd__clkbuf_4_24/X sky130_fd_sc_hd__nand4_1_1/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_43 sky130_fd_sc_hd__clkbuf_4_8/X sky130_fd_sc_hd__clkbuf_4_9/X
+ sky130_fd_sc_hd__clkbuf_1_30/X sky130_fd_sc_hd__a22oi_1_43/A2 sky130_fd_sc_hd__a22oi_1_43/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_167 sky130_fd_sc_hd__a21o_2_7/A2 sky130_fd_sc_hd__a21o_2_7/B1
+ sky130_fd_sc_hd__a21o_2_7/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_54 sky130_fd_sc_hd__nor2_2_2/Y sky130_fd_sc_hd__a22oi_1_82/A1
+ sky130_fd_sc_hd__clkbuf_1_63/X sky130_fd_sc_hd__a22oi_1_54/A2 sky130_fd_sc_hd__nand4_1_7/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_178 sky130_fd_sc_hd__nor3_1_38/A sky130_fd_sc_hd__nor2_1_178/Y
+ sky130_fd_sc_hd__nor2_1_178/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_189 sky130_fd_sc_hd__nor2_1_189/B sky130_fd_sc_hd__nor2_1_189/Y
+ sky130_fd_sc_hd__o21a_1_35/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_65 sky130_fd_sc_hd__a22oi_1_81/B1 sky130_fd_sc_hd__clkbuf_1_99/X
+ sky130_fd_sc_hd__clkbuf_1_39/X sky130_fd_sc_hd__clkbuf_4_14/X sky130_fd_sc_hd__nand4_1_11/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_76 sky130_fd_sc_hd__clkbuf_4_8/X sky130_fd_sc_hd__clkbuf_4_9/X
+ sky130_fd_sc_hd__clkbuf_1_20/X sky130_fd_sc_hd__a22oi_1_76/A2 sky130_fd_sc_hd__a22oi_1_76/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_87 sky130_fd_sc_hd__clkbuf_4_72/X sky130_fd_sc_hd__clkbuf_4_73/X
+ sky130_fd_sc_hd__a22oi_1_87/B2 sky130_fd_sc_hd__buf_2_97/X sky130_fd_sc_hd__buf_2_112/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_98 sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__a22oi_2_12/A1
+ sky130_fd_sc_hd__buf_2_78/X sky130_fd_sc_hd__a22oi_1_98/A2 sky130_fd_sc_hd__a22oi_1_98/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_330 sky130_fd_sc_hd__buf_4_95/X sky130_fd_sc_hd__buf_12_330/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_341 sky130_fd_sc_hd__buf_6_38/X sky130_fd_sc_hd__buf_12_341/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_200 sky130_fd_sc_hd__clkbuf_1_351/X sky130_fd_sc_hd__clkbuf_1_353/X
+ sky130_fd_sc_hd__clkinv_2_8/Y sky130_fd_sc_hd__a22oi_1_200/A2 sky130_fd_sc_hd__nand4_1_45/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_352 sky130_fd_sc_hd__buf_6_48/X sky130_fd_sc_hd__buf_12_352/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_211 sky130_fd_sc_hd__buf_2_166/X sky130_fd_sc_hd__buf_2_167/X
+ sky130_fd_sc_hd__clkbuf_1_438/X sky130_fd_sc_hd__buf_2_183/X sky130_fd_sc_hd__nand4_1_48/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_363 sky130_fd_sc_hd__buf_12_363/A sky130_fd_sc_hd__buf_12_363/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_222 sky130_fd_sc_hd__nor2_4_7/Y sky130_fd_sc_hd__buf_2_165/X
+ sky130_fd_sc_hd__a22oi_1_222/B2 sky130_fd_sc_hd__clkbuf_1_450/X sky130_fd_sc_hd__nand4_1_52/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_374 sky130_fd_sc_hd__buf_12_374/A sky130_fd_sc_hd__buf_12_374/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_233 sky130_fd_sc_hd__buf_2_164/X sky130_fd_sc_hd__nor2_4_8/Y
+ sky130_fd_sc_hd__clkbuf_1_421/X sky130_fd_sc_hd__buf_2_230/X sky130_fd_sc_hd__nand4_1_55/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_385 sky130_fd_sc_hd__inv_2_117/Y sky130_fd_sc_hd__buf_12_427/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_244 sky130_fd_sc_hd__a22oi_2_25/B1 sky130_fd_sc_hd__a22oi_2_25/A1
+ sky130_fd_sc_hd__clkbuf_1_385/X sky130_fd_sc_hd__a22oi_1_244/A2 sky130_fd_sc_hd__a22oi_1_244/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_396 sky130_fd_sc_hd__buf_12_396/A sky130_fd_sc_hd__buf_12_396/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_255 sky130_fd_sc_hd__buf_2_166/X sky130_fd_sc_hd__buf_2_167/X
+ sky130_fd_sc_hd__clkbuf_1_489/X sky130_fd_sc_hd__buf_2_168/X sky130_fd_sc_hd__nand4_1_63/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_266 sky130_fd_sc_hd__clkbuf_1_378/X sky130_fd_sc_hd__clkbuf_1_379/X
+ sky130_fd_sc_hd__clkbuf_4_174/X sky130_fd_sc_hd__buf_2_200/X sky130_fd_sc_hd__nand4_1_66/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_277 sky130_fd_sc_hd__clkbuf_4_165/X sky130_fd_sc_hd__clkinv_2_23/Y
+ sky130_fd_sc_hd__clkbuf_1_408/X sky130_fd_sc_hd__clkbuf_1_532/X sky130_fd_sc_hd__a22oi_1_277/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_288 sky130_fd_sc_hd__clkbuf_1_376/X sky130_fd_sc_hd__nor2_2_5/Y
+ sky130_fd_sc_hd__buf_2_210/X sky130_fd_sc_hd__clkbuf_1_466/X sky130_fd_sc_hd__nand4_1_71/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_530 sky130_fd_sc_hd__a32o_1_0/A3 sky130_fd_sc_hd__nor2_1_89/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_530/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_4_106 VDD VSS sky130_fd_sc_hd__buf_8_185/A sky130_fd_sc_hd__buf_4_106/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__a22oi_1_299 sky130_fd_sc_hd__nor2_2_4/Y sky130_fd_sc_hd__clkbuf_1_377/X
+ sky130_fd_sc_hd__a22oi_1_299/B2 sky130_fd_sc_hd__clkbuf_4_182/X sky130_fd_sc_hd__nand4_1_74/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_541 sky130_fd_sc_hd__o21ai_1_109/A1 sky130_fd_sc_hd__a211o_1_6/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_541/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_4_117 VDD VSS sky130_fd_sc_hd__buf_6_80/A sky130_fd_sc_hd__buf_8_216/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__clkinv_1_552 sky130_fd_sc_hd__o22ai_1_116/A1 sky130_fd_sc_hd__fa_2_984/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_552/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_563 sky130_fd_sc_hd__clkinv_1_563/Y sky130_fd_sc_hd__nand2_1_277/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_563/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_574 sky130_fd_sc_hd__o21ai_1_143/A1 sky130_fd_sc_hd__fa_2_1014/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_574/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_585 sky130_fd_sc_hd__clkinv_1_585/Y sky130_fd_sc_hd__a21oi_1_133/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_585/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_596 sky130_fd_sc_hd__ha_2_171/B sky130_fd_sc_hd__fa_2_1044/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_596/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_4_10 sky130_fd_sc_hd__clkinv_4_10/A sky130_fd_sc_hd__clkinv_8_14/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_10/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_21 sky130_fd_sc_hd__clkinv_8_40/A sky130_fd_sc_hd__clkinv_8_44/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_21/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_32 sky130_fd_sc_hd__clkinv_4_32/A sky130_fd_sc_hd__clkinv_4_32/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_32/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_43 sky130_fd_sc_hd__clkinv_8_84/Y sky130_fd_sc_hd__clkinv_8_85/A
+ VSS VDD VDD VSS VSS sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_54 sky130_fd_sc_hd__clkinv_4_54/A sky130_fd_sc_hd__clkinv_4_54/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_54/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_65 sky130_fd_sc_hd__clkinv_4_70/A sky130_fd_sc_hd__clkinv_4_66/A
+ VSS VDD VDD VSS VSS sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_76 sky130_fd_sc_hd__clkinv_8_17/A sky130_fd_sc_hd__clkinv_4_76/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_76/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__inv_16_6 sky130_fd_sc_hd__inv_16_6/Y sky130_fd_sc_hd__inv_16_6/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__a21oi_1_460 sky130_fd_sc_hd__fa_2_1285/A sky130_fd_sc_hd__o22ai_1_423/Y
+ sky130_fd_sc_hd__a21oi_1_460/Y sky130_fd_sc_hd__nor2_2_18/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_471 sky130_fd_sc_hd__or2_0_12/B sky130_fd_sc_hd__o21ai_1_483/Y
+ sky130_fd_sc_hd__a21oi_1_471/Y sky130_fd_sc_hd__o21ai_1_484/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_482 sky130_fd_sc_hd__nor2_1_312/Y sky130_fd_sc_hd__nand3_1_51/Y
+ sky130_fd_sc_hd__a31oi_1_3/B1 sky130_fd_sc_hd__nand3_1_0/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_493 sky130_fd_sc_hd__nand2_1_569/A sky130_fd_sc_hd__or2_0_0/B
+ sky130_fd_sc_hd__nand2_1_561/A sky130_fd_sc_hd__nor2_1_320/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_8_140 sky130_fd_sc_hd__clkinv_8_140/Y sky130_fd_sc_hd__clkinv_4_77/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_140/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__xor2_1_304 sky130_fd_sc_hd__nor2_4_20/Y sky130_fd_sc_hd__fa_2_1306/B
+ sky130_fd_sc_hd__xor2_1_304/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_315 sky130_fd_sc_hd__nor2_4_20/Y sky130_fd_sc_hd__fa_2_1295/B
+ sky130_fd_sc_hd__xor2_1_315/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_308 VSS VDD sky130_fd_sc_hd__nand4_1_37/D sky130_fd_sc_hd__a22oi_1_167/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_319 VSS VDD sky130_fd_sc_hd__clkinv_1_151/A sky130_fd_sc_hd__and2_1_5/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_12 VDD VSS sky130_fd_sc_hd__dfxtp_1_12/Q sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__a22o_1_9/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_23 VDD VSS sky130_fd_sc_hd__ha_2_110/B sky130_fd_sc_hd__dfxtp_1_26/CLK
+ sky130_fd_sc_hd__buf_2_289/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_34 VDD VSS sky130_fd_sc_hd__fa_2_905/CIN sky130_fd_sc_hd__dfxtp_1_39/CLK
+ sky130_fd_sc_hd__dfxtp_1_66/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_45 VDD VSS sky130_fd_sc_hd__xnor2_1_23/B sky130_fd_sc_hd__clkinv_4_80/Y
+ sky130_fd_sc_hd__dfxtp_1_77/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_56 VDD VSS sky130_fd_sc_hd__ha_2_124/B sky130_fd_sc_hd__dfxtp_1_61/CLK
+ sky130_fd_sc_hd__buf_2_288/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_67 VDD VSS sky130_fd_sc_hd__ha_2_94/B sky130_fd_sc_hd__dfxtp_1_73/CLK
+ sky130_fd_sc_hd__nand4_1_37/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_78 VDD VSS sky130_fd_sc_hd__nor3_1_3/A sky130_fd_sc_hd__dfxtp_1_83/CLK
+ sky130_fd_sc_hd__a21oi_1_1/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_89 VDD VSS sky130_fd_sc_hd__a22o_1_5/B2 sky130_fd_sc_hd__dfxtp_1_93/CLK
+ sky130_fd_sc_hd__buf_6_53/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_4_102 sky130_fd_sc_hd__clkbuf_4_102/X sky130_fd_sc_hd__buf_4_56/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_113 sky130_fd_sc_hd__clkbuf_4_113/X sky130_fd_sc_hd__clkbuf_4_113/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_124 sky130_fd_sc_hd__clkbuf_4_124/X sky130_fd_sc_hd__clkbuf_4_124/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_135 sky130_fd_sc_hd__clkbuf_4_135/X sky130_fd_sc_hd__clkbuf_4_135/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_306 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_306/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_306/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_146 sky130_fd_sc_hd__nand4_1_39/B sky130_fd_sc_hd__a22oi_1_177/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_317 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_317/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_317/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_157 sky130_fd_sc_hd__buf_4_69/A sky130_fd_sc_hd__a22o_1_12/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_328 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_328/X sky130_fd_sc_hd__buf_2_263/X
+ sky130_fd_sc_hd__nor3_1_39/C sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_168 sky130_fd_sc_hd__clkbuf_4_168/X sky130_fd_sc_hd__clkbuf_4_168/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_339 VSS VDD VDD VSS sky130_fd_sc_hd__or2_0_13/B sky130_fd_sc_hd__nor2_1_323/B
+ sky130_fd_sc_hd__nor2_1_323/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_179 sky130_fd_sc_hd__clkbuf_4_179/X sky130_fd_sc_hd__clkbuf_4_179/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__inv_2_106 sky130_fd_sc_hd__inv_2_106/A sky130_fd_sc_hd__inv_2_106/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_117 sky130_fd_sc_hd__inv_2_117/A sky130_fd_sc_hd__inv_2_117/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__or2_0_8 sky130_fd_sc_hd__or2_0_8/A sky130_fd_sc_hd__or2_0_8/X sky130_fd_sc_hd__or2_0_8/B
+ VSS VDD VSS VDD sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__inv_2_128 sky130_fd_sc_hd__inv_2_128/A sky130_fd_sc_hd__inv_2_128/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_139 sky130_fd_sc_hd__nor2_8_1/A sky130_fd_sc_hd__inv_2_139/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_12_160 sky130_fd_sc_hd__buf_8_70/X sky130_fd_sc_hd__buf_12_212/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_171 sky130_fd_sc_hd__buf_8_96/X sky130_fd_sc_hd__buf_12_219/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_182 sky130_fd_sc_hd__buf_8_106/X sky130_fd_sc_hd__buf_12_182/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_193 sky130_fd_sc_hd__inv_16_4/Y sky130_fd_sc_hd__buf_12_193/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_360 sky130_fd_sc_hd__fa_2_829/A sky130_fd_sc_hd__ha_2_145/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_360/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_371 sky130_fd_sc_hd__fa_2_877/B sky130_fd_sc_hd__dfxtp_1_277/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_371/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_382 sky130_fd_sc_hd__fa_2_866/B sky130_fd_sc_hd__dfxtp_1_266/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_382/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_393 sky130_fd_sc_hd__fa_2_879/B sky130_fd_sc_hd__nor2_1_21/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_393/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a211o_1_7 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_77/A sky130_fd_sc_hd__a211o_1_7/A2
+ sky130_fd_sc_hd__nor2_1_76/Y sky130_fd_sc_hd__a211o_1_8/A2 sky130_fd_sc_hd__o22ai_1_95/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o21a_1_12 sky130_fd_sc_hd__o21a_1_12/X sky130_fd_sc_hd__o21a_1_12/A1
+ sky130_fd_sc_hd__o21a_1_12/B1 sky130_fd_sc_hd__fa_2_1060/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21ai_1_307 VSS VDD sky130_fd_sc_hd__o22ai_1_261/A2 sky130_fd_sc_hd__nor2_1_147/B
+ sky130_fd_sc_hd__a21oi_1_279/Y sky130_fd_sc_hd__o21ai_1_307/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_318 VSS VDD sky130_fd_sc_hd__a21oi_1_296/Y sky130_fd_sc_hd__nor2_1_182/A
+ sky130_fd_sc_hd__a21oi_1_287/Y sky130_fd_sc_hd__xor2_1_155/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_23 sky130_fd_sc_hd__o21a_1_23/X sky130_fd_sc_hd__o21a_1_23/A1
+ sky130_fd_sc_hd__xnor2_1_92/B sky130_fd_sc_hd__fa_2_1156/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_34 sky130_fd_sc_hd__o21a_1_34/X sky130_fd_sc_hd__o21a_1_34/A1
+ sky130_fd_sc_hd__o21a_1_34/B1 sky130_fd_sc_hd__fa_2_1181/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21ai_1_329 VSS VDD sky130_fd_sc_hd__o22ai_1_261/A2 sky130_fd_sc_hd__nor2_1_155/B
+ sky130_fd_sc_hd__a21oi_1_298/Y sky130_fd_sc_hd__o21ai_1_329/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_45 sky130_fd_sc_hd__o21a_1_45/X sky130_fd_sc_hd__o21a_1_45/A1
+ sky130_fd_sc_hd__o21a_1_45/B1 sky130_fd_sc_hd__fa_2_1236/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_56 sky130_fd_sc_hd__o21a_1_56/X sky130_fd_sc_hd__o21a_1_56/A1
+ sky130_fd_sc_hd__o21a_1_56/B1 sky130_fd_sc_hd__fa_2_1291/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_67 sky130_fd_sc_hd__o21a_1_67/X sky130_fd_sc_hd__o21a_1_67/A1
+ sky130_fd_sc_hd__o21a_1_67/B1 sky130_fd_sc_hd__fa_2_1298/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__a21oi_1_290 sky130_fd_sc_hd__fa_2_1157/A sky130_fd_sc_hd__nor2_1_178/Y
+ sky130_fd_sc_hd__a21oi_1_290/Y sky130_fd_sc_hd__nor3_1_38/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_220 sky130_fd_sc_hd__buf_8_220/A sky130_fd_sc_hd__buf_8_220/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xor2_1_101 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1056/B
+ sky130_fd_sc_hd__xor2_1_101/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_112 sky130_fd_sc_hd__xor2_1_112/B sky130_fd_sc_hd__xor2_1_112/X
+ sky130_fd_sc_hd__xor2_1_113/X VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_123 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1083/B
+ sky130_fd_sc_hd__xor2_1_123/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_134 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1072/B
+ sky130_fd_sc_hd__xor2_1_134/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_145 sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__fa_2_1138/B
+ sky130_fd_sc_hd__xor2_1_145/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_156 sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__fa_2_1127/B
+ sky130_fd_sc_hd__xor2_1_156/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_507 VDD VSS sky130_fd_sc_hd__nor4_1_12/D sky130_fd_sc_hd__edfxtp_1_0/CLK
+ sky130_fd_sc_hd__a22o_1_64/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_167 sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__fa_2_1155/B
+ sky130_fd_sc_hd__xor2_1_167/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_518 VDD VSS sky130_fd_sc_hd__nor4_1_10/C sky130_fd_sc_hd__dfxtp_1_520/CLK
+ sky130_fd_sc_hd__a22o_1_53/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_178 sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__fa_2_1144/B
+ sky130_fd_sc_hd__xor2_1_178/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_189 sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__fa_2_1190/B
+ sky130_fd_sc_hd__xor2_1_189/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_529 VDD VSS sky130_fd_sc_hd__fa_2_962/A sky130_fd_sc_hd__dfxtp_1_533/CLK
+ sky130_fd_sc_hd__and2_0_261/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_105 VSS VDD sky130_fd_sc_hd__clkinv_1_54/A sky130_fd_sc_hd__inv_2_29/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_116 VSS VDD sky130_fd_sc_hd__buf_6_9/A sky130_fd_sc_hd__buf_4_12/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_127 VSS VDD sky130_fd_sc_hd__clkbuf_1_127/X sky130_fd_sc_hd__clkbuf_4_4/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_138 VSS VDD sky130_fd_sc_hd__a22oi_1_96/A1 sky130_fd_sc_hd__nor3_1_9/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_149 VSS VDD sky130_fd_sc_hd__clkbuf_1_149/X sky130_fd_sc_hd__clkbuf_1_149/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_7 VDD VSS sky130_fd_sc_hd__dfxtp_1_7/Q sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__a22o_1_4/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand3_1_16 sky130_fd_sc_hd__nand3_1_16/Y sky130_fd_sc_hd__nand3_1_16/A
+ sky130_fd_sc_hd__nor3_2_1/A sky130_fd_sc_hd__buf_2_278/X VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_27 sky130_fd_sc_hd__nand3_1_27/Y sky130_fd_sc_hd__nand2_2_0/B
+ sky130_fd_sc_hd__nand3_1_31/B sky130_fd_sc_hd__xor2_1_4/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_38 sky130_fd_sc_hd__nand3_1_38/Y sky130_fd_sc_hd__or2_1_1/X
+ sky130_fd_sc_hd__a22o_1_27/X sky130_fd_sc_hd__a22o_1_28/X VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_49 sky130_fd_sc_hd__nand3_1_49/Y sky130_fd_sc_hd__nand3_1_49/A
+ sky130_fd_sc_hd__nand3_1_49/C sky130_fd_sc_hd__nand3_1_49/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__dfxtp_1_1403 VDD VSS sky130_fd_sc_hd__mux2_2_235/A0 sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__o22ai_1_386/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1414 VDD VSS sky130_fd_sc_hd__mux2_2_264/A0 sky130_fd_sc_hd__clkinv_8_102/Y
+ sky130_fd_sc_hd__dfxtp_1_429/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1425 VDD VSS sky130_fd_sc_hd__mux2_2_260/A0 sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__nor2_1_286/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1436 VDD VSS sky130_fd_sc_hd__mux2_2_230/A1 sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__o22ai_1_397/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1447 VDD VSS sky130_fd_sc_hd__nor2_1_315/A sky130_fd_sc_hd__clkinv_8_116/Y
+ sky130_fd_sc_hd__nor2b_1_135/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1458 VDD VSS sky130_fd_sc_hd__dfxtp_1_1458/Q sky130_fd_sc_hd__dfxtp_1_1458/CLK
+ sky130_fd_sc_hd__and2_0_346/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1469 VDD VSS sky130_fd_sc_hd__nor2_1_319/A sky130_fd_sc_hd__clkinv_2_41/Y
+ sky130_fd_sc_hd__nor2b_1_141/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_103 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_103/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_916/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_11 sky130_fd_sc_hd__ha_2_24/A sky130_fd_sc_hd__inv_2_8/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_11/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_114 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_114/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_837/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_22 sky130_fd_sc_hd__inv_2_11/A sky130_fd_sc_hd__inv_2_3/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_22/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_125 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_125/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_920/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_33 sky130_fd_sc_hd__inv_2_22/A sky130_fd_sc_hd__ha_2_21/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_33/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_136 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_136/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__fa_2_869/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_44 sky130_fd_sc_hd__inv_2_33/A sky130_fd_sc_hd__buf_8_9/A
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_147 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_147/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_896/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_55 sky130_fd_sc_hd__clkinv_1_55/Y sky130_fd_sc_hd__buf_8_19/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_55/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_158 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_158/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__ha_2_158/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_66 sky130_fd_sc_hd__nand3_2_2/C sky130_fd_sc_hd__ha_2_30/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_66/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_169 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_169/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__fa_2_861/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_77 sky130_fd_sc_hd__buf_8_94/A sky130_fd_sc_hd__inv_2_51/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_77/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_88 sky130_fd_sc_hd__buf_2_48/A sky130_fd_sc_hd__clkinv_1_88/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_88/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_99 sky130_fd_sc_hd__inv_2_63/A sky130_fd_sc_hd__buf_8_81/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_99/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_902 sky130_fd_sc_hd__fa_2_901/CIN sky130_fd_sc_hd__fa_2_902/SUM
+ sky130_fd_sc_hd__fa_2_902/A sky130_fd_sc_hd__fa_2_902/B sky130_fd_sc_hd__fa_2_902/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_913 sky130_fd_sc_hd__fa_2_889/A sky130_fd_sc_hd__fa_2_890/B
+ sky130_fd_sc_hd__fa_2_913/A sky130_fd_sc_hd__fa_2_913/B sky130_fd_sc_hd__fa_2_913/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_924 sky130_fd_sc_hd__fa_2_923/CIN sky130_fd_sc_hd__fa_2_924/SUM
+ sky130_fd_sc_hd__fa_2_924/A sky130_fd_sc_hd__fa_2_924/B sky130_fd_sc_hd__fa_2_924/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_935 sky130_fd_sc_hd__fa_2_923/A sky130_fd_sc_hd__fa_2_924/B
+ sky130_fd_sc_hd__fa_2_935/A sky130_fd_sc_hd__fa_2_935/B sky130_fd_sc_hd__ha_2_123/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_946 sky130_fd_sc_hd__fa_2_945/CIN sky130_fd_sc_hd__fa_2_946/SUM
+ sky130_fd_sc_hd__fa_2_946/A sky130_fd_sc_hd__fa_2_946/B sky130_fd_sc_hd__fa_2_946/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_957 sky130_fd_sc_hd__fa_2_956/CIN sky130_fd_sc_hd__fa_2_957/SUM
+ sky130_fd_sc_hd__fa_2_957/A sky130_fd_sc_hd__fa_2_957/B sky130_fd_sc_hd__fa_2_957/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_968 sky130_fd_sc_hd__fa_2_967/CIN sky130_fd_sc_hd__fa_2_968/SUM
+ sky130_fd_sc_hd__fa_2_968/A sky130_fd_sc_hd__fa_2_968/B sky130_fd_sc_hd__fa_2_968/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_979 sky130_fd_sc_hd__fa_2_980/CIN sky130_fd_sc_hd__mux2_2_31/A1
+ sky130_fd_sc_hd__fa_2_979/A sky130_fd_sc_hd__fa_2_979/B sky130_fd_sc_hd__fa_2_979/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__mux2_2_202 VSS VDD sky130_fd_sc_hd__mux2_2_202/A1 sky130_fd_sc_hd__mux2_2_202/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_202/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_213 VSS VDD sky130_fd_sc_hd__mux2_2_213/A1 sky130_fd_sc_hd__mux2_2_213/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_213/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_224 VSS VDD sky130_fd_sc_hd__mux2_2_224/A1 sky130_fd_sc_hd__mux2_2_224/A0
+ sky130_fd_sc_hd__nor2_8_2/A sky130_fd_sc_hd__mux2_2_224/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_235 VSS VDD sky130_fd_sc_hd__mux2_2_235/A1 sky130_fd_sc_hd__mux2_2_235/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_235/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_246 VSS VDD sky130_fd_sc_hd__mux2_2_246/A1 sky130_fd_sc_hd__mux2_2_246/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_246/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_257 VSS VDD sky130_fd_sc_hd__mux2_2_257/A1 sky130_fd_sc_hd__mux2_2_257/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_257/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__buf_8_0 sky130_fd_sc_hd__buf_8_0/A sky130_fd_sc_hd__buf_8_0/X VSS
+ VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__a22o_1_2 sig_frequency[3] sky130_fd_sc_hd__nor2_1_1/Y sky130_fd_sc_hd__a22o_1_2/X
+ sky130_fd_sc_hd__a22o_1_2/B2 sky130_fd_sc_hd__nor2_1_0/Y VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_190 sky130_fd_sc_hd__nor2_2_4/A sky130_fd_sc_hd__nor2_2_5/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_190/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_70 sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__fa_2_996/A
+ sky130_fd_sc_hd__a22o_1_70/X sky130_fd_sc_hd__fa_2_994/A sky130_fd_sc_hd__nor2_2_7/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__inv_12_0 sky130_fd_sc_hd__inv_2_45/Y sky130_fd_sc_hd__inv_12_0/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_12
Xsky130_fd_sc_hd__o21ai_1_104 VSS VDD sky130_fd_sc_hd__o22ai_1_99/A2 sky130_fd_sc_hd__nor2_1_77/A
+ sky130_fd_sc_hd__nand2_1_264/Y sky130_fd_sc_hd__o21ai_1_104/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_115 VSS VDD sky130_fd_sc_hd__o22ai_1_130/B1 sky130_fd_sc_hd__nand4_1_85/A
+ sky130_fd_sc_hd__a21oi_1_100/Y sky130_fd_sc_hd__o21ai_1_115/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_126 VSS VDD sky130_fd_sc_hd__nor2_1_77/A sky130_fd_sc_hd__a21oi_1_119/Y
+ sky130_fd_sc_hd__a21oi_1_107/Y sky130_fd_sc_hd__xor2_1_42/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_137 VSS VDD sky130_fd_sc_hd__nor2_1_86/A sky130_fd_sc_hd__o22ai_1_132/B1
+ sky130_fd_sc_hd__a22oi_1_334/Y sky130_fd_sc_hd__o21ai_1_137/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_148 VSS VDD sky130_fd_sc_hd__o21ai_1_153/A2 sky130_fd_sc_hd__o22ai_1_132/B1
+ sky130_fd_sc_hd__a22oi_1_339/Y sky130_fd_sc_hd__a21o_2_3/B1 VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_159 VSS VDD sky130_fd_sc_hd__o21ai_1_171/A2 sky130_fd_sc_hd__xnor2_1_65/Y
+ sky130_fd_sc_hd__a21oi_1_136/Y sky130_fd_sc_hd__o21ai_1_159/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21bai_1_5 sky130_fd_sc_hd__buf_2_263/X sky130_fd_sc_hd__o21bai_1_5/Y
+ sky130_fd_sc_hd__buf_2_262/A sky130_fd_sc_hd__o21bai_1_5/A2 VDD VSS VDD VSS sky130_fd_sc_hd__o21bai_1
Xsky130_fd_sc_hd__maj3_1_10 sky130_fd_sc_hd__maj3_1_11/X sky130_fd_sc_hd__maj3_1_9/C
+ sky130_fd_sc_hd__maj3_1_10/B sky130_fd_sc_hd__maj3_1_10/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_21 sky130_fd_sc_hd__maj3_1_22/X sky130_fd_sc_hd__maj3_1_21/X
+ sky130_fd_sc_hd__maj3_1_21/B sky130_fd_sc_hd__maj3_1_21/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_400 sky130_fd_sc_hd__nand2_1_516/Y sky130_fd_sc_hd__nand2_1_515/Y
+ sky130_fd_sc_hd__o22ai_1_400/Y sky130_fd_sc_hd__nand2_1_526/B sky130_fd_sc_hd__o21ai_1_442/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_32 sky130_fd_sc_hd__maj3_1_33/X sky130_fd_sc_hd__maj3_1_32/X
+ sky130_fd_sc_hd__maj3_1_32/B sky130_fd_sc_hd__maj3_1_32/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_411 sky130_fd_sc_hd__o32ai_1_9/B2 sky130_fd_sc_hd__nor2_1_309/A
+ sky130_fd_sc_hd__o22ai_1_411/Y sky130_fd_sc_hd__o22ai_1_433/A1 sky130_fd_sc_hd__a222oi_1_35/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_43 sky130_fd_sc_hd__maj3_1_44/X sky130_fd_sc_hd__maj3_1_43/X
+ sky130_fd_sc_hd__maj3_1_43/B sky130_fd_sc_hd__maj3_1_43/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_422 sky130_fd_sc_hd__o32ai_1_11/A3 sky130_fd_sc_hd__nor2_1_273/B
+ sky130_fd_sc_hd__o22ai_1_422/Y sky130_fd_sc_hd__o22ai_1_422/A1 sky130_fd_sc_hd__o21a_1_68/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__inv_8_0 sky130_fd_sc_hd__inv_8_0/A sky130_fd_sc_hd__inv_8_0/Y VSS
+ VDD VSS VDD sky130_fd_sc_hd__inv_8
Xsky130_fd_sc_hd__maj3_1_54 sky130_fd_sc_hd__maj3_1_55/X sky130_fd_sc_hd__maj3_1_54/X
+ sky130_fd_sc_hd__maj3_1_54/B sky130_fd_sc_hd__maj3_1_54/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_433 sky130_fd_sc_hd__nor2_1_284/B sky130_fd_sc_hd__nor2_1_309/A
+ sky130_fd_sc_hd__o22ai_1_433/Y sky130_fd_sc_hd__o22ai_1_433/A1 sky130_fd_sc_hd__a222oi_1_43/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_65 sky130_fd_sc_hd__maj3_1_66/X sky130_fd_sc_hd__maj3_1_65/X
+ sky130_fd_sc_hd__maj3_1_65/B sky130_fd_sc_hd__maj3_1_65/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_508 sky130_fd_sc_hd__o21a_1_65/B1 sky130_fd_sc_hd__fa_2_1303/A
+ sky130_fd_sc_hd__o21a_1_65/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_76 sky130_fd_sc_hd__maj3_1_77/X sky130_fd_sc_hd__maj3_1_76/X
+ sky130_fd_sc_hd__maj3_1_76/B sky130_fd_sc_hd__maj3_1_76/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_519 sky130_fd_sc_hd__nand2_1_519/Y sky130_fd_sc_hd__nand2_1_520/Y
+ sky130_fd_sc_hd__nand2_1_521/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_87 sky130_fd_sc_hd__maj3_1_88/X sky130_fd_sc_hd__maj3_1_87/X
+ sky130_fd_sc_hd__maj3_1_87/B sky130_fd_sc_hd__maj3_1_87/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_98 sky130_fd_sc_hd__maj3_1_99/X sky130_fd_sc_hd__maj3_1_98/X
+ sky130_fd_sc_hd__maj3_1_98/B sky130_fd_sc_hd__maj3_1_98/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_60 sky130_fd_sc_hd__nand2_1_60/Y sky130_fd_sc_hd__nand2_1_61/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_71 sky130_fd_sc_hd__nand2_1_71/Y sky130_fd_sc_hd__nand4_1_69/Y
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_82 sky130_fd_sc_hd__nand2_1_82/Y sky130_fd_sc_hd__nand2_1_83/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_93 sky130_fd_sc_hd__nand2_1_93/Y sky130_fd_sc_hd__nand2_1_93/B
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_304 VDD VSS sky130_fd_sc_hd__a22o_1_45/A1 sky130_fd_sc_hd__dfxtp_1_304/CLK
+ sky130_fd_sc_hd__and2_0_94/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_315 VDD VSS sky130_fd_sc_hd__xor2_1_9/B sky130_fd_sc_hd__dfxtp_1_347/CLK
+ sky130_fd_sc_hd__and2_0_205/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_326 VDD VSS sky130_fd_sc_hd__a22o_1_27/B2 sky130_fd_sc_hd__clkinv_4_27/Y
+ sky130_fd_sc_hd__o21ai_1_18/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_337 VDD VSS sky130_fd_sc_hd__a22o_1_32/B2 sky130_fd_sc_hd__clkinv_4_27/Y
+ sky130_fd_sc_hd__nor2b_1_54/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_348 VDD VSS sky130_fd_sc_hd__a22o_1_24/B2 sky130_fd_sc_hd__dfxtp_1_360/CLK
+ sky130_fd_sc_hd__ha_2_153/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_359 VDD VSS sky130_fd_sc_hd__ha_2_148/A sky130_fd_sc_hd__dfxtp_1_361/CLK
+ sky130_fd_sc_hd__o2bb2ai_1_9/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_209 sky130_fd_sc_hd__fa_2_210/B sky130_fd_sc_hd__fa_2_202/A
+ sky130_fd_sc_hd__fa_2_2/A sky130_fd_sc_hd__fa_2_209/B sky130_fd_sc_hd__fa_2_261/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_12 sky130_fd_sc_hd__fa_2_11/B sky130_fd_sc_hd__fa_2_9/CIN sky130_fd_sc_hd__ha_2_97/A
+ sky130_fd_sc_hd__ha_2_95/B sky130_fd_sc_hd__fa_2_86/A VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_23 sky130_fd_sc_hd__fa_2_20/CIN sky130_fd_sc_hd__fa_2_25/CIN
+ sky130_fd_sc_hd__fa_2_81/B sky130_fd_sc_hd__fa_2_66/B sky130_fd_sc_hd__fa_2_23/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_34 sky130_fd_sc_hd__maj3_1_25/B sky130_fd_sc_hd__maj3_1_26/A
+ sky130_fd_sc_hd__fa_2_87/A sky130_fd_sc_hd__fa_2_34/B sky130_fd_sc_hd__fa_2_35/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_45 sky130_fd_sc_hd__fa_2_47/B sky130_fd_sc_hd__fa_2_45/SUM
+ sky130_fd_sc_hd__fa_2_45/A sky130_fd_sc_hd__fa_2_45/B sky130_fd_sc_hd__fa_2_45/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_56 sky130_fd_sc_hd__fa_2_60/CIN sky130_fd_sc_hd__fa_2_54/B
+ sky130_fd_sc_hd__fa_2_56/A sky130_fd_sc_hd__fa_2_56/B sky130_fd_sc_hd__fa_2_65/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_67 sky130_fd_sc_hd__fa_2_68/B sky130_fd_sc_hd__fa_2_60/A sky130_fd_sc_hd__fa_2_2/A
+ sky130_fd_sc_hd__fa_2_67/B sky130_fd_sc_hd__fa_2_80/B VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_78 sky130_fd_sc_hd__maj3_1_13/B sky130_fd_sc_hd__maj3_1_14/A
+ sky130_fd_sc_hd__fa_2_78/A sky130_fd_sc_hd__fa_2_78/B sky130_fd_sc_hd__fa_2_79/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_89 sky130_fd_sc_hd__maj3_1_11/B sky130_fd_sc_hd__maj3_1_12/A
+ sky130_fd_sc_hd__fa_2_89/A sky130_fd_sc_hd__fa_2_89/B sky130_fd_sc_hd__fa_2_90/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_204 VDD VSS sky130_fd_sc_hd__buf_2_204/X sky130_fd_sc_hd__buf_2_204/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_215 VDD VSS sky130_fd_sc_hd__buf_2_215/X sky130_fd_sc_hd__buf_2_247/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_226 VDD VSS sky130_fd_sc_hd__buf_2_226/X sky130_fd_sc_hd__buf_2_226/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_237 VDD VSS sky130_fd_sc_hd__or2_1_2/A sky130_fd_sc_hd__nor2_4_4/Y
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_248 VDD VSS sky130_fd_sc_hd__buf_2_248/X sky130_fd_sc_hd__buf_2_248/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_259 VDD VSS sky130_fd_sc_hd__fa_2_2/A sky130_fd_sc_hd__buf_2_259/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1200 VDD VSS sky130_fd_sc_hd__fa_2_1249/A sky130_fd_sc_hd__clkinv_8_75/Y
+ sky130_fd_sc_hd__mux2_2_197/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1211 VDD VSS sky130_fd_sc_hd__xor2_1_253/A sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__mux2_2_172/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1222 VDD VSS sky130_fd_sc_hd__fa_2_1234/A sky130_fd_sc_hd__clkinv_8_78/Y
+ sky130_fd_sc_hd__mux2_2_190/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1233 VDD VSS sky130_fd_sc_hd__fa_2_1262/A sky130_fd_sc_hd__clkinv_8_63/Y
+ sky130_fd_sc_hd__mux2_2_217/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1244 VDD VSS sky130_fd_sc_hd__fa_2_1273/A sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__nand2_1_465/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1255 VDD VSS sky130_fd_sc_hd__mux2_2_207/A0 sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__o22ai_1_336/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1266 VDD VSS sky130_fd_sc_hd__mux2_2_179/A1 sky130_fd_sc_hd__clkinv_8_116/Y
+ sky130_fd_sc_hd__o22ai_1_325/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1277 VDD VSS sky130_fd_sc_hd__mux2_2_208/A0 sky130_fd_sc_hd__clkinv_8_65/Y
+ sky130_fd_sc_hd__dfxtp_1_433/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1288 VDD VSS sky130_fd_sc_hd__mux2_2_200/A0 sky130_fd_sc_hd__clkinv_8_75/Y
+ sky130_fd_sc_hd__o22ai_1_347/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_860 VDD VSS sky130_fd_sc_hd__mux2_2_74/A0 sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__a22o_1_73/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1299 VDD VSS sky130_fd_sc_hd__mux2_2_174/A1 sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__o31ai_1_9/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_871 VDD VSS sky130_fd_sc_hd__mux2_2_50/A1 sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__o21ai_1_185/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_882 VDD VSS sky130_fd_sc_hd__fa_2_860/A sky130_fd_sc_hd__dfxtp_1_902/CLK
+ sky130_fd_sc_hd__dfxtp_1_882/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_893 VDD VSS sky130_fd_sc_hd__xnor2_1_8/B sky130_fd_sc_hd__clkinv_4_22/Y
+ sky130_fd_sc_hd__xnor2_1_92/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__or3_1_3 sky130_fd_sc_hd__or3_1_3/A sky130_fd_sc_hd__or3_1_3/X sky130_fd_sc_hd__or3_1_3/B
+ sky130_fd_sc_hd__or3_1_3/C VDD VSS VDD VSS sky130_fd_sc_hd__or3_1
Xsky130_fd_sc_hd__clkbuf_1_480 VSS VDD sky130_fd_sc_hd__nand4_1_49/B sky130_fd_sc_hd__a22oi_1_215/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a21oi_1_17 sky130_fd_sc_hd__nor3_1_30/Y sky130_fd_sc_hd__dfxtp_1_568/Q
+ sky130_fd_sc_hd__nor2_1_24/B sky130_fd_sc_hd__or4_1_2/C VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkbuf_1_491 VSS VDD sky130_fd_sc_hd__nand4_1_52/D sky130_fd_sc_hd__a22oi_2_19/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a21oi_1_28 sky130_fd_sc_hd__nor2_1_41/Y sky130_fd_sc_hd__o22ai_1_61/Y
+ sky130_fd_sc_hd__a21oi_1_28/Y sky130_fd_sc_hd__fa_2_1031/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__fa_2_710 sky130_fd_sc_hd__fa_2_709/CIN sky130_fd_sc_hd__fa_2_710/SUM
+ sky130_fd_sc_hd__fa_2_710/A sky130_fd_sc_hd__fa_2_710/B sky130_fd_sc_hd__fa_2_710/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a21oi_1_39 sky130_fd_sc_hd__nor2_1_41/Y sky130_fd_sc_hd__o22ai_1_72/Y
+ sky130_fd_sc_hd__a21oi_1_39/Y sky130_fd_sc_hd__fa_2_1042/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__fa_2_721 sky130_fd_sc_hd__fa_2_722/B sky130_fd_sc_hd__fa_2_721/SUM
+ sky130_fd_sc_hd__ha_2_144/A sky130_fd_sc_hd__ha_2_141/A sky130_fd_sc_hd__ha_2_142/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_732 sky130_fd_sc_hd__maj3_1_151/B sky130_fd_sc_hd__maj3_1_152/A
+ sky130_fd_sc_hd__fa_2_732/A sky130_fd_sc_hd__fa_2_732/B sky130_fd_sc_hd__fa_2_733/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_743 sky130_fd_sc_hd__fa_2_742/A sky130_fd_sc_hd__fa_2_743/SUM
+ sky130_fd_sc_hd__fa_2_801/B sky130_fd_sc_hd__ha_2_138/A sky130_fd_sc_hd__ha_2_136/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_754 sky130_fd_sc_hd__fa_2_755/CIN sky130_fd_sc_hd__fa_2_749/B
+ sky130_fd_sc_hd__fa_2_832/A sky130_fd_sc_hd__fa_2_834/B sky130_fd_sc_hd__ha_2_138/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_765 sky130_fd_sc_hd__fa_2_766/A sky130_fd_sc_hd__fa_2_761/B
+ sky130_fd_sc_hd__fa_2_820/B sky130_fd_sc_hd__fa_2_811/A sky130_fd_sc_hd__ha_2_141/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_776 sky130_fd_sc_hd__fa_2_779/B sky130_fd_sc_hd__fa_2_776/SUM
+ sky130_fd_sc_hd__fa_2_776/A sky130_fd_sc_hd__fa_2_776/B sky130_fd_sc_hd__fa_2_781/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_787 sky130_fd_sc_hd__fa_2_790/A sky130_fd_sc_hd__fa_2_787/SUM
+ sky130_fd_sc_hd__fa_2_787/A sky130_fd_sc_hd__fa_2_787/B sky130_fd_sc_hd__fa_2_793/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_798 sky130_fd_sc_hd__fa_2_800/CIN sky130_fd_sc_hd__fa_2_794/A
+ sky130_fd_sc_hd__ha_2_139/B sky130_fd_sc_hd__fa_2_798/B sky130_fd_sc_hd__fa_2_798/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor3_1_9 sky130_fd_sc_hd__nor3_2_4/B sky130_fd_sc_hd__nor3_1_9/Y
+ sky130_fd_sc_hd__nor3_2_4/A sky130_fd_sc_hd__nor3_1_9/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor2b_1_140 sky130_fd_sc_hd__a21oi_1_501/Y sky130_fd_sc_hd__nor2b_1_140/Y
+ sky130_fd_sc_hd__nor2b_1_142/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__bufbuf_8_0 sky130_fd_sc_hd__inv_2_79/A sky130_fd_sc_hd__bufbuf_8_0/X
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufbuf_8
Xsky130_fd_sc_hd__buf_6_13 VDD VSS sky130_fd_sc_hd__buf_6_16/A sky130_fd_sc_hd__buf_6_13/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_24 VDD VSS sky130_fd_sc_hd__buf_6_24/X sky130_fd_sc_hd__buf_6_24/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_35 VDD VSS sky130_fd_sc_hd__buf_6_35/X sky130_fd_sc_hd__buf_6_35/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_46 VDD VSS sky130_fd_sc_hd__buf_6_46/X sky130_fd_sc_hd__buf_6_46/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_57 VDD VSS sky130_fd_sc_hd__buf_6_57/X sky130_fd_sc_hd__buf_6_57/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_68 VDD VSS sky130_fd_sc_hd__buf_6_68/X sky130_fd_sc_hd__buf_6_68/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_79 VDD VSS sky130_fd_sc_hd__buf_6_79/X sky130_fd_sc_hd__buf_6_79/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_15 sky130_fd_sc_hd__buf_2_123/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_26 sky130_fd_sc_hd__dfxtp_1_253/Q VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_37 sky130_fd_sc_hd__buf_2_76/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_48 sky130_fd_sc_hd__buf_2_78/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_59 sky130_fd_sc_hd__nand4_1_25/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__o22ai_1_230 sky130_fd_sc_hd__nand2_1_360/Y sky130_fd_sc_hd__nand2_1_359/Y
+ sky130_fd_sc_hd__o22ai_1_230/Y sky130_fd_sc_hd__o22ai_1_230/A1 sky130_fd_sc_hd__a21o_2_9/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_241 sky130_fd_sc_hd__nor2_1_172/A sky130_fd_sc_hd__nor2_1_183/A
+ sky130_fd_sc_hd__o22ai_1_241/Y sky130_fd_sc_hd__a21boi_1_1/Y sky130_fd_sc_hd__a222oi_1_6/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_305 sky130_fd_sc_hd__nand2_1_305/Y sky130_fd_sc_hd__nor2_1_101/B
+ sky130_fd_sc_hd__fa_2_1115/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_904 sky130_fd_sc_hd__nor2_1_215/A sky130_fd_sc_hd__xor2_1_209/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_904/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_252 sky130_fd_sc_hd__o22ai_1_265/A2 sky130_fd_sc_hd__o22ai_1_252/B1
+ sky130_fd_sc_hd__o22ai_1_252/Y sky130_fd_sc_hd__nor2_1_145/B sky130_fd_sc_hd__o32ai_1_2/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_316 sky130_fd_sc_hd__nand2_1_316/Y sky130_fd_sc_hd__nor2_2_12/Y
+ sky130_fd_sc_hd__nor2_1_139/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_915 sky130_fd_sc_hd__o21ai_1_360/A1 sky130_fd_sc_hd__o21ai_1_362/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_915/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_263 sky130_fd_sc_hd__o22ai_1_265/A2 sky130_fd_sc_hd__nor2_1_181/A
+ sky130_fd_sc_hd__o22ai_1_263/Y sky130_fd_sc_hd__nor2_1_151/B sky130_fd_sc_hd__o32ai_1_2/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_327 sky130_fd_sc_hd__nand2_1_327/Y sky130_fd_sc_hd__nand2_1_333/B
+ sky130_fd_sc_hd__o21ai_1_235/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_274 sky130_fd_sc_hd__nand2_1_410/Y sky130_fd_sc_hd__nand2_1_409/Y
+ sky130_fd_sc_hd__o22ai_1_274/Y sky130_fd_sc_hd__o22ai_1_287/A1 sky130_fd_sc_hd__a21o_2_15/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_926 sky130_fd_sc_hd__nor2_1_192/B sky130_fd_sc_hd__fa_2_1206/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_926/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__bufinv_8_0 sky130_fd_sc_hd__bufinv_8_0/A sky130_fd_sc_hd__buf_12_61/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufinv_8
Xsky130_fd_sc_hd__nand2_1_338 sky130_fd_sc_hd__a22o_1_73/B1 sky130_fd_sc_hd__nand2_2_5/Y
+ sky130_fd_sc_hd__nand2_1_338/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_937 sky130_fd_sc_hd__nor2_1_197/B sky130_fd_sc_hd__fa_2_1197/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_937/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_285 sky130_fd_sc_hd__nand2_1_412/Y sky130_fd_sc_hd__nand2_1_411/Y
+ sky130_fd_sc_hd__o22ai_1_285/Y sky130_fd_sc_hd__o22ai_1_285/A1 sky130_fd_sc_hd__a21o_2_14/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_349 sky130_fd_sc_hd__xnor2_1_92/B sky130_fd_sc_hd__fa_2_1156/A
+ sky130_fd_sc_hd__o21a_1_23/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_296 sky130_fd_sc_hd__nor2_1_225/A sky130_fd_sc_hd__nor2_1_222/A
+ sky130_fd_sc_hd__o22ai_1_296/Y sky130_fd_sc_hd__a21boi_1_3/Y sky130_fd_sc_hd__nor2_1_207/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_948 sky130_fd_sc_hd__nand2_1_491/B sky130_fd_sc_hd__nor2_1_267/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_948/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_959 sky130_fd_sc_hd__o32ai_1_7/A2 sky130_fd_sc_hd__fa_2_1242/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_959/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_101 VDD VSS sky130_fd_sc_hd__ha_2_3/A sky130_fd_sc_hd__dfxtp_1_95/CLK
+ sky130_fd_sc_hd__and2_0_8/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_112 VDD VSS sky130_fd_sc_hd__nand2_1_35/A sky130_fd_sc_hd__dfxtp_1_117/CLK
+ sky130_fd_sc_hd__ha_2_4/SUM VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_123 VDD VSS sky130_fd_sc_hd__ha_2_17/A sky130_fd_sc_hd__dfxtp_1_129/CLK
+ sky130_fd_sc_hd__and2_0_22/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_134 VDD VSS sky130_fd_sc_hd__ha_2_28/A sky130_fd_sc_hd__dfxtp_1_138/CLK
+ sky130_fd_sc_hd__nor2b_1_12/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_145 VDD VSS sky130_fd_sc_hd__nor3_2_2/B sky130_fd_sc_hd__clkinv_4_2/Y
+ sky130_fd_sc_hd__ha_2_20/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_156 VDD VSS sky130_fd_sc_hd__ha_2_31/A sky130_fd_sc_hd__dfxtp_1_158/CLK
+ sky130_fd_sc_hd__and2_0_30/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_167 VDD VSS sky130_fd_sc_hd__ha_2_42/A sky130_fd_sc_hd__clkinv_8_14/Y
+ sky130_fd_sc_hd__nor2b_1_20/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_178 VDD VSS sky130_fd_sc_hd__ha_2_56/A sky130_fd_sc_hd__dfxtp_1_182/CLK
+ sky130_fd_sc_hd__and2_0_58/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_189 VDD VSS sky130_fd_sc_hd__ha_2_67/A sky130_fd_sc_hd__dfxtp_1_197/CLK
+ sky130_fd_sc_hd__nor2b_1_36/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_490 VSS VDD sky130_fd_sc_hd__o22ai_1_432/A2 sky130_fd_sc_hd__o21ai_1_490/A1
+ sky130_fd_sc_hd__a21oi_1_477/Y sky130_fd_sc_hd__o21ai_1_490/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_1200 sky130_fd_sc_hd__fa_2_1201/CIN sky130_fd_sc_hd__mux2_2_143/A1
+ sky130_fd_sc_hd__fa_2_1200/A sky130_fd_sc_hd__fa_2_1200/B sky130_fd_sc_hd__fa_2_1200/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1211 sky130_fd_sc_hd__fa_2_1212/CIN sky130_fd_sc_hd__mux2_2_169/A1
+ sky130_fd_sc_hd__fa_2_1211/A sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__fa_2_1211/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1222 sky130_fd_sc_hd__fa_2_1223/CIN sky130_fd_sc_hd__nand2_1_414/A
+ sky130_fd_sc_hd__fa_2_1222/A sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__fa_2_1222/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1233 sky130_fd_sc_hd__fa_2_1234/CIN sky130_fd_sc_hd__mux2_2_192/A1
+ sky130_fd_sc_hd__fa_2_1233/A sky130_fd_sc_hd__fa_2_1233/B sky130_fd_sc_hd__fa_2_1233/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1244 sky130_fd_sc_hd__fa_2_1245/CIN sky130_fd_sc_hd__mux2_2_212/A1
+ sky130_fd_sc_hd__fa_2_1244/A sky130_fd_sc_hd__fa_2_1244/B sky130_fd_sc_hd__fa_2_1244/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1255 sky130_fd_sc_hd__fa_2_1256/CIN sky130_fd_sc_hd__mux2_2_182/A0
+ sky130_fd_sc_hd__fa_2_1255/A sky130_fd_sc_hd__fa_2_1255/B sky130_fd_sc_hd__fa_2_1255/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1266 sky130_fd_sc_hd__fa_2_1267/CIN sky130_fd_sc_hd__mux2_2_211/A1
+ sky130_fd_sc_hd__fa_2_1266/A sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1266/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1277 sky130_fd_sc_hd__fa_2_1278/CIN sky130_fd_sc_hd__mux2_2_261/A1
+ sky130_fd_sc_hd__fa_2_1277/A sky130_fd_sc_hd__fa_2_1277/B sky130_fd_sc_hd__fa_2_1277/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1030 VDD VSS sky130_fd_sc_hd__fa_2_839/A sky130_fd_sc_hd__dfxtp_1_1038/CLK
+ sky130_fd_sc_hd__a21oi_1_310/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_1288 sky130_fd_sc_hd__fa_2_1289/CIN sky130_fd_sc_hd__mux2_2_231/A0
+ sky130_fd_sc_hd__fa_2_1288/A sky130_fd_sc_hd__fa_2_1288/B sky130_fd_sc_hd__fa_2_1288/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1041 VDD VSS sky130_fd_sc_hd__fa_2_907/B sky130_fd_sc_hd__dfxtp_1_1047/CLK
+ sky130_fd_sc_hd__o21a_1_34/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_1299 sky130_fd_sc_hd__fa_2_1300/CIN sky130_fd_sc_hd__mux2_2_248/A1
+ sky130_fd_sc_hd__fa_2_1299/A sky130_fd_sc_hd__fa_2_1299/B sky130_fd_sc_hd__fa_2_1299/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o21ai_1_50 VSS VDD sky130_fd_sc_hd__o21ai_1_53/A2 sky130_fd_sc_hd__xnor2_1_54/Y
+ sky130_fd_sc_hd__a21oi_1_38/Y sky130_fd_sc_hd__o21ai_1_50/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1052 VDD VSS sky130_fd_sc_hd__fa_2_1191/B sky130_fd_sc_hd__clkinv_4_23/Y
+ sky130_fd_sc_hd__and2_0_325/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_61 VSS VDD sky130_fd_sc_hd__nand2_2_3/Y sky130_fd_sc_hd__xnor2_1_42/Y
+ sky130_fd_sc_hd__a21oi_1_47/Y sky130_fd_sc_hd__o21ai_1_61/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1063 VDD VSS sky130_fd_sc_hd__fa_2_1202/A sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__mux2_2_138/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_72 VSS VDD sky130_fd_sc_hd__o21ai_1_72/A2 sky130_fd_sc_hd__o22ai_1_88/B1
+ sky130_fd_sc_hd__a21oi_1_58/Y sky130_fd_sc_hd__o21ai_1_72/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1074 VDD VSS sky130_fd_sc_hd__fa_2_1176/A sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__mux2_2_162/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_83 VSS VDD sky130_fd_sc_hd__xnor2_1_51/A sky130_fd_sc_hd__nor2_1_60/Y
+ sky130_fd_sc_hd__o21ai_1_83/B1 sky130_fd_sc_hd__xnor2_1_53/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1085 VDD VSS sky130_fd_sc_hd__fa_2_1187/A sky130_fd_sc_hd__clkinv_8_70/Y
+ sky130_fd_sc_hd__mux2_2_133/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_94 VSS VDD sky130_fd_sc_hd__a222oi_1_0/Y sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__o21ai_1_96/B1 sky130_fd_sc_hd__xor2_1_62/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1096 VDD VSS sky130_fd_sc_hd__fa_2_1215/A sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__mux2_2_163/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_690 VDD VSS sky130_fd_sc_hd__fa_2_1029/A sky130_fd_sc_hd__clkinv_4_26/Y
+ sky130_fd_sc_hd__or2_0_5/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o2bb2ai_1_14 sky130_fd_sc_hd__maj3_1_2/A sky130_fd_sc_hd__nand2_1_204/B
+ sky130_fd_sc_hd__nor4_1_4/Y sky130_fd_sc_hd__nor4_1_4/Y sky130_fd_sc_hd__nand2_1_204/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__o2bb2ai_1_25 sky130_fd_sc_hd__and2_0_245/A sky130_fd_sc_hd__nand2_1_212/B
+ sky130_fd_sc_hd__nor2_1_30/Y sky130_fd_sc_hd__nor2_1_30/Y sky130_fd_sc_hd__nand2_1_212/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_540 sky130_fd_sc_hd__fa_2_537/B sky130_fd_sc_hd__fa_2_540/SUM
+ sky130_fd_sc_hd__ha_2_125/A sky130_fd_sc_hd__ha_2_125/B sky130_fd_sc_hd__ha_2_124/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_551 sky130_fd_sc_hd__fa_2_553/CIN sky130_fd_sc_hd__fa_2_548/A
+ sky130_fd_sc_hd__fa_2_551/A sky130_fd_sc_hd__fa_2_551/B sky130_fd_sc_hd__fa_2_551/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_562 sky130_fd_sc_hd__fa_2_561/B sky130_fd_sc_hd__fa_2_562/SUM
+ sky130_fd_sc_hd__fa_2_562/A sky130_fd_sc_hd__fa_2_562/B sky130_fd_sc_hd__fa_2_567/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_573 sky130_fd_sc_hd__fa_2_572/CIN sky130_fd_sc_hd__and2_0_91/A
+ sky130_fd_sc_hd__fa_2_573/A sky130_fd_sc_hd__fa_2_573/B sky130_fd_sc_hd__fa_2_573/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_584 sky130_fd_sc_hd__maj3_1_131/B sky130_fd_sc_hd__maj3_1_132/A
+ sky130_fd_sc_hd__ha_2_132/A sky130_fd_sc_hd__ha_2_132/B sky130_fd_sc_hd__ha_2_127/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_595 sky130_fd_sc_hd__maj3_1_125/B sky130_fd_sc_hd__maj3_1_126/A
+ sky130_fd_sc_hd__fa_2_595/A sky130_fd_sc_hd__fa_2_595/B sky130_fd_sc_hd__fa_2_596/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a21oi_1_108 sky130_fd_sc_hd__a211o_1_3/A1 sky130_fd_sc_hd__o21ai_1_128/Y
+ sky130_fd_sc_hd__a21oi_1_108/Y sky130_fd_sc_hd__o21ai_1_136/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_119 sky130_fd_sc_hd__fa_2_1012/A sky130_fd_sc_hd__o21ai_1_143/Y
+ sky130_fd_sc_hd__a21oi_1_119/Y sky130_fd_sc_hd__nor2_4_10/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nor2_1_305 sky130_fd_sc_hd__nor3_1_41/A sky130_fd_sc_hd__nor2_1_305/Y
+ sky130_fd_sc_hd__nor2_1_305/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_316 sky130_fd_sc_hd__or2_0_0/B sky130_fd_sc_hd__nor2_1_316/Y
+ sky130_fd_sc_hd__nor2_1_316/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_501 sky130_fd_sc_hd__buf_12_501/A sky130_fd_sc_hd__buf_12_501/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_512 sky130_fd_sc_hd__buf_12_512/A sky130_fd_sc_hd__buf_12_513/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_404 sky130_fd_sc_hd__nor2_1_315/Y sky130_fd_sc_hd__nor2_1_313/Y
+ sky130_fd_sc_hd__nand3_1_6/Y sky130_fd_sc_hd__nand3_1_7/Y sky130_fd_sc_hd__a31oi_1_3/A2
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkbuf_8_4 sky130_fd_sc_hd__buf_2_149/A sky130_fd_sc_hd__dfxtp_1_91/D
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkbuf_8
Xsky130_fd_sc_hd__nand2_1_102 sky130_fd_sc_hd__nand2_1_102/Y sky130_fd_sc_hd__nand2_1_103/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_701 sky130_fd_sc_hd__nor2_1_113/B sky130_fd_sc_hd__fa_2_1065/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_701/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_113 sky130_fd_sc_hd__nand2_1_113/Y sky130_fd_sc_hd__nand2_1_113/B
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_712 sky130_fd_sc_hd__nor2_1_115/B sky130_fd_sc_hd__fa_2_1061/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_712/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_124 sky130_fd_sc_hd__nand2_1_124/Y sky130_fd_sc_hd__fa_2_705/SUM
+ sky130_fd_sc_hd__and2_0_235/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_723 sky130_fd_sc_hd__nor2_1_120/B sky130_fd_sc_hd__fa_2_1052/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_723/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_135 sky130_fd_sc_hd__nand2_1_135/Y sky130_fd_sc_hd__nand2_1_136/Y
+ sky130_fd_sc_hd__buf_2_264/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_734 sky130_fd_sc_hd__o21a_1_16/A1 sky130_fd_sc_hd__fa_2_1091/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_734/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_146 sky130_fd_sc_hd__nand2_1_146/Y sky130_fd_sc_hd__fa_2_716/SUM
+ sky130_fd_sc_hd__buf_2_257/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_745 sky130_fd_sc_hd__o21ai_1_273/A1 sky130_fd_sc_hd__fa_2_1083/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_745/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_157 sky130_fd_sc_hd__fa_2_137/B sky130_fd_sc_hd__fa_2_91/B
+ sky130_fd_sc_hd__ha_2_97/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_756 sky130_fd_sc_hd__ha_2_188/B sky130_fd_sc_hd__fa_2_1119/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_756/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_168 sky130_fd_sc_hd__fa_2_327/B sky130_fd_sc_hd__fa_2_401/A
+ sky130_fd_sc_hd__fa_2_395/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_767 sky130_fd_sc_hd__ha_2_200/B sky130_fd_sc_hd__fa_2_1107/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_767/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_179 sky130_fd_sc_hd__fa_2_497/A sky130_fd_sc_hd__fa_2_564/B
+ sky130_fd_sc_hd__fa_2_567/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_778 sky130_fd_sc_hd__nand2_1_367/B sky130_fd_sc_hd__fa_2_427/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_778/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_789 sky130_fd_sc_hd__nor2_1_146/A sky130_fd_sc_hd__nor2_1_147/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_789/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor2_1_6 sky130_fd_sc_hd__xor2_1_6/B sky130_fd_sc_hd__xor2_1_6/X
+ sky130_fd_sc_hd__xor2_1_6/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand3_2_7 sky130_fd_sc_hd__nor2_1_7/A sky130_fd_sc_hd__nand3_2_7/Y
+ sky130_fd_sc_hd__or2_1_2/A sky130_fd_sc_hd__nor2_1_6/B VSS VDD VSS VDD sky130_fd_sc_hd__nand3_2
Xsky130_fd_sc_hd__clkinv_8_4 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__clkinv_8_5/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_4/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__nor3_1_12 sky130_fd_sc_hd__nor3_1_13/C sky130_fd_sc_hd__nor3_1_12/Y
+ sky130_fd_sc_hd__nor3_1_9/B sky130_fd_sc_hd__nor2_4_6/A VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_23 sky130_fd_sc_hd__nor3_1_25/C sky130_fd_sc_hd__nor3_1_23/Y
+ sky130_fd_sc_hd__nor3_2_10/A sky130_fd_sc_hd__nor2_2_4/A VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_34 sky130_fd_sc_hd__nor3_1_34/C sky130_fd_sc_hd__nor3_1_34/Y
+ sky130_fd_sc_hd__nor3_1_34/A sky130_fd_sc_hd__fa_2_946/A VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__fa_2_1030 sky130_fd_sc_hd__xor2_1_84/B sky130_fd_sc_hd__mux2_2_30/A0
+ sky130_fd_sc_hd__fa_2_1030/A sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_1030/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1041 sky130_fd_sc_hd__fa_2_1042/CIN sky130_fd_sc_hd__fa_2_1041/SUM
+ sky130_fd_sc_hd__fa_2_1041/A sky130_fd_sc_hd__nor2_1_50/A sky130_fd_sc_hd__fa_2_1041/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1052 sky130_fd_sc_hd__fa_2_1053/CIN sky130_fd_sc_hd__mux2_2_75/A1
+ sky130_fd_sc_hd__fa_2_1052/A sky130_fd_sc_hd__fa_2_1052/B sky130_fd_sc_hd__fa_2_1052/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1063 sky130_fd_sc_hd__fa_2_1064/CIN sky130_fd_sc_hd__mux2_2_51/A0
+ sky130_fd_sc_hd__fa_2_1063/A sky130_fd_sc_hd__xor2_1_94/X sky130_fd_sc_hd__fa_2_1063/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1074 sky130_fd_sc_hd__fa_2_1075/CIN sky130_fd_sc_hd__and2_0_318/A
+ sky130_fd_sc_hd__fa_2_1074/A sky130_fd_sc_hd__fa_2_1074/B sky130_fd_sc_hd__fa_2_1074/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1085 sky130_fd_sc_hd__fa_2_1086/CIN sky130_fd_sc_hd__mux2_2_52/A0
+ sky130_fd_sc_hd__fa_2_1085/A sky130_fd_sc_hd__fa_2_1085/B sky130_fd_sc_hd__fa_2_1085/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1096 sky130_fd_sc_hd__fa_2_1097/CIN sky130_fd_sc_hd__and2_0_298/A
+ sky130_fd_sc_hd__fa_2_1096/A sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1096/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_50 sky130_fd_sc_hd__inv_2_50/A sky130_fd_sc_hd__inv_2_50/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_61 sky130_fd_sc_hd__inv_2_61/A sky130_fd_sc_hd__inv_2_61/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_72 sky130_fd_sc_hd__inv_2_72/A sky130_fd_sc_hd__inv_2_72/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_83 sky130_fd_sc_hd__inv_2_83/A sky130_fd_sc_hd__inv_2_83/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_94 sky130_fd_sc_hd__inv_2_94/A sky130_fd_sc_hd__inv_2_94/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__ha_2_15 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_15/A sky130_fd_sc_hd__ha_2_14/B
+ sky130_fd_sc_hd__ha_2_15/SUM sky130_fd_sc_hd__ha_2_15/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_26 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_26/A sky130_fd_sc_hd__ha_2_25/B
+ sky130_fd_sc_hd__ha_2_26/SUM sky130_fd_sc_hd__ha_2_26/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_37 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_37/A sky130_fd_sc_hd__ha_2_36/B
+ sky130_fd_sc_hd__ha_2_37/SUM sky130_fd_sc_hd__ha_2_37/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_48 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_48/A sky130_fd_sc_hd__ha_2_47/B
+ sky130_fd_sc_hd__ha_2_48/SUM sky130_fd_sc_hd__ha_2_48/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_59 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_59/A sky130_fd_sc_hd__ha_2_58/B
+ sky130_fd_sc_hd__ha_2_59/SUM sky130_fd_sc_hd__ha_2_59/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_370 sky130_fd_sc_hd__fa_2_372/CIN sky130_fd_sc_hd__fa_2_366/A
+ sky130_fd_sc_hd__fa_2_370/A sky130_fd_sc_hd__fa_2_370/B sky130_fd_sc_hd__fa_2_370/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_11 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__clkinv_4_53/Y
+ sky130_fd_sc_hd__dfxtp_1_95/CLK sky130_fd_sc_hd__or2_0_0/X VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_381 sky130_fd_sc_hd__fa_2_383/CIN sky130_fd_sc_hd__fa_2_377/A
+ sky130_fd_sc_hd__fa_2_381/A sky130_fd_sc_hd__fa_2_381/B sky130_fd_sc_hd__fa_2_381/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_22 sky130_fd_sc_hd__conb_1_14/LO sky130_fd_sc_hd__clkinv_4_51/A
+ sky130_fd_sc_hd__dfxtp_1_207/CLK sky130_fd_sc_hd__nand3_1_36/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_392 sky130_fd_sc_hd__fa_2_396/B sky130_fd_sc_hd__fa_2_392/SUM
+ sky130_fd_sc_hd__fa_2_392/A sky130_fd_sc_hd__fa_2_392/B sky130_fd_sc_hd__fa_2_392/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22oi_2_3 sky130_fd_sc_hd__nor3_2_0/A sky130_fd_sc_hd__buf_2_281/X
+ sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__dfxtp_1_62/D sky130_fd_sc_hd__a22oi_2_3/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__sdlclkp_4_33 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_58/A
+ sky130_fd_sc_hd__dfxtp_1_313/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__clkbuf_16_15 sky130_fd_sc_hd__buf_12_506/A sky130_fd_sc_hd__inv_2_130/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__sdlclkp_4_44 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_68/Y
+ sky130_fd_sc_hd__dfxtp_1_411/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__diode_2_220 sig_amplitude[3] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__sdlclkp_4_55 sky130_fd_sc_hd__conb_1_20/LO sky130_fd_sc_hd__clkinv_8_62/Y
+ sky130_fd_sc_hd__dfxtp_1_538/CLK sky130_fd_sc_hd__o21ai_1_32/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__diode_2_231 sig_frequency[1] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__sdlclkp_4_66 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__clkinv_8_61/Y
+ sky130_fd_sc_hd__dfxtp_1_488/CLK sky130_fd_sc_hd__nand2b_1_5/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_77 sky130_fd_sc_hd__conb_1_24/LO sky130_fd_sc_hd__clkinv_8_96/A
+ sky130_fd_sc_hd__dfxtp_1_747/CLK sky130_fd_sc_hd__or2_0_8/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_88 sky130_fd_sc_hd__conb_1_28/LO sky130_fd_sc_hd__clkinv_8_47/A
+ sky130_fd_sc_hd__dfxtp_1_1329/CLK sky130_fd_sc_hd__or2_0_12/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_102 sky130_fd_sc_hd__nor2_1_102/B sky130_fd_sc_hd__nor2_1_95/A
+ sky130_fd_sc_hd__fa_2_1113/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_113 sky130_fd_sc_hd__nor2_1_113/B sky130_fd_sc_hd__o21a_1_9/A1
+ sky130_fd_sc_hd__o21a_1_10/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_124 sky130_fd_sc_hd__nor2_1_135/Y sky130_fd_sc_hd__nor2_1_124/Y
+ sky130_fd_sc_hd__nand2_2_6/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_135 sky130_fd_sc_hd__nor2_1_135/B sky130_fd_sc_hd__nor2_1_135/Y
+ sky130_fd_sc_hd__nor2_1_135/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_11 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__a22oi_1_9/A1
+ sky130_fd_sc_hd__buf_2_288/X sky130_fd_sc_hd__a22oi_1_11/A2 sky130_fd_sc_hd__nand3_1_5/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_22 sky130_fd_sc_hd__nor2_2_0/Y sky130_fd_sc_hd__clkinv_1_4/Y
+ sky130_fd_sc_hd__nand4_1_20/Y sky130_fd_sc_hd__nand4_1_4/Y sky130_fd_sc_hd__a22oi_1_22/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_146 sky130_fd_sc_hd__nor2_1_146/B sky130_fd_sc_hd__o21a_1_21/A1
+ sky130_fd_sc_hd__nor2_1_146/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_33 sky130_fd_sc_hd__nor2_2_2/Y sky130_fd_sc_hd__a22oi_1_82/A1
+ sky130_fd_sc_hd__clkbuf_1_69/X sky130_fd_sc_hd__a22oi_1_33/A2 sky130_fd_sc_hd__nand4_1_1/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_157 sky130_fd_sc_hd__nor2_1_157/B sky130_fd_sc_hd__nor2_1_157/Y
+ sky130_fd_sc_hd__nor2_1_157/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_44 sky130_fd_sc_hd__a22oi_1_81/B1 sky130_fd_sc_hd__clkbuf_1_99/X
+ sky130_fd_sc_hd__clkbuf_1_46/X sky130_fd_sc_hd__clkbuf_4_21/X sky130_fd_sc_hd__nand4_1_4/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_168 sky130_fd_sc_hd__a21o_2_8/A2 sky130_fd_sc_hd__a21o_2_8/B1
+ sky130_fd_sc_hd__a21o_2_8/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_55 sky130_fd_sc_hd__clkbuf_4_8/X sky130_fd_sc_hd__clkbuf_4_9/X
+ sky130_fd_sc_hd__clkbuf_1_26/X sky130_fd_sc_hd__a22oi_1_55/A2 sky130_fd_sc_hd__a22oi_1_55/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_179 sky130_fd_sc_hd__nor2_1_179/B sky130_fd_sc_hd__nor2_1_179/Y
+ sky130_fd_sc_hd__nor2_1_182/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_66 sky130_fd_sc_hd__nor2_2_2/Y sky130_fd_sc_hd__a22oi_1_82/A1
+ sky130_fd_sc_hd__clkbuf_1_59/X sky130_fd_sc_hd__a22oi_1_66/A2 sky130_fd_sc_hd__nand4_1_11/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_77 sky130_fd_sc_hd__a22oi_1_81/B1 sky130_fd_sc_hd__clkbuf_1_99/X
+ sky130_fd_sc_hd__clkbuf_1_36/X sky130_fd_sc_hd__clkbuf_4_11/X sky130_fd_sc_hd__nand4_1_14/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_88 sky130_fd_sc_hd__a22oi_1_96/B1 sky130_fd_sc_hd__a22oi_1_96/A1
+ sky130_fd_sc_hd__a22oi_1_88/B2 sky130_fd_sc_hd__a22oi_1_88/A2 sky130_fd_sc_hd__nand4_1_17/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_99 sky130_fd_sc_hd__clkbuf_4_72/X sky130_fd_sc_hd__clkbuf_4_73/X
+ sky130_fd_sc_hd__a22oi_1_99/B2 sky130_fd_sc_hd__buf_2_94/X sky130_fd_sc_hd__buf_2_109/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_320 sky130_fd_sc_hd__buf_4_74/X sky130_fd_sc_hd__buf_8_173/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_331 sky130_fd_sc_hd__buf_4_71/X sky130_fd_sc_hd__buf_12_331/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_342 sky130_fd_sc_hd__buf_6_43/X sky130_fd_sc_hd__buf_12_342/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_201 sky130_fd_sc_hd__clkbuf_4_111/X sky130_fd_sc_hd__clkbuf_4_112/X
+ sky130_fd_sc_hd__a22oi_1_201/B2 sky130_fd_sc_hd__clkbuf_1_284/X sky130_fd_sc_hd__a22oi_1_201/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_353 sky130_fd_sc_hd__buf_12_353/A sky130_fd_sc_hd__buf_12_353/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_212 sky130_fd_sc_hd__nor2_4_7/Y sky130_fd_sc_hd__buf_2_165/X
+ sky130_fd_sc_hd__a22oi_1_212/B2 sky130_fd_sc_hd__clkbuf_1_454/X sky130_fd_sc_hd__a22oi_1_212/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_364 sky130_fd_sc_hd__buf_12_364/A sky130_fd_sc_hd__buf_12_364/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_223 sky130_fd_sc_hd__buf_2_164/X sky130_fd_sc_hd__nor2_4_8/Y
+ sky130_fd_sc_hd__buf_2_186/X sky130_fd_sc_hd__clkbuf_1_457/X sky130_fd_sc_hd__nand4_1_52/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_375 sky130_fd_sc_hd__buf_12_375/A sky130_fd_sc_hd__buf_12_375/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_234 sky130_fd_sc_hd__buf_2_166/X sky130_fd_sc_hd__buf_2_167/X
+ sky130_fd_sc_hd__clkbuf_1_432/X sky130_fd_sc_hd__buf_2_175/X sky130_fd_sc_hd__nand4_1_56/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_386 sky130_fd_sc_hd__buf_12_386/A sky130_fd_sc_hd__buf_12_437/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_245 sky130_fd_sc_hd__buf_2_166/X sky130_fd_sc_hd__buf_2_167/X
+ sky130_fd_sc_hd__clkbuf_1_429/X sky130_fd_sc_hd__buf_2_171/X sky130_fd_sc_hd__nand4_1_60/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_397 sky130_fd_sc_hd__buf_12_397/A sky130_fd_sc_hd__buf_12_484/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_256 sky130_fd_sc_hd__buf_2_164/X sky130_fd_sc_hd__nor2_4_8/Y
+ sky130_fd_sc_hd__clkbuf_1_414/X sky130_fd_sc_hd__buf_2_223/X sky130_fd_sc_hd__nand4_1_63/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_267 sky130_fd_sc_hd__nor2_2_4/Y sky130_fd_sc_hd__clkbuf_1_377/X
+ sky130_fd_sc_hd__a22oi_1_267/B2 sky130_fd_sc_hd__clkbuf_4_190/X sky130_fd_sc_hd__nand4_1_66/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_278 sky130_fd_sc_hd__clkbuf_1_378/X sky130_fd_sc_hd__clkbuf_1_379/X
+ sky130_fd_sc_hd__clkbuf_4_171/X sky130_fd_sc_hd__buf_2_197/X sky130_fd_sc_hd__nand4_1_69/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_520 sky130_fd_sc_hd__nor2_1_52/B sky130_fd_sc_hd__fa_2_1037/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_520/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22oi_1_289 sky130_fd_sc_hd__clkbuf_4_165/X sky130_fd_sc_hd__clkinv_2_23/Y
+ sky130_fd_sc_hd__clkbuf_1_405/X sky130_fd_sc_hd__a22oi_1_289/A2 sky130_fd_sc_hd__a22oi_1_289/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_531 sky130_fd_sc_hd__o21ai_1_91/A2 sky130_fd_sc_hd__fa_2_998/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_531/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_4_107 VDD VSS sky130_fd_sc_hd__buf_4_112/A sky130_fd_sc_hd__buf_4_107/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__clkinv_1_542 sky130_fd_sc_hd__o22ai_1_99/A2 sky130_fd_sc_hd__nand3_1_49/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_542/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_4_118 VDD VSS sky130_fd_sc_hd__buf_4_118/X sky130_fd_sc_hd__buf_8_216/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__clkinv_1_553 sky130_fd_sc_hd__o22ai_1_117/A1 sky130_fd_sc_hd__fa_2_982/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_553/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_564 sky130_fd_sc_hd__clkinv_1_564/Y sky130_fd_sc_hd__a222oi_1_1/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_564/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_575 sky130_fd_sc_hd__nor2_1_86/A sky130_fd_sc_hd__fa_2_1012/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_575/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_586 sky130_fd_sc_hd__o21ai_1_156/A2 sky130_fd_sc_hd__fa_2_1000/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_586/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_597 sky130_fd_sc_hd__ha_2_172/B sky130_fd_sc_hd__fa_2_1043/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_597/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_4_11 sky130_fd_sc_hd__clkinv_2_7/A sky130_fd_sc_hd__clkinv_4_11/Y
+ VSS VDD VDD VSS VSS sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_22 sky130_fd_sc_hd__clkinv_4_22/A sky130_fd_sc_hd__clkinv_4_22/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_22/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_33 sky130_fd_sc_hd__clkinv_4_75/Y sky130_fd_sc_hd__clkinv_4_33/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_33/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_44 sky130_fd_sc_hd__clkinv_8_99/Y sky130_fd_sc_hd__clkinv_4_45/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_44/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_55 sky130_fd_sc_hd__clkinv_4_55/A sky130_fd_sc_hd__clkinv_8_68/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_55/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_66 sky130_fd_sc_hd__clkinv_4_66/A sky130_fd_sc_hd__clkinv_4_67/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_66/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_77 sky130_fd_sc_hd__clkinv_4_78/A sky130_fd_sc_hd__clkinv_4_77/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_77/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__inv_16_7 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__a21oi_1_450 sky130_fd_sc_hd__nor2_1_309/Y sky130_fd_sc_hd__nor2_1_300/Y
+ sky130_fd_sc_hd__a21oi_1_450/Y sky130_fd_sc_hd__fa_2_1283/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_461 sky130_fd_sc_hd__a21oi_1_464/A1 sky130_fd_sc_hd__a21oi_1_461/B1
+ sky130_fd_sc_hd__a21oi_1_461/Y sky130_fd_sc_hd__nand2_1_543/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_472 sky130_fd_sc_hd__nor3_1_41/A sky130_fd_sc_hd__o22ai_1_427/Y
+ sky130_fd_sc_hd__a21oi_1_472/Y sky130_fd_sc_hd__fa_2_1308/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_483 sky130_fd_sc_hd__nor2_1_314/Y sky130_fd_sc_hd__nand3_1_52/B
+ sky130_fd_sc_hd__a31oi_1_3/A1 sky130_fd_sc_hd__nand3_1_5/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_494 sky130_fd_sc_hd__or2_0_13/B sky130_fd_sc_hd__or2_0_0/B
+ sky130_fd_sc_hd__nand2_1_562/A sky130_fd_sc_hd__nor2_1_320/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_8_130 sky130_fd_sc_hd__clkinv_8_131/A sky130_fd_sc_hd__clkinv_4_72/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_130/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__xor2_1_305 sky130_fd_sc_hd__nor2_4_20/Y sky130_fd_sc_hd__fa_2_1305/B
+ sky130_fd_sc_hd__xor2_1_305/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_316 sky130_fd_sc_hd__nor2_4_20/Y sky130_fd_sc_hd__fa_2_1294/B
+ sky130_fd_sc_hd__xor2_1_316/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nor2b_1_90 sky130_fd_sc_hd__buf_2_263/X sky130_fd_sc_hd__nor2b_1_90/Y
+ sky130_fd_sc_hd__a32o_1_0/A3 VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1090 sky130_fd_sc_hd__o21ai_1_473/A2 sky130_fd_sc_hd__o21ai_1_484/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1090/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkbuf_1_309 VSS VDD sky130_fd_sc_hd__nand4_1_36/D sky130_fd_sc_hd__a22oi_1_163/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_13 VDD VSS sky130_fd_sc_hd__or2_1_1/A sky130_fd_sc_hd__dfxtp_1_8/CLK
+ sky130_fd_sc_hd__nor3_1_1/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_24 VDD VSS sky130_fd_sc_hd__ha_2_115/B sky130_fd_sc_hd__dfxtp_1_29/CLK
+ sky130_fd_sc_hd__buf_2_288/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_35 VDD VSS sky130_fd_sc_hd__fa_2_906/CIN sky130_fd_sc_hd__dfxtp_1_39/CLK
+ sky130_fd_sc_hd__nand4_1_37/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_46 VDD VSS sky130_fd_sc_hd__ha_2_119/A sky130_fd_sc_hd__dfxtp_1_60/CLK
+ sky130_fd_sc_hd__dfxtp_1_62/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_57 VDD VSS sky130_fd_sc_hd__ha_2_125/B sky130_fd_sc_hd__dfxtp_1_61/CLK
+ sky130_fd_sc_hd__buf_2_287/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_68 VDD VSS sky130_fd_sc_hd__ha_2_95/A sky130_fd_sc_hd__dfxtp_1_73/CLK
+ sky130_fd_sc_hd__nand4_1_38/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_79 VDD VSS sky130_fd_sc_hd__o21ai_1_0/A1 sky130_fd_sc_hd__dfxtp_1_83/CLK
+ sky130_fd_sc_hd__a31oi_1_0/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_4_103 sky130_fd_sc_hd__clkbuf_4_103/X sky130_fd_sc_hd__dfxtp_1_1463/Q
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_114 sky130_fd_sc_hd__clkbuf_4_114/X sky130_fd_sc_hd__clkbuf_4_114/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_125 sky130_fd_sc_hd__clkbuf_4_125/X sky130_fd_sc_hd__clkbuf_4_125/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_136 sky130_fd_sc_hd__clkbuf_4_136/X sky130_fd_sc_hd__clkbuf_4_136/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_307 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_307/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_307/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_147 sky130_fd_sc_hd__nand4_1_38/B sky130_fd_sc_hd__a22oi_1_173/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_318 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_318/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_318/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_158 sky130_fd_sc_hd__buf_6_35/A sky130_fd_sc_hd__buf_4_69/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_329 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_329/X sky130_fd_sc_hd__inv_2_139/Y
+ sky130_fd_sc_hd__and2_0_329/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_169 sky130_fd_sc_hd__clkbuf_4_169/X sky130_fd_sc_hd__clkbuf_4_169/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__inv_2_107 sky130_fd_sc_hd__inv_2_107/A sky130_fd_sc_hd__inv_2_107/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_4_90 VDD VSS sky130_fd_sc_hd__buf_4_90/X sky130_fd_sc_hd__buf_6_33/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__inv_2_118 sky130_fd_sc_hd__inv_2_118/A sky130_fd_sc_hd__inv_2_118/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__or2_0_9 sky130_fd_sc_hd__or2_0_9/A sky130_fd_sc_hd__or2_0_9/X sky130_fd_sc_hd__or2_0_9/B
+ VSS VDD VSS VDD sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__inv_2_129 sky130_fd_sc_hd__inv_2_129/A sky130_fd_sc_hd__inv_2_129/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_12_150 sky130_fd_sc_hd__buf_12_150/A sky130_fd_sc_hd__buf_12_228/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_161 sky130_fd_sc_hd__buf_8_81/X sky130_fd_sc_hd__buf_12_213/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_172 sky130_fd_sc_hd__buf_12_172/A sky130_fd_sc_hd__buf_12_172/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_183 sky130_fd_sc_hd__buf_12_183/A sky130_fd_sc_hd__buf_12_183/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_194 sky130_fd_sc_hd__buf_4_55/X sky130_fd_sc_hd__buf_12_226/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_350 sky130_fd_sc_hd__ha_2_128/A sky130_fd_sc_hd__ha_2_133/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_350/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_361 sky130_fd_sc_hd__fa_2_826/A sky130_fd_sc_hd__fa_2_834/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_361/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_372 sky130_fd_sc_hd__fa_2_876/B sky130_fd_sc_hd__dfxtp_1_276/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_372/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_383 sky130_fd_sc_hd__fa_2_865/B sky130_fd_sc_hd__dfxtp_1_265/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_383/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_394 sky130_fd_sc_hd__fa_2_878/B sky130_fd_sc_hd__nand2_1_33/A
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a211o_1_8 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_76/A sky130_fd_sc_hd__a211o_1_8/A2
+ sky130_fd_sc_hd__o22ai_1_96/Y sky130_fd_sc_hd__a211o_1_8/A1 sky130_fd_sc_hd__nor2_1_77/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o21a_1_13 sky130_fd_sc_hd__o21a_1_13/X sky130_fd_sc_hd__o21a_1_13/A1
+ sky130_fd_sc_hd__o21a_1_13/B1 sky130_fd_sc_hd__fa_2_1058/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21ai_1_308 VSS VDD sky130_fd_sc_hd__nor2_1_144/B sky130_fd_sc_hd__o21a_1_29/A1
+ sky130_fd_sc_hd__a21oi_1_280/Y sky130_fd_sc_hd__o21ai_1_308/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_319 VSS VDD sky130_fd_sc_hd__a211oi_1_16/Y sky130_fd_sc_hd__nor2_1_172/A
+ sky130_fd_sc_hd__a21oi_1_288/Y sky130_fd_sc_hd__o21ai_1_319/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_24 sky130_fd_sc_hd__o21a_1_24/X sky130_fd_sc_hd__o21a_1_24/A1
+ sky130_fd_sc_hd__o21a_1_24/B1 sky130_fd_sc_hd__fa_2_1154/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_35 sky130_fd_sc_hd__o21a_1_35/X sky130_fd_sc_hd__o21a_1_35/A1
+ sky130_fd_sc_hd__o21a_1_35/B1 sky130_fd_sc_hd__fa_2_1178/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_46 sky130_fd_sc_hd__o21a_1_46/X sky130_fd_sc_hd__o21a_1_46/A1
+ sky130_fd_sc_hd__o21a_1_46/B1 sky130_fd_sc_hd__fa_2_1234/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_57 sky130_fd_sc_hd__o21a_1_57/X sky130_fd_sc_hd__o21a_1_57/A1
+ sky130_fd_sc_hd__o21a_1_57/B1 sky130_fd_sc_hd__fa_2_1289/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_68 sky130_fd_sc_hd__o21a_1_68/X sky130_fd_sc_hd__o21a_1_68/A1
+ sky130_fd_sc_hd__o21a_1_68/B1 sky130_fd_sc_hd__o21a_1_68/A2 VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__a21oi_1_280 sky130_fd_sc_hd__fa_2_1132/A sky130_fd_sc_hd__o22ai_1_252/Y
+ sky130_fd_sc_hd__a21oi_1_280/Y sky130_fd_sc_hd__nor2_2_15/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_291 sky130_fd_sc_hd__or2_0_9/B sky130_fd_sc_hd__o21ai_1_321/Y
+ sky130_fd_sc_hd__a21oi_1_291/Y sky130_fd_sc_hd__o21ai_1_322/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_210 sky130_fd_sc_hd__buf_8_210/A sky130_fd_sc_hd__buf_8_210/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_221 sky130_fd_sc_hd__buf_8_221/A sky130_fd_sc_hd__buf_8_221/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xor2_1_102 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1055/B
+ sky130_fd_sc_hd__xor2_1_102/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_113 sky130_fd_sc_hd__xor2_1_114/X sky130_fd_sc_hd__xor2_1_113/X
+ sky130_fd_sc_hd__xor2_1_88/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_124 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1082/B
+ sky130_fd_sc_hd__xor2_1_124/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_135 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1071/B
+ sky130_fd_sc_hd__xor2_1_135/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_146 sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__fa_2_1137/B
+ sky130_fd_sc_hd__xor2_1_146/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_157 sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__fa_2_1126/B
+ sky130_fd_sc_hd__xor2_1_157/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_508 VDD VSS sky130_fd_sc_hd__nor4_1_12/C sky130_fd_sc_hd__edfxtp_1_0/CLK
+ sky130_fd_sc_hd__a22o_1_63/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_168 sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__fa_2_1154/B
+ sky130_fd_sc_hd__xor2_1_168/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_519 VDD VSS sky130_fd_sc_hd__nor4_1_9/C sky130_fd_sc_hd__dfxtp_1_520/CLK
+ sky130_fd_sc_hd__a22o_1_52/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_179 sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__fa_2_1143/B
+ sky130_fd_sc_hd__xor2_1_179/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_106 VSS VDD sky130_fd_sc_hd__buf_8_33/A sky130_fd_sc_hd__buf_12_91/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_117 VSS VDD sky130_fd_sc_hd__clkbuf_1_118/A sky130_fd_sc_hd__buf_8_18/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_128 VSS VDD sky130_fd_sc_hd__inv_16_1/A sky130_fd_sc_hd__inv_2_44/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_139 VSS VDD sky130_fd_sc_hd__clkbuf_1_139/X sky130_fd_sc_hd__clkbuf_1_139/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_8 VDD VSS sky130_fd_sc_hd__dfxtp_1_8/Q sky130_fd_sc_hd__dfxtp_1_8/CLK
+ sky130_fd_sc_hd__a22o_1_5/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand3_1_17 sky130_fd_sc_hd__nand3_1_17/Y sky130_fd_sc_hd__nor3_1_4/A
+ sky130_fd_sc_hd__nand3_1_17/C sky130_fd_sc_hd__nor3_2_1/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_28 sky130_fd_sc_hd__nand3_1_28/Y sky130_fd_sc_hd__ha_2_30/A
+ sky130_fd_sc_hd__nand3_1_30/C sky130_fd_sc_hd__nand3_2_2/A VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_39 sky130_fd_sc_hd__nand3_1_39/Y sky130_fd_sc_hd__or2_1_1/X
+ sky130_fd_sc_hd__nand3_2_8/B sky130_fd_sc_hd__a22o_1_27/X VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__dfxtp_1_1404 VDD VSS sky130_fd_sc_hd__mux2_2_233/A0 sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__o22ai_1_385/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1415 VDD VSS sky130_fd_sc_hd__mux2_2_263/A0 sky130_fd_sc_hd__clkinv_8_102/Y
+ sky130_fd_sc_hd__dfxtp_1_430/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1426 VDD VSS sky130_fd_sc_hd__mux2_2_257/A0 sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__a21oi_1_439/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1437 VDD VSS sky130_fd_sc_hd__mux2_2_228/A1 sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__o22ai_1_396/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1448 VDD VSS sky130_fd_sc_hd__nor2_1_314/A sky130_fd_sc_hd__clkinv_8_116/Y
+ sky130_fd_sc_hd__nor2b_1_133/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1459 VDD VSS sky130_fd_sc_hd__buf_6_88/A sky130_fd_sc_hd__dfxtp_1_1461/CLK
+ sky130_fd_sc_hd__and2_0_342/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_104 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_104/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_888/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_12 sky130_fd_sc_hd__nand3_1_25/C sky130_fd_sc_hd__xor2_1_1/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_12/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_115 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_115/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_918/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_23 sky130_fd_sc_hd__inv_2_12/A sky130_fd_sc_hd__inv_2_11/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_23/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_126 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_126/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__fa_2_867/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_34 sky130_fd_sc_hd__inv_2_23/A sky130_fd_sc_hd__inv_2_4/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_34/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_137 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_137/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_894/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_45 sky130_fd_sc_hd__inv_2_34/A sky130_fd_sc_hd__buf_8_1/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_45/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_148 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_148/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_844/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_56 sky130_fd_sc_hd__bufinv_8_0/A sky130_fd_sc_hd__buf_8_4/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_56/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_159 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_159/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_898/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_67 sky130_fd_sc_hd__nand3_1_31/C sky130_fd_sc_hd__xor2_1_4/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_67/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_78 sky130_fd_sc_hd__buf_8_88/A sky130_fd_sc_hd__clkinv_2_4/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_78/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_89 sky130_fd_sc_hd__inv_2_55/A sky130_fd_sc_hd__ha_2_43/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_89/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_903 sky130_fd_sc_hd__fa_2_899/A sky130_fd_sc_hd__fa_2_900/B
+ sky130_fd_sc_hd__fa_2_903/A sky130_fd_sc_hd__fa_2_903/B sky130_fd_sc_hd__fa_2_903/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_914 sky130_fd_sc_hd__fa_2_888/A sky130_fd_sc_hd__fa_2_889/B
+ sky130_fd_sc_hd__fa_2_914/A sky130_fd_sc_hd__fa_2_914/B sky130_fd_sc_hd__fa_2_914/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_925 sky130_fd_sc_hd__fa_2_924/CIN sky130_fd_sc_hd__fa_2_925/SUM
+ sky130_fd_sc_hd__fa_2_925/A sky130_fd_sc_hd__fa_2_925/B sky130_fd_sc_hd__fa_2_925/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_936 sky130_fd_sc_hd__fa_2_922/A sky130_fd_sc_hd__fa_2_923/B
+ sky130_fd_sc_hd__fa_2_936/A sky130_fd_sc_hd__fa_2_936/B sky130_fd_sc_hd__fa_2_535/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_947 sky130_fd_sc_hd__fa_2_946/CIN sky130_fd_sc_hd__fa_2_947/SUM
+ sky130_fd_sc_hd__fa_2_947/A sky130_fd_sc_hd__fa_2_947/B sky130_fd_sc_hd__fa_2_947/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_958 sky130_fd_sc_hd__fa_2_957/CIN sky130_fd_sc_hd__fa_2_958/SUM
+ sky130_fd_sc_hd__or3_1_1/B sky130_fd_sc_hd__fa_2_958/B sky130_fd_sc_hd__fa_2_958/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_969 sky130_fd_sc_hd__fa_2_968/CIN sky130_fd_sc_hd__fa_2_969/SUM
+ sky130_fd_sc_hd__fa_2_969/A sky130_fd_sc_hd__fa_2_969/B sky130_fd_sc_hd__fa_2_969/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__mux2_2_203 VSS VDD sky130_fd_sc_hd__mux2_2_203/A1 sky130_fd_sc_hd__mux2_2_203/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_203/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_214 VSS VDD sky130_fd_sc_hd__mux2_2_214/A1 sky130_fd_sc_hd__mux2_2_214/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_214/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_225 VSS VDD sky130_fd_sc_hd__mux2_2_225/A1 sky130_fd_sc_hd__mux2_2_225/A0
+ sky130_fd_sc_hd__nor2_8_2/A sky130_fd_sc_hd__mux2_2_225/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_236 VSS VDD sky130_fd_sc_hd__xor2_1_318/X sky130_fd_sc_hd__nand2_1_520/B
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_236/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_247 VSS VDD sky130_fd_sc_hd__mux2_2_247/A1 sky130_fd_sc_hd__mux2_2_247/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_247/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_258 VSS VDD sky130_fd_sc_hd__mux2_2_258/A1 sky130_fd_sc_hd__mux2_2_258/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_258/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__buf_8_1 sky130_fd_sc_hd__buf_8_1/A sky130_fd_sc_hd__buf_8_1/X VSS
+ VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__a22o_1_3 sky130_fd_sc_hd__a22o_1_3/A1 sky130_fd_sc_hd__nor2_1_1/Y
+ sky130_fd_sc_hd__a22o_1_3/X sky130_fd_sc_hd__a22o_1_3/B2 sky130_fd_sc_hd__nor2_1_0/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_180 sky130_fd_sc_hd__bufinv_8_8/A sky130_fd_sc_hd__buf_8_131/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_180/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_191 sky130_fd_sc_hd__nor3_1_24/C sky130_fd_sc_hd__nor3_2_10/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_191/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_60 sky130_fd_sc_hd__a22o_1_60/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_60/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__nor4_1_11/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_71 sky130_fd_sc_hd__a22o_1_73/A1 sky130_fd_sc_hd__a22o_1_73/B2
+ sky130_fd_sc_hd__a22o_1_71/X sky130_fd_sc_hd__ha_2_201/SUM sky130_fd_sc_hd__a22o_1_73/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__o21ai_1_105 VSS VDD sky130_fd_sc_hd__nor2_1_79/Y sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__a21oi_1_89/Y sky130_fd_sc_hd__xor2_1_72/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_116 VSS VDD sky130_fd_sc_hd__nor2_1_69/B sky130_fd_sc_hd__o21a_1_8/A2
+ sky130_fd_sc_hd__a21oi_1_101/Y sky130_fd_sc_hd__a211o_1_7/A2 VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_127 VSS VDD sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__a21oi_1_108/Y sky130_fd_sc_hd__xor2_1_43/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_138 VSS VDD sky130_fd_sc_hd__nor2_1_88/A sky130_fd_sc_hd__o21ai_1_92/A1
+ sky130_fd_sc_hd__a22oi_1_335/Y sky130_fd_sc_hd__o21ai_1_138/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_149 VSS VDD sky130_fd_sc_hd__o22ai_1_123/B2 sky130_fd_sc_hd__o21ai_1_92/A1
+ sky130_fd_sc_hd__a22oi_1_340/Y sky130_fd_sc_hd__o21ai_1_149/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__maj3_1_11 sky130_fd_sc_hd__maj3_1_12/X sky130_fd_sc_hd__maj3_1_11/X
+ sky130_fd_sc_hd__maj3_1_11/B sky130_fd_sc_hd__maj3_1_11/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_22 sky130_fd_sc_hd__maj3_1_23/X sky130_fd_sc_hd__maj3_1_22/X
+ sky130_fd_sc_hd__maj3_1_22/B sky130_fd_sc_hd__maj3_1_22/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_401 sky130_fd_sc_hd__nand2_1_516/Y sky130_fd_sc_hd__nand2_1_515/Y
+ sky130_fd_sc_hd__o22ai_1_401/Y sky130_fd_sc_hd__o22ai_1_401/A1 sky130_fd_sc_hd__a21o_2_27/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_33 sky130_fd_sc_hd__maj3_1_34/X sky130_fd_sc_hd__maj3_1_33/X
+ sky130_fd_sc_hd__maj3_1_33/B sky130_fd_sc_hd__maj3_1_33/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_412 sky130_fd_sc_hd__nor2_1_299/A sky130_fd_sc_hd__nor2_1_310/A
+ sky130_fd_sc_hd__o22ai_1_412/Y sky130_fd_sc_hd__a21boi_1_7/Y sky130_fd_sc_hd__a222oi_1_36/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_44 sky130_fd_sc_hd__maj3_1_45/X sky130_fd_sc_hd__maj3_1_44/X
+ sky130_fd_sc_hd__maj3_1_44/B sky130_fd_sc_hd__maj3_1_44/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_423 sky130_fd_sc_hd__o22ai_1_436/A2 sky130_fd_sc_hd__o22ai_1_423/B1
+ sky130_fd_sc_hd__o22ai_1_423/Y sky130_fd_sc_hd__nor2_1_272/B sky130_fd_sc_hd__o32ai_1_11/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__inv_8_1 sky130_fd_sc_hd__inv_8_1/A sky130_fd_sc_hd__inv_8_1/Y VSS
+ VDD VSS VDD sky130_fd_sc_hd__inv_8
Xsky130_fd_sc_hd__maj3_1_55 sky130_fd_sc_hd__maj3_1_55/C sky130_fd_sc_hd__maj3_1_55/X
+ sky130_fd_sc_hd__maj3_1_55/B sky130_fd_sc_hd__maj3_1_55/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_434 sky130_fd_sc_hd__o22ai_1_436/A2 sky130_fd_sc_hd__nor2_1_308/A
+ sky130_fd_sc_hd__o22ai_1_434/Y sky130_fd_sc_hd__nor2_1_278/B sky130_fd_sc_hd__o32ai_1_11/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_66 sky130_fd_sc_hd__maj3_1_67/X sky130_fd_sc_hd__maj3_1_66/X
+ sky130_fd_sc_hd__maj3_1_66/B sky130_fd_sc_hd__maj3_1_66/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_509 sky130_fd_sc_hd__o21a_1_66/B1 sky130_fd_sc_hd__fa_2_1301/A
+ sky130_fd_sc_hd__o21a_1_66/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_77 sky130_fd_sc_hd__maj3_1_78/X sky130_fd_sc_hd__maj3_1_77/X
+ sky130_fd_sc_hd__maj3_1_77/B sky130_fd_sc_hd__maj3_1_77/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_88 sky130_fd_sc_hd__maj3_1_89/X sky130_fd_sc_hd__maj3_1_88/X
+ sky130_fd_sc_hd__maj3_1_88/B sky130_fd_sc_hd__maj3_1_88/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_99 sky130_fd_sc_hd__maj3_1_99/C sky130_fd_sc_hd__maj3_1_99/X
+ sky130_fd_sc_hd__maj3_1_99/B sky130_fd_sc_hd__maj3_1_99/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_50 sky130_fd_sc_hd__nand2_1_50/Y sky130_fd_sc_hd__nand2_1_51/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_61 sky130_fd_sc_hd__nand2_1_61/Y sky130_fd_sc_hd__nand2_1_5/B
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_72 sky130_fd_sc_hd__nand2_1_72/Y sky130_fd_sc_hd__nand2_1_73/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_83 sky130_fd_sc_hd__nand2_1_83/Y sky130_fd_sc_hd__nand2_1_83/B
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_94 sky130_fd_sc_hd__nand2_1_94/Y sky130_fd_sc_hd__nand2_1_95/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_305 VDD VSS sky130_fd_sc_hd__a22o_1_44/A1 sky130_fd_sc_hd__dfxtp_1_313/CLK
+ sky130_fd_sc_hd__and2_0_93/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_316 VDD VSS sky130_fd_sc_hd__or4_1_1/D sky130_fd_sc_hd__dfxtp_1_325/CLK
+ sky130_fd_sc_hd__and2_0_204/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_327 VDD VSS sky130_fd_sc_hd__a22o_1_28/B2 sky130_fd_sc_hd__clkinv_4_27/Y
+ sky130_fd_sc_hd__o21ai_1_19/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_338 VDD VSS sky130_fd_sc_hd__a22o_1_22/B2 sky130_fd_sc_hd__dfxtp_1_354/CLK
+ sky130_fd_sc_hd__ha_2_157/B VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_349 VDD VSS sky130_fd_sc_hd__ha_2_153/A sky130_fd_sc_hd__dfxtp_1_361/CLK
+ sky130_fd_sc_hd__o2bb2ai_1_1/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_13 sky130_fd_sc_hd__fa_2_9/B sky130_fd_sc_hd__fa_2_13/SUM sky130_fd_sc_hd__fa_2_2/A
+ sky130_fd_sc_hd__fa_2_87/A sky130_fd_sc_hd__fa_2_81/B VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_24 sky130_fd_sc_hd__fa_2_20/A sky130_fd_sc_hd__fa_2_25/A sky130_fd_sc_hd__fa_2_67/B
+ sky130_fd_sc_hd__fa_2_5/A sky130_fd_sc_hd__fa_2_2/B VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_35 sky130_fd_sc_hd__fa_2_36/A sky130_fd_sc_hd__fa_2_35/SUM
+ sky130_fd_sc_hd__ha_2_95/B sky130_fd_sc_hd__ha_2_94/B sky130_fd_sc_hd__fa_2_91/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_46 sky130_fd_sc_hd__fa_2_48/B sky130_fd_sc_hd__fa_2_44/A sky130_fd_sc_hd__fa_2_82/A
+ sky130_fd_sc_hd__ha_2_97/B sky130_fd_sc_hd__fa_2_92/B VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_57 sky130_fd_sc_hd__fa_2_56/A sky130_fd_sc_hd__fa_2_51/B sky130_fd_sc_hd__fa_2_57/A
+ sky130_fd_sc_hd__ha_2_97/A sky130_fd_sc_hd__fa_2_66/B VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_68 sky130_fd_sc_hd__fa_2_70/CIN sky130_fd_sc_hd__fa_2_63/A
+ sky130_fd_sc_hd__fa_2_68/A sky130_fd_sc_hd__fa_2_68/B sky130_fd_sc_hd__fa_2_75/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_79 sky130_fd_sc_hd__fa_2_84/B sky130_fd_sc_hd__fa_2_79/SUM
+ sky130_fd_sc_hd__fa_2_79/A sky130_fd_sc_hd__fa_2_79/B sky130_fd_sc_hd__fa_2_79/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_205 VDD VSS sky130_fd_sc_hd__buf_2_205/X sky130_fd_sc_hd__buf_2_205/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_216 VDD VSS sky130_fd_sc_hd__buf_2_216/X sky130_fd_sc_hd__buf_2_216/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_227 VDD VSS sky130_fd_sc_hd__buf_2_227/X sky130_fd_sc_hd__buf_2_227/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_238 VDD VSS sky130_fd_sc_hd__buf_8_203/A sky130_fd_sc_hd__buf_2_238/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_249 VDD VSS sky130_fd_sc_hd__buf_2_249/X sky130_fd_sc_hd__buf_2_249/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1201 VDD VSS sky130_fd_sc_hd__fa_2_1250/A sky130_fd_sc_hd__clkinv_8_75/Y
+ sky130_fd_sc_hd__mux2_2_194/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1212 VDD VSS sky130_fd_sc_hd__fa_2_1224/B sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__and2_0_329/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1223 VDD VSS sky130_fd_sc_hd__fa_2_1235/A sky130_fd_sc_hd__clkinv_8_78/Y
+ sky130_fd_sc_hd__mux2_2_187/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1234 VDD VSS sky130_fd_sc_hd__fa_2_1263/A sky130_fd_sc_hd__clkinv_8_63/Y
+ sky130_fd_sc_hd__mux2_2_216/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1245 VDD VSS sky130_fd_sc_hd__fa_2_1274/A sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__nand2_1_467/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1256 VDD VSS sky130_fd_sc_hd__mux2_2_204/A0 sky130_fd_sc_hd__clkinv_8_75/Y
+ sky130_fd_sc_hd__o22ai_1_335/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1267 VDD VSS sky130_fd_sc_hd__mux2_2_177/A1 sky130_fd_sc_hd__clkinv_8_116/Y
+ sky130_fd_sc_hd__o22ai_1_324/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1278 VDD VSS sky130_fd_sc_hd__mux2_2_205/A0 sky130_fd_sc_hd__clkinv_8_65/Y
+ sky130_fd_sc_hd__dfxtp_1_434/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_850 VDD VSS sky130_fd_sc_hd__mux2_2_53/A1 sky130_fd_sc_hd__clkinv_4_25/Y
+ sky130_fd_sc_hd__o21ai_1_167/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1289 VDD VSS sky130_fd_sc_hd__mux2_2_197/A0 sky130_fd_sc_hd__clkinv_8_75/Y
+ sky130_fd_sc_hd__o22ai_1_346/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_861 VDD VSS sky130_fd_sc_hd__mux2_2_72/A0 sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__o21ai_1_175/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_872 VDD VSS sky130_fd_sc_hd__mux2_2_48/A1 sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__o21ai_1_186/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_883 VDD VSS sky130_fd_sc_hd__fa_2_859/A sky130_fd_sc_hd__dfxtp_1_904/CLK
+ sky130_fd_sc_hd__dfxtp_1_883/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_894 VDD VSS sky130_fd_sc_hd__fa_2_930/CIN sky130_fd_sc_hd__dfxtp_1_899/CLK
+ sky130_fd_sc_hd__o32ai_1_0/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__or3_1_4 sky130_fd_sc_hd__or3_1_4/A sky130_fd_sc_hd__or3_1_4/X sky130_fd_sc_hd__or3_1_4/B
+ sky130_fd_sc_hd__or3_1_4/C VDD VSS VDD VSS sky130_fd_sc_hd__or3_1
Xsky130_fd_sc_hd__clkbuf_1_470 VSS VDD sky130_fd_sc_hd__clkbuf_1_470/X sky130_fd_sc_hd__clkbuf_1_470/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_481 VSS VDD sky130_fd_sc_hd__nand4_1_48/B sky130_fd_sc_hd__a22oi_1_212/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a21oi_1_18 sky130_fd_sc_hd__nor2_1_26/Y sky130_fd_sc_hd__dfxtp_1_572/Q
+ sky130_fd_sc_hd__nor2_1_25/B sky130_fd_sc_hd__or4_1_2/C VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkbuf_1_492 VSS VDD sky130_fd_sc_hd__clkbuf_1_492/X sky130_fd_sc_hd__clkbuf_1_492/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_700 sky130_fd_sc_hd__fa_2_570/A sky130_fd_sc_hd__fa_2_571/B
+ sky130_fd_sc_hd__fa_2_700/A sky130_fd_sc_hd__fa_2_700/B sky130_fd_sc_hd__fa_2_700/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a21oi_1_29 sky130_fd_sc_hd__nor2_1_41/Y sky130_fd_sc_hd__o22ai_1_62/Y
+ sky130_fd_sc_hd__a21oi_1_29/Y sky130_fd_sc_hd__fa_2_1032/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__fa_2_711 sky130_fd_sc_hd__fa_2_710/CIN sky130_fd_sc_hd__fa_2_711/SUM
+ sky130_fd_sc_hd__fa_2_711/A sky130_fd_sc_hd__fa_2_711/B sky130_fd_sc_hd__fa_2_711/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_722 sky130_fd_sc_hd__maj3_1_155/B sky130_fd_sc_hd__maj3_1_156/A
+ sky130_fd_sc_hd__fa_2_722/A sky130_fd_sc_hd__fa_2_722/B sky130_fd_sc_hd__fa_2_723/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_733 sky130_fd_sc_hd__fa_2_735/B sky130_fd_sc_hd__fa_2_733/SUM
+ sky130_fd_sc_hd__fa_2_733/A sky130_fd_sc_hd__fa_2_733/B sky130_fd_sc_hd__fa_2_733/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_744 sky130_fd_sc_hd__maj3_1_147/B sky130_fd_sc_hd__maj3_1_148/A
+ sky130_fd_sc_hd__fa_2_744/A sky130_fd_sc_hd__fa_2_744/B sky130_fd_sc_hd__fa_2_745/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_755 sky130_fd_sc_hd__fa_2_757/CIN sky130_fd_sc_hd__fa_2_752/A
+ sky130_fd_sc_hd__ha_2_140/B sky130_fd_sc_hd__fa_2_755/B sky130_fd_sc_hd__fa_2_755/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_766 sky130_fd_sc_hd__fa_2_767/B sky130_fd_sc_hd__fa_2_764/B
+ sky130_fd_sc_hd__fa_2_766/A sky130_fd_sc_hd__fa_2_766/B sky130_fd_sc_hd__fa_2_769/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_777 sky130_fd_sc_hd__fa_2_776/B sky130_fd_sc_hd__fa_2_777/SUM
+ sky130_fd_sc_hd__fa_2_829/A sky130_fd_sc_hd__ha_2_141/B sky130_fd_sc_hd__ha_2_141/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_788 sky130_fd_sc_hd__fa_2_787/B sky130_fd_sc_hd__fa_2_788/SUM
+ sky130_fd_sc_hd__ha_2_139/B sky130_fd_sc_hd__ha_2_141/B sky130_fd_sc_hd__ha_2_141/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_799 sky130_fd_sc_hd__fa_2_714/A sky130_fd_sc_hd__fa_2_715/B
+ sky130_fd_sc_hd__fa_2_799/A sky130_fd_sc_hd__fa_2_799/B sky130_fd_sc_hd__fa_2_805/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor2b_1_130 sky130_fd_sc_hd__o32ai_1_11/Y sky130_fd_sc_hd__nor2b_1_130/Y
+ sky130_fd_sc_hd__buf_2_262/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_141 sky130_fd_sc_hd__nor2_1_323/B sky130_fd_sc_hd__nor2b_1_141/Y
+ sky130_fd_sc_hd__nor2b_1_142/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__bufbuf_8_1 sky130_fd_sc_hd__inv_2_113/Y sky130_fd_sc_hd__buf_6_64/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufbuf_8
Xsky130_fd_sc_hd__buf_6_14 VDD VSS sky130_fd_sc_hd__buf_6_14/X sky130_fd_sc_hd__buf_6_14/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_25 VDD VSS sky130_fd_sc_hd__buf_6_25/X sky130_fd_sc_hd__buf_6_25/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_36 VDD VSS sky130_fd_sc_hd__buf_6_36/X sky130_fd_sc_hd__buf_6_36/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_47 VDD VSS sky130_fd_sc_hd__buf_6_47/X sky130_fd_sc_hd__buf_6_47/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_58 VDD VSS sky130_fd_sc_hd__buf_6_58/X sky130_fd_sc_hd__buf_6_58/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_69 VDD VSS sky130_fd_sc_hd__buf_6_69/X sky130_fd_sc_hd__buf_6_69/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_16 sky130_fd_sc_hd__buf_2_123/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_27 sky130_fd_sc_hd__buf_2_73/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_38 sky130_fd_sc_hd__buf_2_112/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_49 sky130_fd_sc_hd__buf_2_78/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__o22ai_1_220 sky130_fd_sc_hd__nand2_1_358/Y sky130_fd_sc_hd__nand2_1_357/Y
+ sky130_fd_sc_hd__o22ai_1_220/Y sky130_fd_sc_hd__nand2_1_372/B sky130_fd_sc_hd__o21ai_1_282/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_231 sky130_fd_sc_hd__nand2_1_360/Y sky130_fd_sc_hd__nand2_1_359/Y
+ sky130_fd_sc_hd__o22ai_1_231/Y sky130_fd_sc_hd__nand2_1_371/B sky130_fd_sc_hd__o21ai_1_281/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_242 sky130_fd_sc_hd__o22ai_1_261/A2 sky130_fd_sc_hd__nor2_1_144/B
+ sky130_fd_sc_hd__o22ai_1_242/Y sky130_fd_sc_hd__nor2_1_145/B sky130_fd_sc_hd__o32ai_1_2/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_306 sky130_fd_sc_hd__nand2_1_306/Y sky130_fd_sc_hd__nor2_1_100/B
+ sky130_fd_sc_hd__fa_2_1117/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_905 sky130_fd_sc_hd__clkinv_1_905/Y sky130_fd_sc_hd__nor2_1_214/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_905/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_253 sky130_fd_sc_hd__o22ai_1_261/A2 sky130_fd_sc_hd__o21a_1_29/A2
+ sky130_fd_sc_hd__o22ai_1_253/Y sky130_fd_sc_hd__nor2_1_153/B sky130_fd_sc_hd__o32ai_1_2/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_317 sky130_fd_sc_hd__nand2_1_317/Y sky130_fd_sc_hd__xor2_1_87/A
+ sky130_fd_sc_hd__nand2_2_6/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_916 sky130_fd_sc_hd__o22ai_1_309/B1 sky130_fd_sc_hd__fa_2_1185/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_916/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_264 sky130_fd_sc_hd__o32ai_1_2/A3 sky130_fd_sc_hd__nor2_1_154/B
+ sky130_fd_sc_hd__o22ai_1_264/Y sky130_fd_sc_hd__o22ai_1_264/A1 sky130_fd_sc_hd__o21a_1_29/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_328 sky130_fd_sc_hd__nand2_1_328/Y sky130_fd_sc_hd__nand2_1_333/B
+ sky130_fd_sc_hd__o21ai_1_237/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_275 sky130_fd_sc_hd__nand2_1_410/Y sky130_fd_sc_hd__nand2_1_409/Y
+ sky130_fd_sc_hd__o22ai_1_275/Y sky130_fd_sc_hd__nand2_1_423/B sky130_fd_sc_hd__o21ai_1_335/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_927 sky130_fd_sc_hd__nor2_1_199/B sky130_fd_sc_hd__fa_2_1194/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_927/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__bufinv_8_1 sky130_fd_sc_hd__bufinv_8_1/A sky130_fd_sc_hd__bufinv_8_1/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufinv_8
Xsky130_fd_sc_hd__nand2_1_339 sky130_fd_sc_hd__nor2_2_13/B sky130_fd_sc_hd__nand2_1_339/B
+ sky130_fd_sc_hd__nand2_1_339/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_286 sky130_fd_sc_hd__nand2_1_412/Y sky130_fd_sc_hd__nand2_1_411/Y
+ sky130_fd_sc_hd__o22ai_1_286/Y sky130_fd_sc_hd__nand2_1_422/B sky130_fd_sc_hd__o21ai_1_334/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_938 sky130_fd_sc_hd__o22ai_1_322/B1 sky130_fd_sc_hd__fa_2_1203/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_938/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_297 sky130_fd_sc_hd__o32ai_1_3/B2 sky130_fd_sc_hd__nor2_1_224/A
+ sky130_fd_sc_hd__o22ai_1_297/Y sky130_fd_sc_hd__o22ai_1_319/A1 sky130_fd_sc_hd__a222oi_1_15/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_949 sky130_fd_sc_hd__or2_0_11/B sky130_fd_sc_hd__nor2_1_268/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_949/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_102 VDD VSS sky130_fd_sc_hd__ha_2_2/A sky130_fd_sc_hd__dfxtp_1_95/CLK
+ sky130_fd_sc_hd__and2_0_7/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_113 VDD VSS sky130_fd_sc_hd__nor2_1_22/A sky130_fd_sc_hd__dfxtp_1_117/CLK
+ sky130_fd_sc_hd__ha_2_3/SUM VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_124 VDD VSS sky130_fd_sc_hd__ha_2_16/A sky130_fd_sc_hd__dfxtp_1_129/CLK
+ sky130_fd_sc_hd__and2_0_15/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_135 VDD VSS sky130_fd_sc_hd__ha_2_27/A sky130_fd_sc_hd__dfxtp_1_138/CLK
+ sky130_fd_sc_hd__nor2b_1_6/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_146 VDD VSS sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__clkinv_4_2/Y
+ sky130_fd_sc_hd__xor2_1_2/B VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_157 VDD VSS sky130_fd_sc_hd__ha_2_30/A sky130_fd_sc_hd__dfxtp_1_158/CLK
+ sky130_fd_sc_hd__and2_0_25/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_168 VDD VSS sky130_fd_sc_hd__ha_2_41/A sky130_fd_sc_hd__dfxtp_1_170/CLK
+ sky130_fd_sc_hd__nor2b_1_22/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_179 VDD VSS sky130_fd_sc_hd__ha_2_55/A sky130_fd_sc_hd__dfxtp_1_182/CLK
+ sky130_fd_sc_hd__and2_0_53/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_480 VSS VDD sky130_fd_sc_hd__a21oi_1_476/Y sky130_fd_sc_hd__nor2_1_309/A
+ sky130_fd_sc_hd__a21oi_1_467/Y sky130_fd_sc_hd__xor2_1_290/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_491 VSS VDD sky130_fd_sc_hd__o22ai_1_432/A2 sky130_fd_sc_hd__nor2_1_282/B
+ sky130_fd_sc_hd__a21oi_1_478/Y sky130_fd_sc_hd__o21ai_1_491/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_1201 sky130_fd_sc_hd__fa_2_1202/CIN sky130_fd_sc_hd__mux2_2_141/A1
+ sky130_fd_sc_hd__fa_2_1201/A sky130_fd_sc_hd__fa_2_1201/B sky130_fd_sc_hd__fa_2_1201/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1212 sky130_fd_sc_hd__fa_2_1213/CIN sky130_fd_sc_hd__mux2_2_168/A1
+ sky130_fd_sc_hd__fa_2_1212/A sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__fa_2_1212/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1223 sky130_fd_sc_hd__xor2_1_228/B sky130_fd_sc_hd__nand2_1_417/A
+ sky130_fd_sc_hd__fa_2_1223/A sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__fa_2_1223/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1234 sky130_fd_sc_hd__fa_2_1235/CIN sky130_fd_sc_hd__mux2_2_190/A1
+ sky130_fd_sc_hd__fa_2_1234/A sky130_fd_sc_hd__fa_2_1234/B sky130_fd_sc_hd__fa_2_1234/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1245 sky130_fd_sc_hd__fa_2_1246/CIN sky130_fd_sc_hd__mux2_2_209/A1
+ sky130_fd_sc_hd__fa_2_1245/A sky130_fd_sc_hd__fa_2_1245/B sky130_fd_sc_hd__fa_2_1245/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1256 sky130_fd_sc_hd__fa_2_1257/CIN sky130_fd_sc_hd__mux2_2_180/A0
+ sky130_fd_sc_hd__fa_2_1256/A sky130_fd_sc_hd__fa_2_1256/B sky130_fd_sc_hd__fa_2_1256/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1267 sky130_fd_sc_hd__fa_2_1268/CIN sky130_fd_sc_hd__mux2_2_208/A1
+ sky130_fd_sc_hd__fa_2_1267/A sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1267/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1020 VDD VSS sky130_fd_sc_hd__fa_2_849/A sky130_fd_sc_hd__dfxtp_1_1026/CLK
+ sky130_fd_sc_hd__a21oi_1_316/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_1278 sky130_fd_sc_hd__fa_2_1279/CIN sky130_fd_sc_hd__mux2_2_258/A1
+ sky130_fd_sc_hd__fa_2_1278/A sky130_fd_sc_hd__fa_2_1278/B sky130_fd_sc_hd__fa_2_1278/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1031 VDD VSS sky130_fd_sc_hd__fa_2_838/A sky130_fd_sc_hd__dfxtp_1_1038/CLK
+ sky130_fd_sc_hd__o21a_1_37/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_1289 sky130_fd_sc_hd__fa_2_1290/CIN sky130_fd_sc_hd__mux2_2_229/A0
+ sky130_fd_sc_hd__fa_2_1289/A sky130_fd_sc_hd__fa_2_1289/B sky130_fd_sc_hd__fa_2_1289/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o21ai_1_40 VSS VDD sky130_fd_sc_hd__o21ai_1_53/A2 sky130_fd_sc_hd__xnor2_1_34/Y
+ sky130_fd_sc_hd__a21oi_1_28/Y sky130_fd_sc_hd__o21ai_1_40/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1042 VDD VSS sky130_fd_sc_hd__fa_2_908/B sky130_fd_sc_hd__dfxtp_1_1047/CLK
+ sky130_fd_sc_hd__a21oi_1_304/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_51 VSS VDD sky130_fd_sc_hd__o21ai_1_53/A2 sky130_fd_sc_hd__xnor2_1_56/Y
+ sky130_fd_sc_hd__a21oi_1_39/Y sky130_fd_sc_hd__o21ai_1_51/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1053 VDD VSS sky130_fd_sc_hd__fa_2_1192/A sky130_fd_sc_hd__clkinv_4_23/Y
+ sky130_fd_sc_hd__and2_0_326/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_62 VSS VDD sky130_fd_sc_hd__nand2_2_3/Y sky130_fd_sc_hd__xnor2_1_44/Y
+ sky130_fd_sc_hd__a21oi_1_48/Y sky130_fd_sc_hd__o21ai_1_62/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1064 VDD VSS sky130_fd_sc_hd__fa_2_1203/A sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__mux2_2_136/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_73 VSS VDD sky130_fd_sc_hd__o21ai_1_73/A2 sky130_fd_sc_hd__o22ai_1_88/B1
+ sky130_fd_sc_hd__a21oi_1_58/Y sky130_fd_sc_hd__o21ai_1_73/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1075 VDD VSS sky130_fd_sc_hd__fa_2_1177/A sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__mux2_2_159/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_84 VSS VDD sky130_fd_sc_hd__xnor2_1_47/A sky130_fd_sc_hd__nor2_1_59/Y
+ sky130_fd_sc_hd__o21ai_1_84/B1 sky130_fd_sc_hd__xnor2_1_49/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1086 VDD VSS sky130_fd_sc_hd__fa_2_1188/A sky130_fd_sc_hd__clkinv_8_70/Y
+ sky130_fd_sc_hd__mux2_2_131/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_95 VSS VDD sky130_fd_sc_hd__a21oi_1_97/Y sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__o21ai_1_96/B1 sky130_fd_sc_hd__xor2_1_63/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1097 VDD VSS sky130_fd_sc_hd__fa_2_1216/A sky130_fd_sc_hd__clkinv_8_64/Y
+ sky130_fd_sc_hd__mux2_2_160/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_680 VDD VSS sky130_fd_sc_hd__fa_2_1019/A sky130_fd_sc_hd__clkinv_8_59/Y
+ sky130_fd_sc_hd__and2_0_272/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_691 VDD VSS sky130_fd_sc_hd__fa_2_1030/A sky130_fd_sc_hd__clkinv_4_26/Y
+ sky130_fd_sc_hd__mux2_2_30/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_530 sky130_fd_sc_hd__fa_2_533/B sky130_fd_sc_hd__fa_2_530/SUM
+ sky130_fd_sc_hd__fa_2_530/A sky130_fd_sc_hd__fa_2_530/B sky130_fd_sc_hd__fa_2_530/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o2bb2ai_1_15 sky130_fd_sc_hd__a21oi_1_14/B1 sky130_fd_sc_hd__nor4_1_4/C
+ sky130_fd_sc_hd__xor2_1_9/A sky130_fd_sc_hd__xor2_1_9/A sky130_fd_sc_hd__nor4_1_4/C
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__o2bb2ai_1_26 sky130_fd_sc_hd__and2_0_247/A sky130_fd_sc_hd__or4_1_2/C
+ sky130_fd_sc_hd__or4_1_2/D sky130_fd_sc_hd__or4_1_2/D sky130_fd_sc_hd__or4_1_2/C
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_541 sky130_fd_sc_hd__fa_2_543/CIN sky130_fd_sc_hd__fa_2_534/B
+ sky130_fd_sc_hd__ha_2_117/B sky130_fd_sc_hd__ha_2_119/B sky130_fd_sc_hd__fa_2_427/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_552 sky130_fd_sc_hd__maj3_1_83/B sky130_fd_sc_hd__maj3_1_84/A
+ sky130_fd_sc_hd__fa_2_552/A sky130_fd_sc_hd__fa_2_552/B sky130_fd_sc_hd__fa_2_553/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_563 sky130_fd_sc_hd__fa_2_562/A sky130_fd_sc_hd__fa_2_557/B
+ sky130_fd_sc_hd__ha_2_125/B sky130_fd_sc_hd__ha_2_125/A sky130_fd_sc_hd__fa_2_551/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_574 sky130_fd_sc_hd__fa_2_573/CIN sky130_fd_sc_hd__and2_0_92/A
+ sky130_fd_sc_hd__fa_2_574/A sky130_fd_sc_hd__fa_2_574/B sky130_fd_sc_hd__fa_2_574/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_585 sky130_fd_sc_hd__maj3_1_130/B sky130_fd_sc_hd__maj3_1_131/A
+ sky130_fd_sc_hd__ha_2_126/A sky130_fd_sc_hd__fa_2_585/B sky130_fd_sc_hd__ha_2_128/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_596 sky130_fd_sc_hd__fa_2_598/B sky130_fd_sc_hd__fa_2_596/SUM
+ sky130_fd_sc_hd__fa_2_692/A sky130_fd_sc_hd__fa_2_596/B sky130_fd_sc_hd__fa_2_596/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a21oi_1_109 sky130_fd_sc_hd__clkinv_1_564/Y sky130_fd_sc_hd__o21ai_1_130/Y
+ sky130_fd_sc_hd__a21oi_1_109/Y sky130_fd_sc_hd__a211o_1_3/A1 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nor2_1_306 sky130_fd_sc_hd__nor2_1_306/B sky130_fd_sc_hd__nor2_1_306/Y
+ sky130_fd_sc_hd__nor2_1_309/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_317 sky130_fd_sc_hd__nor2_1_322/B sky130_fd_sc_hd__nor2_1_317/Y
+ sky130_fd_sc_hd__nor2_1_318/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_502 sky130_fd_sc_hd__buf_12_502/A sky130_fd_sc_hd__buf_12_502/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_513 sky130_fd_sc_hd__buf_12_513/A sky130_fd_sc_hd__buf_12_513/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_405 sky130_fd_sc_hd__nor2_1_315/Y sky130_fd_sc_hd__nor2_1_313/Y
+ sky130_fd_sc_hd__nand3_1_10/Y sky130_fd_sc_hd__nand3_1_11/Y sky130_fd_sc_hd__nand3_1_52/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkbuf_8_5 sky130_fd_sc_hd__buf_2_156/A sky130_fd_sc_hd__dfxtp_1_84/D
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkbuf_8
Xsky130_fd_sc_hd__nand2_1_103 sky130_fd_sc_hd__nand2_1_103/Y sky130_fd_sc_hd__buf_2_268/X
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_702 sky130_fd_sc_hd__o21ai_1_227/A1 sky130_fd_sc_hd__o21ai_1_236/Y
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_114 sky130_fd_sc_hd__o21ai_1_31/B1 sky130_fd_sc_hd__ha_2_157/SUM
+ sky130_fd_sc_hd__nor2_1_18/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_713 sky130_fd_sc_hd__o22ai_1_190/A1 sky130_fd_sc_hd__fa_2_1060/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_713/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_125 sky130_fd_sc_hd__nand2_1_125/Y sky130_fd_sc_hd__nand2_1_126/Y
+ sky130_fd_sc_hd__buf_2_264/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_724 sky130_fd_sc_hd__o22ai_1_195/B2 sky130_fd_sc_hd__fa_2_1050/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_724/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_136 sky130_fd_sc_hd__nand2_1_136/Y sky130_fd_sc_hd__fa_2_711/SUM
+ sky130_fd_sc_hd__and2_0_235/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_735 sky130_fd_sc_hd__nand2_1_333/A sky130_fd_sc_hd__a211oi_1_9/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_735/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_147 sky130_fd_sc_hd__nor2_1_17/B sky130_fd_sc_hd__nor3_1_26/C
+ sky130_fd_sc_hd__nor3_1_27/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_746 sky130_fd_sc_hd__nand2_2_6/B sky130_fd_sc_hd__nand2_1_339/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_746/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_158 sky130_fd_sc_hd__fa_2_176/B sky130_fd_sc_hd__fa_2_250/A
+ sky130_fd_sc_hd__fa_2_283/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_757 sky130_fd_sc_hd__ha_2_189/B sky130_fd_sc_hd__fa_2_1118/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_757/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_169 sky130_fd_sc_hd__fa_2_332/CIN sky130_fd_sc_hd__fa_2_413/A
+ sky130_fd_sc_hd__fa_2_409/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_768 sky130_fd_sc_hd__ha_2_200/A sky130_fd_sc_hd__ha_2_201/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_768/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_779 sky130_fd_sc_hd__clkinv_1_779/Y sky130_fd_sc_hd__o21a_1_29/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_779/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor2_1_7 sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__xor2_1_7/X
+ sky130_fd_sc_hd__xor2_1_7/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand3_2_8 sky130_fd_sc_hd__or2_1_1/X sky130_fd_sc_hd__nand3_2_8/Y
+ sky130_fd_sc_hd__nand3_2_8/B sky130_fd_sc_hd__nand3_2_8/C VSS VDD VSS VDD sky130_fd_sc_hd__nand3_2
Xsky130_fd_sc_hd__clkinv_8_5 sky130_fd_sc_hd__clkinv_8_5/Y sky130_fd_sc_hd__clkinv_8_5/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_5/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__nor3_1_13 sky130_fd_sc_hd__nor3_1_13/C sky130_fd_sc_hd__nor3_1_13/Y
+ sky130_fd_sc_hd__nor3_2_4/A sky130_fd_sc_hd__nor3_1_9/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_24 sky130_fd_sc_hd__nor3_1_24/C sky130_fd_sc_hd__nor3_1_24/Y
+ sky130_fd_sc_hd__nor2_2_5/A sky130_fd_sc_hd__nor3_2_10/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_35 sky130_fd_sc_hd__nor3_1_35/C sky130_fd_sc_hd__nor3_1_35/Y
+ sky130_fd_sc_hd__nor3_1_35/A sky130_fd_sc_hd__fa_2_954/A VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__fa_2_1020 sky130_fd_sc_hd__fa_2_1021/CIN sky130_fd_sc_hd__and2_0_273/A
+ sky130_fd_sc_hd__fa_2_1020/A sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_1020/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1031 sky130_fd_sc_hd__fa_2_1032/CIN sky130_fd_sc_hd__fa_2_1031/SUM
+ sky130_fd_sc_hd__fa_2_1031/A sky130_fd_sc_hd__nor2_1_55/A sky130_fd_sc_hd__ha_2_185/COUT
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1042 sky130_fd_sc_hd__fa_2_1043/CIN sky130_fd_sc_hd__fa_2_1042/SUM
+ sky130_fd_sc_hd__nor2_1_61/A sky130_fd_sc_hd__fa_2_1042/B sky130_fd_sc_hd__fa_2_1042/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1053 sky130_fd_sc_hd__fa_2_1054/CIN sky130_fd_sc_hd__mux2_2_73/A1
+ sky130_fd_sc_hd__fa_2_1053/A sky130_fd_sc_hd__fa_2_1053/B sky130_fd_sc_hd__fa_2_1053/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1064 sky130_fd_sc_hd__fa_2_1065/CIN sky130_fd_sc_hd__mux2_2_49/A0
+ sky130_fd_sc_hd__fa_2_1064/A sky130_fd_sc_hd__xor2_1_93/X sky130_fd_sc_hd__fa_2_1064/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1075 sky130_fd_sc_hd__fa_2_1076/CIN sky130_fd_sc_hd__mux2_2_74/A1
+ sky130_fd_sc_hd__fa_2_1075/A sky130_fd_sc_hd__fa_2_1075/B sky130_fd_sc_hd__fa_2_1075/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1086 sky130_fd_sc_hd__fa_2_1087/CIN sky130_fd_sc_hd__mux2_2_50/A0
+ sky130_fd_sc_hd__fa_2_1086/A sky130_fd_sc_hd__fa_2_1086/B sky130_fd_sc_hd__fa_2_1086/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1097 sky130_fd_sc_hd__fa_2_1098/CIN sky130_fd_sc_hd__and2_0_299/A
+ sky130_fd_sc_hd__fa_2_1097/A sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1097/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_40 sky130_fd_sc_hd__inv_2_40/A sky130_fd_sc_hd__inv_2_40/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_51 sky130_fd_sc_hd__ha_2_33/A sky130_fd_sc_hd__inv_2_51/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_62 sky130_fd_sc_hd__inv_2_62/A sky130_fd_sc_hd__inv_2_62/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_73 sky130_fd_sc_hd__inv_2_73/A sky130_fd_sc_hd__inv_2_73/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_84 sky130_fd_sc_hd__inv_2_84/A sky130_fd_sc_hd__inv_2_84/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_95 sky130_fd_sc_hd__inv_2_95/A sky130_fd_sc_hd__inv_2_95/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__o32ai_1_10 sky130_fd_sc_hd__o32ai_1_10/A2 sky130_fd_sc_hd__o32ai_1_10/Y
+ sky130_fd_sc_hd__fa_2_1295/A sky130_fd_sc_hd__o32ai_1_10/A3 sky130_fd_sc_hd__o32ai_1_10/B2
+ sky130_fd_sc_hd__fa_2_1294/A VDD VSS VSS VDD sky130_fd_sc_hd__o32ai_1
Xsky130_fd_sc_hd__ha_2_16 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_16/A sky130_fd_sc_hd__ha_2_15/B
+ sky130_fd_sc_hd__ha_2_16/SUM sky130_fd_sc_hd__ha_2_16/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_27 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_27/A sky130_fd_sc_hd__ha_2_26/B
+ sky130_fd_sc_hd__ha_2_27/SUM sky130_fd_sc_hd__ha_2_27/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_38 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_38/A sky130_fd_sc_hd__ha_2_37/B
+ sky130_fd_sc_hd__ha_2_38/SUM sky130_fd_sc_hd__ha_2_38/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_49 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_49/A sky130_fd_sc_hd__ha_2_48/B
+ sky130_fd_sc_hd__ha_2_49/SUM sky130_fd_sc_hd__ha_2_49/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_360 sky130_fd_sc_hd__fa_2_361/B sky130_fd_sc_hd__fa_2_353/A
+ sky130_fd_sc_hd__ha_2_115/A sky130_fd_sc_hd__fa_2_360/B sky130_fd_sc_hd__fa_2_412/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_371 sky130_fd_sc_hd__maj3_1_65/B sky130_fd_sc_hd__maj3_1_66/A
+ sky130_fd_sc_hd__fa_2_371/A sky130_fd_sc_hd__fa_2_371/B sky130_fd_sc_hd__fa_2_372/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_12 sky130_fd_sc_hd__conb_1_7/LO sky130_fd_sc_hd__clkinv_8_100/Y
+ sky130_fd_sc_hd__dfxtp_1_117/CLK sky130_fd_sc_hd__a21oi_1_0/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_382 sky130_fd_sc_hd__maj3_1_63/B sky130_fd_sc_hd__maj3_1_64/A
+ sky130_fd_sc_hd__fa_2_382/A sky130_fd_sc_hd__fa_2_382/B sky130_fd_sc_hd__fa_2_383/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_23 sky130_fd_sc_hd__conb_1_14/LO sky130_fd_sc_hd__clkinv_4_51/A
+ sky130_fd_sc_hd__dfxtp_1_212/CLK sky130_fd_sc_hd__nand3_1_36/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_393 sky130_fd_sc_hd__fa_2_390/B sky130_fd_sc_hd__fa_2_386/B
+ sky130_fd_sc_hd__fa_2_393/A sky130_fd_sc_hd__ha_2_115/B sky130_fd_sc_hd__fa_2_425/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22oi_2_4 sky130_fd_sc_hd__nor2_4_5/Y sky130_fd_sc_hd__a22oi_2_4/A2
+ sky130_fd_sc_hd__a22oi_2_9/B1 sky130_fd_sc_hd__a22oi_2_4/B2 sky130_fd_sc_hd__a22oi_2_4/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__sdlclkp_4_34 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_62/Y
+ sky130_fd_sc_hd__dfxtp_1_304/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__clkbuf_16_16 sky130_fd_sc_hd__buf_12_507/A sky130_fd_sc_hd__buf_6_63/X
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__diode_2_210 sig_frequency[7] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__sdlclkp_4_45 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_68/Y
+ sky130_fd_sc_hd__dfxtp_1_424/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__diode_2_221 sig_amplitude[3] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__sdlclkp_4_56 sky130_fd_sc_hd__conb_1_20/LO sky130_fd_sc_hd__clkinv_8_62/Y
+ sky130_fd_sc_hd__dfxtp_1_533/CLK sky130_fd_sc_hd__o21ai_1_32/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__diode_2_232 sig_frequency[1] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__sdlclkp_4_67 sky130_fd_sc_hd__conb_1_22/LO sky130_fd_sc_hd__clkinv_8_61/Y
+ sky130_fd_sc_hd__dfxtp_1_571/CLK sky130_fd_sc_hd__nor4_1_5/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_78 sky130_fd_sc_hd__conb_1_25/LO sky130_fd_sc_hd__clkinv_8_72/A
+ sky130_fd_sc_hd__dfxtp_1_902/CLK sky130_fd_sc_hd__or2_0_9/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_89 sky130_fd_sc_hd__conb_1_28/LO sky130_fd_sc_hd__clkinv_8_47/A
+ sky130_fd_sc_hd__dfxtp_1_1332/CLK sky130_fd_sc_hd__or2_0_12/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_103 sky130_fd_sc_hd__nor2_1_103/B sky130_fd_sc_hd__nor2_1_94/A
+ sky130_fd_sc_hd__fa_2_1111/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_114 sky130_fd_sc_hd__nor2_1_114/B sky130_fd_sc_hd__o21a_1_10/A1
+ sky130_fd_sc_hd__o21a_1_11/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_125 sky130_fd_sc_hd__nor2_1_132/Y sky130_fd_sc_hd__nor2_1_125/Y
+ sky130_fd_sc_hd__nor2_1_126/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_12 sky130_fd_sc_hd__nor2_2_0/Y sky130_fd_sc_hd__clkinv_1_4/Y
+ sky130_fd_sc_hd__nand4_1_25/Y sky130_fd_sc_hd__nand4_1_9/Y sky130_fd_sc_hd__a22oi_1_12/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_136 sky130_fd_sc_hd__o21a_1_16/A2 sky130_fd_sc_hd__nor2_1_136/Y
+ sky130_fd_sc_hd__nor2_1_136/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_23 sky130_fd_sc_hd__nor2_2_0/Y sky130_fd_sc_hd__clkinv_1_4/Y
+ sky130_fd_sc_hd__nand4_1_19/Y sky130_fd_sc_hd__nand4_1_3/Y sky130_fd_sc_hd__a22oi_1_23/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_147 sky130_fd_sc_hd__nor2_1_147/B sky130_fd_sc_hd__nor2_1_147/Y
+ sky130_fd_sc_hd__o21a_1_22/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_34 sky130_fd_sc_hd__a22oi_2_9/B1 sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__clkbuf_4_40/X sky130_fd_sc_hd__a22oi_1_34/A2 sky130_fd_sc_hd__a22oi_1_34/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_158 sky130_fd_sc_hd__nor2_1_158/B sky130_fd_sc_hd__nor2_1_158/Y
+ sky130_fd_sc_hd__nor2_2_14/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_45 sky130_fd_sc_hd__nor2_2_2/Y sky130_fd_sc_hd__a22oi_1_82/A1
+ sky130_fd_sc_hd__clkbuf_1_66/X sky130_fd_sc_hd__a22oi_1_45/A2 sky130_fd_sc_hd__nand4_1_4/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_169 sky130_fd_sc_hd__a21o_2_9/A2 sky130_fd_sc_hd__a21o_2_9/B1
+ sky130_fd_sc_hd__a21o_2_9/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_56 sky130_fd_sc_hd__a22oi_1_81/B1 sky130_fd_sc_hd__clkbuf_1_99/X
+ sky130_fd_sc_hd__clkbuf_1_42/X sky130_fd_sc_hd__clkbuf_4_17/X sky130_fd_sc_hd__nand4_1_8/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_67 sky130_fd_sc_hd__a22oi_2_9/B1 sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__clkbuf_4_30/X sky130_fd_sc_hd__a22oi_1_67/A2 sky130_fd_sc_hd__a22oi_1_67/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_78 sky130_fd_sc_hd__nor2_2_2/Y sky130_fd_sc_hd__a22oi_1_82/A1
+ sky130_fd_sc_hd__clkbuf_1_56/X sky130_fd_sc_hd__clkbuf_1_52/X sky130_fd_sc_hd__nand4_1_14/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_89 sky130_fd_sc_hd__a22oi_1_97/B1 sky130_fd_sc_hd__a22oi_1_97/A1
+ sky130_fd_sc_hd__buf_2_64/X sky130_fd_sc_hd__clkbuf_4_88/X sky130_fd_sc_hd__nand4_1_17/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_310 sky130_fd_sc_hd__inv_16_6/Y sky130_fd_sc_hd__buf_12_310/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_321 sky130_fd_sc_hd__buf_4_73/X sky130_fd_sc_hd__buf_12_321/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_332 sky130_fd_sc_hd__buf_4_86/X sky130_fd_sc_hd__buf_12_354/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_343 sky130_fd_sc_hd__buf_6_37/X sky130_fd_sc_hd__buf_12_343/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_202 sky130_fd_sc_hd__clkbuf_1_264/X sky130_fd_sc_hd__nor2_2_3/Y
+ sky130_fd_sc_hd__a22oi_1_202/B2 sky130_fd_sc_hd__clkbuf_4_124/X sky130_fd_sc_hd__nand4_1_45/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_354 sky130_fd_sc_hd__buf_12_354/A sky130_fd_sc_hd__buf_12_354/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_213 sky130_fd_sc_hd__buf_2_164/X sky130_fd_sc_hd__nor2_4_8/Y
+ sky130_fd_sc_hd__clkbuf_1_426/X sky130_fd_sc_hd__buf_2_235/X sky130_fd_sc_hd__nand4_1_48/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_365 sky130_fd_sc_hd__buf_12_365/A sky130_fd_sc_hd__buf_12_365/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_224 sky130_fd_sc_hd__nor3_2_8/Y sky130_fd_sc_hd__nor3_2_7/Y
+ sky130_fd_sc_hd__clkbuf_1_392/X sky130_fd_sc_hd__a22oi_1_224/A2 sky130_fd_sc_hd__a22oi_1_224/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_376 sky130_fd_sc_hd__buf_2_274/X sky130_fd_sc_hd__buf_2_140/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_235 sky130_fd_sc_hd__buf_2_164/X sky130_fd_sc_hd__nor2_4_8/Y
+ sky130_fd_sc_hd__clkbuf_1_420/X sky130_fd_sc_hd__buf_2_229/X sky130_fd_sc_hd__nand4_1_56/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_387 sky130_fd_sc_hd__inv_2_125/Y sky130_fd_sc_hd__buf_12_489/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_246 sky130_fd_sc_hd__buf_2_164/X sky130_fd_sc_hd__nor2_4_8/Y
+ sky130_fd_sc_hd__clkbuf_1_416/X sky130_fd_sc_hd__buf_2_225/X sky130_fd_sc_hd__nand4_1_60/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_398 sky130_fd_sc_hd__buf_12_398/A sky130_fd_sc_hd__buf_12_497/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_257 sky130_fd_sc_hd__clkbuf_4_165/X sky130_fd_sc_hd__clkinv_2_23/Y
+ sky130_fd_sc_hd__clkbuf_1_413/X sky130_fd_sc_hd__a22oi_1_257/A2 sky130_fd_sc_hd__a22oi_1_257/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_268 sky130_fd_sc_hd__clkbuf_1_376/X sky130_fd_sc_hd__nor2_2_5/Y
+ sky130_fd_sc_hd__buf_2_215/X sky130_fd_sc_hd__clkbuf_1_471/X sky130_fd_sc_hd__nand4_1_66/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_510 sky130_fd_sc_hd__a21oi_1_60/A1 sky130_fd_sc_hd__nor2_1_50/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_510/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22oi_1_279 sky130_fd_sc_hd__nor2_2_4/Y sky130_fd_sc_hd__clkbuf_1_377/X
+ sky130_fd_sc_hd__a22oi_1_279/B2 sky130_fd_sc_hd__clkbuf_4_187/X sky130_fd_sc_hd__nand4_1_69/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_521 sky130_fd_sc_hd__nor2_1_59/B sky130_fd_sc_hd__fa_2_1038/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_521/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_532 sky130_fd_sc_hd__o21ai_1_92/A2 sky130_fd_sc_hd__fa_2_1002/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_532/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_4_108 VDD VSS sky130_fd_sc_hd__buf_6_63/A sky130_fd_sc_hd__buf_6_79/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__clkinv_1_543 sky130_fd_sc_hd__o21ai_1_111/A2 sky130_fd_sc_hd__a211o_1_5/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_543/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_4_119 VDD VSS sky130_fd_sc_hd__buf_4_119/X sky130_fd_sc_hd__buf_4_119/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__clkinv_1_554 sky130_fd_sc_hd__nand4_1_85/C sky130_fd_sc_hd__fa_2_971/A
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_565 sky130_fd_sc_hd__clkinv_1_565/Y sky130_fd_sc_hd__a21oi_1_132/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_565/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_576 sky130_fd_sc_hd__nor2_1_88/A sky130_fd_sc_hd__fa_2_1010/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_576/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_587 sky130_fd_sc_hd__nand2_2_4/A sky130_fd_sc_hd__o22ai_1_90/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_587/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_598 sky130_fd_sc_hd__ha_2_173/B sky130_fd_sc_hd__fa_2_1042/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_598/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_4_12 sky130_fd_sc_hd__clkinv_4_13/A sky130_fd_sc_hd__clkinv_4_12/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_12/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_23 sky130_fd_sc_hd__clkinv_8_49/A sky130_fd_sc_hd__clkinv_4_23/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_23/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_34 sky130_fd_sc_hd__buf_6_86/X sky130_fd_sc_hd__or2_0_0/B
+ VSS VDD VDD VSS VSS sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_90 sky130_fd_sc_hd__nor2_1_90/B sky130_fd_sc_hd__nor2_1_90/Y
+ sky130_fd_sc_hd__or2_0_5/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_45 sky130_fd_sc_hd__clkinv_4_45/A sky130_fd_sc_hd__clkinv_8_0/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_45/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_56 sky130_fd_sc_hd__clkinv_4_56/A sky130_fd_sc_hd__clkinv_4_56/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_56/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_67 sky130_fd_sc_hd__clkinv_4_67/A sky130_fd_sc_hd__clkinv_2_6/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_67/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_78 sky130_fd_sc_hd__clkinv_4_78/A sky130_fd_sc_hd__clkinv_4_78/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_78/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__a21oi_1_440 sky130_fd_sc_hd__nor2_2_18/Y sky130_fd_sc_hd__o21ai_1_447/Y
+ sky130_fd_sc_hd__nor2_1_291/B sky130_fd_sc_hd__fa_2_1298/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_451 sky130_fd_sc_hd__nand2_1_543/B sky130_fd_sc_hd__o22ai_1_415/Y
+ sky130_fd_sc_hd__a21oi_1_451/Y sky130_fd_sc_hd__o21ai_1_469/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_462 sky130_fd_sc_hd__nor2b_2_5/Y sky130_fd_sc_hd__o21ai_1_477/Y
+ sky130_fd_sc_hd__a21oi_1_462/Y sky130_fd_sc_hd__o21ai_1_490/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_473 sky130_fd_sc_hd__fa_2_1307/A sky130_fd_sc_hd__o22ai_1_428/Y
+ sky130_fd_sc_hd__a21oi_1_473/Y sky130_fd_sc_hd__nor3_1_41/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_484 sky130_fd_sc_hd__nor2_1_312/Y sky130_fd_sc_hd__nand3_1_52/Y
+ sky130_fd_sc_hd__a31oi_1_4/B1 sky130_fd_sc_hd__nand3_1_8/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_495 sky130_fd_sc_hd__or2_0_13/A sky130_fd_sc_hd__or2_0_0/B
+ sky130_fd_sc_hd__nand2_1_563/A sky130_fd_sc_hd__nor2_1_320/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_8_120 sky130_fd_sc_hd__clkinv_8_7/A sky130_fd_sc_hd__clkinv_8_120/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_131 sky130_fd_sc_hd__clkinv_8_13/A sky130_fd_sc_hd__clkinv_8_131/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__o21a_1_0 sky130_fd_sc_hd__o21a_1_0/X sky130_fd_sc_hd__nor2_1_2/Y
+ sky130_fd_sc_hd__buf_6_86/X sky130_fd_sc_hd__o21a_1_0/A2 VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__xor2_1_306 sky130_fd_sc_hd__nor2_4_20/Y sky130_fd_sc_hd__fa_2_1304/B
+ sky130_fd_sc_hd__xor2_1_306/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_317 sky130_fd_sc_hd__nor2_4_20/Y sky130_fd_sc_hd__xor2_1_317/X
+ sky130_fd_sc_hd__xor2_1_317/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nor2b_1_80 sky130_fd_sc_hd__xnor2_1_32/A sky130_fd_sc_hd__nor2b_1_80/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_91 sky130_fd_sc_hd__or2_0_6/X sky130_fd_sc_hd__nor2b_1_91/Y
+ sky130_fd_sc_hd__buf_2_262/X VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1080 sky130_fd_sc_hd__o22ai_1_421/B1 sky130_fd_sc_hd__fa_2_1291/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1080/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1091 sky130_fd_sc_hd__a21oi_1_464/A1 sky130_fd_sc_hd__a21boi_1_8/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1091/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_14 VDD VSS sky130_fd_sc_hd__ha_2_110/A sky130_fd_sc_hd__dfxtp_1_26/CLK
+ sky130_fd_sc_hd__nand4_1_32/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_25 VDD VSS sky130_fd_sc_hd__ha_2_116/B sky130_fd_sc_hd__dfxtp_1_26/CLK
+ sky130_fd_sc_hd__buf_2_287/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_36 VDD VSS sky130_fd_sc_hd__fa_2_907/CIN sky130_fd_sc_hd__dfxtp_1_39/CLK
+ sky130_fd_sc_hd__nand4_1_38/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_190 sky130_fd_sc_hd__fa_2_192/A sky130_fd_sc_hd__fa_2_190/SUM
+ sky130_fd_sc_hd__fa_2_190/A sky130_fd_sc_hd__fa_2_190/B sky130_fd_sc_hd__fa_2_195/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_47 VDD VSS sky130_fd_sc_hd__ha_2_169/B sky130_fd_sc_hd__dfxtp_1_60/CLK
+ sky130_fd_sc_hd__dfxtp_1_63/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_58 VDD VSS sky130_fd_sc_hd__fa_2_546/A sky130_fd_sc_hd__dfxtp_1_61/CLK
+ sky130_fd_sc_hd__buf_2_286/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_69 VDD VSS sky130_fd_sc_hd__fa_2_87/A sky130_fd_sc_hd__dfxtp_1_77/CLK
+ sky130_fd_sc_hd__nand4_1_39/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_4_104 sky130_fd_sc_hd__clkbuf_4_104/X sky130_fd_sc_hd__buf_2_274/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_115 sky130_fd_sc_hd__clkbuf_4_115/X sky130_fd_sc_hd__clkbuf_4_115/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_126 sky130_fd_sc_hd__clkbuf_4_126/X sky130_fd_sc_hd__clkbuf_4_126/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_137 sky130_fd_sc_hd__clkbuf_4_137/X sky130_fd_sc_hd__clkbuf_4_137/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_308 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_308/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_308/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_148 sky130_fd_sc_hd__nand4_1_37/B sky130_fd_sc_hd__a22oi_1_169/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_319 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_319/X sky130_fd_sc_hd__mux2_2_99/S
+ sky130_fd_sc_hd__and2_0_319/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_159 sky130_fd_sc_hd__buf_12_290/A sky130_fd_sc_hd__buf_8_156/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_4_80 VDD VSS sky130_fd_sc_hd__buf_4_80/X sky130_fd_sc_hd__buf_4_80/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__inv_2_108 sky130_fd_sc_hd__inv_2_108/A sky130_fd_sc_hd__inv_2_108/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_4_91 VDD VSS sky130_fd_sc_hd__buf_4_91/X sky130_fd_sc_hd__buf_4_91/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__inv_2_119 sky130_fd_sc_hd__inv_2_119/A sky130_fd_sc_hd__inv_2_119/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_12_140 sky130_fd_sc_hd__inv_2_50/Y sky130_fd_sc_hd__buf_12_140/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_151 sky130_fd_sc_hd__buf_8_82/X sky130_fd_sc_hd__buf_12_263/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_162 sky130_fd_sc_hd__buf_8_94/X sky130_fd_sc_hd__buf_6_28/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_173 sky130_fd_sc_hd__buf_8_98/X sky130_fd_sc_hd__buf_12_173/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_184 sky130_fd_sc_hd__buf_8_110/X sky130_fd_sc_hd__buf_12_214/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_195 sky130_fd_sc_hd__buf_4_49/X sky130_fd_sc_hd__buf_12_195/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_340 sky130_fd_sc_hd__ha_2_129/B sky130_fd_sc_hd__ha_2_134/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_340/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_351 sky130_fd_sc_hd__ha_2_131/A sky130_fd_sc_hd__ha_2_133/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_351/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_362 sky130_fd_sc_hd__ha_2_142/B sky130_fd_sc_hd__fa_2_806/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_362/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_373 sky130_fd_sc_hd__fa_2_875/B sky130_fd_sc_hd__dfxtp_1_275/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_373/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_384 sky130_fd_sc_hd__fa_2_864/B sky130_fd_sc_hd__dfxtp_1_264/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_384/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_395 sky130_fd_sc_hd__o22ai_1_57/B2 sky130_fd_sc_hd__a21oi_1_14/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_395/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a211o_1_9 VSS VDD VSS VDD sky130_fd_sc_hd__a211o_1_9/X sky130_fd_sc_hd__a211o_1_9/A2
+ sky130_fd_sc_hd__nor2_1_122/Y sky130_fd_sc_hd__a211o_1_9/A1 sky130_fd_sc_hd__a211o_1_9/C1
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o21a_1_14 sky130_fd_sc_hd__o21a_1_14/X sky130_fd_sc_hd__o21a_1_14/A1
+ sky130_fd_sc_hd__o21a_1_14/B1 sky130_fd_sc_hd__fa_2_1055/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21ai_1_309 VSS VDD sky130_fd_sc_hd__a21oi_1_290/Y sky130_fd_sc_hd__nor2_1_182/A
+ sky130_fd_sc_hd__nand2_1_382/Y sky130_fd_sc_hd__xor2_1_144/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_25 sky130_fd_sc_hd__o21a_1_25/X sky130_fd_sc_hd__o21a_1_25/A1
+ sky130_fd_sc_hd__o21a_1_25/B1 sky130_fd_sc_hd__fa_2_1152/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_36 sky130_fd_sc_hd__o21a_1_36/X sky130_fd_sc_hd__o21a_1_36/A1
+ sky130_fd_sc_hd__xnor2_1_95/B sky130_fd_sc_hd__fa_2_1207/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_47 sky130_fd_sc_hd__o21a_1_47/X sky130_fd_sc_hd__o21a_1_47/A1
+ sky130_fd_sc_hd__o21a_1_47/B1 sky130_fd_sc_hd__fa_2_1232/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_58 sky130_fd_sc_hd__o21a_1_58/X sky130_fd_sc_hd__o21a_1_58/A1
+ sky130_fd_sc_hd__o21a_1_58/B1 sky130_fd_sc_hd__fa_2_1287/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__a21oi_1_270 sky130_fd_sc_hd__nor2_1_182/Y sky130_fd_sc_hd__nor2_1_173/Y
+ sky130_fd_sc_hd__a21oi_1_270/Y sky130_fd_sc_hd__fa_2_1130/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_281 sky130_fd_sc_hd__clkinv_1_838/Y sky130_fd_sc_hd__clkinv_1_836/Y
+ sky130_fd_sc_hd__a21oi_1_281/Y sky130_fd_sc_hd__nand2_1_387/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_292 sky130_fd_sc_hd__nor3_1_38/A sky130_fd_sc_hd__o22ai_1_256/Y
+ sky130_fd_sc_hd__a21oi_1_292/Y sky130_fd_sc_hd__fa_2_1155/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_200 sky130_fd_sc_hd__buf_8_200/A sky130_fd_sc_hd__buf_8_200/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_211 sky130_fd_sc_hd__buf_8_211/A sky130_fd_sc_hd__buf_8_211/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_222 sky130_fd_sc_hd__buf_8_222/A sky130_fd_sc_hd__buf_6_73/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xor2_1_103 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1054/B
+ sky130_fd_sc_hd__xor2_1_103/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_114 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__xor2_1_114/X
+ sky130_fd_sc_hd__xor2_1_87/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_125 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1081/B
+ sky130_fd_sc_hd__xor2_1_125/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_136 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1070/B
+ sky130_fd_sc_hd__xor2_1_136/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_147 sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__fa_2_1136/B
+ sky130_fd_sc_hd__xor2_1_147/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_158 sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__fa_2_1125/B
+ sky130_fd_sc_hd__xor2_1_158/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_509 VDD VSS sky130_fd_sc_hd__nor4_1_12/A sky130_fd_sc_hd__edfxtp_1_0/CLK
+ sky130_fd_sc_hd__a22o_1_62/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_169 sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__fa_2_1153/B
+ sky130_fd_sc_hd__xor2_1_169/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_107 VSS VDD sky130_fd_sc_hd__buf_8_32/A sky130_fd_sc_hd__clkbuf_1_122/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_118 VSS VDD sky130_fd_sc_hd__buf_8_41/A sky130_fd_sc_hd__clkbuf_1_118/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_129 VSS VDD sky130_fd_sc_hd__ha_2_14/A sky130_fd_sc_hd__dfxtp_1_126/Q
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_9 VDD VSS sky130_fd_sc_hd__dfxtp_1_9/Q sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__a22o_1_6/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand3_1_18 sky130_fd_sc_hd__nor2_4_3/A sky130_fd_sc_hd__nor4_1_0/A
+ sky130_fd_sc_hd__nor3_1_0/A sky130_fd_sc_hd__nor4_1_0/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_29 sky130_fd_sc_hd__nand3_1_29/Y sky130_fd_sc_hd__ha_2_40/A
+ sky130_fd_sc_hd__nand3_1_31/C sky130_fd_sc_hd__nand2_2_0/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__dfxtp_1_1405 VDD VSS sky130_fd_sc_hd__mux2_2_231/A1 sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__o22ai_1_384/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1416 VDD VSS sky130_fd_sc_hd__mux2_2_262/A0 sky130_fd_sc_hd__clkinv_8_63/Y
+ sky130_fd_sc_hd__dfxtp_1_431/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1427 VDD VSS sky130_fd_sc_hd__mux2_2_254/A0 sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__o22ai_1_406/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1438 VDD VSS sky130_fd_sc_hd__mux2_2_226/A1 sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__o22ai_1_395/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1449 VDD VSS sky130_fd_sc_hd__nand2_1_568/B sky130_fd_sc_hd__dfxtp_1_1458/CLK
+ sky130_fd_sc_hd__and2_0_352/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_105 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_105/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__xnor2_1_8/Y sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_13 sky130_fd_sc_hd__nor3_2_2/C sky130_fd_sc_hd__nor3_2_3/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_13/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_116 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_116/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__fa_2_865/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_24 sky130_fd_sc_hd__inv_2_13/A sky130_fd_sc_hd__buf_8_54/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_24/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_127 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_127/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_892/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_35 sky130_fd_sc_hd__inv_2_24/A sky130_fd_sc_hd__buf_2_16/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_35/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_138 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_138/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_842/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_46 sky130_fd_sc_hd__inv_2_35/A sky130_fd_sc_hd__inv_2_18/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_46/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_149 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_149/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_858/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_57 sky130_fd_sc_hd__buf_8_29/A sky130_fd_sc_hd__bufinv_8_0/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_57/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_0 sky130_fd_sc_hd__fa_2_6/CIN sky130_fd_sc_hd__fa_2_0/SUM sky130_fd_sc_hd__fa_2_0/A
+ sky130_fd_sc_hd__fa_2_0/B sky130_fd_sc_hd__fa_2_0/CIN VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_1_68 sky130_fd_sc_hd__nand3_1_31/B sky130_fd_sc_hd__ha_2_40/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_68/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_79 sky130_fd_sc_hd__buf_8_68/A sky130_fd_sc_hd__clkinv_2_4/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_79/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_904 sky130_fd_sc_hd__fa_2_898/A sky130_fd_sc_hd__fa_2_899/B
+ sky130_fd_sc_hd__fa_2_904/A sky130_fd_sc_hd__fa_2_904/B sky130_fd_sc_hd__fa_2_904/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_915 sky130_fd_sc_hd__xnor2_1_23/A sky130_fd_sc_hd__fa_2_888/B
+ sky130_fd_sc_hd__fa_2_915/A sky130_fd_sc_hd__fa_2_915/B sky130_fd_sc_hd__fa_2_915/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_926 sky130_fd_sc_hd__fa_2_925/CIN sky130_fd_sc_hd__fa_2_926/SUM
+ sky130_fd_sc_hd__fa_2_926/A sky130_fd_sc_hd__fa_2_926/B sky130_fd_sc_hd__fa_2_926/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_937 sky130_fd_sc_hd__fa_2_921/A sky130_fd_sc_hd__fa_2_922/B
+ sky130_fd_sc_hd__fa_2_937/A sky130_fd_sc_hd__fa_2_937/B sky130_fd_sc_hd__ha_2_123/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_948 sky130_fd_sc_hd__fa_2_947/CIN sky130_fd_sc_hd__fa_2_948/SUM
+ sky130_fd_sc_hd__fa_2_948/A sky130_fd_sc_hd__fa_2_948/B sky130_fd_sc_hd__fa_2_948/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_959 sky130_fd_sc_hd__fa_2_958/CIN sky130_fd_sc_hd__fa_2_959/SUM
+ sky130_fd_sc_hd__fa_2_959/A sky130_fd_sc_hd__fa_2_959/B sky130_fd_sc_hd__fa_2_959/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__mux2_2_204 VSS VDD sky130_fd_sc_hd__mux2_2_204/A1 sky130_fd_sc_hd__mux2_2_204/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_204/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_215 VSS VDD sky130_fd_sc_hd__mux2_2_215/A1 sky130_fd_sc_hd__mux2_2_215/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_215/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_226 VSS VDD sky130_fd_sc_hd__mux2_2_226/A1 sky130_fd_sc_hd__mux2_2_226/A0
+ sky130_fd_sc_hd__nor2_8_2/A sky130_fd_sc_hd__mux2_2_226/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_237 VSS VDD sky130_fd_sc_hd__mux2_2_237/A1 sky130_fd_sc_hd__mux2_2_237/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_237/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_248 VSS VDD sky130_fd_sc_hd__mux2_2_248/A1 sky130_fd_sc_hd__mux2_2_248/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_248/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_259 VSS VDD sky130_fd_sc_hd__mux2_2_259/A1 sky130_fd_sc_hd__mux2_2_259/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_259/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__clkinv_1_170 sky130_fd_sc_hd__buf_8_158/A sky130_fd_sc_hd__clkinv_1_170/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_170/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_2 sky130_fd_sc_hd__buf_8_2/A sky130_fd_sc_hd__buf_8_2/X VSS
+ VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__a22o_1_4 sig_frequency[5] sky130_fd_sc_hd__nor2_1_1/Y sky130_fd_sc_hd__a22o_1_4/X
+ sky130_fd_sc_hd__a22o_1_4/B2 sky130_fd_sc_hd__nor2_1_0/Y VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_181 sky130_fd_sc_hd__buf_8_153/A sky130_fd_sc_hd__bufinv_8_8/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_181/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_192 sky130_fd_sc_hd__nor3_1_25/C sky130_fd_sc_hd__nor3_2_10/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_192/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_50 sky130_fd_sc_hd__a22o_1_50/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_50/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__fa_2_956/SUM
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_61 sky130_fd_sc_hd__a22o_1_61/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_61/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__nor4_1_11/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_72 sky130_fd_sc_hd__nor2_2_10/Y sky130_fd_sc_hd__a22o_1_72/A2
+ sky130_fd_sc_hd__a22o_1_72/X sky130_fd_sc_hd__a22o_1_72/B2 sky130_fd_sc_hd__nor2_2_11/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__nand4_1_0 sky130_fd_sc_hd__nand4_1_0/C sky130_fd_sc_hd__nand4_1_0/B
+ sky130_fd_sc_hd__nand4_1_0/Y sky130_fd_sc_hd__nand4_1_0/D sky130_fd_sc_hd__nand4_1_0/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__o21ai_1_106 VSS VDD sky130_fd_sc_hd__a21oi_1_90/Y sky130_fd_sc_hd__nor2_1_76/A
+ sky130_fd_sc_hd__nand2_1_264/Y sky130_fd_sc_hd__o21ai_1_106/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_117 VSS VDD sky130_fd_sc_hd__o22ai_1_130/B1 sky130_fd_sc_hd__nand4_1_85/B
+ sky130_fd_sc_hd__a21oi_1_102/Y sky130_fd_sc_hd__o21ai_1_117/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_128 VSS VDD sky130_fd_sc_hd__o22ai_1_92/A1 sky130_fd_sc_hd__nor2_1_77/A
+ sky130_fd_sc_hd__nand2b_1_13/Y sky130_fd_sc_hd__o21ai_1_128/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_139 VSS VDD sky130_fd_sc_hd__o21ai_1_153/A2 sky130_fd_sc_hd__o21a_1_8/A2
+ sky130_fd_sc_hd__a21oi_1_115/Y sky130_fd_sc_hd__a211o_1_4/A2 VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__maj3_1_12 sky130_fd_sc_hd__maj3_1_13/X sky130_fd_sc_hd__maj3_1_12/X
+ sky130_fd_sc_hd__maj3_1_12/B sky130_fd_sc_hd__maj3_1_12/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_23 sky130_fd_sc_hd__maj3_1_24/X sky130_fd_sc_hd__maj3_1_23/X
+ sky130_fd_sc_hd__maj3_1_23/B sky130_fd_sc_hd__maj3_1_23/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_402 sky130_fd_sc_hd__nand2_1_516/Y sky130_fd_sc_hd__nand2_1_515/Y
+ sky130_fd_sc_hd__o22ai_1_402/Y sky130_fd_sc_hd__nand2_1_527/B sky130_fd_sc_hd__o21ai_1_443/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_34 sky130_fd_sc_hd__maj3_1_35/X sky130_fd_sc_hd__maj3_1_34/X
+ sky130_fd_sc_hd__maj3_1_34/B sky130_fd_sc_hd__maj3_1_34/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_413 sky130_fd_sc_hd__o22ai_1_432/A2 sky130_fd_sc_hd__nor2_1_271/B
+ sky130_fd_sc_hd__o22ai_1_413/Y sky130_fd_sc_hd__nor2_1_272/B sky130_fd_sc_hd__o32ai_1_11/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_45 sky130_fd_sc_hd__maj3_1_46/X sky130_fd_sc_hd__maj3_1_45/X
+ sky130_fd_sc_hd__maj3_1_45/B sky130_fd_sc_hd__maj3_1_45/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_424 sky130_fd_sc_hd__o22ai_1_432/A2 sky130_fd_sc_hd__o21a_1_68/A2
+ sky130_fd_sc_hd__o22ai_1_424/Y sky130_fd_sc_hd__nor2_1_280/B sky130_fd_sc_hd__o32ai_1_11/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_56 sky130_fd_sc_hd__maj3_1_57/X sky130_fd_sc_hd__maj3_1_56/X
+ sky130_fd_sc_hd__maj3_1_56/B sky130_fd_sc_hd__maj3_1_56/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_435 sky130_fd_sc_hd__o32ai_1_11/A3 sky130_fd_sc_hd__nor2_1_281/B
+ sky130_fd_sc_hd__o22ai_1_435/Y sky130_fd_sc_hd__o22ai_1_435/A1 sky130_fd_sc_hd__o21a_1_68/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_67 sky130_fd_sc_hd__maj3_1_68/X sky130_fd_sc_hd__maj3_1_67/X
+ sky130_fd_sc_hd__maj3_1_67/B sky130_fd_sc_hd__maj3_1_67/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_78 sky130_fd_sc_hd__maj3_1_79/X sky130_fd_sc_hd__maj3_1_78/X
+ sky130_fd_sc_hd__maj3_1_78/B sky130_fd_sc_hd__maj3_1_78/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_89 sky130_fd_sc_hd__maj3_1_90/X sky130_fd_sc_hd__maj3_1_89/X
+ sky130_fd_sc_hd__maj3_1_89/B sky130_fd_sc_hd__maj3_1_89/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_40 sky130_fd_sc_hd__nand2_1_40/Y sky130_fd_sc_hd__nand2_1_40/B
+ sky130_fd_sc_hd__a21oi_2_0/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_51 sky130_fd_sc_hd__nand2_1_51/Y sky130_fd_sc_hd__nand2_1_0/B
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_62 sky130_fd_sc_hd__nand2_1_62/Y sky130_fd_sc_hd__nand2_1_63/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_73 sky130_fd_sc_hd__nand2_1_73/Y sky130_fd_sc_hd__nand4_1_68/Y
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_84 sky130_fd_sc_hd__nand2_1_84/Y sky130_fd_sc_hd__nand2_1_85/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_95 sky130_fd_sc_hd__nand2_1_95/Y sky130_fd_sc_hd__nand2_1_95/B
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_306 VDD VSS sky130_fd_sc_hd__a22o_1_43/A1 sky130_fd_sc_hd__dfxtp_1_313/CLK
+ sky130_fd_sc_hd__and2_0_92/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_317 VDD VSS sky130_fd_sc_hd__nor4_1_2/B sky130_fd_sc_hd__dfxtp_1_325/CLK
+ sky130_fd_sc_hd__and2_0_199/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_328 VDD VSS sky130_fd_sc_hd__a22o_2_7/B2 sky130_fd_sc_hd__clkinv_4_27/Y
+ sky130_fd_sc_hd__o21ai_1_20/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_339 VDD VSS sky130_fd_sc_hd__ha_2_157/B sky130_fd_sc_hd__dfxtp_1_347/CLK
+ sky130_fd_sc_hd__dfxtp_1_339/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_14 sky130_fd_sc_hd__fa_2_7/B sky130_fd_sc_hd__fa_2_6/B sky130_fd_sc_hd__fa_2_2/A
+ sky130_fd_sc_hd__ha_2_96/B sky130_fd_sc_hd__fa_2_14/CIN VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_25 sky130_fd_sc_hd__fa_2_19/A sky130_fd_sc_hd__fa_2_22/B sky130_fd_sc_hd__fa_2_25/A
+ sky130_fd_sc_hd__fa_2_25/B sky130_fd_sc_hd__fa_2_25/CIN VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_36 sky130_fd_sc_hd__maj3_1_24/B sky130_fd_sc_hd__maj3_1_25/A
+ sky130_fd_sc_hd__fa_2_36/A sky130_fd_sc_hd__fa_2_36/B sky130_fd_sc_hd__o22ai_1_3/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_47 sky130_fd_sc_hd__maj3_1_20/B sky130_fd_sc_hd__maj3_1_21/A
+ sky130_fd_sc_hd__fa_2_47/A sky130_fd_sc_hd__fa_2_47/B sky130_fd_sc_hd__fa_2_48/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_58 sky130_fd_sc_hd__fa_2_56/B sky130_fd_sc_hd__fa_2_51/A sky130_fd_sc_hd__fa_2_2/A
+ sky130_fd_sc_hd__ha_2_93/A sky130_fd_sc_hd__fa_2_45/A VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_69 sky130_fd_sc_hd__maj3_1_15/B sky130_fd_sc_hd__maj3_1_16/A
+ sky130_fd_sc_hd__fa_2_69/A sky130_fd_sc_hd__fa_2_69/B sky130_fd_sc_hd__fa_2_70/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_206 VDD VSS sky130_fd_sc_hd__buf_2_206/X sky130_fd_sc_hd__buf_2_206/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_217 VDD VSS sky130_fd_sc_hd__buf_2_217/X sky130_fd_sc_hd__buf_2_217/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_228 VDD VSS sky130_fd_sc_hd__buf_2_228/X sky130_fd_sc_hd__buf_2_228/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_239 VDD VSS sky130_fd_sc_hd__buf_8_187/A sky130_fd_sc_hd__buf_8_203/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_sram_2kbyte_1rw1r_32x512_8_10 sky130_fd_sc_hd__clkbuf_4_102/X sky130_fd_sc_hd__clkbuf_4_103/X
+ sky130_fd_sc_hd__clkbuf_4_104/X sky130_fd_sc_hd__clkbuf_4_105/X sky130_fd_sc_hd__inv_8_0/Y
+ sky130_fd_sc_hd__buf_6_88/X sky130_fd_sc_hd__buf_2_285/X sky130_fd_sc_hd__buf_6_89/X
+ sky130_fd_sc_hd__clkbuf_4_227/X sky130_fd_sc_hd__buf_6_84/X sky130_fd_sc_hd__buf_4_122/X
+ sky130_fd_sc_hd__buf_4_121/X sky130_fd_sc_hd__buf_6_85/X sky130_fd_sc_hd__nand2_1_566/B
+ sky130_fd_sc_hd__nand2_1_567/B sky130_fd_sc_hd__clkbuf_4_109/X sky130_fd_sc_hd__clkbuf_4_102/X
+ sky130_fd_sc_hd__clkbuf_4_103/X sky130_fd_sc_hd__clkbuf_4_104/X sky130_fd_sc_hd__clkbuf_4_105/X
+ sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__buf_6_88/X sky130_fd_sc_hd__buf_2_285/X
+ sky130_fd_sc_hd__buf_6_89/X sky130_fd_sc_hd__clkbuf_4_227/X sky130_fd_sc_hd__buf_6_84/X
+ sky130_fd_sc_hd__buf_4_122/X sky130_fd_sc_hd__buf_4_121/X sky130_fd_sc_hd__buf_6_85/X
+ sky130_fd_sc_hd__nand2_1_566/B sky130_fd_sc_hd__nand2_1_567/B sky130_fd_sc_hd__clkbuf_4_109/X
+ sky130_fd_sc_hd__buf_8_179/X sky130_fd_sc_hd__buf_12_363/X sky130_fd_sc_hd__buf_12_305/X
+ sky130_fd_sc_hd__buf_12_298/X sky130_fd_sc_hd__buf_12_287/X sky130_fd_sc_hd__buf_12_270/X
+ sky130_fd_sc_hd__buf_12_272/X sky130_fd_sc_hd__buf_12_319/X sky130_fd_sc_hd__buf_12_374/X
+ sky130_fd_sc_hd__buf_12_266/X sky130_fd_sc_hd__buf_12_303/X sky130_fd_sc_hd__buf_12_338/X
+ sky130_fd_sc_hd__buf_12_293/X sky130_fd_sc_hd__buf_12_294/X sky130_fd_sc_hd__buf_12_318/X
+ sky130_fd_sc_hd__buf_12_282/X sky130_fd_sc_hd__buf_12_350/X sky130_fd_sc_hd__buf_12_308/X
+ sky130_fd_sc_hd__buf_2_132/X sky130_fd_sc_hd__clkbuf_1_263/X sky130_fd_sc_hd__buf_2_132/X
+ sky130_fd_sc_hd__clkinv_8_140/Y sky130_fd_sc_hd__clkinv_8_16/Y sky130_fd_sc_hd__buf_8_175/X
+ sky130_fd_sc_hd__buf_8_173/X sky130_fd_sc_hd__buf_12_330/X sky130_fd_sc_hd__buf_8_176/X
+ sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[0] sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[1]
+ sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[2] sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[3]
+ sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[4] sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[5]
+ sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[6] sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[7]
+ sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[8] sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[9]
+ sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[10] sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[11]
+ sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[12] sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[13]
+ sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[14] sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[15]
+ sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[16] sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[17]
+ sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[18] sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[19]
+ sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[20] sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[21]
+ sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[22] sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[23]
+ sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[24] sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[25]
+ sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[26] sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[27]
+ sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[28] sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[29]
+ sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[30] sky130_sram_2kbyte_1rw1r_32x512_8_10/dout0[31]
+ sky130_fd_sc_hd__a22oi_1_208/A2 sky130_fd_sc_hd__a22oi_1_204/A2 sky130_fd_sc_hd__a22oi_1_200/A2
+ sky130_fd_sc_hd__a22oi_1_196/A2 sky130_fd_sc_hd__a22oi_1_192/A2 sky130_fd_sc_hd__a22oi_1_188/A2
+ sky130_fd_sc_hd__a22oi_1_184/A2 sky130_fd_sc_hd__a22oi_1_180/A2 sky130_fd_sc_hd__a22oi_1_176/A2
+ sky130_fd_sc_hd__a22oi_1_172/A2 sky130_fd_sc_hd__a22oi_1_168/A2 sky130_fd_sc_hd__a22oi_1_164/A2
+ sky130_fd_sc_hd__a22oi_1_160/A2 sky130_fd_sc_hd__a22oi_1_156/A2 sky130_fd_sc_hd__a22oi_1_152/A2
+ sky130_fd_sc_hd__a22oi_1_148/A2 sky130_fd_sc_hd__a22oi_1_210/B2 sky130_fd_sc_hd__a22oi_1_206/B2
+ sky130_fd_sc_hd__a22oi_1_202/B2 sky130_fd_sc_hd__a22oi_1_198/B2 sky130_fd_sc_hd__a22oi_1_194/B2
+ sky130_fd_sc_hd__a22oi_1_190/B2 sky130_fd_sc_hd__a22oi_1_186/B2 sky130_fd_sc_hd__a22oi_1_182/B2
+ sky130_fd_sc_hd__a22oi_1_178/B2 sky130_fd_sc_hd__a22oi_1_174/B2 sky130_fd_sc_hd__a22oi_1_170/B2
+ sky130_fd_sc_hd__a22oi_1_166/B2 sky130_fd_sc_hd__a22oi_1_162/B2 sky130_fd_sc_hd__a22oi_1_158/B2
+ sky130_fd_sc_hd__a22oi_1_154/B2 sky130_fd_sc_hd__a22oi_1_150/B2 VDD VSS sky130_sram_2kbyte_1rw1r_32x512_8
Xsky130_fd_sc_hd__dfxtp_1_1202 VDD VSS sky130_fd_sc_hd__fa_2_1251/A sky130_fd_sc_hd__clkinv_8_75/Y
+ sky130_fd_sc_hd__mux2_2_191/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1213 VDD VSS sky130_fd_sc_hd__fa_2_1225/A sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__and2_0_331/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1224 VDD VSS sky130_fd_sc_hd__fa_2_1236/A sky130_fd_sc_hd__clkinv_8_78/Y
+ sky130_fd_sc_hd__mux2_2_185/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1235 VDD VSS sky130_fd_sc_hd__fa_2_1264/A sky130_fd_sc_hd__clkinv_8_63/Y
+ sky130_fd_sc_hd__mux2_2_215/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1246 VDD VSS sky130_fd_sc_hd__nor2_8_1/B sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__mux2_2_188/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1257 VDD VSS sky130_fd_sc_hd__mux2_2_201/A0 sky130_fd_sc_hd__clkinv_8_78/Y
+ sky130_fd_sc_hd__o22ai_1_334/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1268 VDD VSS sky130_fd_sc_hd__mux2_2_175/A1 sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__o31ai_1_10/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_840 VDD VSS sky130_fd_sc_hd__mux2_2_75/A0 sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__a22o_1_71/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1279 VDD VSS sky130_fd_sc_hd__mux2_2_202/A0 sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__dfxtp_1_435/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_851 VDD VSS sky130_fd_sc_hd__mux2_2_51/A1 sky130_fd_sc_hd__clkinv_4_25/Y
+ sky130_fd_sc_hd__o21ai_1_168/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_862 VDD VSS sky130_fd_sc_hd__mux2_2_70/A0 sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__o21ai_1_176/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_873 VDD VSS sky130_fd_sc_hd__mux2_2_46/A1 sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__o21ai_1_187/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_884 VDD VSS sky130_fd_sc_hd__fa_2_858/A sky130_fd_sc_hd__dfxtp_1_904/CLK
+ sky130_fd_sc_hd__o21a_1_27/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_895 VDD VSS sky130_fd_sc_hd__fa_2_929/A sky130_fd_sc_hd__dfxtp_1_899/CLK
+ sky130_fd_sc_hd__dfxtp_1_895/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_460 VSS VDD sky130_fd_sc_hd__clkbuf_1_460/X sky130_fd_sc_hd__clkbuf_1_460/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__or3_1_5 sky130_fd_sc_hd__or3_1_5/A sky130_fd_sc_hd__or3_1_5/X sky130_fd_sc_hd__or3_1_5/B
+ sky130_fd_sc_hd__or3_1_5/C VDD VSS VDD VSS sky130_fd_sc_hd__or3_1
Xsky130_fd_sc_hd__clkbuf_1_471 VSS VDD sky130_fd_sc_hd__clkbuf_1_471/X sky130_fd_sc_hd__clkbuf_1_471/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_482 VSS VDD sky130_fd_sc_hd__buf_8_188/A sky130_fd_sc_hd__inv_2_113/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a21oi_1_19 sky130_fd_sc_hd__nor3_1_31/Y sky130_fd_sc_hd__dfxtp_1_576/Q
+ sky130_fd_sc_hd__nor2_1_27/B sky130_fd_sc_hd__or4_1_2/C VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkbuf_1_493 VSS VDD sky130_fd_sc_hd__a22oi_2_23/B2 sky130_fd_sc_hd__clkbuf_1_493/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_701 sky130_fd_sc_hd__fa_2_569/A sky130_fd_sc_hd__fa_2_570/B
+ sky130_fd_sc_hd__ha_2_135/A sky130_fd_sc_hd__fa_2_701/B sky130_fd_sc_hd__fa_2_698/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_712 sky130_fd_sc_hd__fa_2_711/CIN sky130_fd_sc_hd__fa_2_712/SUM
+ sky130_fd_sc_hd__fa_2_712/A sky130_fd_sc_hd__fa_2_712/B sky130_fd_sc_hd__fa_2_712/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_723 sky130_fd_sc_hd__fa_2_724/B sky130_fd_sc_hd__fa_2_723/SUM
+ sky130_fd_sc_hd__fa_2_817/B sky130_fd_sc_hd__ha_2_136/A sky130_fd_sc_hd__ha_2_142/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_734 sky130_fd_sc_hd__fa_2_736/CIN sky130_fd_sc_hd__fa_2_732/A
+ sky130_fd_sc_hd__ha_2_139/B sky130_fd_sc_hd__fa_2_823/B sky130_fd_sc_hd__fa_2_829/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_745 sky130_fd_sc_hd__fa_2_748/A sky130_fd_sc_hd__fa_2_745/SUM
+ sky130_fd_sc_hd__fa_2_745/A sky130_fd_sc_hd__fa_2_745/B sky130_fd_sc_hd__fa_2_751/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_756 sky130_fd_sc_hd__maj3_1_144/B sky130_fd_sc_hd__maj3_1_145/A
+ sky130_fd_sc_hd__fa_2_756/A sky130_fd_sc_hd__fa_2_756/B sky130_fd_sc_hd__fa_2_757/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_767 sky130_fd_sc_hd__maj3_1_141/B sky130_fd_sc_hd__maj3_1_142/A
+ sky130_fd_sc_hd__fa_2_767/A sky130_fd_sc_hd__fa_2_767/B sky130_fd_sc_hd__fa_2_768/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_778 sky130_fd_sc_hd__fa_2_780/B sky130_fd_sc_hd__fa_2_775/A
+ sky130_fd_sc_hd__fa_2_834/B sky130_fd_sc_hd__ha_2_142/B sky130_fd_sc_hd__ha_2_142/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_789 sky130_fd_sc_hd__fa_2_791/A sky130_fd_sc_hd__fa_2_786/A
+ sky130_fd_sc_hd__ha_2_145/B sky130_fd_sc_hd__ha_2_142/A sky130_fd_sc_hd__ha_2_142/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor2b_1_120 sky130_fd_sc_hd__or2_0_11/X sky130_fd_sc_hd__nor2b_1_120/Y
+ sky130_fd_sc_hd__buf_2_262/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_131 sky130_fd_sc_hd__and2_0_338/X sky130_fd_sc_hd__nor2b_1_131/Y
+ sky130_fd_sc_hd__buf_2_262/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_142 sky130_fd_sc_hd__or2_0_13/X sky130_fd_sc_hd__nor2b_1_142/Y
+ sky130_fd_sc_hd__nor2b_1_142/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__bufbuf_8_2 sky130_fd_sc_hd__buf_2_159/X sky130_fd_sc_hd__buf_6_65/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufbuf_8
Xsky130_fd_sc_hd__buf_6_15 VDD VSS sky130_fd_sc_hd__buf_6_15/X sky130_fd_sc_hd__buf_6_15/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_26 VDD VSS sky130_fd_sc_hd__buf_6_26/X sky130_fd_sc_hd__buf_6_26/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_37 VDD VSS sky130_fd_sc_hd__buf_6_37/X sky130_fd_sc_hd__buf_6_37/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_48 VDD VSS sky130_fd_sc_hd__buf_6_48/X sky130_fd_sc_hd__buf_6_48/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_59 VDD VSS sky130_fd_sc_hd__buf_6_59/X sky130_fd_sc_hd__buf_6_59/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_17 sky130_fd_sc_hd__buf_2_123/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_28 sky130_fd_sc_hd__buf_2_73/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_39 sky130_fd_sc_hd__buf_2_112/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__o22ai_1_210 sky130_fd_sc_hd__nand2_1_358/Y sky130_fd_sc_hd__o21ai_1_277/Y
+ sky130_fd_sc_hd__o22ai_1_210/Y sky130_fd_sc_hd__nand2_1_367/B sky130_fd_sc_hd__nand2_1_357/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_221 sky130_fd_sc_hd__nand2_1_358/Y sky130_fd_sc_hd__nand2_1_357/Y
+ sky130_fd_sc_hd__o22ai_1_221/Y sky130_fd_sc_hd__o22ai_1_234/A1 sky130_fd_sc_hd__a21o_2_11/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_232 sky130_fd_sc_hd__nand2_1_360/Y sky130_fd_sc_hd__nand2_1_359/Y
+ sky130_fd_sc_hd__o22ai_1_232/Y sky130_fd_sc_hd__o22ai_1_232/A1 sky130_fd_sc_hd__a21o_2_10/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_243 sky130_fd_sc_hd__o22ai_1_265/A2 sky130_fd_sc_hd__nor2_1_176/A
+ sky130_fd_sc_hd__o22ai_1_243/Y sky130_fd_sc_hd__o22ai_1_252/B1 sky130_fd_sc_hd__o32ai_1_2/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_307 sky130_fd_sc_hd__nand2_1_307/Y sky130_fd_sc_hd__nor2_1_99/B
+ sky130_fd_sc_hd__nor2_1_99/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_906 sky130_fd_sc_hd__o21ai_1_358/A2 sky130_fd_sc_hd__fa_2_1187/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_906/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_254 sky130_fd_sc_hd__o22ai_1_265/A2 sky130_fd_sc_hd__nor2_1_150/B
+ sky130_fd_sc_hd__o22ai_1_254/Y sky130_fd_sc_hd__o22ai_1_265/B1 sky130_fd_sc_hd__o32ai_1_2/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_1_0 sky130_fd_sc_hd__nor3_1_0/A sky130_fd_sc_hd__nor2_1_0/Y
+ sky130_fd_sc_hd__nor2_1_1/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nand2_1_318 sky130_fd_sc_hd__nand2_1_318/Y sky130_fd_sc_hd__nand2_1_333/B
+ sky130_fd_sc_hd__nand2_1_318/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_917 sky130_fd_sc_hd__nor2_1_187/B sky130_fd_sc_hd__fa_2_1182/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_917/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_265 sky130_fd_sc_hd__o22ai_1_265/A2 sky130_fd_sc_hd__o22ai_1_265/B1
+ sky130_fd_sc_hd__o22ai_1_265/Y sky130_fd_sc_hd__nor2_1_153/B sky130_fd_sc_hd__o32ai_1_2/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_329 sky130_fd_sc_hd__nand2_1_329/Y sky130_fd_sc_hd__a211o_1_9/A1
+ sky130_fd_sc_hd__o21ai_1_239/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_276 sky130_fd_sc_hd__nand2_1_410/Y sky130_fd_sc_hd__nand2_1_409/Y
+ sky130_fd_sc_hd__o22ai_1_276/Y sky130_fd_sc_hd__o22ai_1_289/A1 sky130_fd_sc_hd__a21o_2_16/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_928 sky130_fd_sc_hd__o22ai_1_319/A1 sky130_fd_sc_hd__nor2_1_224/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_928/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__bufinv_8_2 sky130_fd_sc_hd__bufinv_8_2/A sky130_fd_sc_hd__bufinv_8_2/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufinv_8
Xsky130_fd_sc_hd__o22ai_1_287 sky130_fd_sc_hd__nand2_1_412/Y sky130_fd_sc_hd__nand2_1_411/Y
+ sky130_fd_sc_hd__o22ai_1_287/Y sky130_fd_sc_hd__o22ai_1_287/A1 sky130_fd_sc_hd__a21o_2_15/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_939 sky130_fd_sc_hd__nor2_1_195/B sky130_fd_sc_hd__fa_2_1200/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_939/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_298 sky130_fd_sc_hd__nor2_1_214/A sky130_fd_sc_hd__nor2_1_225/A
+ sky130_fd_sc_hd__o22ai_1_298/Y sky130_fd_sc_hd__a21boi_1_3/Y sky130_fd_sc_hd__a222oi_1_16/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__dfxtp_1_103 VDD VSS sky130_fd_sc_hd__ha_2_1/A sky130_fd_sc_hd__dfxtp_1_95/CLK
+ sky130_fd_sc_hd__and2_0_6/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_114 VDD VSS sky130_fd_sc_hd__nand2_1_34/A sky130_fd_sc_hd__dfxtp_1_117/CLK
+ sky130_fd_sc_hd__ha_2_2/SUM VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_125 VDD VSS sky130_fd_sc_hd__ha_2_15/A sky130_fd_sc_hd__dfxtp_1_129/CLK
+ sky130_fd_sc_hd__and2_0_18/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_136 VDD VSS sky130_fd_sc_hd__ha_2_26/A sky130_fd_sc_hd__dfxtp_1_138/CLK
+ sky130_fd_sc_hd__nor2b_1_7/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_147 VDD VSS sky130_fd_sc_hd__ha_2_39/B sky130_fd_sc_hd__dfxtp_1_155/CLK
+ sky130_fd_sc_hd__and2_0_34/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_158 VDD VSS sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__dfxtp_1_158/CLK
+ sky130_fd_sc_hd__and2_0_29/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_169 VDD VSS sky130_fd_sc_hd__ha_2_40/A sky130_fd_sc_hd__dfxtp_1_170/CLK
+ sky130_fd_sc_hd__nor2b_1_14/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_470 VSS VDD sky130_fd_sc_hd__nor2_1_271/B sky130_fd_sc_hd__o21a_1_68/A1
+ sky130_fd_sc_hd__a21oi_1_460/Y sky130_fd_sc_hd__o21ai_1_470/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_481 VSS VDD sky130_fd_sc_hd__a211oi_1_37/Y sky130_fd_sc_hd__nor2_1_299/A
+ sky130_fd_sc_hd__a21oi_1_468/Y sky130_fd_sc_hd__o21ai_1_481/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_492 VSS VDD sky130_fd_sc_hd__nor2_1_316/Y sky130_fd_sc_hd__o21ai_1_507/A1
+ sky130_fd_sc_hd__nand2_1_553/Y sky130_fd_sc_hd__and2_0_340/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_1202 sky130_fd_sc_hd__fa_2_1203/CIN sky130_fd_sc_hd__mux2_2_138/A1
+ sky130_fd_sc_hd__fa_2_1202/A sky130_fd_sc_hd__fa_2_1202/B sky130_fd_sc_hd__fa_2_1202/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1213 sky130_fd_sc_hd__fa_2_1214/CIN sky130_fd_sc_hd__mux2_2_167/A1
+ sky130_fd_sc_hd__fa_2_1213/A sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__fa_2_1213/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1224 sky130_fd_sc_hd__fa_2_1225/CIN sky130_fd_sc_hd__and2_0_329/A
+ sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1224/B sky130_fd_sc_hd__xor2_1_251/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1235 sky130_fd_sc_hd__fa_2_1236/CIN sky130_fd_sc_hd__mux2_2_187/A1
+ sky130_fd_sc_hd__fa_2_1235/A sky130_fd_sc_hd__fa_2_1235/B sky130_fd_sc_hd__fa_2_1235/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1246 sky130_fd_sc_hd__fa_2_1247/CIN sky130_fd_sc_hd__mux2_2_206/A1
+ sky130_fd_sc_hd__fa_2_1246/A sky130_fd_sc_hd__fa_2_1246/B sky130_fd_sc_hd__fa_2_1246/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1257 sky130_fd_sc_hd__fa_2_1258/CIN sky130_fd_sc_hd__mux2_2_178/A0
+ sky130_fd_sc_hd__fa_2_1257/A sky130_fd_sc_hd__fa_2_1257/B sky130_fd_sc_hd__fa_2_1257/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1010 VDD VSS sky130_fd_sc_hd__mux2_2_93/A0 sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__o22ai_1_229/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_1268 sky130_fd_sc_hd__fa_2_1269/CIN sky130_fd_sc_hd__mux2_2_205/A1
+ sky130_fd_sc_hd__fa_2_1268/A sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1268/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1021 VDD VSS sky130_fd_sc_hd__fa_2_848/A sky130_fd_sc_hd__dfxtp_1_1026/CLK
+ sky130_fd_sc_hd__a21oi_1_315/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_1279 sky130_fd_sc_hd__fa_2_1280/CIN sky130_fd_sc_hd__mux2_2_255/A1
+ sky130_fd_sc_hd__fa_2_1279/A sky130_fd_sc_hd__fa_2_1279/B sky130_fd_sc_hd__fa_2_1279/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o21ai_1_30 VSS VDD sky130_fd_sc_hd__inv_4_1/A sky130_fd_sc_hd__nor4_1_2/Y
+ sky130_fd_sc_hd__o21ai_1_3/B1 sky130_fd_sc_hd__o21ai_1_30/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1032 VDD VSS sky130_fd_sc_hd__fa_2_837/A sky130_fd_sc_hd__dfxtp_1_1038/CLK
+ sky130_fd_sc_hd__a21oi_1_309/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_41 VSS VDD sky130_fd_sc_hd__o21ai_1_53/A2 sky130_fd_sc_hd__xnor2_1_36/Y
+ sky130_fd_sc_hd__a21oi_1_29/Y sky130_fd_sc_hd__o21ai_1_41/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1043 VDD VSS sky130_fd_sc_hd__fa_2_909/B sky130_fd_sc_hd__dfxtp_1_1050/CLK
+ sky130_fd_sc_hd__o21a_1_33/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_52 VSS VDD sky130_fd_sc_hd__o21ai_1_53/A2 sky130_fd_sc_hd__xnor2_1_58/Y
+ sky130_fd_sc_hd__a21oi_1_40/Y sky130_fd_sc_hd__o21ai_1_52/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1054 VDD VSS sky130_fd_sc_hd__fa_2_1193/A sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__mux2_2_164/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_63 VSS VDD sky130_fd_sc_hd__nand2_2_3/Y sky130_fd_sc_hd__xnor2_1_46/Y
+ sky130_fd_sc_hd__a21oi_1_49/Y sky130_fd_sc_hd__o21ai_1_63/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1065 VDD VSS sky130_fd_sc_hd__fa_2_1204/A sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__mux2_2_134/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_74 VSS VDD sky130_fd_sc_hd__xnor2_1_60/A sky130_fd_sc_hd__o21ai_1_74/A1
+ sky130_fd_sc_hd__o21ai_1_74/B1 sky130_fd_sc_hd__o21ai_1_74/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1076 VDD VSS sky130_fd_sc_hd__fa_2_1178/A sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__mux2_2_156/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_85 VSS VDD sky130_fd_sc_hd__xnor2_1_43/A sky130_fd_sc_hd__nor2_1_58/Y
+ sky130_fd_sc_hd__o21ai_1_85/B1 sky130_fd_sc_hd__xnor2_1_45/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1087 VDD VSS sky130_fd_sc_hd__fa_2_1189/A sky130_fd_sc_hd__clkinv_8_70/Y
+ sky130_fd_sc_hd__mux2_2_129/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_96 VSS VDD sky130_fd_sc_hd__a21oi_1_90/Y sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__o21ai_1_96/B1 sky130_fd_sc_hd__xor2_1_64/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1098 VDD VSS sky130_fd_sc_hd__fa_2_1217/A sky130_fd_sc_hd__clkinv_8_65/Y
+ sky130_fd_sc_hd__mux2_2_157/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_670 VDD VSS sky130_fd_sc_hd__fa_2_987/A sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__mux2_2_13/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_681 VDD VSS sky130_fd_sc_hd__fa_2_1020/A sky130_fd_sc_hd__clkinv_8_59/Y
+ sky130_fd_sc_hd__and2_0_273/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_692 VDD VSS sky130_fd_sc_hd__xor2_1_85/A sky130_fd_sc_hd__clkinv_4_26/Y
+ sky130_fd_sc_hd__mux2_2_28/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_290 VSS VDD sky130_fd_sc_hd__clkbuf_1_290/X sky130_fd_sc_hd__clkbuf_1_290/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_520 sky130_fd_sc_hd__fa_2_524/B sky130_fd_sc_hd__fa_2_520/SUM
+ sky130_fd_sc_hd__fa_2_520/A sky130_fd_sc_hd__fa_2_520/B sky130_fd_sc_hd__fa_2_520/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o2bb2ai_1_16 sky130_fd_sc_hd__xor2_1_19/B sky130_fd_sc_hd__nand2_1_203/B
+ sky130_fd_sc_hd__nor2_1_23/Y sky130_fd_sc_hd__nor2_1_23/Y sky130_fd_sc_hd__nand2_1_203/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_531 sky130_fd_sc_hd__fa_2_530/B sky130_fd_sc_hd__fa_2_525/B
+ sky130_fd_sc_hd__fa_2_559/A sky130_fd_sc_hd__fa_2_531/B sky130_fd_sc_hd__fa_2_531/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o2bb2ai_1_27 sky130_fd_sc_hd__and2_0_246/A sky130_fd_sc_hd__nand2_1_216/B
+ sky130_fd_sc_hd__nor2_1_35/Y sky130_fd_sc_hd__nor2_1_35/Y sky130_fd_sc_hd__nand2_1_216/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_542 sky130_fd_sc_hd__fa_2_539/A sky130_fd_sc_hd__fa_2_534/A
+ sky130_fd_sc_hd__fa_2_546/A sky130_fd_sc_hd__ha_2_125/B sky130_fd_sc_hd__fa_2_559/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_553 sky130_fd_sc_hd__fa_2_556/B sky130_fd_sc_hd__fa_2_553/SUM
+ sky130_fd_sc_hd__fa_2_553/A sky130_fd_sc_hd__fa_2_553/B sky130_fd_sc_hd__fa_2_553/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_564 sky130_fd_sc_hd__fa_2_462/B sky130_fd_sc_hd__fa_2_565/CIN
+ sky130_fd_sc_hd__fa_2_567/B sky130_fd_sc_hd__fa_2_564/B sky130_fd_sc_hd__fa_2_537/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_575 sky130_fd_sc_hd__fa_2_574/CIN sky130_fd_sc_hd__and2_0_93/A
+ sky130_fd_sc_hd__fa_2_575/A sky130_fd_sc_hd__fa_2_575/B sky130_fd_sc_hd__fa_2_575/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_586 sky130_fd_sc_hd__maj3_1_129/B sky130_fd_sc_hd__maj3_1_130/A
+ sky130_fd_sc_hd__fa_2_624/B sky130_fd_sc_hd__fa_2_586/B sky130_fd_sc_hd__fa_2_587/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_597 sky130_fd_sc_hd__fa_2_599/CIN sky130_fd_sc_hd__fa_2_595/A
+ sky130_fd_sc_hd__ha_2_128/A sky130_fd_sc_hd__ha_2_126/A sky130_fd_sc_hd__fa_2_683/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor2_1_307 sky130_fd_sc_hd__o21a_1_68/A1 sky130_fd_sc_hd__nor2_1_307/Y
+ sky130_fd_sc_hd__nor2_1_307/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_318 sky130_fd_sc_hd__nor2_1_320/A sky130_fd_sc_hd__nor2_1_318/Y
+ sky130_fd_sc_hd__nor2_1_318/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_503 sky130_fd_sc_hd__buf_12_503/A sky130_fd_sc_hd__buf_12_503/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_514 sky130_fd_sc_hd__buf_12_514/A sky130_fd_sc_hd__buf_12_514/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_406 sky130_fd_sc_hd__nor2_1_315/Y sky130_fd_sc_hd__nor2_1_313/Y
+ sky130_fd_sc_hd__nand3_1_14/Y sky130_fd_sc_hd__nand3_1_15/Y sky130_fd_sc_hd__a31oi_1_4/A2
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nand2_1_104 sky130_fd_sc_hd__nand2_1_104/Y sky130_fd_sc_hd__nand2_1_105/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_703 sky130_fd_sc_hd__o22ai_1_173/A2 sky130_fd_sc_hd__nand3_1_50/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_703/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_115 sky130_fd_sc_hd__nand2_1_115/Y sky130_fd_sc_hd__nand2_1_116/Y
+ sky130_fd_sc_hd__buf_2_264/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_714 sky130_fd_sc_hd__nor2_1_116/B sky130_fd_sc_hd__fa_2_1059/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_714/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_126 sky130_fd_sc_hd__nand2_1_126/Y sky130_fd_sc_hd__fa_2_706/SUM
+ sky130_fd_sc_hd__and2_0_235/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_725 sky130_fd_sc_hd__nor2_1_120/A sky130_fd_sc_hd__fa_2_1051/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_725/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_137 sky130_fd_sc_hd__nand2_1_137/Y sky130_fd_sc_hd__nand2_1_138/Y
+ sky130_fd_sc_hd__buf_2_264/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_736 sky130_fd_sc_hd__o21ai_1_261/A1 sky130_fd_sc_hd__fa_2_1090/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_736/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_148 sky130_fd_sc_hd__o21ai_1_31/A1 sky130_fd_sc_hd__nor3_1_28/Y
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_747 sky130_fd_sc_hd__clkinv_1_747/Y sky130_fd_sc_hd__a21oi_1_239/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_747/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_159 sky130_fd_sc_hd__fa_2_181/CIN sky130_fd_sc_hd__fa_2_281/B
+ sky130_fd_sc_hd__fa_2_258/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_758 sky130_fd_sc_hd__ha_2_190/B sky130_fd_sc_hd__fa_2_1117/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_758/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_769 sky130_fd_sc_hd__nor2_1_141/B sky130_fd_sc_hd__fa_2_1121/COUT
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_769/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor2_1_8 sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__xor2_1_8/X
+ sky130_fd_sc_hd__xor2_1_8/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkinv_8_6 sky130_fd_sc_hd__clkinv_8_6/Y sky130_fd_sc_hd__clkinv_8_6/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_6/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__nor3_1_14 sky130_fd_sc_hd__nor3_2_6/C sky130_fd_sc_hd__nor3_1_14/Y
+ sky130_fd_sc_hd__nor3_2_6/B sky130_fd_sc_hd__nor3_1_16/C VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_25 sky130_fd_sc_hd__nor3_1_25/C sky130_fd_sc_hd__nor3_1_25/Y
+ sky130_fd_sc_hd__nor2_2_5/A sky130_fd_sc_hd__nor3_2_10/A VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_36 sky130_fd_sc_hd__nor3_1_36/C sky130_fd_sc_hd__nor3_1_36/Y
+ sky130_fd_sc_hd__nor3_1_36/A sky130_fd_sc_hd__fa_2_962/A VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__fa_2_1010 sky130_fd_sc_hd__fa_2_1011/CIN sky130_fd_sc_hd__mux2_2_12/A0
+ sky130_fd_sc_hd__fa_2_1010/A sky130_fd_sc_hd__xor2_1_66/X sky130_fd_sc_hd__fa_2_1010/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1021 sky130_fd_sc_hd__fa_2_1022/CIN sky130_fd_sc_hd__and2_0_274/A
+ sky130_fd_sc_hd__fa_2_1021/A sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_1021/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1032 sky130_fd_sc_hd__fa_2_1033/CIN sky130_fd_sc_hd__fa_2_1032/SUM
+ sky130_fd_sc_hd__nor2_1_56/A sky130_fd_sc_hd__fa_2_1032/B sky130_fd_sc_hd__fa_2_1032/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1043 sky130_fd_sc_hd__fa_2_1044/CIN sky130_fd_sc_hd__fa_2_1043/SUM
+ sky130_fd_sc_hd__fa_2_1043/A sky130_fd_sc_hd__nor2_1_49/A sky130_fd_sc_hd__fa_2_1043/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1054 sky130_fd_sc_hd__fa_2_1055/CIN sky130_fd_sc_hd__mux2_2_71/A1
+ sky130_fd_sc_hd__fa_2_1054/A sky130_fd_sc_hd__fa_2_1054/B sky130_fd_sc_hd__fa_2_1054/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1065 sky130_fd_sc_hd__fa_2_1066/CIN sky130_fd_sc_hd__mux2_2_47/A0
+ sky130_fd_sc_hd__fa_2_1065/A sky130_fd_sc_hd__xor2_1_92/X sky130_fd_sc_hd__fa_2_1065/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1076 sky130_fd_sc_hd__fa_2_1077/CIN sky130_fd_sc_hd__mux2_2_72/A1
+ sky130_fd_sc_hd__fa_2_1076/A sky130_fd_sc_hd__fa_2_1076/B sky130_fd_sc_hd__fa_2_1076/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1087 sky130_fd_sc_hd__fa_2_1088/CIN sky130_fd_sc_hd__mux2_2_48/A0
+ sky130_fd_sc_hd__fa_2_1087/A sky130_fd_sc_hd__fa_2_1087/B sky130_fd_sc_hd__fa_2_1087/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1098 sky130_fd_sc_hd__fa_2_1099/CIN sky130_fd_sc_hd__and2_0_300/A
+ sky130_fd_sc_hd__fa_2_1098/A sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1098/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_30 sky130_fd_sc_hd__inv_2_30/A sky130_fd_sc_hd__inv_2_30/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_41 sky130_fd_sc_hd__inv_2_41/A sky130_fd_sc_hd__inv_2_41/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_52 sky130_fd_sc_hd__ha_2_36/A sky130_fd_sc_hd__inv_2_53/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_63 sky130_fd_sc_hd__inv_2_63/A sky130_fd_sc_hd__inv_2_63/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_74 sky130_fd_sc_hd__inv_2_74/A sky130_fd_sc_hd__inv_2_74/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_85 sky130_fd_sc_hd__inv_2_85/A sky130_fd_sc_hd__inv_2_85/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_96 sky130_fd_sc_hd__inv_2_96/A sky130_fd_sc_hd__inv_2_97/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__o32ai_1_11 sky130_fd_sc_hd__nor3_1_41/C sky130_fd_sc_hd__o32ai_1_11/Y
+ sky130_fd_sc_hd__o32ai_1_11/A1 sky130_fd_sc_hd__o32ai_1_11/A3 sky130_fd_sc_hd__o32ai_1_11/B2
+ sky130_fd_sc_hd__o32ai_1_11/B1 VDD VSS VSS VDD sky130_fd_sc_hd__o32ai_1
Xsky130_fd_sc_hd__ha_2_17 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_17/A sky130_fd_sc_hd__ha_2_16/B
+ sky130_fd_sc_hd__ha_2_17/SUM sky130_fd_sc_hd__ha_2_17/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_28 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_28/A sky130_fd_sc_hd__ha_2_27/B
+ sky130_fd_sc_hd__ha_2_28/SUM sky130_fd_sc_hd__ha_2_28/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_39 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_39/A sky130_fd_sc_hd__ha_2_38/B
+ sky130_fd_sc_hd__ha_2_39/SUM sky130_fd_sc_hd__ha_2_39/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_350 sky130_fd_sc_hd__fa_2_349/A sky130_fd_sc_hd__fa_2_344/B
+ sky130_fd_sc_hd__ha_2_109/B sky130_fd_sc_hd__ha_2_116/A sky130_fd_sc_hd__fa_2_401/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_361 sky130_fd_sc_hd__fa_2_363/CIN sky130_fd_sc_hd__fa_2_356/A
+ sky130_fd_sc_hd__fa_2_361/A sky130_fd_sc_hd__fa_2_361/B sky130_fd_sc_hd__fa_2_368/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_372 sky130_fd_sc_hd__fa_2_377/B sky130_fd_sc_hd__fa_2_372/SUM
+ sky130_fd_sc_hd__fa_2_372/A sky130_fd_sc_hd__fa_2_372/B sky130_fd_sc_hd__fa_2_372/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_13 sky130_fd_sc_hd__conb_1_8/LO sky130_fd_sc_hd__clkinv_8_9/Y
+ sky130_fd_sc_hd__dfxtp_1_129/CLK sky130_fd_sc_hd__nand2b_1_0/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_383 sky130_fd_sc_hd__fa_2_387/B sky130_fd_sc_hd__fa_2_383/SUM
+ sky130_fd_sc_hd__fa_2_383/A sky130_fd_sc_hd__fa_2_383/B sky130_fd_sc_hd__fa_2_383/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_24 sky130_fd_sc_hd__conb_1_15/LO sky130_fd_sc_hd__clkinv_4_51/A
+ sky130_fd_sc_hd__dfxtp_1_224/CLK sky130_fd_sc_hd__or2_0_3/X VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_394 sky130_fd_sc_hd__fa_2_395/CIN sky130_fd_sc_hd__fa_2_388/A
+ sky130_fd_sc_hd__ha_2_114/B sky130_fd_sc_hd__fa_2_404/B sky130_fd_sc_hd__fa_2_422/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22oi_2_5 sky130_fd_sc_hd__nor2_4_5/Y sky130_fd_sc_hd__a22oi_2_5/A2
+ sky130_fd_sc_hd__a22oi_2_9/B1 sky130_fd_sc_hd__a22oi_2_5/B2 sky130_fd_sc_hd__a22oi_2_5/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__diode_2_200 sky130_fd_sc_hd__buf_2_269/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__sdlclkp_4_35 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_61/Y
+ sky130_fd_sc_hd__clkinv_4_30/A sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__diode_2_211 sig_frequency[7] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__sdlclkp_4_46 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_68/Y
+ sky130_fd_sc_hd__dfxtp_1_425/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__diode_2_222 sig_amplitude[3] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__sdlclkp_4_57 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__clkinv_8_62/Y
+ sky130_fd_sc_hd__edfxtp_1_0/CLK sky130_fd_sc_hd__nand2b_1_5/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__diode_2_233 sky130_fd_sc_hd__a22oi_1_7/A2 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__sdlclkp_4_68 sky130_fd_sc_hd__conb_1_22/LO sky130_fd_sc_hd__clkinv_8_61/Y
+ sky130_fd_sc_hd__dfxtp_1_577/CLK sky130_fd_sc_hd__nor4_1_5/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_79 sky130_fd_sc_hd__conb_1_25/LO sky130_fd_sc_hd__clkinv_8_118/Y
+ sky130_fd_sc_hd__dfxtp_1_904/CLK sky130_fd_sc_hd__or2_0_9/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_104 sky130_fd_sc_hd__nor2_1_104/B sky130_fd_sc_hd__nor2_1_93/A
+ sky130_fd_sc_hd__fa_2_1109/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_115 sky130_fd_sc_hd__nor2_1_115/B sky130_fd_sc_hd__o21a_1_11/A1
+ sky130_fd_sc_hd__o21a_1_12/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_126 sky130_fd_sc_hd__nor2_1_130/Y sky130_fd_sc_hd__nor2_1_126/Y
+ sky130_fd_sc_hd__nor2_1_126/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_13 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__a22oi_1_9/A1
+ sky130_fd_sc_hd__buf_2_289/X sky130_fd_sc_hd__a22oi_1_13/A2 sky130_fd_sc_hd__nand3_1_6/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_137 sky130_fd_sc_hd__o21a_1_16/A2 sky130_fd_sc_hd__nor2_1_137/Y
+ sky130_fd_sc_hd__nor2_1_137/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_24 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__nor3_2_0/A
+ sky130_fd_sc_hd__nand4_1_35/Y sig_frequency[3] sky130_fd_sc_hd__nand3_1_12/A VDD
+ VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_148 sky130_fd_sc_hd__nor2_1_148/B sky130_fd_sc_hd__o21a_1_22/A1
+ sky130_fd_sc_hd__nor2_1_148/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_35 sky130_fd_sc_hd__clkbuf_4_8/X sky130_fd_sc_hd__clkbuf_4_9/X
+ sky130_fd_sc_hd__clkbuf_1_32/X sky130_fd_sc_hd__a22oi_1_35/A2 sky130_fd_sc_hd__a22oi_1_35/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_159 sky130_fd_sc_hd__nor2_1_163/A sky130_fd_sc_hd__nor2_1_159/Y
+ sky130_fd_sc_hd__xnor2_1_93/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_46 sky130_fd_sc_hd__clkbuf_4_8/X sky130_fd_sc_hd__clkbuf_4_9/X
+ sky130_fd_sc_hd__clkbuf_1_29/X sky130_fd_sc_hd__a22oi_1_46/A2 sky130_fd_sc_hd__a22oi_1_46/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_57 sky130_fd_sc_hd__nor2_2_2/Y sky130_fd_sc_hd__a22oi_1_82/A1
+ sky130_fd_sc_hd__clkbuf_1_62/X sky130_fd_sc_hd__a22oi_1_57/A2 sky130_fd_sc_hd__nand4_1_8/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_68 sky130_fd_sc_hd__clkbuf_4_8/X sky130_fd_sc_hd__clkbuf_4_9/X
+ sky130_fd_sc_hd__clkbuf_1_22/X sky130_fd_sc_hd__a22oi_1_68/A2 sky130_fd_sc_hd__a22oi_1_68/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_79 sky130_fd_sc_hd__a22oi_2_9/B1 sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__clkbuf_4_27/X sky130_fd_sc_hd__a22oi_1_79/A2 sky130_fd_sc_hd__a22oi_1_79/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_300 sky130_fd_sc_hd__buf_8_132/X sky130_fd_sc_hd__buf_8_178/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_311 sky130_fd_sc_hd__bufinv_8_8/Y sky130_fd_sc_hd__buf_12_311/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_322 sky130_fd_sc_hd__buf_4_96/X sky130_fd_sc_hd__buf_12_371/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_333 sky130_fd_sc_hd__buf_4_88/X sky130_fd_sc_hd__buf_12_333/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_344 sky130_fd_sc_hd__buf_6_36/X sky130_fd_sc_hd__buf_12_344/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_203 sky130_fd_sc_hd__clkbuf_1_265/X sky130_fd_sc_hd__clkbuf_1_266/X
+ sky130_fd_sc_hd__clkbuf_1_268/X sky130_fd_sc_hd__a22oi_1_203/A2 sky130_fd_sc_hd__a22oi_1_203/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_355 sky130_fd_sc_hd__buf_12_355/A sky130_fd_sc_hd__buf_12_355/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_214 sky130_fd_sc_hd__buf_2_166/X sky130_fd_sc_hd__buf_2_167/X
+ sky130_fd_sc_hd__clkbuf_1_437/X sky130_fd_sc_hd__buf_2_182/X sky130_fd_sc_hd__nand4_1_49/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_366 sky130_fd_sc_hd__buf_12_366/A sky130_fd_sc_hd__buf_12_366/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_225 sky130_fd_sc_hd__buf_2_166/X sky130_fd_sc_hd__buf_2_167/X
+ sky130_fd_sc_hd__a22oi_1_225/B2 sky130_fd_sc_hd__buf_2_178/X sky130_fd_sc_hd__nand4_1_53/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_377 sky130_fd_sc_hd__buf_2_145/X sky130_fd_sc_hd__buf_2_146/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_236 sky130_fd_sc_hd__buf_2_166/X sky130_fd_sc_hd__buf_2_167/X
+ sky130_fd_sc_hd__clkbuf_1_431/X sky130_fd_sc_hd__buf_2_174/X sky130_fd_sc_hd__nand4_1_57/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_388 sky130_fd_sc_hd__inv_2_123/Y sky130_fd_sc_hd__buf_12_388/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_247 sky130_fd_sc_hd__a22oi_2_25/B1 sky130_fd_sc_hd__a22oi_2_25/A1
+ sky130_fd_sc_hd__clkbuf_1_384/X sky130_fd_sc_hd__a22oi_1_247/A2 sky130_fd_sc_hd__a22oi_1_247/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_399 sky130_fd_sc_hd__buf_8_185/X sky130_fd_sc_hd__buf_12_399/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_258 sky130_fd_sc_hd__clkbuf_1_378/X sky130_fd_sc_hd__clkbuf_1_379/X
+ sky130_fd_sc_hd__clkbuf_4_176/X sky130_fd_sc_hd__buf_2_202/X sky130_fd_sc_hd__nand4_1_64/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_500 sky130_fd_sc_hd__a21oi_1_65/A1 sky130_fd_sc_hd__nor2_1_55/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_500/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22oi_1_269 sky130_fd_sc_hd__clkbuf_4_165/X sky130_fd_sc_hd__clkinv_2_23/Y
+ sky130_fd_sc_hd__clkbuf_1_410/X sky130_fd_sc_hd__a22oi_1_269/A2 sky130_fd_sc_hd__a22oi_1_269/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_511 sky130_fd_sc_hd__o21ai_1_75/A1 sky130_fd_sc_hd__o21ai_1_82/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_511/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_522 sky130_fd_sc_hd__nor2_1_51/B sky130_fd_sc_hd__fa_2_1039/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_522/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_4_109 VDD VSS sky130_fd_sc_hd__buf_4_109/X sky130_fd_sc_hd__buf_8_202/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__clkinv_1_533 sky130_fd_sc_hd__a21oi_1_85/B1 sky130_fd_sc_hd__o211ai_1_5/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_533/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_544 sky130_fd_sc_hd__a21oi_1_89/A1 sky130_fd_sc_hd__a21oi_1_99/Y
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_555 sky130_fd_sc_hd__nand4_1_85/A sky130_fd_sc_hd__fa_2_973/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_555/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_566 sky130_fd_sc_hd__clkinv_1_566/Y sky130_fd_sc_hd__a211oi_1_7/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_566/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_577 sky130_fd_sc_hd__nor2_1_87/A sky130_fd_sc_hd__fa_2_1011/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_577/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_588 sky130_fd_sc_hd__o22ai_1_123/A2 sky130_fd_sc_hd__fa_2_1004/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_588/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_599 sky130_fd_sc_hd__ha_2_174/B sky130_fd_sc_hd__fa_2_1041/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_599/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_4_13 sky130_fd_sc_hd__clkinv_4_13/A sky130_fd_sc_hd__clkinv_4_13/Y
+ VSS VDD VDD VSS VSS sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_24 sky130_fd_sc_hd__clkinv_4_24/A sky130_fd_sc_hd__clkinv_4_24/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_24/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_80 sky130_fd_sc_hd__nor2_1_80/B sky130_fd_sc_hd__nor2_1_80/Y
+ sky130_fd_sc_hd__nor2_1_80/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_35 sky130_fd_sc_hd__clkinv_4_35/A sky130_fd_sc_hd__dfxtp_1_92/D
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_35/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_91 sky130_fd_sc_hd__nor2_1_91/B sky130_fd_sc_hd__nor2_1_91/Y
+ sky130_fd_sc_hd__nor2_1_91/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_46 sky130_fd_sc_hd__clkinv_8_99/A sky130_fd_sc_hd__clkinv_4_49/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_46/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_57 sky130_fd_sc_hd__clkinv_4_57/A sky130_fd_sc_hd__clkinv_8_69/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_57/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_68 sky130_fd_sc_hd__clkinv_2_6/A sky130_fd_sc_hd__clkinv_4_69/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_68/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_79 sky130_fd_sc_hd__clkinv_4_79/A sky130_fd_sc_hd__clkinv_4_80/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_79/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__a21oi_1_430 sky130_fd_sc_hd__o21a_1_64/B1 sky130_fd_sc_hd__o21a_1_63/A1
+ sky130_fd_sc_hd__a21oi_1_430/Y sky130_fd_sc_hd__nor2_1_278/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_441 sky130_fd_sc_hd__nor2_2_18/Y sky130_fd_sc_hd__o21ai_1_448/Y
+ sky130_fd_sc_hd__nor2_1_292/B sky130_fd_sc_hd__fa_2_1280/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_452 sky130_fd_sc_hd__or2_0_12/B sky130_fd_sc_hd__o21ai_1_461/Y
+ sky130_fd_sc_hd__a21oi_1_452/Y sky130_fd_sc_hd__a21oi_1_452/A2 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_463 sky130_fd_sc_hd__fa_2_1301/A sky130_fd_sc_hd__o22ai_1_424/Y
+ sky130_fd_sc_hd__a21oi_1_463/Y sky130_fd_sc_hd__nor3_1_41/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_474 sky130_fd_sc_hd__fa_2_1301/A sky130_fd_sc_hd__o22ai_1_429/Y
+ sky130_fd_sc_hd__a21oi_1_474/Y sky130_fd_sc_hd__nor2_2_18/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_485 sky130_fd_sc_hd__nor2_1_314/Y sky130_fd_sc_hd__nand3_1_52/B
+ sky130_fd_sc_hd__a31oi_1_4/A1 sky130_fd_sc_hd__nand3_1_13/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_496 sky130_fd_sc_hd__nor2_1_319/Y sky130_fd_sc_hd__or2_0_0/B
+ sky130_fd_sc_hd__nand2_1_564/A sky130_fd_sc_hd__nor2_1_320/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_8_110 sky130_fd_sc_hd__clkinv_2_47/A sky130_fd_sc_hd__clkinv_4_55/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_121 sky130_fd_sc_hd__clkinv_8_122/A sky130_fd_sc_hd__clkinv_4_61/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_121/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_132 sky130_fd_sc_hd__clkinv_8_132/Y sky130_fd_sc_hd__clkinv_8_13/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_132/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__o21a_1_1 sky130_fd_sc_hd__o21a_1_1/X sky130_fd_sc_hd__o21a_1_1/A1
+ sky130_fd_sc_hd__o21a_1_1/B1 sky130_fd_sc_hd__fa_2_990/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__xor2_1_307 sky130_fd_sc_hd__nor2_4_20/Y sky130_fd_sc_hd__fa_2_1303/B
+ sky130_fd_sc_hd__xor2_1_307/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_490 sky130_fd_sc_hd__nand2_1_490/Y sky130_fd_sc_hd__nor2b_2_4/A
+ sky130_fd_sc_hd__xor2_1_253/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_318 sky130_fd_sc_hd__xor2_1_318/B sky130_fd_sc_hd__xor2_1_318/X
+ sky130_fd_sc_hd__xor2_1_319/X VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nor2b_1_70 sky130_fd_sc_hd__dfxtp_1_489/Q sky130_fd_sc_hd__nor2b_1_70/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_81 sky130_fd_sc_hd__dfxtp_1_480/Q sky130_fd_sc_hd__nor2b_1_81/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_92 sky130_fd_sc_hd__nor2_1_71/Y sky130_fd_sc_hd__nor2b_1_92/Y
+ sky130_fd_sc_hd__buf_2_262/X VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__xnor2_1_0 VSS VDD sky130_fd_sc_hd__xnor2_1_0/B sky130_fd_sc_hd__xnor2_1_0/Y
+ sky130_fd_sc_hd__xnor2_1_0/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_1070 sky130_fd_sc_hd__nand2_1_528/B sky130_fd_sc_hd__fa_2_22/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1070/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1081 sky130_fd_sc_hd__nor2_1_270/B sky130_fd_sc_hd__fa_2_1288/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1081/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1092 sky130_fd_sc_hd__o21ai_1_479/B1 sky130_fd_sc_hd__nor2_1_304/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1092/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_15 VDD VSS sky130_fd_sc_hd__ha_2_112/A sky130_fd_sc_hd__dfxtp_1_26/CLK
+ sky130_fd_sc_hd__nand4_1_33/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_26 VDD VSS sky130_fd_sc_hd__fa_2_404/A sky130_fd_sc_hd__dfxtp_1_26/CLK
+ sky130_fd_sc_hd__buf_2_286/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_180 sky130_fd_sc_hd__maj3_1_49/B sky130_fd_sc_hd__maj3_1_50/A
+ sky130_fd_sc_hd__fa_2_180/A sky130_fd_sc_hd__fa_2_180/B sky130_fd_sc_hd__fa_2_181/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_37 VDD VSS sky130_fd_sc_hd__fa_2_908/CIN sky130_fd_sc_hd__dfxtp_1_39/CLK
+ sky130_fd_sc_hd__nand4_1_39/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_191 sky130_fd_sc_hd__fa_2_193/CIN sky130_fd_sc_hd__fa_2_189/A
+ sky130_fd_sc_hd__fa_2_242/B sky130_fd_sc_hd__fa_2_283/A sky130_fd_sc_hd__fa_2_191/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_48 VDD VSS sky130_fd_sc_hd__ha_2_118/B sky130_fd_sc_hd__dfxtp_1_61/CLK
+ sky130_fd_sc_hd__nand4_1_34/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_59 VDD VSS sky130_fd_sc_hd__ha_2_124/A sky130_fd_sc_hd__dfxtp_1_61/CLK
+ sky130_fd_sc_hd__dfxtp_1_75/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_4_105 sky130_fd_sc_hd__clkbuf_4_105/X sky130_fd_sc_hd__buf_2_275/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_116 sky130_fd_sc_hd__clkbuf_4_116/X sky130_fd_sc_hd__clkbuf_4_116/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o22ai_1_90 sky130_fd_sc_hd__o22ai_1_90/A2 sky130_fd_sc_hd__nand2_2_4/A
+ sky130_fd_sc_hd__o22ai_1_90/Y sky130_fd_sc_hd__o22ai_1_90/A1 sky130_fd_sc_hd__a21oi_1_81/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkbuf_4_127 sky130_fd_sc_hd__clkbuf_4_127/X sky130_fd_sc_hd__clkbuf_4_127/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_138 sky130_fd_sc_hd__nand4_1_47/B sky130_fd_sc_hd__a22oi_1_209/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_309 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_309/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_309/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_149 sky130_fd_sc_hd__nand4_1_36/B sky130_fd_sc_hd__a22oi_1_165/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_4_70 VDD VSS sky130_fd_sc_hd__buf_4_70/X sky130_fd_sc_hd__buf_4_70/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_81 VDD VSS sky130_fd_sc_hd__buf_4_81/X sky130_fd_sc_hd__buf_4_81/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__inv_2_109 sky130_fd_sc_hd__a22o_2_4/X sky130_fd_sc_hd__inv_2_110/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_4_92 VDD VSS sky130_fd_sc_hd__buf_4_93/A sky130_fd_sc_hd__buf_4_92/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_12_130 sky130_fd_sc_hd__buf_12_130/A sky130_fd_sc_hd__buf_12_238/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_141 sky130_fd_sc_hd__inv_2_64/Y sky130_fd_sc_hd__buf_12_152/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_152 sky130_fd_sc_hd__buf_12_152/A sky130_fd_sc_hd__buf_12_232/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_163 sky130_fd_sc_hd__buf_8_68/X sky130_fd_sc_hd__buf_12_207/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_4_0 sky130_fd_sc_hd__clkbuf_4_0/X sky130_fd_sc_hd__buf_2_1/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_12_174 sky130_fd_sc_hd__buf_8_71/X sky130_fd_sc_hd__buf_12_254/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_185 sky130_fd_sc_hd__buf_8_111/X sky130_fd_sc_hd__buf_12_225/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_196 sky130_fd_sc_hd__buf_4_43/X sky130_fd_sc_hd__buf_12_196/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_330 sky130_fd_sc_hd__fa_2_551/A sky130_fd_sc_hd__ha_2_119/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_330/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_341 sky130_fd_sc_hd__fa_2_700/B sky130_fd_sc_hd__fa_2_701/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_341/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_352 sky130_fd_sc_hd__fa_2_689/B sky130_fd_sc_hd__ha_2_134/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_352/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_363 sky130_fd_sc_hd__ha_2_140/A sky130_fd_sc_hd__fa_2_807/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_363/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_374 sky130_fd_sc_hd__fa_2_874/B sky130_fd_sc_hd__dfxtp_1_274/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_374/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_385 sky130_fd_sc_hd__fa_2_887/B sky130_fd_sc_hd__xor2_1_9/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_385/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_396 sky130_fd_sc_hd__nand2_1_201/B sky130_fd_sc_hd__nand2_1_33/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_396/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21a_1_15 sky130_fd_sc_hd__o21a_1_15/X sky130_fd_sc_hd__o21a_1_15/A1
+ sky130_fd_sc_hd__o21a_1_15/B1 sky130_fd_sc_hd__fa_2_1053/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_26 sky130_fd_sc_hd__o21a_1_26/X sky130_fd_sc_hd__o21a_1_26/A1
+ sky130_fd_sc_hd__o21a_1_26/B1 sky130_fd_sc_hd__fa_2_1150/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_37 sky130_fd_sc_hd__o21a_1_37/X sky130_fd_sc_hd__o21a_1_37/A1
+ sky130_fd_sc_hd__o21a_1_37/B1 sky130_fd_sc_hd__fa_2_1205/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_48 sky130_fd_sc_hd__o21a_1_48/X sky130_fd_sc_hd__o21a_1_48/A1
+ sky130_fd_sc_hd__o21a_1_48/B1 sky130_fd_sc_hd__fa_2_1229/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_59 sky130_fd_sc_hd__o21a_1_59/X sky130_fd_sc_hd__o21a_1_59/A1
+ sky130_fd_sc_hd__o21a_1_59/B1 sky130_fd_sc_hd__fa_2_1285/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__a21oi_1_260 sky130_fd_sc_hd__nor2_2_15/Y sky130_fd_sc_hd__o21ai_1_285/Y
+ sky130_fd_sc_hd__nor2_1_164/B sky130_fd_sc_hd__fa_2_1145/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_271 sky130_fd_sc_hd__nand2_1_387/B sky130_fd_sc_hd__o22ai_1_244/Y
+ sky130_fd_sc_hd__a21oi_1_271/Y sky130_fd_sc_hd__o21ai_1_307/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_282 sky130_fd_sc_hd__nor2b_1_104/Y sky130_fd_sc_hd__o21ai_1_315/Y
+ sky130_fd_sc_hd__a21oi_1_282/Y sky130_fd_sc_hd__o21ai_1_328/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_4_0 sky130_fd_sc_hd__clkinv_4_0/A sky130_fd_sc_hd__clkinv_4_1/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_0/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__a21oi_1_293 sky130_fd_sc_hd__fa_2_1154/A sky130_fd_sc_hd__o22ai_1_257/Y
+ sky130_fd_sc_hd__a21oi_1_293/Y sky130_fd_sc_hd__nor3_1_38/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_201 sky130_fd_sc_hd__buf_8_201/A sky130_fd_sc_hd__buf_8_201/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_212 sky130_fd_sc_hd__buf_8_212/A sky130_fd_sc_hd__buf_8_212/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_223 sky130_fd_sc_hd__buf_8_223/A sky130_fd_sc_hd__buf_8_223/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xor2_1_104 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1053/B
+ sky130_fd_sc_hd__xor2_1_104/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_115 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1091/B
+ sky130_fd_sc_hd__xor2_1_115/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_126 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1080/B
+ sky130_fd_sc_hd__xor2_1_126/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_137 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__xor2_1_137/X
+ sky130_fd_sc_hd__xor2_1_137/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_148 sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__fa_2_1135/B
+ sky130_fd_sc_hd__xor2_1_148/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_159 sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__fa_2_1124/B
+ sky130_fd_sc_hd__xor2_1_159/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_108 VSS VDD sky130_fd_sc_hd__buf_8_31/A sky130_fd_sc_hd__clkbuf_1_124/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_119 VSS VDD sky130_fd_sc_hd__clkbuf_1_119/X sky130_fd_sc_hd__buf_8_7/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__nand3_1_19 sky130_fd_sc_hd__buf_2_24/A sky130_fd_sc_hd__nand3_2_2/A
+ sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__ha_2_10/A VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__dfxtp_1_1406 VDD VSS sky130_fd_sc_hd__mux2_2_229/A1 sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__o22ai_1_383/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1417 VDD VSS sky130_fd_sc_hd__mux2_2_259/A0 sky130_fd_sc_hd__clkinv_8_65/Y
+ sky130_fd_sc_hd__dfxtp_1_432/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1428 VDD VSS sky130_fd_sc_hd__mux2_2_251/A0 sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__o22ai_1_405/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1439 VDD VSS sky130_fd_sc_hd__mux2_2_224/A1 sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__o22ai_1_394/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_106 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_106/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__xnor2_1_6/Y sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_14 sky130_fd_sc_hd__nor3_1_8/C sky130_fd_sc_hd__nor3_2_3/B
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_117 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_117/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_890/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_25 sky130_fd_sc_hd__inv_2_14/A sky130_fd_sc_hd__ha_2_29/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_25/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_128 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_128/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_840/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_36 sky130_fd_sc_hd__inv_2_25/A sky130_fd_sc_hd__buf_2_15/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_36/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_139 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_139/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_856/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_47 sky130_fd_sc_hd__inv_2_36/A sky130_fd_sc_hd__inv_2_3/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_47/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_58 sky130_fd_sc_hd__inv_16_2/A sky130_fd_sc_hd__buf_4_30/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_58/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_1 sky130_fd_sc_hd__fa_2_0/CIN sky130_fd_sc_hd__fa_2_1/SUM sky130_fd_sc_hd__fa_2_1/A
+ sky130_fd_sc_hd__fa_2_1/B sky130_fd_sc_hd__fa_2_1/CIN VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_1_69 sky130_fd_sc_hd__buf_8_86/A sky130_fd_sc_hd__buf_8_76/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_69/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_905 sky130_fd_sc_hd__fa_2_897/A sky130_fd_sc_hd__fa_2_898/B
+ sky130_fd_sc_hd__fa_2_905/A sky130_fd_sc_hd__fa_2_905/B sky130_fd_sc_hd__fa_2_905/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_916 sky130_fd_sc_hd__xor2_1_26/A sky130_fd_sc_hd__fa_2_916/SUM
+ sky130_fd_sc_hd__fa_2_916/A sky130_fd_sc_hd__fa_2_916/B sky130_fd_sc_hd__fa_2_916/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_927 sky130_fd_sc_hd__fa_2_926/CIN sky130_fd_sc_hd__fa_2_927/SUM
+ sky130_fd_sc_hd__fa_2_927/A sky130_fd_sc_hd__fa_2_927/B sky130_fd_sc_hd__fa_2_927/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_938 sky130_fd_sc_hd__fa_2_920/A sky130_fd_sc_hd__fa_2_921/B
+ sky130_fd_sc_hd__fa_2_938/A sky130_fd_sc_hd__fa_2_938/B sky130_fd_sc_hd__ha_2_119/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_949 sky130_fd_sc_hd__fa_2_948/CIN sky130_fd_sc_hd__fa_2_949/SUM
+ sky130_fd_sc_hd__fa_2_949/A sky130_fd_sc_hd__fa_2_949/B sky130_fd_sc_hd__fa_2_949/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__mux2_2_205 VSS VDD sky130_fd_sc_hd__mux2_2_205/A1 sky130_fd_sc_hd__mux2_2_205/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_205/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_216 VSS VDD sky130_fd_sc_hd__mux2_2_216/A1 sky130_fd_sc_hd__mux2_2_216/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_216/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_227 VSS VDD sky130_fd_sc_hd__mux2_2_227/A1 sky130_fd_sc_hd__mux2_2_227/A0
+ sky130_fd_sc_hd__nor2_8_2/A sky130_fd_sc_hd__mux2_2_227/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_238 VSS VDD sky130_fd_sc_hd__mux2_2_238/A1 sky130_fd_sc_hd__mux2_2_238/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_238/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_249 VSS VDD sky130_fd_sc_hd__mux2_2_249/A1 sky130_fd_sc_hd__mux2_2_249/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_249/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__clkinv_1_160 sky130_fd_sc_hd__inv_2_91/A sky130_fd_sc_hd__inv_2_83/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_160/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_171 sky130_fd_sc_hd__inv_2_100/A sky130_fd_sc_hd__buf_8_142/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_171/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_3 sky130_fd_sc_hd__buf_8_3/A sky130_fd_sc_hd__buf_8_3/X VSS
+ VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__a22o_1_5 sig_frequency[6] sky130_fd_sc_hd__nor2_1_1/Y sky130_fd_sc_hd__a22o_1_5/X
+ sky130_fd_sc_hd__a22o_1_5/B2 sky130_fd_sc_hd__nor2_1_0/Y VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_182 sky130_fd_sc_hd__inv_16_7/A sky130_fd_sc_hd__buf_6_34/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_182/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_193 sky130_fd_sc_hd__nand3_2_8/C sky130_fd_sc_hd__a22o_1_27/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_193/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_40 sky130_fd_sc_hd__a22o_1_40/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_40/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__fa_2_946/SUM
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_51 sky130_fd_sc_hd__a22o_1_51/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_51/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__fa_2_957/SUM
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_62 sky130_fd_sc_hd__a22o_1_62/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_62/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__nor4_1_11/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_73 sky130_fd_sc_hd__a22o_1_73/A1 sky130_fd_sc_hd__ha_2_201/SUM
+ sky130_fd_sc_hd__a22o_1_73/X sky130_fd_sc_hd__a22o_1_73/B2 sky130_fd_sc_hd__a22o_1_73/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__nand4_1_1 sky130_fd_sc_hd__nand4_1_1/C sky130_fd_sc_hd__nand4_1_1/B
+ sky130_fd_sc_hd__nand4_1_1/Y sky130_fd_sc_hd__nand4_1_1/D sky130_fd_sc_hd__nand4_1_1/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__o21ai_1_107 VSS VDD sky130_fd_sc_hd__o211ai_1_6/A1 sky130_fd_sc_hd__o22ai_1_132/B1
+ sky130_fd_sc_hd__a22oi_1_325/Y sky130_fd_sc_hd__o21ai_1_107/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_118 VSS VDD sky130_fd_sc_hd__nor2_1_67/B sky130_fd_sc_hd__o21a_1_8/A2
+ sky130_fd_sc_hd__a21oi_1_103/Y sky130_fd_sc_hd__a211o_1_6/A2 VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_129 VSS VDD sky130_fd_sc_hd__nor2_1_77/A sky130_fd_sc_hd__a211oi_1_5/Y
+ sky130_fd_sc_hd__a21oi_1_109/Y sky130_fd_sc_hd__xor2_1_44/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__maj3_1_13 sky130_fd_sc_hd__maj3_1_14/X sky130_fd_sc_hd__maj3_1_13/X
+ sky130_fd_sc_hd__maj3_1_13/B sky130_fd_sc_hd__maj3_1_13/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_24 sky130_fd_sc_hd__maj3_1_25/X sky130_fd_sc_hd__maj3_1_24/X
+ sky130_fd_sc_hd__maj3_1_24/B sky130_fd_sc_hd__maj3_1_24/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_403 sky130_fd_sc_hd__nand2_1_516/Y sky130_fd_sc_hd__nand2_1_515/Y
+ sky130_fd_sc_hd__o22ai_1_403/Y sky130_fd_sc_hd__o22ai_1_403/A1 sky130_fd_sc_hd__a21o_2_28/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_35 sky130_fd_sc_hd__maj3_1_36/X sky130_fd_sc_hd__maj3_1_35/X
+ sky130_fd_sc_hd__maj3_1_35/B sky130_fd_sc_hd__maj3_1_35/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_414 sky130_fd_sc_hd__o22ai_1_436/A2 sky130_fd_sc_hd__nor2_1_303/A
+ sky130_fd_sc_hd__o22ai_1_414/Y sky130_fd_sc_hd__o22ai_1_423/B1 sky130_fd_sc_hd__o32ai_1_11/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_46 sky130_fd_sc_hd__maj3_1_47/X sky130_fd_sc_hd__maj3_1_46/X
+ sky130_fd_sc_hd__maj3_1_46/B sky130_fd_sc_hd__maj3_1_46/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_425 sky130_fd_sc_hd__o22ai_1_436/A2 sky130_fd_sc_hd__nor2_1_277/B
+ sky130_fd_sc_hd__o22ai_1_425/Y sky130_fd_sc_hd__o22ai_1_436/B1 sky130_fd_sc_hd__o32ai_1_11/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_57 sky130_fd_sc_hd__maj3_1_58/X sky130_fd_sc_hd__maj3_1_57/X
+ sky130_fd_sc_hd__maj3_1_57/B sky130_fd_sc_hd__maj3_1_57/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_436 sky130_fd_sc_hd__o22ai_1_436/A2 sky130_fd_sc_hd__o22ai_1_436/B1
+ sky130_fd_sc_hd__o22ai_1_436/Y sky130_fd_sc_hd__nor2_1_280/B sky130_fd_sc_hd__o32ai_1_11/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_68 sky130_fd_sc_hd__maj3_1_69/X sky130_fd_sc_hd__maj3_1_68/X
+ sky130_fd_sc_hd__maj3_1_68/B sky130_fd_sc_hd__maj3_1_68/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_79 sky130_fd_sc_hd__maj3_1_80/X sky130_fd_sc_hd__maj3_1_79/X
+ sky130_fd_sc_hd__maj3_1_79/B sky130_fd_sc_hd__maj3_1_79/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_30 sky130_fd_sc_hd__buf_2_242/A sky130_fd_sc_hd__nor2_1_7/Y
+ sky130_fd_sc_hd__or2_1_2/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_41 sky130_fd_sc_hd__nand2_1_41/Y sky130_fd_sc_hd__nand2_1_41/B
+ sky130_fd_sc_hd__a21oi_2_0/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_52 sky130_fd_sc_hd__nand2_1_52/Y sky130_fd_sc_hd__nand2_1_53/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_63 sky130_fd_sc_hd__nand2_1_63/Y sky130_fd_sc_hd__nand2_1_6/B
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_74 sky130_fd_sc_hd__nand2_1_74/Y sky130_fd_sc_hd__nand2_1_75/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_85 sky130_fd_sc_hd__nand2_1_85/Y sky130_fd_sc_hd__buf_2_265/X
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_96 sky130_fd_sc_hd__nand2_1_96/Y sky130_fd_sc_hd__nand2_1_97/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_307 VDD VSS sky130_fd_sc_hd__a22o_1_42/A1 sky130_fd_sc_hd__dfxtp_1_313/CLK
+ sky130_fd_sc_hd__and2_0_91/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_318 VDD VSS sky130_fd_sc_hd__or4_1_1/B sky130_fd_sc_hd__dfxtp_1_325/CLK
+ sky130_fd_sc_hd__and2_0_198/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_329 VDD VSS sky130_fd_sc_hd__a22o_1_29/B2 sky130_fd_sc_hd__clkinv_4_27/Y
+ sky130_fd_sc_hd__o21ai_1_21/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_15 sky130_fd_sc_hd__fa_2_4/A sky130_fd_sc_hd__fa_2_7/A sky130_fd_sc_hd__ha_2_97/A
+ sky130_fd_sc_hd__fa_2_15/B sky130_fd_sc_hd__fa_2_9/A VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_26 sky130_fd_sc_hd__fa_2_22/CIN sky130_fd_sc_hd__fa_2_26/SUM
+ sky130_fd_sc_hd__fa_2_26/A sky130_fd_sc_hd__fa_2_26/B sky130_fd_sc_hd__fa_2_26/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_37 sky130_fd_sc_hd__fa_2_38/A sky130_fd_sc_hd__fa_2_36/B sky130_fd_sc_hd__ha_2_95/A
+ sky130_fd_sc_hd__fa_2_87/B sky130_fd_sc_hd__fa_2_76/A VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_48 sky130_fd_sc_hd__fa_2_50/A sky130_fd_sc_hd__fa_2_48/SUM
+ sky130_fd_sc_hd__fa_2_48/A sky130_fd_sc_hd__fa_2_48/B sky130_fd_sc_hd__fa_2_53/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_59 sky130_fd_sc_hd__maj3_1_17/B sky130_fd_sc_hd__maj3_1_18/A
+ sky130_fd_sc_hd__fa_2_59/A sky130_fd_sc_hd__fa_2_59/B sky130_fd_sc_hd__fa_2_60/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_207 VDD VSS sky130_fd_sc_hd__buf_2_207/X sky130_fd_sc_hd__buf_2_207/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_218 VDD VSS sky130_fd_sc_hd__buf_2_218/X sky130_fd_sc_hd__buf_2_218/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_229 VDD VSS sky130_fd_sc_hd__buf_2_229/X sky130_fd_sc_hd__buf_2_229/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_sram_2kbyte_1rw1r_32x512_8_11 sky130_fd_sc_hd__buf_4_56/X sky130_fd_sc_hd__buf_4_57/X
+ sky130_fd_sc_hd__buf_4_58/X sky130_fd_sc_hd__clkbuf_4_106/X sky130_fd_sc_hd__clkbuf_4_155/X
+ sky130_fd_sc_hd__buf_4_59/X sky130_fd_sc_hd__buf_4_60/X sky130_fd_sc_hd__buf_4_61/X
+ sky130_fd_sc_hd__buf_4_62/X sky130_fd_sc_hd__clkbuf_4_107/X sky130_fd_sc_hd__buf_4_63/X
+ sky130_fd_sc_hd__buf_4_64/X sky130_fd_sc_hd__buf_4_65/X sky130_fd_sc_hd__buf_4_66/X
+ sky130_fd_sc_hd__clkbuf_4_108/X sky130_fd_sc_hd__buf_4_67/X sky130_fd_sc_hd__buf_4_56/X
+ sky130_fd_sc_hd__buf_4_57/X sky130_fd_sc_hd__buf_4_58/X sky130_fd_sc_hd__clkbuf_4_106/X
+ sky130_fd_sc_hd__clkbuf_4_155/X sky130_fd_sc_hd__buf_4_59/X sky130_fd_sc_hd__buf_4_60/X
+ sky130_fd_sc_hd__buf_4_61/X sky130_fd_sc_hd__buf_4_62/X sky130_fd_sc_hd__clkbuf_4_107/X
+ sky130_fd_sc_hd__buf_4_63/X sky130_fd_sc_hd__buf_4_64/X sky130_fd_sc_hd__buf_4_65/X
+ sky130_fd_sc_hd__buf_4_66/X sky130_fd_sc_hd__clkbuf_4_108/X sky130_fd_sc_hd__buf_4_67/X
+ sky130_fd_sc_hd__buf_12_349/X sky130_fd_sc_hd__buf_12_291/X sky130_fd_sc_hd__buf_12_351/X
+ sky130_fd_sc_hd__buf_12_337/X sky130_fd_sc_hd__buf_12_357/X sky130_fd_sc_hd__buf_12_354/X
+ sky130_fd_sc_hd__buf_12_335/X sky130_fd_sc_hd__buf_12_311/X sky130_fd_sc_hd__buf_12_269/X
+ sky130_fd_sc_hd__buf_12_284/X sky130_fd_sc_hd__buf_12_331/X sky130_fd_sc_hd__buf_12_352/X
+ sky130_fd_sc_hd__buf_12_348/X sky130_fd_sc_hd__buf_12_375/X sky130_fd_sc_hd__buf_12_358/X
+ sky130_fd_sc_hd__buf_12_306/X sky130_fd_sc_hd__buf_12_315/X sky130_fd_sc_hd__buf_12_325/X
+ sky130_fd_sc_hd__clkbuf_1_321/X sky130_fd_sc_hd__buf_2_124/X sky130_fd_sc_hd__clkbuf_1_321/X
+ sky130_fd_sc_hd__clkinv_4_13/Y sky130_fd_sc_hd__clkinv_8_15/Y sky130_fd_sc_hd__buf_12_314/X
+ sky130_fd_sc_hd__buf_8_172/X sky130_fd_sc_hd__buf_12_326/X sky130_fd_sc_hd__buf_12_316/X
+ sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[0] sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[1]
+ sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[2] sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[3]
+ sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[4] sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[5]
+ sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[6] sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[7]
+ sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[8] sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[9]
+ sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[10] sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[11]
+ sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[12] sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[13]
+ sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[14] sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[15]
+ sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[16] sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[17]
+ sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[18] sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[19]
+ sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[20] sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[21]
+ sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[22] sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[23]
+ sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[24] sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[25]
+ sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[26] sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[27]
+ sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[28] sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[29]
+ sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[30] sky130_sram_2kbyte_1rw1r_32x512_8_11/dout0[31]
+ sky130_fd_sc_hd__clkbuf_1_267/A sky130_fd_sc_hd__clkbuf_1_268/A sky130_fd_sc_hd__clkbuf_1_269/A
+ sky130_fd_sc_hd__clkbuf_1_270/A sky130_fd_sc_hd__clkbuf_1_271/A sky130_fd_sc_hd__clkbuf_1_272/A
+ sky130_fd_sc_hd__clkbuf_1_273/A sky130_fd_sc_hd__clkbuf_1_274/A sky130_fd_sc_hd__clkbuf_1_275/A
+ sky130_fd_sc_hd__clkbuf_1_276/A sky130_fd_sc_hd__clkbuf_1_277/A sky130_fd_sc_hd__clkbuf_1_278/A
+ sky130_fd_sc_hd__clkbuf_1_336/A sky130_fd_sc_hd__clkbuf_1_279/A sky130_fd_sc_hd__clkbuf_1_280/A
+ sky130_fd_sc_hd__clkbuf_1_281/A sky130_fd_sc_hd__a22oi_1_207/A2 sky130_fd_sc_hd__a22oi_1_203/A2
+ sky130_fd_sc_hd__a22oi_1_199/A2 sky130_fd_sc_hd__a22oi_1_195/A2 sky130_fd_sc_hd__a22oi_1_191/A2
+ sky130_fd_sc_hd__a22oi_1_187/A2 sky130_fd_sc_hd__a22oi_1_183/A2 sky130_fd_sc_hd__a22oi_1_179/A2
+ sky130_fd_sc_hd__a22oi_1_175/A2 sky130_fd_sc_hd__a22oi_1_171/A2 sky130_fd_sc_hd__a22oi_1_167/A2
+ sky130_fd_sc_hd__a22oi_1_163/A2 sky130_fd_sc_hd__a22oi_1_159/A2 sky130_fd_sc_hd__a22oi_1_155/A2
+ sky130_fd_sc_hd__a22oi_1_151/A2 sky130_fd_sc_hd__a22oi_1_147/A2 VDD VSS sky130_sram_2kbyte_1rw1r_32x512_8
Xsky130_fd_sc_hd__dfxtp_1_1203 VDD VSS sky130_fd_sc_hd__fa_2_1252/A sky130_fd_sc_hd__clkinv_8_75/Y
+ sky130_fd_sc_hd__mux2_2_189/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1214 VDD VSS sky130_fd_sc_hd__fa_2_1226/A sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__mux2_2_213/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1225 VDD VSS sky130_fd_sc_hd__fa_2_1237/A sky130_fd_sc_hd__clkinv_8_78/Y
+ sky130_fd_sc_hd__mux2_2_183/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1236 VDD VSS sky130_fd_sc_hd__fa_2_1265/A sky130_fd_sc_hd__clkinv_8_65/Y
+ sky130_fd_sc_hd__mux2_2_214/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1247 VDD VSS sky130_fd_sc_hd__nor2b_2_4/A sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__nor2b_1_125/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1258 VDD VSS sky130_fd_sc_hd__mux2_2_198/A0 sky130_fd_sc_hd__clkinv_8_78/Y
+ sky130_fd_sc_hd__o22ai_1_333/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_830 VDD VSS sky130_fd_sc_hd__fa_2_1104/A sky130_fd_sc_hd__clkinv_8_54/Y
+ sky130_fd_sc_hd__and2_0_317/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1269 VDD VSS sky130_fd_sc_hd__mux2_2_173/A1 sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__a21oi_1_382/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_841 VDD VSS sky130_fd_sc_hd__mux2_2_73/A0 sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__o21ai_1_158/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_852 VDD VSS sky130_fd_sc_hd__mux2_2_49/A1 sky130_fd_sc_hd__clkinv_4_25/Y
+ sky130_fd_sc_hd__o21ai_1_169/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_863 VDD VSS sky130_fd_sc_hd__mux2_2_67/A0 sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__o21ai_1_177/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_874 VDD VSS sky130_fd_sc_hd__mux2_2_44/A1 sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__o21ai_1_188/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_885 VDD VSS sky130_fd_sc_hd__fa_2_857/A sky130_fd_sc_hd__dfxtp_1_902/CLK
+ sky130_fd_sc_hd__dfxtp_1_885/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_896 VDD VSS sky130_fd_sc_hd__fa_2_931/B sky130_fd_sc_hd__dfxtp_1_899/CLK
+ sky130_fd_sc_hd__dfxtp_1_896/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_450 VSS VDD sky130_fd_sc_hd__clkbuf_1_450/X sky130_fd_sc_hd__clkbuf_1_450/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_461 VSS VDD sky130_fd_sc_hd__clkbuf_1_461/X sky130_fd_sc_hd__clkbuf_1_523/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_472 VSS VDD sky130_fd_sc_hd__clkbuf_1_472/X sky130_fd_sc_hd__clkbuf_1_472/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_483 VSS VDD sky130_fd_sc_hd__buf_6_60/A sky130_fd_sc_hd__a22o_1_22/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_702 sky130_fd_sc_hd__xnor2_1_5/B sky130_fd_sc_hd__fa_2_702/SUM
+ sky130_fd_sc_hd__fa_2_832/A sky130_fd_sc_hd__fa_2_702/B sky130_fd_sc_hd__fa_2_702/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_494 VSS VDD sky130_fd_sc_hd__a22oi_2_28/B2 sky130_fd_sc_hd__clkbuf_1_494/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_713 sky130_fd_sc_hd__fa_2_712/CIN sky130_fd_sc_hd__fa_2_713/SUM
+ sky130_fd_sc_hd__fa_2_713/A sky130_fd_sc_hd__fa_2_713/B sky130_fd_sc_hd__fa_2_713/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_724 sky130_fd_sc_hd__maj3_1_154/B sky130_fd_sc_hd__maj3_1_155/A
+ sky130_fd_sc_hd__fa_2_733/B sky130_fd_sc_hd__fa_2_724/B sky130_fd_sc_hd__fa_2_725/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_735 sky130_fd_sc_hd__maj3_1_150/B sky130_fd_sc_hd__maj3_1_151/A
+ sky130_fd_sc_hd__fa_2_735/A sky130_fd_sc_hd__fa_2_735/B sky130_fd_sc_hd__fa_2_736/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_746 sky130_fd_sc_hd__fa_2_745/B sky130_fd_sc_hd__fa_2_746/SUM
+ sky130_fd_sc_hd__ha_2_140/B sky130_fd_sc_hd__ha_2_141/A sky130_fd_sc_hd__ha_2_139/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_757 sky130_fd_sc_hd__fa_2_760/B sky130_fd_sc_hd__fa_2_757/SUM
+ sky130_fd_sc_hd__fa_2_757/A sky130_fd_sc_hd__fa_2_810/B sky130_fd_sc_hd__fa_2_757/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_768 sky130_fd_sc_hd__fa_2_772/B sky130_fd_sc_hd__fa_2_768/SUM
+ sky130_fd_sc_hd__fa_2_768/A sky130_fd_sc_hd__fa_2_768/B sky130_fd_sc_hd__fa_2_774/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_779 sky130_fd_sc_hd__maj3_1_138/B sky130_fd_sc_hd__maj3_1_139/A
+ sky130_fd_sc_hd__fa_2_779/A sky130_fd_sc_hd__fa_2_779/B sky130_fd_sc_hd__fa_2_780/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor2b_1_110 sky130_fd_sc_hd__and2_0_323/X sky130_fd_sc_hd__nor2b_1_110/Y
+ sky130_fd_sc_hd__buf_2_262/X VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_121 sky130_fd_sc_hd__nor3_1_40/Y sky130_fd_sc_hd__nor2b_1_121/Y
+ sky130_fd_sc_hd__buf_2_262/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_132 sky130_fd_sc_hd__o22ai_1_380/Y sky130_fd_sc_hd__nor2b_1_132/Y
+ sky130_fd_sc_hd__buf_2_262/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__buf_6_0 VDD VSS sky130_fd_sc_hd__buf_6_1/A sky130_fd_sc_hd__buf_6_0/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__bufbuf_8_3 sky130_fd_sc_hd__buf_2_238/A sky130_fd_sc_hd__buf_6_72/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufbuf_8
Xsky130_fd_sc_hd__buf_6_16 VDD VSS sky130_fd_sc_hd__buf_6_16/X sky130_fd_sc_hd__buf_6_16/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_27 VDD VSS sky130_fd_sc_hd__buf_6_27/X sky130_fd_sc_hd__buf_6_27/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_38 VDD VSS sky130_fd_sc_hd__buf_6_38/X sky130_fd_sc_hd__buf_6_38/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_49 VDD VSS sky130_fd_sc_hd__buf_6_49/X sky130_fd_sc_hd__buf_6_49/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_18 sky130_fd_sc_hd__buf_2_123/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_29 sky130_fd_sc_hd__buf_2_77/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__o22ai_1_200 sky130_fd_sc_hd__a21oi_1_226/Y sky130_fd_sc_hd__nor2_1_126/A
+ sky130_fd_sc_hd__o22ai_1_200/Y sky130_fd_sc_hd__nor2_2_13/B sky130_fd_sc_hd__a211oi_1_10/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_211 sky130_fd_sc_hd__nand2_1_358/Y sky130_fd_sc_hd__nand2_1_357/Y
+ sky130_fd_sc_hd__o22ai_1_211/Y sky130_fd_sc_hd__o22ai_1_224/A1 sky130_fd_sc_hd__a21o_2_6/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_222 sky130_fd_sc_hd__nand2_1_358/Y sky130_fd_sc_hd__nand2_1_357/Y
+ sky130_fd_sc_hd__o22ai_1_222/Y sky130_fd_sc_hd__o22ai_1_235/A1 sky130_fd_sc_hd__o21ai_1_283/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_233 sky130_fd_sc_hd__nand2_1_360/Y sky130_fd_sc_hd__nand2_1_359/Y
+ sky130_fd_sc_hd__o22ai_1_233/Y sky130_fd_sc_hd__nand2_1_372/B sky130_fd_sc_hd__o21ai_1_282/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_244 sky130_fd_sc_hd__nor2_1_183/A sky130_fd_sc_hd__nor2_1_172/A
+ sky130_fd_sc_hd__o22ai_1_244/Y sky130_fd_sc_hd__o22ai_1_244/A1 sky130_fd_sc_hd__nor2_1_175/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_308 sky130_fd_sc_hd__o21a_1_9/B1 sky130_fd_sc_hd__o21a_1_9/A2
+ sky130_fd_sc_hd__o21a_1_9/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_907 sky130_fd_sc_hd__o22ai_1_304/A1 sky130_fd_sc_hd__fa_2_1183/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_907/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_255 sky130_fd_sc_hd__nor2_1_183/A sky130_fd_sc_hd__nor2_1_172/A
+ sky130_fd_sc_hd__o22ai_1_255/Y sky130_fd_sc_hd__a21oi_1_290/Y sky130_fd_sc_hd__nor2_1_183/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_1_1 sky130_fd_sc_hd__nor2_1_1/B sky130_fd_sc_hd__nor2_1_1/Y
+ sky130_fd_sc_hd__nor3_2_0/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nand2_1_319 sky130_fd_sc_hd__nand2_1_319/Y sky130_fd_sc_hd__nand2_1_331/B
+ sky130_fd_sc_hd__nand2_1_319/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_918 sky130_fd_sc_hd__nor2_1_186/B sky130_fd_sc_hd__fa_2_1184/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_918/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_266 sky130_fd_sc_hd__a21oi_1_317/Y sky130_fd_sc_hd__nand2_1_393/B
+ sky130_fd_sc_hd__o22ai_1_266/Y sky130_fd_sc_hd__nor3_1_39/C sky130_fd_sc_hd__o32ai_1_5/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_277 sky130_fd_sc_hd__nand2_1_410/Y sky130_fd_sc_hd__nand2_1_409/Y
+ sky130_fd_sc_hd__o22ai_1_277/Y sky130_fd_sc_hd__nand2_1_424/B sky130_fd_sc_hd__o21ai_1_336/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_929 sky130_fd_sc_hd__nand2_1_393/B sky130_fd_sc_hd__nor2b_2_3/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_929/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__bufinv_8_3 sky130_fd_sc_hd__bufinv_8_3/A sky130_fd_sc_hd__bufinv_8_3/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufinv_8
Xsky130_fd_sc_hd__o22ai_1_288 sky130_fd_sc_hd__nand2_1_412/Y sky130_fd_sc_hd__nand2_1_411/Y
+ sky130_fd_sc_hd__o22ai_1_288/Y sky130_fd_sc_hd__nand2_1_423/B sky130_fd_sc_hd__o21ai_1_335/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_299 sky130_fd_sc_hd__o22ai_1_318/A2 sky130_fd_sc_hd__nor2_1_186/B
+ sky130_fd_sc_hd__o22ai_1_299/Y sky130_fd_sc_hd__nor2_1_187/B sky130_fd_sc_hd__o32ai_1_5/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__dfxtp_1_104 VDD VSS sky130_fd_sc_hd__ha_2_0/A sky130_fd_sc_hd__dfxtp_1_95/CLK
+ sky130_fd_sc_hd__and2_0_5/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_115 VDD VSS sky130_fd_sc_hd__nor2_1_21/A sky130_fd_sc_hd__dfxtp_1_117/CLK
+ sky130_fd_sc_hd__ha_2_1/SUM VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_126 VDD VSS sky130_fd_sc_hd__dfxtp_1_126/Q sky130_fd_sc_hd__dfxtp_1_126/CLK
+ sky130_fd_sc_hd__and2_1_0/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_137 VDD VSS sky130_fd_sc_hd__ha_2_25/A sky130_fd_sc_hd__dfxtp_1_138/CLK
+ sky130_fd_sc_hd__nor2b_1_4/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_148 VDD VSS sky130_fd_sc_hd__ha_2_39/A sky130_fd_sc_hd__dfxtp_1_155/CLK
+ sky130_fd_sc_hd__and2_0_33/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_159 VDD VSS sky130_fd_sc_hd__ha_2_49/B sky130_fd_sc_hd__dfxtp_1_170/CLK
+ sky130_fd_sc_hd__nor2b_1_16/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_460 VSS VDD sky130_fd_sc_hd__nor3_1_41/A sky130_fd_sc_hd__nor2_1_300/A
+ sky130_fd_sc_hd__nand2_1_536/Y sky130_fd_sc_hd__o21ai_1_460/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_471 VSS VDD sky130_fd_sc_hd__a21oi_1_470/Y sky130_fd_sc_hd__nor2_1_309/A
+ sky130_fd_sc_hd__nand2_1_538/Y sky130_fd_sc_hd__xor2_1_279/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_482 VSS VDD sky130_fd_sc_hd__o21a_1_68/X sky130_fd_sc_hd__nor2_1_307/A
+ sky130_fd_sc_hd__a21oi_1_469/Y sky130_fd_sc_hd__xor2_1_291/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_493 VSS VDD sky130_fd_sc_hd__nand2_1_554/A sky130_fd_sc_hd__o21ai_1_507/A1
+ sky130_fd_sc_hd__nand2_1_554/Y sky130_fd_sc_hd__and2_0_344/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_1203 sky130_fd_sc_hd__fa_2_1204/CIN sky130_fd_sc_hd__mux2_2_136/A1
+ sky130_fd_sc_hd__fa_2_1203/A sky130_fd_sc_hd__fa_2_1203/B sky130_fd_sc_hd__fa_2_1203/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1214 sky130_fd_sc_hd__fa_2_1215/CIN sky130_fd_sc_hd__mux2_2_166/A1
+ sky130_fd_sc_hd__fa_2_1214/A sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__fa_2_1214/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1225 sky130_fd_sc_hd__fa_2_1226/CIN sky130_fd_sc_hd__and2_0_331/A
+ sky130_fd_sc_hd__fa_2_1225/A sky130_fd_sc_hd__fa_2_1225/B sky130_fd_sc_hd__fa_2_1225/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1236 sky130_fd_sc_hd__fa_2_1237/CIN sky130_fd_sc_hd__mux2_2_185/A1
+ sky130_fd_sc_hd__fa_2_1236/A sky130_fd_sc_hd__fa_2_1236/B sky130_fd_sc_hd__fa_2_1236/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1247 sky130_fd_sc_hd__fa_2_1248/CIN sky130_fd_sc_hd__mux2_2_203/A1
+ sky130_fd_sc_hd__fa_2_1247/A sky130_fd_sc_hd__fa_2_1247/B sky130_fd_sc_hd__fa_2_1247/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1000 VDD VSS sky130_fd_sc_hd__mux2_2_97/A0 sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__dfxtp_1_454/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_1258 sky130_fd_sc_hd__fa_2_1259/CIN sky130_fd_sc_hd__mux2_2_176/A0
+ sky130_fd_sc_hd__fa_2_1258/A sky130_fd_sc_hd__fa_2_1258/B sky130_fd_sc_hd__fa_2_1258/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1011 VDD VSS sky130_fd_sc_hd__mux2_2_90/A0 sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__o22ai_1_228/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_20 VSS VDD sky130_fd_sc_hd__a21oi_2_0/Y sky130_fd_sc_hd__o22ai_1_0/B2
+ sky130_fd_sc_hd__nand2_1_39/Y sky130_fd_sc_hd__o21ai_1_20/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_1269 sky130_fd_sc_hd__fa_2_1270/CIN sky130_fd_sc_hd__mux2_2_202/A1
+ sky130_fd_sc_hd__fa_2_1269/A sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1269/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1022 VDD VSS sky130_fd_sc_hd__fa_2_847/A sky130_fd_sc_hd__dfxtp_1_1026/CLK
+ sky130_fd_sc_hd__o21a_1_41/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_31 VSS VDD sky130_fd_sc_hd__nor2_1_13/B sky130_fd_sc_hd__o21ai_1_31/A1
+ sky130_fd_sc_hd__o21ai_1_31/B1 sky130_fd_sc_hd__o21ai_1_31/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1033 VDD VSS sky130_fd_sc_hd__fa_2_836/A sky130_fd_sc_hd__dfxtp_1_1050/CLK
+ sky130_fd_sc_hd__o21a_1_36/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_42 VSS VDD sky130_fd_sc_hd__o21ai_1_53/A2 sky130_fd_sc_hd__xnor2_1_38/Y
+ sky130_fd_sc_hd__a21oi_1_30/Y sky130_fd_sc_hd__o21ai_1_42/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1044 VDD VSS sky130_fd_sc_hd__fa_2_910/B sky130_fd_sc_hd__dfxtp_1_1047/CLK
+ sky130_fd_sc_hd__a21oi_1_303/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_53 VSS VDD sky130_fd_sc_hd__o21ai_1_53/A2 sky130_fd_sc_hd__xnor2_1_60/Y
+ sky130_fd_sc_hd__a21oi_1_41/Y sky130_fd_sc_hd__o21ai_1_53/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1055 VDD VSS sky130_fd_sc_hd__fa_2_1194/A sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__mux2_2_161/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_64 VSS VDD sky130_fd_sc_hd__nand2_2_3/Y sky130_fd_sc_hd__xnor2_1_48/Y
+ sky130_fd_sc_hd__a21oi_1_50/Y sky130_fd_sc_hd__o21ai_1_64/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1066 VDD VSS sky130_fd_sc_hd__fa_2_1205/A sky130_fd_sc_hd__clkinv_8_70/Y
+ sky130_fd_sc_hd__mux2_2_132/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_75 VSS VDD sky130_fd_sc_hd__xnor2_1_56/A sky130_fd_sc_hd__o21ai_1_75/A1
+ sky130_fd_sc_hd__o21ai_1_75/B1 sky130_fd_sc_hd__xnor2_1_58/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1077 VDD VSS sky130_fd_sc_hd__fa_2_1179/A sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__mux2_2_153/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_86 VSS VDD sky130_fd_sc_hd__xnor2_1_39/A sky130_fd_sc_hd__nor2_1_57/Y
+ sky130_fd_sc_hd__o21ai_1_86/B1 sky130_fd_sc_hd__xnor2_1_41/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1088 VDD VSS sky130_fd_sc_hd__fa_2_1190/A sky130_fd_sc_hd__clkinv_8_70/Y
+ sky130_fd_sc_hd__mux2_2_127/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_97 VSS VDD sky130_fd_sc_hd__nor2_1_74/A sky130_fd_sc_hd__o22ai_1_99/A2
+ sky130_fd_sc_hd__a21oi_1_84/Y sky130_fd_sc_hd__xor2_1_67/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_660 VDD VSS sky130_fd_sc_hd__fa_2_977/A sky130_fd_sc_hd__clkinv_8_41/Y
+ sky130_fd_sc_hd__mux2_2_35/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1099 VDD VSS sky130_fd_sc_hd__fa_2_1218/A sky130_fd_sc_hd__clkinv_8_65/Y
+ sky130_fd_sc_hd__mux2_2_154/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_671 VDD VSS sky130_fd_sc_hd__fa_2_988/A sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__mux2_2_11/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_682 VDD VSS sky130_fd_sc_hd__fa_2_1021/A sky130_fd_sc_hd__clkinv_8_59/Y
+ sky130_fd_sc_hd__and2_0_274/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_693 VDD VSS sky130_fd_sc_hd__o22ai_1_90/A1 sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__nor2b_1_95/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_280 VSS VDD sky130_fd_sc_hd__clkbuf_1_280/X sky130_fd_sc_hd__clkbuf_1_280/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_291 VSS VDD sky130_fd_sc_hd__clkbuf_1_291/X sky130_fd_sc_hd__clkbuf_1_291/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_510 sky130_fd_sc_hd__fa_2_507/A sky130_fd_sc_hd__fa_2_510/SUM
+ sky130_fd_sc_hd__ha_2_124/B sky130_fd_sc_hd__ha_2_125/A sky130_fd_sc_hd__fa_2_502/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_521 sky130_fd_sc_hd__fa_2_523/CIN sky130_fd_sc_hd__fa_2_514/B
+ sky130_fd_sc_hd__fa_2_567/B sky130_fd_sc_hd__fa_2_566/B sky130_fd_sc_hd__fa_2_558/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o2bb2ai_1_17 sky130_fd_sc_hd__dfxtp_1_554/D sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__dfxtp_1_554/Q sky130_fd_sc_hd__nor4_1_5/C sky130_fd_sc_hd__nand3_1_44/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_532 sky130_fd_sc_hd__fa_2_534/CIN sky130_fd_sc_hd__fa_2_529/A
+ sky130_fd_sc_hd__fa_2_532/A sky130_fd_sc_hd__fa_2_532/B sky130_fd_sc_hd__fa_2_540/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o2bb2ai_1_28 sky130_fd_sc_hd__and2_0_243/A sky130_fd_sc_hd__nand2_1_215/B
+ sky130_fd_sc_hd__nor2_1_34/Y sky130_fd_sc_hd__nor2_1_34/Y sky130_fd_sc_hd__nand2_1_215/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_543 sky130_fd_sc_hd__fa_2_545/CIN sky130_fd_sc_hd__fa_2_538/A
+ sky130_fd_sc_hd__fa_2_543/A sky130_fd_sc_hd__fa_2_543/B sky130_fd_sc_hd__fa_2_543/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_554 sky130_fd_sc_hd__fa_2_555/CIN sky130_fd_sc_hd__fa_2_549/A
+ sky130_fd_sc_hd__fa_2_554/A sky130_fd_sc_hd__fa_2_567/A sky130_fd_sc_hd__fa_2_543/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_565 sky130_fd_sc_hd__fa_2_463/B sky130_fd_sc_hd__fa_2_565/SUM
+ sky130_fd_sc_hd__fa_2_565/A sky130_fd_sc_hd__fa_2_565/B sky130_fd_sc_hd__fa_2_565/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_576 sky130_fd_sc_hd__fa_2_575/CIN sky130_fd_sc_hd__and2_0_94/A
+ sky130_fd_sc_hd__fa_2_576/A sky130_fd_sc_hd__fa_2_576/B sky130_fd_sc_hd__fa_2_576/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_587 sky130_fd_sc_hd__fa_2_588/B sky130_fd_sc_hd__fa_2_587/SUM
+ sky130_fd_sc_hd__ha_2_134/A sky130_fd_sc_hd__ha_2_131/A sky130_fd_sc_hd__ha_2_132/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_598 sky130_fd_sc_hd__maj3_1_124/B sky130_fd_sc_hd__maj3_1_125/A
+ sky130_fd_sc_hd__fa_2_598/A sky130_fd_sc_hd__fa_2_598/B sky130_fd_sc_hd__fa_2_599/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor2_1_308 sky130_fd_sc_hd__o21a_1_68/A1 sky130_fd_sc_hd__nor2_1_308/Y
+ sky130_fd_sc_hd__nor2_1_308/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_319 sky130_fd_sc_hd__nor2_1_323/A sky130_fd_sc_hd__nor2_1_319/Y
+ sky130_fd_sc_hd__nor2_1_319/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_504 sky130_fd_sc_hd__buf_12_504/A sky130_fd_sc_hd__buf_12_504/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_515 sky130_fd_sc_hd__buf_12_515/A sky130_fd_sc_hd__buf_12_515/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__nand2_1_105 sky130_fd_sc_hd__nand2_1_105/Y sky130_fd_sc_hd__buf_2_269/X
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_704 sky130_fd_sc_hd__o21ai_1_229/A2 sky130_fd_sc_hd__o21ai_1_239/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_704/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_116 sky130_fd_sc_hd__nand2_1_116/Y sky130_fd_sc_hd__xnor2_1_5/Y
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_715 sky130_fd_sc_hd__o22ai_1_191/A1 sky130_fd_sc_hd__fa_2_1058/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_715/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_127 sky130_fd_sc_hd__nand2_1_127/Y sky130_fd_sc_hd__nand2_1_128/Y
+ sky130_fd_sc_hd__buf_2_264/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_726 sky130_fd_sc_hd__clkinv_1_726/Y sky130_fd_sc_hd__nand2_1_334/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_726/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_138 sky130_fd_sc_hd__nand2_1_138/Y sky130_fd_sc_hd__fa_2_712/SUM
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_737 sky130_fd_sc_hd__nor2_1_136/A sky130_fd_sc_hd__fa_2_1088/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_737/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_149 sky130_fd_sc_hd__fa_2_34/B sky130_fd_sc_hd__fa_2_66/B
+ sky130_fd_sc_hd__fa_2_49/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_748 sky130_fd_sc_hd__nor2_4_13/B sky130_fd_sc_hd__nor2_4_12/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_748/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_759 sky130_fd_sc_hd__ha_2_191/B sky130_fd_sc_hd__fa_2_1116/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_759/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor2_1_9 sky130_fd_sc_hd__xor2_1_9/B sky130_fd_sc_hd__xor2_1_9/X
+ sky130_fd_sc_hd__xor2_1_9/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkinv_8_7 sky130_fd_sc_hd__clkinv_8_7/Y sky130_fd_sc_hd__clkinv_8_7/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__o21ai_1_290 VSS VDD sky130_fd_sc_hd__nor2_1_172/B sky130_fd_sc_hd__nor2_1_182/A
+ sky130_fd_sc_hd__nand2_1_373/Y sky130_fd_sc_hd__xor2_1_167/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor3_1_15 sky130_fd_sc_hd__nor3_1_17/C sky130_fd_sc_hd__nor3_1_15/Y
+ sky130_fd_sc_hd__nor3_2_6/A sky130_fd_sc_hd__nor3_2_6/C VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_26 sky130_fd_sc_hd__nor3_1_26/C sky130_fd_sc_hd__nor3_1_26/Y
+ sky130_fd_sc_hd__nor3_1_26/A sky130_fd_sc_hd__nor3_1_27/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_37 sky130_fd_sc_hd__nor3_1_37/C sky130_fd_sc_hd__nor3_1_37/Y
+ sky130_fd_sc_hd__nor3_1_37/A sky130_fd_sc_hd__fa_2_968/A VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__fa_2_1000 sky130_fd_sc_hd__fa_2_1001/CIN sky130_fd_sc_hd__mux2_2_34/A1
+ sky130_fd_sc_hd__fa_2_1000/A sky130_fd_sc_hd__xor2_1_76/X sky130_fd_sc_hd__fa_2_999/COUT
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1011 sky130_fd_sc_hd__fa_2_1012/CIN sky130_fd_sc_hd__mux2_2_10/A0
+ sky130_fd_sc_hd__fa_2_1011/A sky130_fd_sc_hd__xor2_1_65/X sky130_fd_sc_hd__fa_2_1011/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1022 sky130_fd_sc_hd__fa_2_1023/CIN sky130_fd_sc_hd__and2_0_275/A
+ sky130_fd_sc_hd__fa_2_1022/A sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_1022/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1033 sky130_fd_sc_hd__fa_2_1034/CIN sky130_fd_sc_hd__fa_2_1033/SUM
+ sky130_fd_sc_hd__fa_2_1033/A sky130_fd_sc_hd__nor2_1_54/A sky130_fd_sc_hd__fa_2_1033/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1044 sky130_fd_sc_hd__fa_2_1045/CIN sky130_fd_sc_hd__fa_2_1044/SUM
+ sky130_fd_sc_hd__nor2_1_62/A sky130_fd_sc_hd__fa_2_1044/B sky130_fd_sc_hd__fa_2_1044/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1055 sky130_fd_sc_hd__fa_2_1056/CIN sky130_fd_sc_hd__mux2_2_69/A1
+ sky130_fd_sc_hd__fa_2_1055/A sky130_fd_sc_hd__fa_2_1055/B sky130_fd_sc_hd__fa_2_1055/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1066 sky130_fd_sc_hd__fa_2_1067/CIN sky130_fd_sc_hd__mux2_2_45/A0
+ sky130_fd_sc_hd__o21a_1_9/A2 sky130_fd_sc_hd__xor2_1_91/X sky130_fd_sc_hd__fa_2_1066/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1077 sky130_fd_sc_hd__fa_2_1078/CIN sky130_fd_sc_hd__mux2_2_70/A1
+ sky130_fd_sc_hd__fa_2_1077/A sky130_fd_sc_hd__fa_2_1077/B sky130_fd_sc_hd__fa_2_1077/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1088 sky130_fd_sc_hd__fa_2_1089/CIN sky130_fd_sc_hd__mux2_2_46/A0
+ sky130_fd_sc_hd__fa_2_1088/A sky130_fd_sc_hd__fa_2_1088/B sky130_fd_sc_hd__fa_2_1088/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1099 sky130_fd_sc_hd__fa_2_1100/CIN sky130_fd_sc_hd__and2_0_305/A
+ sky130_fd_sc_hd__fa_2_1099/A sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1099/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_20 sky130_fd_sc_hd__inv_2_20/A sky130_fd_sc_hd__inv_2_20/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_31 sky130_fd_sc_hd__inv_2_31/A sky130_fd_sc_hd__buf_8_0/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_42 sky130_fd_sc_hd__inv_2_42/A sky130_fd_sc_hd__inv_2_42/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_53 sky130_fd_sc_hd__inv_2_53/A sky130_fd_sc_hd__inv_2_53/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_64 sky130_fd_sc_hd__inv_2_64/A sky130_fd_sc_hd__inv_2_64/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_75 sky130_fd_sc_hd__inv_2_75/A sky130_fd_sc_hd__inv_2_75/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_86 sky130_fd_sc_hd__inv_2_86/A sky130_fd_sc_hd__inv_2_86/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_490 VDD VSS sky130_fd_sc_hd__dfxtp_1_490/Q sky130_fd_sc_hd__dfxtp_1_496/CLK
+ sky130_fd_sc_hd__nor2b_1_65/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_97 sky130_fd_sc_hd__inv_2_97/A sky130_fd_sc_hd__inv_2_97/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__ha_2_18 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_18/A sky130_fd_sc_hd__ha_2_17/B
+ sky130_fd_sc_hd__ha_2_18/SUM sky130_fd_sc_hd__ha_2_18/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_29 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_29/A sky130_fd_sc_hd__ha_2_28/B
+ sky130_fd_sc_hd__ha_2_29/SUM sky130_fd_sc_hd__ha_2_29/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_340 sky130_fd_sc_hd__maj3_1_72/B sky130_fd_sc_hd__maj3_1_73/A
+ sky130_fd_sc_hd__fa_2_340/A sky130_fd_sc_hd__fa_2_340/B sky130_fd_sc_hd__fa_2_341/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_351 sky130_fd_sc_hd__fa_2_349/B sky130_fd_sc_hd__fa_2_344/A
+ sky130_fd_sc_hd__ha_2_115/A sky130_fd_sc_hd__ha_2_112/A sky130_fd_sc_hd__fa_2_404/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_362 sky130_fd_sc_hd__maj3_1_67/B sky130_fd_sc_hd__maj3_1_68/A
+ sky130_fd_sc_hd__fa_2_362/A sky130_fd_sc_hd__fa_2_362/B sky130_fd_sc_hd__fa_2_363/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_373 sky130_fd_sc_hd__fa_2_370/B sky130_fd_sc_hd__fa_2_373/SUM
+ sky130_fd_sc_hd__ha_2_114/A sky130_fd_sc_hd__fa_2_412/A sky130_fd_sc_hd__fa_2_424/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_14 sky130_fd_sc_hd__conb_1_9/LO sky130_fd_sc_hd__clkinv_8_9/Y
+ sky130_fd_sc_hd__dfxtp_1_138/CLK sky130_fd_sc_hd__or2_0_1/X VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_384 sky130_fd_sc_hd__fa_2_386/CIN sky130_fd_sc_hd__fa_2_378/B
+ sky130_fd_sc_hd__fa_2_424/B sky130_fd_sc_hd__fa_2_417/B sky130_fd_sc_hd__fa_2_384/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_25 sky130_fd_sc_hd__conb_1_17/LO sky130_fd_sc_hd__clkinv_8_100/Y
+ sky130_fd_sc_hd__dfxtp_1_360/CLK sky130_fd_sc_hd__nor2_1_14/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__and2_1_0 VDD VSS sky130_fd_sc_hd__and2_1_0/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__and2_1_0/A VDD VSS sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__fa_2_395 sky130_fd_sc_hd__fa_2_397/CIN sky130_fd_sc_hd__fa_2_391/A
+ sky130_fd_sc_hd__fa_2_395/A sky130_fd_sc_hd__fa_2_395/B sky130_fd_sc_hd__fa_2_395/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22oi_2_6 sky130_fd_sc_hd__nor2_4_5/Y sky130_fd_sc_hd__a22oi_2_6/A2
+ sky130_fd_sc_hd__a22oi_2_9/B1 sky130_fd_sc_hd__a22oi_2_6/B2 sky130_fd_sc_hd__a22oi_2_6/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__diode_2_201 sky130_fd_sc_hd__buf_2_268/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__sdlclkp_4_36 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_100/Y
+ sky130_fd_sc_hd__dfxtp_1_347/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__diode_2_212 amplitude_adc_done VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__sdlclkp_4_47 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_4_53/Y
+ sky130_fd_sc_hd__dfxtp_1_452/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__diode_2_223 sig_amplitude[3] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__sdlclkp_4_58 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__clkinv_8_62/Y
+ sky130_fd_sc_hd__dfxtp_1_502/CLK sky130_fd_sc_hd__nand2b_1_5/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__diode_2_234 sky130_fd_sc_hd__a22oi_1_7/A2 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__sdlclkp_4_69 sky130_fd_sc_hd__conb_1_23/LO sky130_fd_sc_hd__clkinv_8_58/A
+ sky130_fd_sc_hd__dfxtp_1_611/CLK sky130_fd_sc_hd__or2_0_6/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_105 sky130_fd_sc_hd__nor2_1_105/B sky130_fd_sc_hd__nor2_1_92/A
+ sky130_fd_sc_hd__fa_2_1107/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_116 sky130_fd_sc_hd__nor2_1_116/B sky130_fd_sc_hd__o21a_1_12/A1
+ sky130_fd_sc_hd__o21a_1_13/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_127 sky130_fd_sc_hd__nor2_1_129/Y sky130_fd_sc_hd__nor2_1_127/Y
+ sky130_fd_sc_hd__nor2_1_127/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_14 sky130_fd_sc_hd__nor2_2_0/Y sky130_fd_sc_hd__clkinv_1_4/Y
+ sky130_fd_sc_hd__nand4_1_24/Y sky130_fd_sc_hd__nand4_1_8/Y sky130_fd_sc_hd__a22oi_1_14/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_138 sky130_fd_sc_hd__o21a_1_16/A2 sky130_fd_sc_hd__nor2_1_138/Y
+ sky130_fd_sc_hd__nor2_1_138/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_149 sky130_fd_sc_hd__nor2_1_149/B sky130_fd_sc_hd__nor2_1_149/Y
+ sky130_fd_sc_hd__nor2_1_149/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_25 sky130_fd_sc_hd__nor2_2_0/Y sky130_fd_sc_hd__clkinv_1_4/Y
+ sky130_fd_sc_hd__nand4_1_18/Y sky130_fd_sc_hd__nand4_1_2/Y sky130_fd_sc_hd__a22oi_1_25/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_36 sky130_fd_sc_hd__a22oi_1_81/B1 sky130_fd_sc_hd__clkbuf_1_99/X
+ sky130_fd_sc_hd__clkbuf_1_48/X sky130_fd_sc_hd__clkbuf_4_23/X sky130_fd_sc_hd__nand4_1_2/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_47 sky130_fd_sc_hd__a22oi_1_81/B1 sky130_fd_sc_hd__clkbuf_1_99/X
+ sky130_fd_sc_hd__clkbuf_1_45/X sky130_fd_sc_hd__clkbuf_4_20/X sky130_fd_sc_hd__nand4_1_5/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_58 sky130_fd_sc_hd__clkbuf_4_8/X sky130_fd_sc_hd__clkbuf_4_9/X
+ sky130_fd_sc_hd__clkbuf_1_25/X sky130_fd_sc_hd__a22oi_1_58/A2 sky130_fd_sc_hd__a22oi_1_58/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_69 sky130_fd_sc_hd__a22oi_1_81/B1 sky130_fd_sc_hd__clkbuf_1_99/X
+ sky130_fd_sc_hd__clkbuf_1_38/X sky130_fd_sc_hd__clkbuf_4_13/X sky130_fd_sc_hd__nand4_1_12/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_301 sky130_fd_sc_hd__buf_8_137/X sky130_fd_sc_hd__buf_12_301/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_312 sky130_fd_sc_hd__bufinv_8_6/Y sky130_fd_sc_hd__buf_12_312/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_323 sky130_fd_sc_hd__buf_4_83/X sky130_fd_sc_hd__buf_12_323/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_334 sky130_fd_sc_hd__buf_4_77/X sky130_fd_sc_hd__buf_12_334/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_345 sky130_fd_sc_hd__buf_6_42/X sky130_fd_sc_hd__buf_12_345/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_204 sky130_fd_sc_hd__clkbuf_1_351/X sky130_fd_sc_hd__clkbuf_1_353/X
+ sky130_fd_sc_hd__clkbuf_4_114/X sky130_fd_sc_hd__a22oi_1_204/A2 sky130_fd_sc_hd__nand4_1_46/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_356 sky130_fd_sc_hd__buf_12_356/A sky130_fd_sc_hd__buf_12_356/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_215 sky130_fd_sc_hd__nor2_4_7/Y sky130_fd_sc_hd__buf_2_165/X
+ sky130_fd_sc_hd__a22oi_1_215/B2 sky130_fd_sc_hd__clkbuf_1_453/X sky130_fd_sc_hd__a22oi_1_215/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_367 sky130_fd_sc_hd__buf_12_367/A sky130_fd_sc_hd__buf_12_367/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_226 sky130_fd_sc_hd__nor2_4_7/Y sky130_fd_sc_hd__buf_2_165/X
+ sky130_fd_sc_hd__a22oi_1_226/B2 sky130_fd_sc_hd__clkbuf_1_449/X sky130_fd_sc_hd__nand4_1_53/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_378 sky130_fd_sc_hd__dfxtp_1_87/D sky130_fd_sc_hd__buf_2_153/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_237 sky130_fd_sc_hd__nor2_4_7/Y sky130_fd_sc_hd__buf_2_165/X
+ sky130_fd_sc_hd__clkbuf_1_497/X sky130_fd_sc_hd__clkbuf_1_445/X sky130_fd_sc_hd__a22oi_1_237/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_389 sky130_fd_sc_hd__buf_12_389/A sky130_fd_sc_hd__buf_6_75/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_248 sky130_fd_sc_hd__buf_2_166/X sky130_fd_sc_hd__buf_2_167/X
+ sky130_fd_sc_hd__clkbuf_1_428/X sky130_fd_sc_hd__buf_2_170/X sky130_fd_sc_hd__nand4_1_61/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_259 sky130_fd_sc_hd__nor2_2_4/Y sky130_fd_sc_hd__clkbuf_1_377/X
+ sky130_fd_sc_hd__a22oi_1_259/B2 sky130_fd_sc_hd__clkbuf_4_192/X sky130_fd_sc_hd__nand4_1_64/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_501 sky130_fd_sc_hd__o21ai_1_80/A1 sky130_fd_sc_hd__o21ai_1_87/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_501/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_512 sky130_fd_sc_hd__a21oi_1_59/A1 sky130_fd_sc_hd__nor2_1_49/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_512/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_523 sky130_fd_sc_hd__nor2_1_60/B sky130_fd_sc_hd__fa_2_1040/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_523/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_534 sky130_fd_sc_hd__a21oi_1_85/A1 sky130_fd_sc_hd__a21oi_1_90/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_534/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_545 sky130_fd_sc_hd__clkinv_1_545/Y sky130_fd_sc_hd__nor2_1_80/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_545/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_556 sky130_fd_sc_hd__nand4_1_85/D sky130_fd_sc_hd__fa_2_970/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_556/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_567 sky130_fd_sc_hd__o21ai_1_133/A2 sky130_fd_sc_hd__a21o_2_3/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_567/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_578 sky130_fd_sc_hd__o21ai_1_147/A2 sky130_fd_sc_hd__fa_2_999/A
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_589 sky130_fd_sc_hd__nor2_2_8/B sky130_fd_sc_hd__nor2_4_10/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_589/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_4_14 sky130_fd_sc_hd__clkinv_8_17/Y sky130_fd_sc_hd__clkinv_4_14/Y
+ VSS VDD VDD VSS VSS sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_70 sky130_fd_sc_hd__nor2_1_70/B sky130_fd_sc_hd__o21a_1_7/A1
+ sky130_fd_sc_hd__nor2_1_70/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_25 sky130_fd_sc_hd__clkinv_4_26/A sky130_fd_sc_hd__clkinv_4_25/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_25/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_81 sky130_fd_sc_hd__nor2_1_81/B sky130_fd_sc_hd__nor2_1_81/Y
+ sky130_fd_sc_hd__nor2_1_81/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_36 sky130_fd_sc_hd__clkinv_4_36/A sky130_fd_sc_hd__dfxtp_1_91/D
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_36/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_92 sky130_fd_sc_hd__nor2_1_92/B sky130_fd_sc_hd__nor2_1_92/Y
+ sky130_fd_sc_hd__nor2_1_92/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_47 sky130_fd_sc_hd__clkinv_4_49/A sky130_fd_sc_hd__clkinv_4_48/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_47/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_58 sky130_fd_sc_hd__clkinv_8_71/A sky130_fd_sc_hd__clkinv_4_59/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_58/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_69 sky130_fd_sc_hd__clkinv_4_69/A sky130_fd_sc_hd__clkinv_4_69/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_69/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_sram_2kbyte_1rw1r_32x512_8_0 sky130_fd_sc_hd__buf_6_1/X sky130_fd_sc_hd__clkbuf_4_0/X
+ sky130_fd_sc_hd__buf_4_2/X sky130_fd_sc_hd__buf_4_3/X sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__buf_6_4/X sky130_fd_sc_hd__buf_4_7/X sky130_fd_sc_hd__buf_6_6/X
+ sky130_fd_sc_hd__clkbuf_4_1/X sky130_fd_sc_hd__buf_4_8/X sky130_fd_sc_hd__buf_4_9/X
+ sky130_fd_sc_hd__clkbuf_4_5/X sky130_fd_sc_hd__clkbuf_4_6/X sky130_fd_sc_hd__buf_4_11/X
+ sky130_fd_sc_hd__buf_12_0/X sky130_fd_sc_hd__buf_6_9/X sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__clkbuf_4_0/X sky130_fd_sc_hd__buf_4_2/X sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__buf_4_5/X sky130_fd_sc_hd__buf_6_4/X sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__buf_6_6/X sky130_fd_sc_hd__clkbuf_4_1/X sky130_fd_sc_hd__buf_4_8/X
+ sky130_fd_sc_hd__buf_4_9/X sky130_fd_sc_hd__clkbuf_4_5/X sky130_fd_sc_hd__clkbuf_4_6/X
+ sky130_fd_sc_hd__buf_4_11/X sky130_fd_sc_hd__buf_12_0/X sky130_fd_sc_hd__buf_6_9/X
+ sky130_fd_sc_hd__buf_12_35/X sky130_fd_sc_hd__buf_12_48/X sky130_fd_sc_hd__buf_12_53/X
+ sky130_fd_sc_hd__buf_12_52/X sky130_fd_sc_hd__buf_12_33/X sky130_fd_sc_hd__buf_12_89/X
+ sky130_fd_sc_hd__buf_12_84/X sky130_fd_sc_hd__buf_12_50/X sky130_fd_sc_hd__buf_12_49/X
+ sky130_fd_sc_hd__buf_12_74/X sky130_fd_sc_hd__buf_12_110/X sky130_fd_sc_hd__buf_12_93/X
+ sky130_fd_sc_hd__buf_12_15/X sky130_fd_sc_hd__buf_12_106/X sky130_fd_sc_hd__buf_12_62/X
+ sky130_fd_sc_hd__buf_12_109/X sky130_fd_sc_hd__buf_12_72/X sky130_fd_sc_hd__buf_12_6/X
+ sky130_fd_sc_hd__buf_2_24/X sky130_fd_sc_hd__clkbuf_1_91/X sky130_fd_sc_hd__buf_2_24/X
+ sky130_fd_sc_hd__clkinv_8_1/Y sky130_fd_sc_hd__clkinv_8_6/Y sky130_fd_sc_hd__buf_12_114/X
+ sky130_fd_sc_hd__buf_12_44/X sky130_fd_sc_hd__buf_8_60/X sky130_fd_sc_hd__buf_12_41/X
+ sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[0] sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[1]
+ sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[2] sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[3]
+ sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[4] sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[5]
+ sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[6] sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[7]
+ sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[8] sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[9]
+ sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[10] sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[11]
+ sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[12] sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[13]
+ sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[14] sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[15]
+ sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[16] sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[17]
+ sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[18] sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[19]
+ sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[20] sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[21]
+ sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[22] sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[23]
+ sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[24] sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[25]
+ sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[26] sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[27]
+ sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[28] sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[29]
+ sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[30] sky130_sram_2kbyte_1rw1r_32x512_8_0/dout0[31]
+ sky130_fd_sc_hd__clkbuf_1_55/A sky130_fd_sc_hd__clkbuf_1_56/A sky130_fd_sc_hd__clkbuf_1_57/A
+ sky130_fd_sc_hd__clkbuf_1_58/A sky130_fd_sc_hd__clkbuf_1_59/A sky130_fd_sc_hd__clkbuf_1_60/A
+ sky130_fd_sc_hd__clkbuf_1_61/A sky130_fd_sc_hd__clkbuf_1_62/A sky130_fd_sc_hd__clkbuf_1_63/A
+ sky130_fd_sc_hd__clkbuf_1_64/A sky130_fd_sc_hd__clkbuf_1_65/A sky130_fd_sc_hd__clkbuf_1_66/A
+ sky130_fd_sc_hd__clkbuf_1_67/A sky130_fd_sc_hd__clkbuf_1_68/A sky130_fd_sc_hd__clkbuf_1_69/A
+ sky130_fd_sc_hd__clkbuf_1_70/A sky130_fd_sc_hd__a22oi_1_83/A2 sky130_fd_sc_hd__a22oi_1_79/A2
+ sky130_fd_sc_hd__a22oi_1_75/A2 sky130_fd_sc_hd__a22oi_1_71/A2 sky130_fd_sc_hd__a22oi_1_67/A2
+ sky130_fd_sc_hd__a22oi_2_11/A2 sky130_fd_sc_hd__a22oi_2_10/A2 sky130_fd_sc_hd__a22oi_2_9/A2
+ sky130_fd_sc_hd__a22oi_2_8/A2 sky130_fd_sc_hd__a22oi_2_7/A2 sky130_fd_sc_hd__a22oi_2_6/A2
+ sky130_fd_sc_hd__a22oi_2_5/A2 sky130_fd_sc_hd__a22oi_1_42/A2 sky130_fd_sc_hd__a22oi_1_38/A2
+ sky130_fd_sc_hd__a22oi_1_34/A2 sky130_fd_sc_hd__a22oi_2_4/A2 VDD VSS sky130_sram_2kbyte_1rw1r_32x512_8
Xsky130_fd_sc_hd__a21oi_1_420 sky130_fd_sc_hd__or2_0_11/B sky130_fd_sc_hd__nor3_1_40/C
+ sky130_fd_sc_hd__o21bai_1_4/A2 sky130_fd_sc_hd__nor3_1_40/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_431 sky130_fd_sc_hd__o21a_1_65/B1 sky130_fd_sc_hd__o21a_1_64/A1
+ sky130_fd_sc_hd__a21oi_1_431/Y sky130_fd_sc_hd__o21a_1_68/A2 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_442 sky130_fd_sc_hd__xor2_1_275/X sky130_fd_sc_hd__o21ai_1_449/Y
+ sky130_fd_sc_hd__a21oi_1_442/Y sky130_fd_sc_hd__nand2_1_522/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_453 sky130_fd_sc_hd__nor2_2_18/Y sky130_fd_sc_hd__o21ai_1_462/Y
+ sky130_fd_sc_hd__nor2_1_299/B sky130_fd_sc_hd__fa_2_1291/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_464 sky130_fd_sc_hd__a21oi_1_464/A1 sky130_fd_sc_hd__nor2_1_304/Y
+ sky130_fd_sc_hd__a21oi_1_464/Y sky130_fd_sc_hd__nor2b_2_5/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_475 sky130_fd_sc_hd__nor3_1_41/A sky130_fd_sc_hd__o22ai_1_431/Y
+ sky130_fd_sc_hd__a21oi_1_475/Y sky130_fd_sc_hd__fa_2_1303/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_486 sky130_fd_sc_hd__or2_0_13/B sky130_fd_sc_hd__or2_0_0/B
+ sky130_fd_sc_hd__nand2_1_554/A sky130_fd_sc_hd__nor2_1_322/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_8_100 sky130_fd_sc_hd__clkinv_8_100/Y sky130_fd_sc_hd__clkinv_4_48/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_100/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__a21oi_1_497 sky130_fd_sc_hd__nor2_1_318/Y sky130_fd_sc_hd__or2_0_0/B
+ sky130_fd_sc_hd__nand2_1_565/A sky130_fd_sc_hd__nand2_1_569/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_8_111 sky130_fd_sc_hd__clkinv_8_112/A sky130_fd_sc_hd__clkinv_4_56/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_111/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_122 sky130_fd_sc_hd__clkinv_4_0/A sky130_fd_sc_hd__clkinv_8_122/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_122/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_133 sky130_fd_sc_hd__clkinv_8_134/A sky130_fd_sc_hd__clkinv_4_64/Y
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__o21a_1_2 sky130_fd_sc_hd__o21a_1_2/X sky130_fd_sc_hd__o21a_1_2/A1
+ sky130_fd_sc_hd__o21a_1_2/B1 sky130_fd_sc_hd__fa_2_988/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__nand2_1_480 sky130_fd_sc_hd__nand2_1_480/Y sky130_fd_sc_hd__nor2b_2_4/A
+ sky130_fd_sc_hd__xor2_1_254/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_308 sky130_fd_sc_hd__nor2_4_20/Y sky130_fd_sc_hd__fa_2_1302/B
+ sky130_fd_sc_hd__xor2_1_308/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_491 sky130_fd_sc_hd__nand2_1_491/Y sky130_fd_sc_hd__nand2_1_491/B
+ sky130_fd_sc_hd__o21ai_1_424/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_319 sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__xor2_1_319/X
+ sky130_fd_sc_hd__nor2_8_2/B VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nor2b_1_60 sky130_fd_sc_hd__dfxtp_1_494/Q sky130_fd_sc_hd__nor2b_1_60/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_71 sky130_fd_sc_hd__nand3_1_48/C sky130_fd_sc_hd__nor2b_1_71/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_82 sky130_fd_sc_hd__nor2_1_40/B sky130_fd_sc_hd__nor2b_1_82/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_93 sky130_fd_sc_hd__a32o_1_0/X sky130_fd_sc_hd__nor2b_1_93/Y
+ sky130_fd_sc_hd__buf_2_262/X VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1060 sky130_fd_sc_hd__nor2_1_283/B sky130_fd_sc_hd__fa_2_1297/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1060/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_1 VSS VDD sky130_fd_sc_hd__xnor2_1_1/B sky130_fd_sc_hd__xnor2_1_1/Y
+ sky130_fd_sc_hd__xnor2_1_1/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_1071 sky130_fd_sc_hd__a21oi_1_444/B1 sky130_fd_sc_hd__nand2_1_532/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1071/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1082 sky130_fd_sc_hd__nor2_1_273/B sky130_fd_sc_hd__fa_2_1282/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1082/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1093 sky130_fd_sc_hd__nor2_1_305/A sky130_fd_sc_hd__xor2_1_298/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1093/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_16 VDD VSS sky130_fd_sc_hd__ha_2_109/B sky130_fd_sc_hd__dfxtp_1_29/CLK
+ sky130_fd_sc_hd__nand4_1_34/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_170 sky130_fd_sc_hd__fa_2_171/CIN sky130_fd_sc_hd__or3_1_4/B
+ sky130_fd_sc_hd__fa_2_170/A sky130_fd_sc_hd__fa_2_170/B sky130_fd_sc_hd__maj3_1_30/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_27 VDD VSS sky130_fd_sc_hd__ha_2_115/A sky130_fd_sc_hd__dfxtp_1_29/CLK
+ sky130_fd_sc_hd__nand4_1_45/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_181 sky130_fd_sc_hd__fa_2_183/B sky130_fd_sc_hd__fa_2_181/SUM
+ sky130_fd_sc_hd__ha_2_91/B sky130_fd_sc_hd__fa_2_277/B sky130_fd_sc_hd__fa_2_181/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_38 VDD VSS sky130_fd_sc_hd__fa_2_909/CIN sky130_fd_sc_hd__dfxtp_1_39/CLK
+ sky130_fd_sc_hd__buf_2_290/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_192 sky130_fd_sc_hd__maj3_1_45/B sky130_fd_sc_hd__maj3_1_46/A
+ sky130_fd_sc_hd__fa_2_192/A sky130_fd_sc_hd__fa_2_192/B sky130_fd_sc_hd__fa_2_193/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_49 VDD VSS sky130_fd_sc_hd__ha_2_121/B sky130_fd_sc_hd__dfxtp_1_61/CLK
+ sky130_fd_sc_hd__nand4_1_35/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_4_106 sky130_fd_sc_hd__clkbuf_4_106/X sky130_fd_sc_hd__buf_2_275/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o22ai_1_80 sky130_fd_sc_hd__o22ai_1_89/A1 sky130_fd_sc_hd__o22ai_1_88/B1
+ sky130_fd_sc_hd__o22ai_1_80/Y sky130_fd_sc_hd__xnor2_1_43/Y sky130_fd_sc_hd__o22ai_1_80/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkbuf_4_117 sky130_fd_sc_hd__clkbuf_4_117/X sky130_fd_sc_hd__clkbuf_4_117/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o22ai_1_91 sky130_fd_sc_hd__nor2_1_74/A sky130_fd_sc_hd__nor2_1_77/A
+ sky130_fd_sc_hd__o22ai_1_91/Y sky130_fd_sc_hd__a21oi_1_82/Y sky130_fd_sc_hd__a21oi_1_83/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkbuf_4_128 sky130_fd_sc_hd__clkbuf_4_128/X sky130_fd_sc_hd__clkbuf_4_128/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_139 sky130_fd_sc_hd__nand4_1_46/B sky130_fd_sc_hd__a22oi_1_205/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_4_60 VDD VSS sky130_fd_sc_hd__buf_4_60/X sky130_fd_sc_hd__buf_4_60/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_71 VDD VSS sky130_fd_sc_hd__buf_4_71/X sky130_fd_sc_hd__buf_4_71/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_82 VDD VSS sky130_fd_sc_hd__buf_4_82/X sky130_fd_sc_hd__buf_4_82/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_93 VDD VSS sky130_fd_sc_hd__buf_4_93/X sky130_fd_sc_hd__buf_4_93/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_12_120 sky130_fd_sc_hd__buf_12_3/X sky130_fd_sc_hd__buf_12_120/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_131 sky130_fd_sc_hd__buf_12_131/A sky130_fd_sc_hd__buf_12_253/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_142 sky130_fd_sc_hd__inv_2_66/Y sky130_fd_sc_hd__buf_12_142/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_153 sky130_fd_sc_hd__buf_12_153/A sky130_fd_sc_hd__buf_12_153/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_164 sky130_fd_sc_hd__buf_12_164/A sky130_fd_sc_hd__buf_12_237/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_4_1 sky130_fd_sc_hd__clkbuf_4_1/X sky130_fd_sc_hd__buf_2_5/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_12_175 sky130_fd_sc_hd__buf_8_89/X sky130_fd_sc_hd__buf_12_239/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_186 sky130_fd_sc_hd__buf_8_97/X sky130_fd_sc_hd__buf_6_30/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_197 sky130_fd_sc_hd__buf_4_51/X sky130_fd_sc_hd__buf_12_197/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_320 sky130_fd_sc_hd__fa_2_425/A sky130_fd_sc_hd__ha_2_109/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_320/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_331 sky130_fd_sc_hd__fa_2_555/A sky130_fd_sc_hd__ha_2_123/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_331/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_342 sky130_fd_sc_hd__fa_2_698/A sky130_fd_sc_hd__fa_2_699/A
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_353 sky130_fd_sc_hd__ha_2_130/B sky130_fd_sc_hd__ha_2_135/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_353/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_364 sky130_fd_sc_hd__ha_2_141/B sky130_fd_sc_hd__fa_2_812/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_364/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_375 sky130_fd_sc_hd__fa_2_873/B sky130_fd_sc_hd__dfxtp_1_273/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_375/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_386 sky130_fd_sc_hd__fa_2_886/B sky130_fd_sc_hd__nor4_1_4/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_386/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_397 sky130_fd_sc_hd__nand2_1_202/B sky130_fd_sc_hd__nand2_1_34/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_397/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21a_1_16 sky130_fd_sc_hd__o21a_1_16/X sky130_fd_sc_hd__o21a_1_16/A1
+ sky130_fd_sc_hd__o21a_1_16/B1 sky130_fd_sc_hd__o21a_1_16/A2 VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_27 sky130_fd_sc_hd__o21a_1_27/X sky130_fd_sc_hd__o21a_1_27/A1
+ sky130_fd_sc_hd__o21a_1_27/B1 sky130_fd_sc_hd__fa_2_1148/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_38 sky130_fd_sc_hd__o21a_1_38/X sky130_fd_sc_hd__o21a_1_38/A1
+ sky130_fd_sc_hd__o21a_1_38/B1 sky130_fd_sc_hd__fa_2_1203/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_49 sky130_fd_sc_hd__o21a_1_49/X sky130_fd_sc_hd__o21a_1_49/A1
+ sky130_fd_sc_hd__xnor2_1_98/B sky130_fd_sc_hd__fa_2_1258/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__a21oi_1_250 sky130_fd_sc_hd__o21a_1_25/B1 sky130_fd_sc_hd__o21a_1_24/A1
+ sky130_fd_sc_hd__dfxtp_1_889/D sky130_fd_sc_hd__nor2_1_151/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_261 sky130_fd_sc_hd__nor2_2_15/Y sky130_fd_sc_hd__o21ai_1_286/Y
+ sky130_fd_sc_hd__nor2_1_165/B sky130_fd_sc_hd__fa_2_1127/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_272 sky130_fd_sc_hd__or2_0_9/B sky130_fd_sc_hd__o21ai_1_299/Y
+ sky130_fd_sc_hd__a21oi_1_272/Y sky130_fd_sc_hd__clkinv_1_822/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_283 sky130_fd_sc_hd__fa_2_1148/A sky130_fd_sc_hd__o22ai_1_253/Y
+ sky130_fd_sc_hd__a21oi_1_283/Y sky130_fd_sc_hd__nor3_1_38/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_4_1 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkinv_4_1/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_1/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__a21oi_1_294 sky130_fd_sc_hd__fa_2_1148/A sky130_fd_sc_hd__o22ai_1_258/Y
+ sky130_fd_sc_hd__a21oi_1_294/Y sky130_fd_sc_hd__nor2_2_15/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_202 sky130_fd_sc_hd__buf_8_202/A sky130_fd_sc_hd__buf_8_202/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_213 sky130_fd_sc_hd__buf_8_213/A sky130_fd_sc_hd__buf_8_213/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xor2_1_105 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1052/B
+ sky130_fd_sc_hd__xor2_1_105/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_116 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1090/B
+ sky130_fd_sc_hd__xor2_1_116/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_127 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1079/B
+ sky130_fd_sc_hd__xor2_1_127/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_138 sky130_fd_sc_hd__xor2_1_138/B sky130_fd_sc_hd__xor2_1_138/X
+ sky130_fd_sc_hd__xor2_1_139/X VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_149 sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__fa_2_1134/B
+ sky130_fd_sc_hd__xor2_1_149/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_109 VSS VDD sky130_fd_sc_hd__buf_8_35/A sky130_fd_sc_hd__buf_12_90/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_1407 VDD VSS sky130_fd_sc_hd__mux2_2_227/A1 sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__o22ai_1_382/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1418 VDD VSS sky130_fd_sc_hd__mux2_2_256/A0 sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__dfxtp_1_433/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1429 VDD VSS sky130_fd_sc_hd__mux2_2_248/A0 sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__o22ai_1_404/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_107 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_107/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__xnor2_1_10/Y sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_15 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__nor3_2_2/B
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_118 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_118/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_838/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_26 sky130_fd_sc_hd__inv_2_15/A sky130_fd_sc_hd__ha_2_28/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_26/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_129 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_129/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_854/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_37 sky130_fd_sc_hd__inv_2_26/A sky130_fd_sc_hd__buf_2_14/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_37/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_48 sky130_fd_sc_hd__inv_2_37/A sky130_fd_sc_hd__buf_2_13/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_48/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_59 sky130_fd_sc_hd__inv_2_8/A sky130_fd_sc_hd__dfxtp_1_138/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_59/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_2 sky130_fd_sc_hd__xnor2_1_0/A sky130_fd_sc_hd__fa_2_2/SUM
+ sky130_fd_sc_hd__fa_2_2/A sky130_fd_sc_hd__fa_2_2/B sky130_fd_sc_hd__fa_2_2/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_200 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_200/A sky130_fd_sc_hd__ha_2_199/A
+ sky130_fd_sc_hd__ha_2_200/SUM sky130_fd_sc_hd__ha_2_200/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_906 sky130_fd_sc_hd__fa_2_896/A sky130_fd_sc_hd__fa_2_897/B
+ sky130_fd_sc_hd__fa_2_906/A sky130_fd_sc_hd__fa_2_906/B sky130_fd_sc_hd__fa_2_906/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_917 sky130_fd_sc_hd__fa_2_916/CIN sky130_fd_sc_hd__fa_2_917/SUM
+ sky130_fd_sc_hd__fa_2_917/A sky130_fd_sc_hd__fa_2_917/B sky130_fd_sc_hd__fa_2_917/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_928 sky130_fd_sc_hd__fa_2_927/CIN sky130_fd_sc_hd__fa_2_928/SUM
+ sky130_fd_sc_hd__fa_2_928/A sky130_fd_sc_hd__fa_2_928/B sky130_fd_sc_hd__fa_2_928/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_939 sky130_fd_sc_hd__fa_2_919/A sky130_fd_sc_hd__fa_2_920/B
+ sky130_fd_sc_hd__fa_2_939/A sky130_fd_sc_hd__fa_2_939/B sky130_fd_sc_hd__ha_2_124/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a211o_1_30 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_313/A sky130_fd_sc_hd__o21ai_1_456/Y
+ sky130_fd_sc_hd__nor2_1_292/Y sky130_fd_sc_hd__nor2b_2_5/Y sky130_fd_sc_hd__o22ai_1_412/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__mux2_2_206 VSS VDD sky130_fd_sc_hd__mux2_2_206/A1 sky130_fd_sc_hd__mux2_2_206/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_206/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_217 VSS VDD sky130_fd_sc_hd__mux2_2_217/A1 sky130_fd_sc_hd__mux2_2_217/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_217/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_228 VSS VDD sky130_fd_sc_hd__mux2_2_228/A1 sky130_fd_sc_hd__mux2_2_228/A0
+ sky130_fd_sc_hd__nor2_8_2/A sky130_fd_sc_hd__mux2_2_228/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_239 VSS VDD sky130_fd_sc_hd__mux2_2_239/A1 sky130_fd_sc_hd__mux2_2_239/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_239/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__clkinv_1_150 sky130_fd_sc_hd__buf_8_117/A sky130_fd_sc_hd__clkinv_1_150/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_150/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_161 sky130_fd_sc_hd__inv_2_92/A sky130_fd_sc_hd__inv_2_82/Y
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_172 sky130_fd_sc_hd__inv_2_101/A sky130_fd_sc_hd__inv_2_97/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_172/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_4 sky130_fd_sc_hd__buf_8_4/A sky130_fd_sc_hd__buf_8_4/X VSS
+ VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__a22o_1_6 sky130_fd_sc_hd__buf_2_291/X sky130_fd_sc_hd__nor2_1_1/Y
+ sky130_fd_sc_hd__a22o_1_6/X sky130_fd_sc_hd__a22o_1_6/B2 sky130_fd_sc_hd__nor2_1_0/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_183 sky130_fd_sc_hd__a22o_2_6/B1 sky130_fd_sc_hd__nor2_4_4/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_183/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_194 sky130_fd_sc_hd__nand3_2_8/B sky130_fd_sc_hd__a22o_1_28/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_194/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_30 sky130_fd_sc_hd__or2_1_1/B sky130_fd_sc_hd__ha_2_83/A
+ sky130_fd_sc_hd__a22o_1_30/X sky130_fd_sc_hd__a22o_1_30/B2 sky130_fd_sc_hd__a22o_4_0/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_41 sky130_fd_sc_hd__a22o_1_41/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_41/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__fa_2_947/SUM
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_52 sky130_fd_sc_hd__a22o_1_52/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_52/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__nor4_1_10/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_63 sky130_fd_sc_hd__a22o_1_63/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_63/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__nor4_1_12/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_74 sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__fa_2_1071/A
+ sky130_fd_sc_hd__a22o_1_74/X sky130_fd_sc_hd__fa_2_1073/A sky130_fd_sc_hd__nor2_2_12/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__nand4_1_2 sky130_fd_sc_hd__nand4_1_2/C sky130_fd_sc_hd__nand4_1_2/B
+ sky130_fd_sc_hd__nand4_1_2/Y sky130_fd_sc_hd__nand4_1_2/D sky130_fd_sc_hd__nand4_1_2/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__o21ai_1_108 VSS VDD sky130_fd_sc_hd__nor2_1_77/A sky130_fd_sc_hd__nor2_1_80/Y
+ sky130_fd_sc_hd__a21oi_1_91/Y sky130_fd_sc_hd__xor2_1_73/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_119 VSS VDD sky130_fd_sc_hd__o22ai_1_130/B1 sky130_fd_sc_hd__nand4_1_85/C
+ sky130_fd_sc_hd__a21oi_1_104/Y sky130_fd_sc_hd__o21ai_1_119/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__maj3_1_14 sky130_fd_sc_hd__maj3_1_15/X sky130_fd_sc_hd__maj3_1_14/X
+ sky130_fd_sc_hd__maj3_1_14/B sky130_fd_sc_hd__maj3_1_14/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_25 sky130_fd_sc_hd__maj3_1_26/X sky130_fd_sc_hd__maj3_1_25/X
+ sky130_fd_sc_hd__maj3_1_25/B sky130_fd_sc_hd__maj3_1_25/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_404 sky130_fd_sc_hd__nand2_1_516/Y sky130_fd_sc_hd__nand2_1_515/Y
+ sky130_fd_sc_hd__o22ai_1_404/Y sky130_fd_sc_hd__nand2_1_528/B sky130_fd_sc_hd__o21ai_1_444/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_36 sky130_fd_sc_hd__maj3_1_37/X sky130_fd_sc_hd__maj3_1_36/X
+ sky130_fd_sc_hd__maj3_1_36/B sky130_fd_sc_hd__maj3_1_36/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_415 sky130_fd_sc_hd__nor2_1_310/A sky130_fd_sc_hd__nor2_1_299/A
+ sky130_fd_sc_hd__o22ai_1_415/Y sky130_fd_sc_hd__o22ai_1_415/A1 sky130_fd_sc_hd__nor2_1_302/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_47 sky130_fd_sc_hd__maj3_1_48/X sky130_fd_sc_hd__maj3_1_47/X
+ sky130_fd_sc_hd__maj3_1_47/B sky130_fd_sc_hd__maj3_1_47/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_426 sky130_fd_sc_hd__nor2_1_310/A sky130_fd_sc_hd__nor2_1_299/A
+ sky130_fd_sc_hd__o22ai_1_426/Y sky130_fd_sc_hd__a21oi_1_470/Y sky130_fd_sc_hd__nor2_1_310/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_58 sky130_fd_sc_hd__maj3_1_59/X sky130_fd_sc_hd__maj3_1_58/X
+ sky130_fd_sc_hd__maj3_1_58/B sky130_fd_sc_hd__maj3_1_58/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_437 sky130_fd_sc_hd__a31oi_1_4/Y sky130_fd_sc_hd__nor4_1_13/B
+ sky130_fd_sc_hd__nor2_2_19/B sky130_fd_sc_hd__o22ai_1_437/A1 sky130_fd_sc_hd__a31oi_1_3/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_69 sky130_fd_sc_hd__maj3_1_70/X sky130_fd_sc_hd__maj3_1_69/X
+ sky130_fd_sc_hd__maj3_1_69/B sky130_fd_sc_hd__maj3_1_69/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_20 sky130_fd_sc_hd__nor2_2_0/B sky130_fd_sc_hd__nor3_1_0/A
+ sky130_fd_sc_hd__nor4_1_0/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_31 sky130_fd_sc_hd__nand2_1_31/Y sky130_fd_sc_hd__or4_1_0/D
+ sky130_fd_sc_hd__o21ai_1_14/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_42 sky130_fd_sc_hd__nand2_1_42/Y sky130_fd_sc_hd__nand2_1_42/B
+ sky130_fd_sc_hd__a21oi_2_0/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_53 sky130_fd_sc_hd__nand2_1_53/Y sky130_fd_sc_hd__nand2_1_1/B
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_64 sky130_fd_sc_hd__nand2_1_64/Y sky130_fd_sc_hd__nand2_1_65/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_75 sky130_fd_sc_hd__nand2_1_75/Y sky130_fd_sc_hd__nand4_1_67/Y
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_86 sky130_fd_sc_hd__nand2_1_86/Y sky130_fd_sc_hd__nand2_1_87/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_97 sky130_fd_sc_hd__nand2_1_97/Y sky130_fd_sc_hd__buf_2_266/X
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_308 VDD VSS sky130_fd_sc_hd__a22o_1_41/A1 sky130_fd_sc_hd__dfxtp_1_313/CLK
+ sky130_fd_sc_hd__and2_0_90/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_319 VDD VSS sky130_fd_sc_hd__or4_1_1/C sky130_fd_sc_hd__dfxtp_1_325/CLK
+ sky130_fd_sc_hd__and2_0_197/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_16 sky130_fd_sc_hd__fa_2_8/CIN sky130_fd_sc_hd__fa_2_16/SUM
+ sky130_fd_sc_hd__fa_2_16/A sky130_fd_sc_hd__fa_2_16/B sky130_fd_sc_hd__fa_2_16/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_27 sky130_fd_sc_hd__fa_2_26/CIN sky130_fd_sc_hd__or3_1_5/A
+ sky130_fd_sc_hd__fa_2_27/A sky130_fd_sc_hd__fa_2_27/B sky130_fd_sc_hd__fa_2_27/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_38 sky130_fd_sc_hd__maj3_1_23/B sky130_fd_sc_hd__maj3_1_24/A
+ sky130_fd_sc_hd__fa_2_38/A sky130_fd_sc_hd__fa_2_38/B sky130_fd_sc_hd__fa_2_39/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_49 sky130_fd_sc_hd__fa_2_51/CIN sky130_fd_sc_hd__fa_2_47/A
+ sky130_fd_sc_hd__ha_2_96/B sky130_fd_sc_hd__fa_2_49/B sky130_fd_sc_hd__fa_2_49/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_208 VDD VSS sky130_fd_sc_hd__buf_2_208/X sky130_fd_sc_hd__buf_2_208/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_219 VDD VSS sky130_fd_sc_hd__buf_2_219/X sky130_fd_sc_hd__buf_2_219/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_sram_2kbyte_1rw1r_32x512_8_12 sky130_fd_sc_hd__buf_6_49/X sky130_fd_sc_hd__buf_6_50/X
+ sky130_fd_sc_hd__buf_2_140/A sky130_fd_sc_hd__buf_6_51/X sky130_fd_sc_hd__buf_2_144/A
+ sky130_fd_sc_hd__buf_2_146/A sky130_fd_sc_hd__buf_2_147/A sky130_fd_sc_hd__buf_2_148/A
+ sky130_fd_sc_hd__buf_2_149/A sky130_fd_sc_hd__buf_6_52/X sky130_fd_sc_hd__buf_6_53/X
+ sky130_fd_sc_hd__buf_6_55/X sky130_fd_sc_hd__buf_2_153/A sky130_fd_sc_hd__buf_6_56/X
+ sky130_fd_sc_hd__buf_6_57/X sky130_fd_sc_hd__buf_2_156/A sky130_fd_sc_hd__buf_6_49/X
+ sky130_fd_sc_hd__buf_6_50/X sky130_fd_sc_hd__buf_2_140/A sky130_fd_sc_hd__buf_6_51/X
+ sky130_fd_sc_hd__buf_2_144/A sky130_fd_sc_hd__buf_2_146/A sky130_fd_sc_hd__buf_2_147/A
+ sky130_fd_sc_hd__clkbuf_8_3/X sky130_fd_sc_hd__buf_2_149/A sky130_fd_sc_hd__buf_6_52/X
+ sky130_fd_sc_hd__buf_6_53/X sky130_fd_sc_hd__buf_6_55/X sky130_fd_sc_hd__buf_2_153/A
+ sky130_fd_sc_hd__buf_6_56/X sky130_fd_sc_hd__buf_6_57/X sky130_fd_sc_hd__buf_2_156/A
+ sky130_fd_sc_hd__buf_12_420/X sky130_fd_sc_hd__buf_12_454/X sky130_fd_sc_hd__buf_12_409/X
+ sky130_fd_sc_hd__buf_12_449/X sky130_fd_sc_hd__buf_12_381/X sky130_fd_sc_hd__buf_12_502/X
+ sky130_fd_sc_hd__buf_12_498/X sky130_fd_sc_hd__buf_12_458/X sky130_fd_sc_hd__buf_12_517/X
+ sky130_fd_sc_hd__buf_12_415/X sky130_fd_sc_hd__buf_12_504/X sky130_fd_sc_hd__buf_12_393/X
+ sky130_fd_sc_hd__buf_12_497/X sky130_fd_sc_hd__buf_12_468/X sky130_fd_sc_hd__buf_12_481/X
+ sky130_fd_sc_hd__buf_12_488/X sky130_fd_sc_hd__buf_12_442/X sky130_fd_sc_hd__buf_12_509/X
+ sky130_fd_sc_hd__clkbuf_1_519/X sky130_fd_sc_hd__clkbuf_1_375/X sky130_fd_sc_hd__nand3_2_5/Y
+ sky130_fd_sc_hd__clkinv_8_38/Y sky130_fd_sc_hd__dfxtp_1_83/CLK sky130_fd_sc_hd__buf_12_460/X
+ sky130_fd_sc_hd__buf_12_421/X sky130_fd_sc_hd__buf_12_440/X sky130_fd_sc_hd__buf_12_518/X
+ sky130_fd_sc_hd__clkbuf_1_490/A sky130_fd_sc_hd__clkbuf_1_492/A sky130_fd_sc_hd__a22oi_2_29/B2
+ sky130_fd_sc_hd__clkbuf_1_494/A sky130_fd_sc_hd__clkbuf_1_496/A sky130_fd_sc_hd__clkbuf_1_498/A
+ sky130_fd_sc_hd__clkbuf_1_497/A sky130_fd_sc_hd__clkbuf_1_493/A sky130_fd_sc_hd__clkbuf_1_495/A
+ sky130_fd_sc_hd__a22oi_1_229/B2 sky130_fd_sc_hd__a22oi_1_226/B2 sky130_fd_sc_hd__a22oi_1_222/B2
+ sky130_fd_sc_hd__a22oi_2_18/B2 sky130_fd_sc_hd__a22oi_2_16/B2 sky130_fd_sc_hd__a22oi_1_215/B2
+ sky130_fd_sc_hd__a22oi_1_212/B2 sky130_fd_sc_hd__buf_2_223/A sky130_fd_sc_hd__clkbuf_1_455/A
+ sky130_fd_sc_hd__buf_2_224/A sky130_fd_sc_hd__clkbuf_1_534/A sky130_fd_sc_hd__buf_2_226/A
+ sky130_fd_sc_hd__buf_2_227/A sky130_fd_sc_hd__buf_2_228/A sky130_fd_sc_hd__buf_2_229/A
+ sky130_fd_sc_hd__buf_2_230/A sky130_fd_sc_hd__buf_2_231/A sky130_fd_sc_hd__clkbuf_1_456/A
+ sky130_fd_sc_hd__clkbuf_1_457/A sky130_fd_sc_hd__buf_2_232/A sky130_fd_sc_hd__clkbuf_1_533/A
+ sky130_fd_sc_hd__buf_2_234/A sky130_fd_sc_hd__buf_2_235/A sky130_fd_sc_hd__a22oi_1_319/B2
+ sky130_fd_sc_hd__a22oi_1_315/B2 sky130_fd_sc_hd__a22oi_1_311/B2 sky130_fd_sc_hd__a22oi_1_307/B2
+ sky130_fd_sc_hd__a22oi_1_303/B2 sky130_fd_sc_hd__a22oi_1_299/B2 sky130_fd_sc_hd__a22oi_1_295/B2
+ sky130_fd_sc_hd__a22oi_1_291/B2 sky130_fd_sc_hd__a22oi_1_287/B2 sky130_fd_sc_hd__a22oi_1_283/B2
+ sky130_fd_sc_hd__a22oi_1_279/B2 sky130_fd_sc_hd__a22oi_1_275/B2 sky130_fd_sc_hd__a22oi_1_271/B2
+ sky130_fd_sc_hd__a22oi_1_267/B2 sky130_fd_sc_hd__a22oi_1_263/B2 sky130_fd_sc_hd__a22oi_1_259/B2
+ sky130_fd_sc_hd__clkbuf_1_458/A sky130_fd_sc_hd__clkbuf_1_459/A sky130_fd_sc_hd__clkbuf_1_460/A
+ sky130_fd_sc_hd__clkbuf_1_523/A sky130_fd_sc_hd__clkbuf_1_525/A sky130_fd_sc_hd__clkbuf_1_463/A
+ sky130_fd_sc_hd__clkbuf_1_464/A sky130_fd_sc_hd__clkbuf_1_465/A sky130_fd_sc_hd__clkbuf_1_466/A
+ sky130_fd_sc_hd__clkbuf_1_467/A sky130_fd_sc_hd__clkbuf_1_468/A sky130_fd_sc_hd__clkbuf_1_469/A
+ sky130_fd_sc_hd__clkbuf_1_470/A sky130_fd_sc_hd__clkbuf_1_471/A sky130_fd_sc_hd__clkbuf_1_472/A
+ sky130_fd_sc_hd__clkbuf_1_473/A VDD VSS sky130_sram_2kbyte_1rw1r_32x512_8
Xsky130_fd_sc_hd__dfxtp_1_1204 VDD VSS sky130_fd_sc_hd__fa_2_1253/A sky130_fd_sc_hd__clkinv_8_75/Y
+ sky130_fd_sc_hd__mux2_2_186/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1215 VDD VSS sky130_fd_sc_hd__fa_2_1227/A sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__mux2_2_210/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1226 VDD VSS sky130_fd_sc_hd__fa_2_1238/A sky130_fd_sc_hd__clkinv_8_116/Y
+ sky130_fd_sc_hd__mux2_2_181/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1237 VDD VSS sky130_fd_sc_hd__fa_2_1266/A sky130_fd_sc_hd__clkinv_8_65/Y
+ sky130_fd_sc_hd__mux2_2_211/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1248 VDD VSS sky130_fd_sc_hd__o32ai_1_8/A1 sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__nor2b_1_123/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_820 VDD VSS sky130_fd_sc_hd__fa_2_1094/A sky130_fd_sc_hd__clkinv_8_59/Y
+ sky130_fd_sc_hd__and2_0_296/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1259 VDD VSS sky130_fd_sc_hd__mux2_2_195/A0 sky130_fd_sc_hd__clkinv_8_78/Y
+ sky130_fd_sc_hd__o22ai_1_332/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_831 VDD VSS sky130_fd_sc_hd__fa_2_1105/A sky130_fd_sc_hd__clkinv_4_26/Y
+ sky130_fd_sc_hd__or2_0_7/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_842 VDD VSS sky130_fd_sc_hd__mux2_2_71/A0 sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__o21ai_1_159/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_853 VDD VSS sky130_fd_sc_hd__mux2_2_47/A1 sky130_fd_sc_hd__clkinv_4_25/Y
+ sky130_fd_sc_hd__o21ai_1_170/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_864 VDD VSS sky130_fd_sc_hd__mux2_2_64/A1 sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__o21ai_1_178/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_875 VDD VSS sky130_fd_sc_hd__mux2_2_42/A1 sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__o21ai_1_189/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_886 VDD VSS sky130_fd_sc_hd__fa_2_856/A sky130_fd_sc_hd__dfxtp_1_902/CLK
+ sky130_fd_sc_hd__o21a_1_26/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_897 VDD VSS sky130_fd_sc_hd__fa_2_932/B sky130_fd_sc_hd__dfxtp_1_899/CLK
+ sky130_fd_sc_hd__o21a_1_22/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_440 VSS VDD sky130_fd_sc_hd__clkbuf_1_440/X sky130_fd_sc_hd__clkbuf_1_440/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_451 VSS VDD sky130_fd_sc_hd__a22oi_2_18/A2 sky130_fd_sc_hd__clkbuf_1_451/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_462 VSS VDD sky130_fd_sc_hd__clkbuf_1_462/X sky130_fd_sc_hd__clkbuf_1_525/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_473 VSS VDD sky130_fd_sc_hd__clkbuf_1_473/X sky130_fd_sc_hd__clkbuf_1_473/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_484 VSS VDD sky130_fd_sc_hd__clkbuf_1_484/X sky130_fd_sc_hd__nand3_2_6/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_495 VSS VDD sky130_fd_sc_hd__a22oi_2_21/B2 sky130_fd_sc_hd__clkbuf_1_495/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_703 sky130_fd_sc_hd__fa_2_702/CIN sky130_fd_sc_hd__fa_2_703/SUM
+ sky130_fd_sc_hd__fa_2_703/A sky130_fd_sc_hd__fa_2_703/B sky130_fd_sc_hd__fa_2_703/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_714 sky130_fd_sc_hd__fa_2_713/CIN sky130_fd_sc_hd__fa_2_714/SUM
+ sky130_fd_sc_hd__fa_2_714/A sky130_fd_sc_hd__fa_2_714/B sky130_fd_sc_hd__fa_2_714/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_725 sky130_fd_sc_hd__fa_2_726/B sky130_fd_sc_hd__fa_2_725/SUM
+ sky130_fd_sc_hd__fa_2_823/B sky130_fd_sc_hd__ha_2_138/A sky130_fd_sc_hd__fa_2_725/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_736 sky130_fd_sc_hd__fa_2_738/B sky130_fd_sc_hd__fa_2_736/SUM
+ sky130_fd_sc_hd__fa_2_736/A sky130_fd_sc_hd__fa_2_736/B sky130_fd_sc_hd__fa_2_736/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_747 sky130_fd_sc_hd__fa_2_749/A sky130_fd_sc_hd__fa_2_744/A
+ sky130_fd_sc_hd__fa_2_826/A sky130_fd_sc_hd__ha_2_142/A sky130_fd_sc_hd__fa_2_817/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_758 sky130_fd_sc_hd__fa_2_759/CIN sky130_fd_sc_hd__fa_2_753/A
+ sky130_fd_sc_hd__fa_2_834/B sky130_fd_sc_hd__fa_2_758/B sky130_fd_sc_hd__ha_2_139/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_769 sky130_fd_sc_hd__fa_2_768/B sky130_fd_sc_hd__fa_2_769/SUM
+ sky130_fd_sc_hd__ha_2_142/B sky130_fd_sc_hd__ha_2_140/B sky130_fd_sc_hd__fa_2_834/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor2b_1_100 sky130_fd_sc_hd__a32o_1_1/X sky130_fd_sc_hd__nor2b_1_100/Y
+ sky130_fd_sc_hd__buf_2_262/X VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_111 sky130_fd_sc_hd__o22ai_1_209/Y sky130_fd_sc_hd__nor2b_1_111/Y
+ sky130_fd_sc_hd__buf_2_262/X VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_122 sky130_fd_sc_hd__nor2_1_243/Y sky130_fd_sc_hd__nor2b_1_122/Y
+ sky130_fd_sc_hd__buf_2_262/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_133 sky130_fd_sc_hd__nor2_1_315/B sky130_fd_sc_hd__nor2b_1_133/Y
+ sky130_fd_sc_hd__nor4_1_13/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__buf_6_1 VDD VSS sky130_fd_sc_hd__buf_6_1/X sky130_fd_sc_hd__buf_6_1/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__bufbuf_8_4 sky130_fd_sc_hd__a22o_1_23/X sky130_fd_sc_hd__buf_6_71/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufbuf_8
Xsky130_fd_sc_hd__buf_6_17 VDD VSS sky130_fd_sc_hd__buf_6_17/X sky130_fd_sc_hd__buf_6_17/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_28 VDD VSS sky130_fd_sc_hd__buf_6_28/X sky130_fd_sc_hd__buf_6_28/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_39 VDD VSS sky130_fd_sc_hd__buf_6_39/X sky130_fd_sc_hd__buf_6_39/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_19 sky130_fd_sc_hd__buf_2_123/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__o22ai_1_201 sky130_fd_sc_hd__nor2_1_126/A sky130_fd_sc_hd__nor2_2_13/B
+ sky130_fd_sc_hd__o22ai_1_201/Y sky130_fd_sc_hd__a21oi_1_234/Y sky130_fd_sc_hd__a211oi_1_8/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_212 sky130_fd_sc_hd__nand2_1_358/Y sky130_fd_sc_hd__nand2_1_357/Y
+ sky130_fd_sc_hd__o22ai_1_212/Y sky130_fd_sc_hd__nand2_1_368/B sky130_fd_sc_hd__o21ai_1_278/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_223 sky130_fd_sc_hd__nand2_1_360/Y sky130_fd_sc_hd__o21ai_1_277/Y
+ sky130_fd_sc_hd__o22ai_1_223/Y sky130_fd_sc_hd__nand2_1_367/B sky130_fd_sc_hd__nand2_1_359/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_234 sky130_fd_sc_hd__nand2_1_360/Y sky130_fd_sc_hd__nand2_1_359/Y
+ sky130_fd_sc_hd__o22ai_1_234/Y sky130_fd_sc_hd__o22ai_1_234/A1 sky130_fd_sc_hd__a21o_2_11/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_245 sky130_fd_sc_hd__o22ai_1_265/A2 sky130_fd_sc_hd__o22ai_1_252/B1
+ sky130_fd_sc_hd__o22ai_1_245/Y sky130_fd_sc_hd__nor2_1_144/B sky130_fd_sc_hd__o22ai_1_261/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_309 sky130_fd_sc_hd__o21a_1_10/B1 sky130_fd_sc_hd__fa_2_1064/A
+ sky130_fd_sc_hd__o21a_1_10/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_908 sky130_fd_sc_hd__nor2_1_191/B sky130_fd_sc_hd__fa_2_1176/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_908/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_256 sky130_fd_sc_hd__o32ai_1_2/A3 sky130_fd_sc_hd__o22ai_1_259/B1
+ sky130_fd_sc_hd__o22ai_1_256/Y sky130_fd_sc_hd__nor2_1_178/A sky130_fd_sc_hd__o21a_1_29/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_1_2 sky130_fd_sc_hd__nor3_1_1/B sky130_fd_sc_hd__nor2_1_2/Y
+ sky130_fd_sc_hd__nor2_1_2/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_1_919 sky130_fd_sc_hd__clkinv_1_919/Y sky130_fd_sc_hd__nand2_1_438/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_919/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_267 sky130_fd_sc_hd__nand2_1_410/Y sky130_fd_sc_hd__o21ai_1_331/Y
+ sky130_fd_sc_hd__o22ai_1_267/Y sky130_fd_sc_hd__nand2_1_419/B sky130_fd_sc_hd__nand2_1_409/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_278 sky130_fd_sc_hd__nand2_1_410/Y sky130_fd_sc_hd__nand2_1_409/Y
+ sky130_fd_sc_hd__o22ai_1_278/Y sky130_fd_sc_hd__o22ai_1_291/A1 sky130_fd_sc_hd__a21o_2_17/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__bufinv_8_4 sky130_fd_sc_hd__bufinv_8_4/A sky130_fd_sc_hd__buf_6_45/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufinv_8
Xsky130_fd_sc_hd__o22ai_1_289 sky130_fd_sc_hd__nand2_1_412/Y sky130_fd_sc_hd__nand2_1_411/Y
+ sky130_fd_sc_hd__o22ai_1_289/Y sky130_fd_sc_hd__o22ai_1_289/A1 sky130_fd_sc_hd__a21o_2_16/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__dfxtp_1_105 VDD VSS sky130_fd_sc_hd__xor2_1_0/B sky130_fd_sc_hd__dfxtp_1_95/CLK
+ sky130_fd_sc_hd__and2_0_4/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_116 VDD VSS sky130_fd_sc_hd__nand2_1_33/A sky130_fd_sc_hd__dfxtp_1_117/CLK
+ sky130_fd_sc_hd__ha_2_0/SUM VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_127 VDD VSS sky130_fd_sc_hd__ha_2_13/A sky130_fd_sc_hd__dfxtp_1_129/CLK
+ sky130_fd_sc_hd__and2_0_16/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_138 VDD VSS sky130_fd_sc_hd__dfxtp_1_138/Q sky130_fd_sc_hd__dfxtp_1_138/CLK
+ sky130_fd_sc_hd__nor2b_1_13/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_149 VDD VSS sky130_fd_sc_hd__ha_2_38/A sky130_fd_sc_hd__dfxtp_1_155/CLK
+ sky130_fd_sc_hd__and2_0_32/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_450 VSS VDD sky130_fd_sc_hd__o22ai_1_415/A1 sky130_fd_sc_hd__nor2_1_309/A
+ sky130_fd_sc_hd__nand2_1_529/Y sky130_fd_sc_hd__xor2_1_300/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_461 VSS VDD sky130_fd_sc_hd__a222oi_1_37/Y sky130_fd_sc_hd__nor2_1_309/A
+ sky130_fd_sc_hd__a22oi_1_397/Y sky130_fd_sc_hd__o21ai_1_461/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_472 VSS VDD sky130_fd_sc_hd__a222oi_1_40/Y sky130_fd_sc_hd__nor2_1_309/A
+ sky130_fd_sc_hd__nand2_1_538/Y sky130_fd_sc_hd__xor2_1_280/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_483 VSS VDD sky130_fd_sc_hd__a222oi_1_41/Y sky130_fd_sc_hd__nor2_1_309/A
+ sky130_fd_sc_hd__a22oi_1_401/Y sky130_fd_sc_hd__o21ai_1_483/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_494 VSS VDD sky130_fd_sc_hd__nand2_1_555/A sky130_fd_sc_hd__o21ai_1_507/A1
+ sky130_fd_sc_hd__nand2_1_555/Y sky130_fd_sc_hd__and2_0_343/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_1204 sky130_fd_sc_hd__fa_2_1205/CIN sky130_fd_sc_hd__mux2_2_134/A0
+ sky130_fd_sc_hd__fa_2_1204/A sky130_fd_sc_hd__fa_2_1204/B sky130_fd_sc_hd__fa_2_1204/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1215 sky130_fd_sc_hd__fa_2_1216/CIN sky130_fd_sc_hd__mux2_2_163/A1
+ sky130_fd_sc_hd__fa_2_1215/A sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__fa_2_1215/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1226 sky130_fd_sc_hd__fa_2_1227/CIN sky130_fd_sc_hd__mux2_2_213/A1
+ sky130_fd_sc_hd__fa_2_1226/A sky130_fd_sc_hd__fa_2_1226/B sky130_fd_sc_hd__fa_2_1226/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1237 sky130_fd_sc_hd__fa_2_1238/CIN sky130_fd_sc_hd__mux2_2_183/A0
+ sky130_fd_sc_hd__fa_2_1237/A sky130_fd_sc_hd__fa_2_1237/B sky130_fd_sc_hd__fa_2_1237/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1248 sky130_fd_sc_hd__fa_2_1249/CIN sky130_fd_sc_hd__mux2_2_200/A1
+ sky130_fd_sc_hd__fa_2_1248/A sky130_fd_sc_hd__fa_2_1248/B sky130_fd_sc_hd__fa_2_1248/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1001 VDD VSS sky130_fd_sc_hd__mux2_2_92/A0 sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__xnor2_1_96/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_1259 sky130_fd_sc_hd__xor2_1_252/B sky130_fd_sc_hd__mux2_2_174/A0
+ sky130_fd_sc_hd__fa_2_1259/A sky130_fd_sc_hd__fa_2_1259/B sky130_fd_sc_hd__fa_2_1259/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o21ai_1_10 VSS VDD sky130_fd_sc_hd__nor2b_1_52/A sky130_fd_sc_hd__or4_1_1/C
+ sky130_fd_sc_hd__nor2_1_23/A sky130_fd_sc_hd__o21ai_1_10/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1012 VDD VSS sky130_fd_sc_hd__mux2_2_88/A0 sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__o22ai_1_227/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_21 VSS VDD sky130_fd_sc_hd__a21oi_2_0/Y sky130_fd_sc_hd__o22ai_1_0/A2
+ sky130_fd_sc_hd__nand2_1_40/Y sky130_fd_sc_hd__o21ai_1_21/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1023 VDD VSS sky130_fd_sc_hd__fa_2_846/A sky130_fd_sc_hd__dfxtp_1_1026/CLK
+ sky130_fd_sc_hd__a21oi_1_314/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_32 VSS VDD sky130_fd_sc_hd__nor3_1_32/C sky130_fd_sc_hd__nor2_1_29/A
+ sky130_fd_sc_hd__o21ai_1_32/B1 sky130_fd_sc_hd__o21ai_1_32/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1034 VDD VSS sky130_fd_sc_hd__xnor2_1_6/B sky130_fd_sc_hd__dfxtp_1_1050/CLK
+ sky130_fd_sc_hd__xnor2_1_95/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_43 VSS VDD sky130_fd_sc_hd__o21ai_1_53/A2 sky130_fd_sc_hd__xnor2_1_40/Y
+ sky130_fd_sc_hd__a21oi_1_31/Y sky130_fd_sc_hd__o21ai_1_43/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1045 VDD VSS sky130_fd_sc_hd__fa_2_911/B sky130_fd_sc_hd__dfxtp_1_1050/CLK
+ sky130_fd_sc_hd__o21a_1_32/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_54 VSS VDD sky130_fd_sc_hd__o21ai_1_71/A2 sky130_fd_sc_hd__nand2_2_3/Y
+ sky130_fd_sc_hd__a21oi_1_42/Y sky130_fd_sc_hd__o21ai_1_54/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1056 VDD VSS sky130_fd_sc_hd__fa_2_1195/A sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__mux2_2_158/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_65 VSS VDD sky130_fd_sc_hd__nand2_2_3/Y sky130_fd_sc_hd__xnor2_1_50/Y
+ sky130_fd_sc_hd__a21oi_1_51/Y sky130_fd_sc_hd__o21ai_1_65/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1067 VDD VSS sky130_fd_sc_hd__fa_2_1206/A sky130_fd_sc_hd__clkinv_8_70/Y
+ sky130_fd_sc_hd__mux2_2_130/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_76 VSS VDD sky130_fd_sc_hd__xnor2_1_52/A sky130_fd_sc_hd__o21ai_1_76/A1
+ sky130_fd_sc_hd__o21ai_1_76/B1 sky130_fd_sc_hd__xnor2_1_54/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1078 VDD VSS sky130_fd_sc_hd__fa_2_1180/A sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__mux2_2_150/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_650 VDD VSS sky130_fd_sc_hd__fa_2_1014/A sky130_fd_sc_hd__clkinv_8_44/Y
+ sky130_fd_sc_hd__mux2_2_4/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_87 VSS VDD sky130_fd_sc_hd__xnor2_1_35/A sky130_fd_sc_hd__nor2_1_56/Y
+ sky130_fd_sc_hd__o21ai_1_87/B1 sky130_fd_sc_hd__xnor2_1_37/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1089 VDD VSS sky130_fd_sc_hd__xor2_1_209/A sky130_fd_sc_hd__clkinv_8_70/Y
+ sky130_fd_sc_hd__mux2_2_125/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_98 VSS VDD sky130_fd_sc_hd__nor2_1_74/A sky130_fd_sc_hd__a21oi_1_99/Y
+ sky130_fd_sc_hd__a21oi_1_85/Y sky130_fd_sc_hd__xor2_1_68/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_661 VDD VSS sky130_fd_sc_hd__fa_2_978/A sky130_fd_sc_hd__clkinv_8_41/Y
+ sky130_fd_sc_hd__mux2_2_33/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_672 VDD VSS sky130_fd_sc_hd__fa_2_989/A sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__mux2_2_9/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_683 VDD VSS sky130_fd_sc_hd__fa_2_1022/A sky130_fd_sc_hd__clkinv_8_59/Y
+ sky130_fd_sc_hd__and2_0_275/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_694 VDD VSS sky130_fd_sc_hd__nor2_2_7/A sky130_fd_sc_hd__clkinv_8_41/Y
+ sky130_fd_sc_hd__nor2b_1_93/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_270 VSS VDD sky130_fd_sc_hd__clkbuf_1_270/X sky130_fd_sc_hd__clkbuf_1_270/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_281 VSS VDD sky130_fd_sc_hd__clkbuf_1_281/X sky130_fd_sc_hd__clkbuf_1_281/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_292 VSS VDD sky130_fd_sc_hd__clkbuf_1_292/X sky130_fd_sc_hd__clkbuf_1_292/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_500 sky130_fd_sc_hd__fa_2_497/B sky130_fd_sc_hd__fa_2_500/SUM
+ sky130_fd_sc_hd__fa_2_546/A sky130_fd_sc_hd__ha_2_125/A sky130_fd_sc_hd__fa_2_537/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_511 sky130_fd_sc_hd__fa_2_512/CIN sky130_fd_sc_hd__fa_2_505/A
+ sky130_fd_sc_hd__fa_2_558/B sky130_fd_sc_hd__fa_2_551/A sky130_fd_sc_hd__fa_2_567/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_522 sky130_fd_sc_hd__fa_2_523/B sky130_fd_sc_hd__fa_2_514/A
+ sky130_fd_sc_hd__fa_2_535/A sky130_fd_sc_hd__fa_2_567/A sky130_fd_sc_hd__fa_2_531/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o2bb2ai_1_18 sky130_fd_sc_hd__dfxtp_1_556/D sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__dfxtp_1_556/Q sky130_fd_sc_hd__nand2_1_210/Y sky130_fd_sc_hd__nand3_1_44/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_533 sky130_fd_sc_hd__maj3_1_87/B sky130_fd_sc_hd__maj3_1_88/A
+ sky130_fd_sc_hd__fa_2_533/A sky130_fd_sc_hd__fa_2_533/B sky130_fd_sc_hd__fa_2_534/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o2bb2ai_1_29 sky130_fd_sc_hd__and2_0_252/A sky130_fd_sc_hd__nand2_1_214/B
+ sky130_fd_sc_hd__nor2_1_33/Y sky130_fd_sc_hd__nor2_1_33/Y sky130_fd_sc_hd__nand2_1_214/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_544 sky130_fd_sc_hd__maj3_1_85/B sky130_fd_sc_hd__maj3_1_86/A
+ sky130_fd_sc_hd__fa_2_544/A sky130_fd_sc_hd__fa_2_544/B sky130_fd_sc_hd__fa_2_545/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_555 sky130_fd_sc_hd__fa_2_557/CIN sky130_fd_sc_hd__fa_2_552/A
+ sky130_fd_sc_hd__fa_2_555/A sky130_fd_sc_hd__fa_2_555/B sky130_fd_sc_hd__fa_2_555/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_566 sky130_fd_sc_hd__fa_2_565/B sky130_fd_sc_hd__fa_2_562/B
+ sky130_fd_sc_hd__fa_2_566/A sky130_fd_sc_hd__fa_2_566/B sky130_fd_sc_hd__fa_2_554/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_577 sky130_fd_sc_hd__fa_2_576/CIN sky130_fd_sc_hd__and2_0_95/A
+ sky130_fd_sc_hd__fa_2_577/A sky130_fd_sc_hd__fa_2_577/B sky130_fd_sc_hd__fa_2_577/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_588 sky130_fd_sc_hd__maj3_1_128/B sky130_fd_sc_hd__maj3_1_129/A
+ sky130_fd_sc_hd__fa_2_588/A sky130_fd_sc_hd__fa_2_588/B sky130_fd_sc_hd__fa_2_589/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_599 sky130_fd_sc_hd__fa_2_601/B sky130_fd_sc_hd__fa_2_599/SUM
+ sky130_fd_sc_hd__fa_2_599/A sky130_fd_sc_hd__fa_2_599/B sky130_fd_sc_hd__fa_2_599/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor2_1_309 sky130_fd_sc_hd__o21a_1_68/A1 sky130_fd_sc_hd__nor2_1_309/Y
+ sky130_fd_sc_hd__nor2_1_309/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__and2_0_290 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_290/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__and2_0_290/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_505 sky130_fd_sc_hd__buf_12_505/A sky130_fd_sc_hd__buf_12_505/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_516 sky130_fd_sc_hd__buf_12_516/A sky130_fd_sc_hd__buf_12_516/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__nand2_1_106 sky130_fd_sc_hd__nand2_1_106/Y sky130_fd_sc_hd__nand2_1_107/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_705 sky130_fd_sc_hd__clkinv_1_705/Y sky130_fd_sc_hd__a21oi_1_206/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_705/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_117 sky130_fd_sc_hd__nand2_1_117/Y sky130_fd_sc_hd__nand2_1_118/Y
+ sky130_fd_sc_hd__buf_2_264/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_716 sky130_fd_sc_hd__nand4_1_86/C sky130_fd_sc_hd__fa_2_1047/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_716/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_128 sky130_fd_sc_hd__nand2_1_128/Y sky130_fd_sc_hd__fa_2_707/SUM
+ sky130_fd_sc_hd__and2_0_235/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_727 sky130_fd_sc_hd__clkinv_1_727/Y sky130_fd_sc_hd__a222oi_1_3/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_727/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_139 sky130_fd_sc_hd__nand2_1_139/Y sky130_fd_sc_hd__nand2_1_140/Y
+ sky130_fd_sc_hd__buf_2_264/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_738 sky130_fd_sc_hd__nor2_1_138/A sky130_fd_sc_hd__fa_2_1086/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_738/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_749 sky130_fd_sc_hd__a22o_1_73/A1 sky130_fd_sc_hd__a22o_1_73/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_749/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_280 VSS VDD sky130_fd_sc_hd__nand2_1_370/B sky130_fd_sc_hd__a21o_2_9/B1
+ sky130_fd_sc_hd__a21o_2_8/A2 sky130_fd_sc_hd__o21ai_1_280/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkinv_8_8 sky130_fd_sc_hd__clkinv_8_8/Y sky130_fd_sc_hd__clkinv_8_8/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__o21ai_1_291 VSS VDD sky130_fd_sc_hd__nor2_1_174/B sky130_fd_sc_hd__nor2_1_182/A
+ sky130_fd_sc_hd__nand2_1_373/Y sky130_fd_sc_hd__xor2_1_168/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor3_1_16 sky130_fd_sc_hd__nor3_1_16/C sky130_fd_sc_hd__nor3_1_16/Y
+ sky130_fd_sc_hd__nor3_2_5/A sky130_fd_sc_hd__nor3_2_6/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_27 sky130_fd_sc_hd__nor3_1_27/C sky130_fd_sc_hd__or2_0_4/A
+ sky130_fd_sc_hd__nor3_1_27/A sky130_fd_sc_hd__nor3_1_27/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_38 sky130_fd_sc_hd__nor3_1_38/C sky130_fd_sc_hd__nor3_1_38/Y
+ sky130_fd_sc_hd__nor3_1_38/A sky130_fd_sc_hd__nor3_1_38/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__fa_2_1001 sky130_fd_sc_hd__fa_2_1002/CIN sky130_fd_sc_hd__mux2_2_32/A1
+ sky130_fd_sc_hd__fa_2_1001/A sky130_fd_sc_hd__xor2_1_75/X sky130_fd_sc_hd__fa_2_1001/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1012 sky130_fd_sc_hd__fa_2_1013/CIN sky130_fd_sc_hd__mux2_2_8/A0
+ sky130_fd_sc_hd__fa_2_1012/A sky130_fd_sc_hd__xor2_1_64/X sky130_fd_sc_hd__fa_2_1012/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1023 sky130_fd_sc_hd__fa_2_1024/CIN sky130_fd_sc_hd__and2_0_280/A
+ sky130_fd_sc_hd__fa_2_1023/A sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_1023/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1034 sky130_fd_sc_hd__fa_2_1035/CIN sky130_fd_sc_hd__fa_2_1034/SUM
+ sky130_fd_sc_hd__nor2_1_57/A sky130_fd_sc_hd__fa_2_1034/B sky130_fd_sc_hd__fa_2_1034/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1045 sky130_fd_sc_hd__fa_2_1045/COUT sky130_fd_sc_hd__a22o_1_67/A2
+ sky130_fd_sc_hd__nor2_2_6/B sky130_fd_sc_hd__fa_2_1045/B sky130_fd_sc_hd__fa_2_1045/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1056 sky130_fd_sc_hd__fa_2_1057/CIN sky130_fd_sc_hd__mux2_2_65/A0
+ sky130_fd_sc_hd__fa_2_1056/A sky130_fd_sc_hd__fa_2_1056/B sky130_fd_sc_hd__fa_2_1056/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1067 sky130_fd_sc_hd__fa_2_1068/CIN sky130_fd_sc_hd__mux2_2_43/A0
+ sky130_fd_sc_hd__fa_2_1067/A sky130_fd_sc_hd__xor2_1_90/X sky130_fd_sc_hd__fa_2_1067/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1078 sky130_fd_sc_hd__fa_2_1079/CIN sky130_fd_sc_hd__mux2_2_67/A1
+ sky130_fd_sc_hd__fa_2_1078/A sky130_fd_sc_hd__fa_2_1078/B sky130_fd_sc_hd__fa_2_1078/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1089 sky130_fd_sc_hd__fa_2_1090/CIN sky130_fd_sc_hd__mux2_2_44/A0
+ sky130_fd_sc_hd__fa_2_1089/A sky130_fd_sc_hd__fa_2_1089/B sky130_fd_sc_hd__fa_2_1089/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_10 sky130_fd_sc_hd__inv_2_10/A sky130_fd_sc_hd__inv_2_10/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_21 sky130_fd_sc_hd__inv_2_21/A sky130_fd_sc_hd__inv_2_21/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_32 sky130_fd_sc_hd__inv_2_32/A sky130_fd_sc_hd__buf_8_5/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_43 sky130_fd_sc_hd__inv_2_43/A sky130_fd_sc_hd__inv_2_43/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_54 sky130_fd_sc_hd__ha_2_37/A sky130_fd_sc_hd__inv_2_54/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_65 sky130_fd_sc_hd__inv_2_65/A sky130_fd_sc_hd__inv_2_65/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_76 sky130_fd_sc_hd__inv_2_76/A sky130_fd_sc_hd__inv_2_78/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_480 VDD VSS sky130_fd_sc_hd__dfxtp_1_480/Q sky130_fd_sc_hd__dfxtp_1_483/CLK
+ sky130_fd_sc_hd__nor2b_1_82/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_2_0 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__nand2_2_0/A
+ sky130_fd_sc_hd__nand2_2_0/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__inv_2_87 sky130_fd_sc_hd__inv_2_87/A sky130_fd_sc_hd__inv_2_87/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_491 VDD VSS sky130_fd_sc_hd__nor2b_1_89/A sky130_fd_sc_hd__dfxtp_1_496/CLK
+ sky130_fd_sc_hd__nor2b_1_66/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_98 sky130_fd_sc_hd__inv_2_98/A sky130_fd_sc_hd__inv_2_98/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__ha_2_19 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_19/A sky130_fd_sc_hd__ha_2_18/B
+ sky130_fd_sc_hd__ha_2_19/SUM sky130_fd_sc_hd__inv_2_3/A sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_330 sky130_fd_sc_hd__fa_2_331/A sky130_fd_sc_hd__fa_2_329/B
+ sky130_fd_sc_hd__ha_2_114/A sky130_fd_sc_hd__fa_2_425/A sky130_fd_sc_hd__fa_2_416/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_341 sky130_fd_sc_hd__fa_2_343/A sky130_fd_sc_hd__fa_2_341/SUM
+ sky130_fd_sc_hd__fa_2_341/A sky130_fd_sc_hd__fa_2_341/B sky130_fd_sc_hd__fa_2_346/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_352 sky130_fd_sc_hd__maj3_1_69/B sky130_fd_sc_hd__maj3_1_70/A
+ sky130_fd_sc_hd__fa_2_352/A sky130_fd_sc_hd__fa_2_352/B sky130_fd_sc_hd__fa_2_353/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_363 sky130_fd_sc_hd__fa_2_366/B sky130_fd_sc_hd__fa_2_363/SUM
+ sky130_fd_sc_hd__fa_2_363/A sky130_fd_sc_hd__fa_2_363/B sky130_fd_sc_hd__fa_2_363/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_374 sky130_fd_sc_hd__fa_2_376/CIN sky130_fd_sc_hd__fa_2_367/B
+ sky130_fd_sc_hd__fa_2_393/A sky130_fd_sc_hd__fa_2_424/A sky130_fd_sc_hd__fa_2_417/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_15 sky130_fd_sc_hd__conb_1_9/LO sky130_fd_sc_hd__clkinv_8_9/Y
+ sky130_fd_sc_hd__dfxtp_1_140/CLK sky130_fd_sc_hd__or2_0_1/X VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_385 sky130_fd_sc_hd__fa_2_386/A sky130_fd_sc_hd__fa_2_378/A
+ sky130_fd_sc_hd__ha_2_110/B sky130_fd_sc_hd__fa_2_422/B sky130_fd_sc_hd__fa_2_286/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_26 sky130_fd_sc_hd__conb_1_17/LO sky130_fd_sc_hd__clkinv_4_51/A
+ sky130_fd_sc_hd__dfxtp_1_354/CLK sky130_fd_sc_hd__nor2_1_14/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__and2_1_1 VDD VSS sky130_fd_sc_hd__and2_1_1/X sky130_fd_sc_hd__ha_2_51/A
+ sky130_fd_sc_hd__nor2_4_2/Y VDD VSS sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__fa_2_396 sky130_fd_sc_hd__maj3_1_60/B sky130_fd_sc_hd__maj3_1_61/A
+ sky130_fd_sc_hd__fa_2_396/A sky130_fd_sc_hd__fa_2_396/B sky130_fd_sc_hd__fa_2_397/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22oi_2_7 sky130_fd_sc_hd__nor2_4_5/Y sky130_fd_sc_hd__a22oi_2_7/A2
+ sky130_fd_sc_hd__a22oi_2_9/B1 sky130_fd_sc_hd__a22oi_2_7/B2 sky130_fd_sc_hd__a22oi_2_7/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__diode_2_202 sky130_fd_sc_hd__buf_2_265/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__sdlclkp_4_37 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_4_51/A
+ sky130_fd_sc_hd__dfxtp_1_433/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__diode_2_213 amplitude_adc_done VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__sdlclkp_4_48 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_104/A
+ sky130_fd_sc_hd__dfxtp_1_454/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__diode_2_224 sig_amplitude[0] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__sdlclkp_4_59 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__clkinv_8_62/Y
+ sky130_fd_sc_hd__dfxtp_1_496/CLK sky130_fd_sc_hd__nand2b_1_5/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__diode_2_235 sky130_fd_sc_hd__a22oi_1_9/A2 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkinv_8_90 sky130_fd_sc_hd__clkinv_8_91/A sky130_fd_sc_hd__clkinv_8_90/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_90/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__nor2_1_106 sky130_fd_sc_hd__nor2_1_106/B sky130_fd_sc_hd__nor2_1_106/Y
+ sky130_fd_sc_hd__fa_2_1108/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_117 sky130_fd_sc_hd__nor2_1_117/B sky130_fd_sc_hd__o21a_1_13/A1
+ sky130_fd_sc_hd__nor2_1_117/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_128 sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__nor2_1_128/Y
+ sky130_fd_sc_hd__nor2_1_128/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_15 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__a22oi_1_9/A1
+ sky130_fd_sc_hd__buf_2_290/X sky130_fd_sc_hd__buf_2_282/X sky130_fd_sc_hd__nand3_1_7/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_139 sky130_fd_sc_hd__or2_0_8/B sky130_fd_sc_hd__nor2_1_139/Y
+ sky130_fd_sc_hd__nor2_1_139/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_26 sky130_fd_sc_hd__nor2_2_0/Y sky130_fd_sc_hd__clkinv_1_4/Y
+ sky130_fd_sc_hd__nand4_1_17/Y sky130_fd_sc_hd__nand4_1_1/Y sky130_fd_sc_hd__a22oi_1_26/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_37 sky130_fd_sc_hd__nor2_2_2/Y sky130_fd_sc_hd__a22oi_1_82/A1
+ sky130_fd_sc_hd__clkbuf_1_68/X sky130_fd_sc_hd__a22oi_1_37/A2 sky130_fd_sc_hd__nand4_1_2/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_48 sky130_fd_sc_hd__nor2_2_2/Y sky130_fd_sc_hd__a22oi_1_82/A1
+ sky130_fd_sc_hd__clkbuf_1_65/X sky130_fd_sc_hd__a22oi_1_48/A2 sky130_fd_sc_hd__nand4_1_5/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_59 sky130_fd_sc_hd__a22oi_1_81/B1 sky130_fd_sc_hd__clkbuf_1_99/X
+ sky130_fd_sc_hd__clkbuf_1_41/X sky130_fd_sc_hd__clkbuf_4_16/X sky130_fd_sc_hd__nand4_1_9/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_302 sky130_fd_sc_hd__buf_8_123/X sky130_fd_sc_hd__buf_12_302/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_313 sky130_fd_sc_hd__bufinv_8_7/Y sky130_fd_sc_hd__buf_12_313/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_324 sky130_fd_sc_hd__buf_4_93/X sky130_fd_sc_hd__buf_8_176/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_335 sky130_fd_sc_hd__buf_4_85/X sky130_fd_sc_hd__buf_12_335/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_346 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__buf_12_346/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_205 sky130_fd_sc_hd__clkbuf_4_111/X sky130_fd_sc_hd__clkbuf_4_112/X
+ sky130_fd_sc_hd__a22oi_1_205/B2 sky130_fd_sc_hd__clkbuf_1_283/X sky130_fd_sc_hd__a22oi_1_205/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_357 sky130_fd_sc_hd__buf_12_357/A sky130_fd_sc_hd__buf_12_357/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_216 sky130_fd_sc_hd__buf_2_164/X sky130_fd_sc_hd__nor2_4_8/Y
+ sky130_fd_sc_hd__clkbuf_1_425/X sky130_fd_sc_hd__buf_2_234/X sky130_fd_sc_hd__nand4_1_49/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_368 sky130_fd_sc_hd__buf_12_368/A sky130_fd_sc_hd__buf_12_373/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_227 sky130_fd_sc_hd__buf_2_164/X sky130_fd_sc_hd__nor2_4_8/Y
+ sky130_fd_sc_hd__buf_2_185/X sky130_fd_sc_hd__clkbuf_1_456/X sky130_fd_sc_hd__nand4_1_53/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_379 sky130_fd_sc_hd__inv_2_115/Y sky130_fd_sc_hd__buf_12_501/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_238 sky130_fd_sc_hd__buf_2_164/X sky130_fd_sc_hd__nor2_4_8/Y
+ sky130_fd_sc_hd__clkbuf_1_419/X sky130_fd_sc_hd__buf_2_228/X sky130_fd_sc_hd__nand4_1_57/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_249 sky130_fd_sc_hd__buf_2_164/X sky130_fd_sc_hd__nor2_4_8/Y
+ sky130_fd_sc_hd__clkbuf_1_415/X sky130_fd_sc_hd__buf_2_224/X sky130_fd_sc_hd__nand4_1_61/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_502 sky130_fd_sc_hd__a21oi_1_64/A1 sky130_fd_sc_hd__nor2_1_54/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_502/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_513 sky130_fd_sc_hd__o21ai_1_74/A1 sky130_fd_sc_hd__o21ai_1_81/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_513/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_524 sky130_fd_sc_hd__nor2_1_50/B sky130_fd_sc_hd__fa_2_1041/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_524/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_535 sky130_fd_sc_hd__nand2_1_261/A sky130_fd_sc_hd__a21oi_1_92/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_535/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_546 sky130_fd_sc_hd__nor2_1_64/B sky130_fd_sc_hd__fa_2_987/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_546/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_557 sky130_fd_sc_hd__o22ai_1_119/A1 sky130_fd_sc_hd__fa_2_979/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_557/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_568 sky130_fd_sc_hd__o22ai_1_122/B1 sky130_fd_sc_hd__o21ai_1_136/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_568/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_579 sky130_fd_sc_hd__o22ai_1_123/B2 sky130_fd_sc_hd__fa_2_1003/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_579/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_60 sky130_fd_sc_hd__nor2_1_60/B sky130_fd_sc_hd__nor2_1_60/Y
+ sky130_fd_sc_hd__nor2_1_60/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_15 sky130_fd_sc_hd__bufinv_8_4/A sky130_fd_sc_hd__clkinv_4_15/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_15/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_71 sky130_fd_sc_hd__nor2_1_71/B sky130_fd_sc_hd__nor2_1_71/Y
+ sky130_fd_sc_hd__nor2_4_10/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_26 sky130_fd_sc_hd__clkinv_4_26/A sky130_fd_sc_hd__clkinv_4_26/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_26/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_82 sky130_fd_sc_hd__nor2_1_82/B sky130_fd_sc_hd__nor2_1_82/Y
+ sky130_fd_sc_hd__nor2_1_82/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_37 sky130_fd_sc_hd__clkinv_4_37/A sky130_fd_sc_hd__buf_6_53/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_37/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_93 sky130_fd_sc_hd__nor2_1_93/B sky130_fd_sc_hd__nor2_1_93/Y
+ sky130_fd_sc_hd__nor2_1_93/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_48 sky130_fd_sc_hd__clkinv_4_48/A sky130_fd_sc_hd__clkinv_4_48/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_48/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_59 sky130_fd_sc_hd__clkinv_4_59/A sky130_fd_sc_hd__clkinv_8_75/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_59/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_sram_2kbyte_1rw1r_32x512_8_1 sky130_fd_sc_hd__buf_6_1/A sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__buf_4_1/X sky130_fd_sc_hd__buf_6_2/X sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__buf_6_3/X sky130_fd_sc_hd__buf_4_6/X sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__buf_6_7/X sky130_fd_sc_hd__clkbuf_4_2/X sky130_fd_sc_hd__clkbuf_4_3/X
+ sky130_fd_sc_hd__clkbuf_1_127/X sky130_fd_sc_hd__buf_4_10/X sky130_fd_sc_hd__clkbuf_4_7/X
+ sky130_fd_sc_hd__buf_6_8/X sky130_fd_sc_hd__buf_4_12/X sky130_fd_sc_hd__buf_6_1/A
+ sky130_fd_sc_hd__buf_4_0/X sky130_fd_sc_hd__buf_4_1/X sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__buf_4_4/X sky130_fd_sc_hd__buf_6_3/X sky130_fd_sc_hd__buf_4_6/X
+ sky130_fd_sc_hd__buf_6_5/X sky130_fd_sc_hd__buf_6_7/X sky130_fd_sc_hd__clkbuf_4_2/X
+ sky130_fd_sc_hd__clkbuf_4_3/X sky130_fd_sc_hd__clkbuf_4_4/X sky130_fd_sc_hd__buf_4_10/X
+ sky130_fd_sc_hd__clkbuf_4_7/X sky130_fd_sc_hd__buf_6_8/X sky130_fd_sc_hd__buf_4_12/X
+ sky130_fd_sc_hd__buf_12_45/X sky130_fd_sc_hd__buf_12_21/X sky130_fd_sc_hd__buf_12_57/X
+ sky130_fd_sc_hd__buf_12_43/X sky130_fd_sc_hd__buf_12_40/X sky130_fd_sc_hd__buf_12_80/X
+ sky130_fd_sc_hd__buf_12_19/X sky130_fd_sc_hd__buf_12_68/X sky130_fd_sc_hd__buf_12_75/X
+ sky130_fd_sc_hd__buf_12_1/X sky130_fd_sc_hd__buf_12_4/X sky130_fd_sc_hd__buf_12_16/X
+ sky130_fd_sc_hd__buf_12_54/X sky130_fd_sc_hd__buf_12_115/X sky130_fd_sc_hd__buf_12_67/X
+ sky130_fd_sc_hd__buf_12_8/X sky130_fd_sc_hd__buf_12_100/X sky130_fd_sc_hd__buf_12_46/X
+ sky130_fd_sc_hd__buf_2_23/X sky130_fd_sc_hd__clkbuf_1_126/X sky130_fd_sc_hd__buf_2_23/X
+ sky130_fd_sc_hd__clkinv_8_0/Y sky130_fd_sc_hd__clkinv_4_2/Y sky130_fd_sc_hd__buf_8_59/X
+ sky130_fd_sc_hd__buf_12_105/X sky130_fd_sc_hd__buf_12_103/X sky130_fd_sc_hd__buf_12_7/X
+ sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[0] sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[1]
+ sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[2] sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[3]
+ sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[4] sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[5]
+ sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[6] sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[7]
+ sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[8] sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[9]
+ sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[10] sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[11]
+ sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[12] sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[13]
+ sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[14] sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[15]
+ sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[16] sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[17]
+ sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[18] sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[19]
+ sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[20] sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[21]
+ sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[22] sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[23]
+ sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[24] sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[25]
+ sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[26] sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[27]
+ sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[28] sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[29]
+ sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[30] sky130_sram_2kbyte_1rw1r_32x512_8_1/dout0[31]
+ sky130_fd_sc_hd__clkbuf_1_35/A sky130_fd_sc_hd__clkbuf_1_36/A sky130_fd_sc_hd__clkbuf_1_37/A
+ sky130_fd_sc_hd__clkbuf_1_38/A sky130_fd_sc_hd__clkbuf_1_39/A sky130_fd_sc_hd__clkbuf_1_40/A
+ sky130_fd_sc_hd__clkbuf_1_41/A sky130_fd_sc_hd__clkbuf_1_42/A sky130_fd_sc_hd__clkbuf_1_43/A
+ sky130_fd_sc_hd__clkbuf_1_44/A sky130_fd_sc_hd__clkbuf_1_45/A sky130_fd_sc_hd__clkbuf_1_46/A
+ sky130_fd_sc_hd__clkbuf_1_47/A sky130_fd_sc_hd__clkbuf_1_48/A sky130_fd_sc_hd__clkbuf_1_49/A
+ sky130_fd_sc_hd__clkbuf_1_50/A sky130_fd_sc_hd__clkbuf_1_51/A sky130_fd_sc_hd__clkbuf_1_52/A
+ sky130_fd_sc_hd__clkbuf_1_53/A sky130_fd_sc_hd__clkbuf_1_54/A sky130_fd_sc_hd__a22oi_1_66/A2
+ sky130_fd_sc_hd__a22oi_1_63/A2 sky130_fd_sc_hd__a22oi_1_60/A2 sky130_fd_sc_hd__a22oi_1_57/A2
+ sky130_fd_sc_hd__a22oi_1_54/A2 sky130_fd_sc_hd__a22oi_1_51/A2 sky130_fd_sc_hd__a22oi_1_48/A2
+ sky130_fd_sc_hd__a22oi_1_45/A2 sky130_fd_sc_hd__a22oi_1_41/A2 sky130_fd_sc_hd__a22oi_1_37/A2
+ sky130_fd_sc_hd__a22oi_1_33/A2 sky130_fd_sc_hd__a22oi_1_30/A2 VDD VSS sky130_sram_2kbyte_1rw1r_32x512_8
Xsky130_fd_sc_hd__a21oi_1_410 sky130_fd_sc_hd__fa_2_1259/A sky130_fd_sc_hd__nor2_1_263/Y
+ sky130_fd_sc_hd__a21oi_1_410/Y sky130_fd_sc_hd__nor3_1_40/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_421 sky130_fd_sc_hd__o21a_1_57/B1 sky130_fd_sc_hd__o21a_1_56/A1
+ sky130_fd_sc_hd__a21oi_1_421/Y sky130_fd_sc_hd__nor2_1_303/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_432 sky130_fd_sc_hd__o21a_1_66/B1 sky130_fd_sc_hd__o21a_1_65/A1
+ sky130_fd_sc_hd__a21oi_1_432/Y sky130_fd_sc_hd__nor2_1_280/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_443 sky130_fd_sc_hd__o21ai_1_460/Y sky130_fd_sc_hd__a21oi_1_444/B1
+ sky130_fd_sc_hd__a21oi_1_443/Y sky130_fd_sc_hd__nor2b_2_5/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_454 sky130_fd_sc_hd__fa_2_1289/A sky130_fd_sc_hd__o22ai_1_416/Y
+ sky130_fd_sc_hd__a21oi_1_454/Y sky130_fd_sc_hd__nor3_1_41/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_465 sky130_fd_sc_hd__fa_2_1307/A sky130_fd_sc_hd__o22ai_1_425/Y
+ sky130_fd_sc_hd__a21oi_1_465/Y sky130_fd_sc_hd__a22oi_1_400/B1 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_476 sky130_fd_sc_hd__fa_2_1299/A sky130_fd_sc_hd__o22ai_1_432/Y
+ sky130_fd_sc_hd__a21oi_1_476/Y sky130_fd_sc_hd__nor3_1_41/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_487 sky130_fd_sc_hd__or2_0_13/A sky130_fd_sc_hd__or2_0_0/B
+ sky130_fd_sc_hd__nand2_1_555/A sky130_fd_sc_hd__nor2_1_322/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_8_101 sky130_fd_sc_hd__clkinv_4_51/A sky130_fd_sc_hd__clkinv_4_50/Y
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__a21oi_1_498 sky130_fd_sc_hd__nor2_1_318/Y sky130_fd_sc_hd__or2_0_0/B
+ sky130_fd_sc_hd__nand2_1_566/A sky130_fd_sc_hd__or2_0_13/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_8_112 sky130_fd_sc_hd__clkinv_8_15/A sky130_fd_sc_hd__clkinv_8_112/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_123 sky130_fd_sc_hd__clkinv_8_6/A sky130_fd_sc_hd__clkinv_4_63/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_123/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_134 sky130_fd_sc_hd__clkinv_8_135/A sky130_fd_sc_hd__clkinv_8_134/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__o21a_1_3 sky130_fd_sc_hd__o21a_1_3/X sky130_fd_sc_hd__o21a_1_3/A1
+ sky130_fd_sc_hd__o21a_1_3/B1 sky130_fd_sc_hd__fa_2_986/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__nand2_1_470 sky130_fd_sc_hd__nand2_1_470/Y sky130_fd_sc_hd__o31ai_1_9/A3
+ sky130_fd_sc_hd__o31ai_1_9/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_481 sky130_fd_sc_hd__nand2_1_481/Y sky130_fd_sc_hd__nand2_1_491/B
+ sky130_fd_sc_hd__o21ai_1_416/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_309 sky130_fd_sc_hd__nor2_4_20/Y sky130_fd_sc_hd__fa_2_1301/B
+ sky130_fd_sc_hd__xor2_1_309/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_492 sky130_fd_sc_hd__nand2_1_492/Y sky130_fd_sc_hd__nor2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_431/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_50 sky130_fd_sc_hd__nor2_1_21/A sky130_fd_sc_hd__nor2b_1_50/Y
+ sky130_fd_sc_hd__xor2_1_11/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_61 sky130_fd_sc_hd__dfxtp_1_502/Q sky130_fd_sc_hd__nor2b_1_61/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_72 sky130_fd_sc_hd__nor2_1_37/B sky130_fd_sc_hd__nor2b_1_72/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_83 sky130_fd_sc_hd__nor2b_1_87/A sky130_fd_sc_hd__nor2b_1_83/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1050 sky130_fd_sc_hd__o22ai_1_395/A1 sky130_fd_sc_hd__fa_2_3/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1050/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_94 sky130_fd_sc_hd__nor2b_1_90/Y sky130_fd_sc_hd__nor2b_1_94/Y
+ sky130_fd_sc_hd__buf_2_262/X VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1061 sky130_fd_sc_hd__o32ai_1_9/B2 sky130_fd_sc_hd__fa_2_1277/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1061/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_2 VSS VDD sky130_fd_sc_hd__xnor2_1_2/B sky130_fd_sc_hd__xnor2_1_2/Y
+ sky130_fd_sc_hd__xnor2_1_2/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_1072 sky130_fd_sc_hd__a21oi_1_447/A1 sky130_fd_sc_hd__a21boi_1_7/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1072/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1083 sky130_fd_sc_hd__o22ai_1_422/A1 sky130_fd_sc_hd__fa_2_1283/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1083/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1094 sky130_fd_sc_hd__o22ai_1_429/B1 sky130_fd_sc_hd__fa_2_1303/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1094/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_160 sky130_fd_sc_hd__fa_2_150/A sky130_fd_sc_hd__fa_2_158/A
+ sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__fa_2_160/B sky130_fd_sc_hd__fa_2_160/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_17 VDD VSS sky130_fd_sc_hd__ha_2_112/B sky130_fd_sc_hd__dfxtp_1_29/CLK
+ sky130_fd_sc_hd__nand4_1_35/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_171 sky130_fd_sc_hd__fa_2_169/CIN sky130_fd_sc_hd__or3_1_4/C
+ sky130_fd_sc_hd__fa_2_171/A sky130_fd_sc_hd__fa_2_171/B sky130_fd_sc_hd__fa_2_171/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_28 VDD VSS sky130_fd_sc_hd__ha_2_116/A sky130_fd_sc_hd__dfxtp_1_29/CLK
+ sky130_fd_sc_hd__nand4_1_46/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_182 sky130_fd_sc_hd__fa_2_184/CIN sky130_fd_sc_hd__fa_2_180/B
+ sky130_fd_sc_hd__fa_2_242/B sky130_fd_sc_hd__fa_2_242/A sky130_fd_sc_hd__fa_2_266/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_39 VDD VSS sky130_fd_sc_hd__fa_2_910/CIN sky130_fd_sc_hd__dfxtp_1_39/CLK
+ sky130_fd_sc_hd__buf_2_289/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_193 sky130_fd_sc_hd__fa_2_196/A sky130_fd_sc_hd__fa_2_193/SUM
+ sky130_fd_sc_hd__fa_2_193/A sky130_fd_sc_hd__fa_2_193/B sky130_fd_sc_hd__fa_2_193/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o22ai_1_70 sky130_fd_sc_hd__o22ai_1_88/B1 sky130_fd_sc_hd__nand2_2_3/Y
+ sky130_fd_sc_hd__o22ai_1_70/Y sky130_fd_sc_hd__xnor2_1_51/Y sky130_fd_sc_hd__o22ai_1_84/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkbuf_4_107 sky130_fd_sc_hd__clkbuf_4_107/X sky130_fd_sc_hd__buf_6_84/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o22ai_1_81 sky130_fd_sc_hd__o22ai_1_89/A1 sky130_fd_sc_hd__o22ai_1_88/B1
+ sky130_fd_sc_hd__o22ai_1_81/Y sky130_fd_sc_hd__xnor2_1_45/Y sky130_fd_sc_hd__o22ai_1_81/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkbuf_4_118 sky130_fd_sc_hd__clkbuf_4_118/X sky130_fd_sc_hd__clkbuf_4_118/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o22ai_1_92 sky130_fd_sc_hd__nor2_2_9/B sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__o22ai_1_92/Y sky130_fd_sc_hd__o22ai_1_92/A1 sky130_fd_sc_hd__a21oi_1_83/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkbuf_4_129 sky130_fd_sc_hd__clkbuf_4_129/X sky130_fd_sc_hd__clkbuf_4_129/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_4_50 VDD VSS sky130_fd_sc_hd__buf_4_50/X sky130_fd_sc_hd__buf_8_90/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_61 VDD VSS sky130_fd_sc_hd__buf_4_61/X sky130_fd_sc_hd__buf_6_89/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_72 VDD VSS sky130_fd_sc_hd__buf_4_72/X sky130_fd_sc_hd__buf_6_31/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_83 VDD VSS sky130_fd_sc_hd__buf_4_83/X sky130_fd_sc_hd__buf_4_83/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_94 VDD VSS sky130_fd_sc_hd__buf_4_96/A sky130_fd_sc_hd__buf_4_95/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_12_110 sky130_fd_sc_hd__buf_12_69/X sky130_fd_sc_hd__buf_12_110/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_121 sky130_fd_sc_hd__buf_4_34/X sky130_fd_sc_hd__buf_12_121/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_132 sky130_fd_sc_hd__buf_12_132/A sky130_fd_sc_hd__buf_12_167/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_143 sky130_fd_sc_hd__inv_2_72/Y sky130_fd_sc_hd__buf_12_143/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_154 sky130_fd_sc_hd__buf_8_92/X sky130_fd_sc_hd__buf_12_154/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_165 sky130_fd_sc_hd__buf_8_86/X sky130_fd_sc_hd__buf_12_233/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_4_2 sky130_fd_sc_hd__clkbuf_4_2/X sky130_fd_sc_hd__buf_2_6/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_12_176 sky130_fd_sc_hd__buf_8_100/X sky130_fd_sc_hd__buf_12_176/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_187 sky130_fd_sc_hd__buf_4_41/X sky130_fd_sc_hd__buf_12_187/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_198 sky130_fd_sc_hd__buf_4_47/X sky130_fd_sc_hd__buf_12_198/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_310 sky130_fd_sc_hd__fa_2_389/B sky130_fd_sc_hd__ha_2_115/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_310/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_321 sky130_fd_sc_hd__fa_2_424/A sky130_fd_sc_hd__ha_2_115/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_321/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_332 sky130_fd_sc_hd__fa_2_543/A sky130_fd_sc_hd__fa_2_535/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_332/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_343 sky130_fd_sc_hd__fa_2_695/A sky130_fd_sc_hd__ha_2_135/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_343/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_354 sky130_fd_sc_hd__fa_2_624/B sky130_fd_sc_hd__fa_2_667/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_354/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_365 sky130_fd_sc_hd__ha_2_136/A sky130_fd_sc_hd__fa_2_811/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_365/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_376 sky130_fd_sc_hd__fa_2_872/B sky130_fd_sc_hd__dfxtp_1_272/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_376/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_387 sky130_fd_sc_hd__fa_2_885/B sky130_fd_sc_hd__nor4_1_4/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_387/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_398 sky130_fd_sc_hd__nand2_1_203/B sky130_fd_sc_hd__nand2_1_35/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_398/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21a_1_17 sky130_fd_sc_hd__o21a_1_17/X sky130_fd_sc_hd__o21a_1_17/A1
+ sky130_fd_sc_hd__xnor2_1_91/B sky130_fd_sc_hd__fa_2_1138/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_28 sky130_fd_sc_hd__o21a_1_28/X sky130_fd_sc_hd__o21a_1_28/A1
+ sky130_fd_sc_hd__o21a_1_28/B1 sky130_fd_sc_hd__fa_2_1145/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_39 sky130_fd_sc_hd__o21a_1_39/X sky130_fd_sc_hd__o21a_1_39/A1
+ sky130_fd_sc_hd__o21a_1_39/B1 sky130_fd_sc_hd__fa_2_1201/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__a21oi_1_240 sky130_fd_sc_hd__a21o_2_5/A2 sky130_fd_sc_hd__o21ai_1_275/Y
+ sky130_fd_sc_hd__a21oi_1_240/Y sky130_fd_sc_hd__fa_2_1079/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_251 sky130_fd_sc_hd__o21a_1_26/B1 sky130_fd_sc_hd__o21a_1_25/A1
+ sky130_fd_sc_hd__dfxtp_1_887/D sky130_fd_sc_hd__o21a_1_29/A2 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_262 sky130_fd_sc_hd__xor2_1_140/X sky130_fd_sc_hd__o21ai_1_287/Y
+ sky130_fd_sc_hd__dfxtp_1_987/D sky130_fd_sc_hd__nand2_1_366/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_273 sky130_fd_sc_hd__nor2_2_15/Y sky130_fd_sc_hd__o21ai_1_300/Y
+ sky130_fd_sc_hd__nor2_1_172/B sky130_fd_sc_hd__fa_2_1138/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_284 sky130_fd_sc_hd__clkinv_1_838/Y sky130_fd_sc_hd__nor2_1_177/Y
+ sky130_fd_sc_hd__a21oi_1_284/Y sky130_fd_sc_hd__nor2b_1_104/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_4_2 sky130_fd_sc_hd__clkinv_4_2/A sky130_fd_sc_hd__clkinv_4_2/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_2/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__a21oi_1_295 sky130_fd_sc_hd__nor3_1_38/A sky130_fd_sc_hd__o22ai_1_260/Y
+ sky130_fd_sc_hd__a21oi_1_295/Y sky130_fd_sc_hd__fa_2_1150/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_203 sky130_fd_sc_hd__buf_8_203/A sky130_fd_sc_hd__buf_8_203/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_214 sky130_fd_sc_hd__buf_8_214/A sky130_fd_sc_hd__buf_8_214/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xor2_1_106 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1051/B
+ sky130_fd_sc_hd__xor2_1_106/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_117 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1089/B
+ sky130_fd_sc_hd__xor2_1_117/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_128 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1078/B
+ sky130_fd_sc_hd__xor2_1_128/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_139 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__xor2_1_139/X
+ sky130_fd_sc_hd__xor2_1_139/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_1408 VDD VSS sky130_fd_sc_hd__mux2_2_225/A1 sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__o22ai_1_381/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1419 VDD VSS sky130_fd_sc_hd__mux2_2_253/A0 sky130_fd_sc_hd__clkinv_8_65/Y
+ sky130_fd_sc_hd__dfxtp_1_434/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_108 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_108/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_836/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_16 sky130_fd_sc_hd__nand3_1_25/B sky130_fd_sc_hd__ha_2_10/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_16/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_119 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_119/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_852/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_27 sky130_fd_sc_hd__inv_2_16/A sky130_fd_sc_hd__ha_2_27/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_27/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_38 sky130_fd_sc_hd__inv_2_27/A sky130_fd_sc_hd__buf_2_13/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_38/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_49 sky130_fd_sc_hd__inv_2_38/A sky130_fd_sc_hd__ha_2_23/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_49/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_3 sky130_fd_sc_hd__fa_2_2/CIN sky130_fd_sc_hd__fa_2_3/SUM sky130_fd_sc_hd__fa_2_9/A
+ sky130_fd_sc_hd__fa_2_3/B sky130_fd_sc_hd__fa_2_3/CIN VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_201 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_201/A sky130_fd_sc_hd__ha_2_201/COUT
+ sky130_fd_sc_hd__ha_2_201/SUM sky130_fd_sc_hd__ha_2_201/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_907 sky130_fd_sc_hd__fa_2_895/A sky130_fd_sc_hd__fa_2_896/B
+ sky130_fd_sc_hd__fa_2_907/A sky130_fd_sc_hd__fa_2_907/B sky130_fd_sc_hd__fa_2_907/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_918 sky130_fd_sc_hd__fa_2_917/CIN sky130_fd_sc_hd__fa_2_918/SUM
+ sky130_fd_sc_hd__fa_2_918/A sky130_fd_sc_hd__fa_2_918/B sky130_fd_sc_hd__fa_2_918/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_929 sky130_fd_sc_hd__fa_2_928/CIN sky130_fd_sc_hd__fa_2_929/SUM
+ sky130_fd_sc_hd__fa_2_929/A sky130_fd_sc_hd__fa_2_929/B sky130_fd_sc_hd__fa_2_929/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a211o_1_20 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_202/A sky130_fd_sc_hd__o21ai_1_370/Y
+ sky130_fd_sc_hd__nor2_1_206/Y sky130_fd_sc_hd__nor2b_2_3/Y sky130_fd_sc_hd__o22ai_1_295/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__mux2_2_207 VSS VDD sky130_fd_sc_hd__mux2_2_207/A1 sky130_fd_sc_hd__mux2_2_207/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_207/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_218 VSS VDD sky130_fd_sc_hd__mux2_2_218/A1 sky130_fd_sc_hd__mux2_2_218/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_218/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_229 VSS VDD sky130_fd_sc_hd__mux2_2_229/A1 sky130_fd_sc_hd__mux2_2_229/A0
+ sky130_fd_sc_hd__nor2_8_2/A sky130_fd_sc_hd__mux2_2_229/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__clkinv_1_140 sky130_fd_sc_hd__clkinv_1_141/A sky130_fd_sc_hd__buf_2_126/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_140/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_151 sky130_fd_sc_hd__inv_2_84/A sky130_fd_sc_hd__clkinv_1_151/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_151/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_162 sky130_fd_sc_hd__inv_2_93/A sky130_fd_sc_hd__inv_2_80/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_162/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_173 sky130_fd_sc_hd__inv_2_102/A sky130_fd_sc_hd__inv_2_94/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_173/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_5 sky130_fd_sc_hd__buf_8_5/A sky130_fd_sc_hd__buf_8_5/X VSS
+ VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__a22o_1_7 sky130_fd_sc_hd__a22o_1_7/A1 sky130_fd_sc_hd__nor2_1_1/Y
+ sky130_fd_sc_hd__a22o_1_7/X sky130_fd_sc_hd__a22o_1_7/B2 sky130_fd_sc_hd__nor2_1_0/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_184 sky130_fd_sc_hd__a22o_4_0/B1 sky130_fd_sc_hd__or2_1_1/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_184/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_195 sky130_fd_sc_hd__buf_6_59/A sky130_fd_sc_hd__buf_2_240/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_195/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_20 sky130_fd_sc_hd__nor2_4_4/Y sky130_fd_sc_hd__ha_2_77/A
+ sky130_fd_sc_hd__inv_4_0/A sky130_fd_sc_hd__a22o_1_20/B2 sky130_fd_sc_hd__a22o_2_6/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_31 sky130_fd_sc_hd__or2_1_1/B sky130_fd_sc_hd__ha_2_85/A
+ sky130_fd_sc_hd__a22o_1_31/X sky130_fd_sc_hd__a22o_1_31/B2 sky130_fd_sc_hd__a22o_4_0/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_42 sky130_fd_sc_hd__a22o_1_42/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_42/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__fa_2_948/SUM
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_53 sky130_fd_sc_hd__a22o_1_53/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_53/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__nor4_1_9/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_64 sky130_fd_sc_hd__a22o_1_64/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_64/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__nor4_1_12/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_75 sky130_fd_sc_hd__nor2_2_12/Y sky130_fd_sc_hd__fa_2_1072/A
+ sky130_fd_sc_hd__a22o_1_75/X sky130_fd_sc_hd__fa_2_1070/A sky130_fd_sc_hd__nor2_4_13/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__nand4_1_3 sky130_fd_sc_hd__nand4_1_3/C sky130_fd_sc_hd__nand4_1_3/B
+ sky130_fd_sc_hd__nand4_1_3/Y sky130_fd_sc_hd__nand4_1_3/D sky130_fd_sc_hd__nand4_1_3/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__o21ai_1_109 VSS VDD sky130_fd_sc_hd__nor2_1_74/A sky130_fd_sc_hd__o21ai_1_109/A1
+ sky130_fd_sc_hd__a21oi_1_94/Y sky130_fd_sc_hd__xor2_1_74/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__maj3_1_15 sky130_fd_sc_hd__maj3_1_16/X sky130_fd_sc_hd__maj3_1_15/X
+ sky130_fd_sc_hd__maj3_1_15/B sky130_fd_sc_hd__maj3_1_15/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_26 sky130_fd_sc_hd__maj3_1_27/X sky130_fd_sc_hd__maj3_1_26/X
+ sky130_fd_sc_hd__maj3_1_26/B sky130_fd_sc_hd__maj3_1_26/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_405 sky130_fd_sc_hd__nand2_1_516/Y sky130_fd_sc_hd__nand2_1_515/Y
+ sky130_fd_sc_hd__o22ai_1_405/Y sky130_fd_sc_hd__o22ai_1_405/A1 sky130_fd_sc_hd__a21o_2_29/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_37 sky130_fd_sc_hd__maj3_1_38/X sky130_fd_sc_hd__maj3_1_37/X
+ sky130_fd_sc_hd__maj3_1_37/B sky130_fd_sc_hd__maj3_1_37/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_416 sky130_fd_sc_hd__o22ai_1_436/A2 sky130_fd_sc_hd__o22ai_1_423/B1
+ sky130_fd_sc_hd__o22ai_1_416/Y sky130_fd_sc_hd__nor2_1_271/B sky130_fd_sc_hd__o22ai_1_432/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_48 sky130_fd_sc_hd__maj3_1_49/X sky130_fd_sc_hd__maj3_1_48/X
+ sky130_fd_sc_hd__maj3_1_48/B sky130_fd_sc_hd__maj3_1_48/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_427 sky130_fd_sc_hd__o32ai_1_11/A3 sky130_fd_sc_hd__o22ai_1_430/B1
+ sky130_fd_sc_hd__o22ai_1_427/Y sky130_fd_sc_hd__nor2_1_305/A sky130_fd_sc_hd__o21a_1_68/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_59 sky130_fd_sc_hd__maj3_1_60/X sky130_fd_sc_hd__maj3_1_59/X
+ sky130_fd_sc_hd__maj3_1_59/B sky130_fd_sc_hd__maj3_1_59/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_10 sky130_fd_sc_hd__nand3_1_10/C sky130_fd_sc_hd__nand4_1_69/Y
+ sky130_fd_sc_hd__nand2_1_9/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_21 sky130_fd_sc_hd__or2_0_1/B sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__inv_8_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_32 sky130_fd_sc_hd__nand2_1_32/Y sky130_fd_sc_hd__xor2_1_10/X
+ sky130_fd_sc_hd__o31ai_1_1/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_43 sky130_fd_sc_hd__nand2_1_43/Y sky130_fd_sc_hd__nand2_1_43/B
+ sky130_fd_sc_hd__a21oi_2_0/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_54 sky130_fd_sc_hd__nand2_1_54/Y sky130_fd_sc_hd__nand2_1_55/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_65 sky130_fd_sc_hd__nand2_1_65/Y sky130_fd_sc_hd__nand2_1_7/B
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_76 sky130_fd_sc_hd__nand2_1_76/Y sky130_fd_sc_hd__nand2_1_77/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_87 sky130_fd_sc_hd__nand2_1_87/Y sky130_fd_sc_hd__nand2_1_87/B
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_98 sky130_fd_sc_hd__nand2_1_98/Y sky130_fd_sc_hd__nand2_1_99/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_309 VDD VSS sky130_fd_sc_hd__a22o_1_40/A1 sky130_fd_sc_hd__dfxtp_1_313/CLK
+ sky130_fd_sc_hd__and2_0_89/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_17 sky130_fd_sc_hd__fa_2_10/B sky130_fd_sc_hd__fa_2_18/CIN
+ sky130_fd_sc_hd__fa_2_82/A sky130_fd_sc_hd__ha_2_95/A sky130_fd_sc_hd__fa_2_76/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_28 sky130_fd_sc_hd__fa_2_29/CIN sky130_fd_sc_hd__or3_1_5/B
+ sky130_fd_sc_hd__fa_2_28/A sky130_fd_sc_hd__fa_2_28/B sky130_fd_sc_hd__maj3_1_4/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_39 sky130_fd_sc_hd__fa_2_41/B sky130_fd_sc_hd__fa_2_39/SUM
+ sky130_fd_sc_hd__ha_2_91/B sky130_fd_sc_hd__fa_2_92/B sky130_fd_sc_hd__fa_2_39/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_209 VDD VSS sky130_fd_sc_hd__buf_2_209/X sky130_fd_sc_hd__buf_2_209/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_sram_2kbyte_1rw1r_32x512_8_13 sky130_fd_sc_hd__buf_6_49/X sky130_fd_sc_hd__buf_6_50/X
+ sky130_fd_sc_hd__buf_2_140/A sky130_fd_sc_hd__buf_6_51/X sky130_fd_sc_hd__buf_2_144/A
+ sky130_fd_sc_hd__buf_2_146/A sky130_fd_sc_hd__buf_2_147/A sky130_fd_sc_hd__clkbuf_8_3/X
+ sky130_fd_sc_hd__buf_2_149/A sky130_fd_sc_hd__buf_6_52/X sky130_fd_sc_hd__buf_6_53/X
+ sky130_fd_sc_hd__buf_6_55/X sky130_fd_sc_hd__buf_2_153/A sky130_fd_sc_hd__buf_6_56/X
+ sky130_fd_sc_hd__buf_6_57/X sky130_fd_sc_hd__buf_2_156/A sky130_fd_sc_hd__buf_6_49/X
+ sky130_fd_sc_hd__buf_6_50/X sky130_fd_sc_hd__buf_2_140/A sky130_fd_sc_hd__buf_6_51/X
+ sky130_fd_sc_hd__buf_2_144/A sky130_fd_sc_hd__buf_2_146/A sky130_fd_sc_hd__buf_2_147/A
+ sky130_fd_sc_hd__clkbuf_8_3/X sky130_fd_sc_hd__buf_2_149/A sky130_fd_sc_hd__buf_6_52/X
+ sky130_fd_sc_hd__buf_6_53/X sky130_fd_sc_hd__buf_6_55/X sky130_fd_sc_hd__buf_2_153/A
+ sky130_fd_sc_hd__buf_6_56/X sky130_fd_sc_hd__buf_6_57/X sky130_fd_sc_hd__buf_2_156/A
+ sky130_fd_sc_hd__buf_12_459/X sky130_fd_sc_hd__buf_12_486/X sky130_fd_sc_hd__buf_12_473/X
+ sky130_fd_sc_hd__buf_12_443/X sky130_fd_sc_hd__buf_12_476/X sky130_fd_sc_hd__buf_12_515/X
+ sky130_fd_sc_hd__buf_12_501/X sky130_fd_sc_hd__buf_12_477/X sky130_fd_sc_hd__buf_12_427/X
+ sky130_fd_sc_hd__buf_12_407/X sky130_fd_sc_hd__buf_12_456/X sky130_fd_sc_hd__buf_12_489/X
+ sky130_fd_sc_hd__buf_12_448/X sky130_fd_sc_hd__buf_12_445/X sky130_fd_sc_hd__buf_12_493/X
+ sky130_fd_sc_hd__buf_12_499/X sky130_fd_sc_hd__buf_12_485/X sky130_fd_sc_hd__buf_12_410/X
+ sky130_fd_sc_hd__nand2_2_1/Y sky130_fd_sc_hd__clkinv_1_208/Y sky130_fd_sc_hd__buf_2_244/X
+ sky130_fd_sc_hd__clkinv_8_38/Y sky130_fd_sc_hd__clkinv_8_31/Y sky130_fd_sc_hd__buf_12_432/X
+ sky130_fd_sc_hd__buf_12_513/X sky130_fd_sc_hd__buf_6_83/X sky130_fd_sc_hd__buf_12_510/X
+ sky130_fd_sc_hd__clkbuf_1_540/A sky130_fd_sc_hd__a22oi_1_251/B2 sky130_fd_sc_hd__clkbuf_1_428/A
+ sky130_fd_sc_hd__clkbuf_1_429/A sky130_fd_sc_hd__clkbuf_1_430/A sky130_fd_sc_hd__clkbuf_1_499/A
+ sky130_fd_sc_hd__clkbuf_1_431/A sky130_fd_sc_hd__clkbuf_1_432/A sky130_fd_sc_hd__clkbuf_1_433/A
+ sky130_fd_sc_hd__clkbuf_1_434/A sky130_fd_sc_hd__a22oi_1_225/B2 sky130_fd_sc_hd__clkbuf_1_521/A
+ sky130_fd_sc_hd__clkbuf_1_435/A sky130_fd_sc_hd__clkbuf_1_436/A sky130_fd_sc_hd__clkbuf_1_437/A
+ sky130_fd_sc_hd__clkbuf_1_438/A sky130_fd_sc_hd__clkbuf_1_439/A sky130_fd_sc_hd__clkbuf_1_440/A
+ sky130_fd_sc_hd__clkbuf_1_441/A sky130_fd_sc_hd__clkbuf_1_442/A sky130_fd_sc_hd__clkbuf_1_443/A
+ sky130_fd_sc_hd__clkbuf_1_444/A sky130_fd_sc_hd__clkbuf_1_445/A sky130_fd_sc_hd__clkbuf_1_446/A
+ sky130_fd_sc_hd__clkbuf_1_447/A sky130_fd_sc_hd__clkbuf_1_448/A sky130_fd_sc_hd__clkbuf_1_449/A
+ sky130_fd_sc_hd__clkbuf_1_450/A sky130_fd_sc_hd__clkbuf_1_451/A sky130_fd_sc_hd__clkbuf_1_539/A
+ sky130_fd_sc_hd__clkbuf_1_453/A sky130_fd_sc_hd__clkbuf_1_454/A sky130_fd_sc_hd__buf_2_218/A
+ sky130_fd_sc_hd__buf_2_219/A sky130_fd_sc_hd__buf_2_220/A sky130_fd_sc_hd__clkbuf_4_166/A
+ sky130_fd_sc_hd__clkbuf_4_167/A sky130_fd_sc_hd__clkbuf_4_168/A sky130_fd_sc_hd__clkbuf_4_169/A
+ sky130_fd_sc_hd__clkbuf_1_538/A sky130_fd_sc_hd__buf_2_221/A sky130_fd_sc_hd__buf_2_222/A
+ sky130_fd_sc_hd__clkbuf_4_171/A sky130_fd_sc_hd__clkbuf_4_172/A sky130_fd_sc_hd__clkbuf_4_173/A
+ sky130_fd_sc_hd__clkbuf_4_174/A sky130_fd_sc_hd__clkbuf_4_175/A sky130_fd_sc_hd__clkbuf_4_176/A
+ sky130_fd_sc_hd__clkbuf_4_177/A sky130_fd_sc_hd__clkbuf_4_178/A sky130_fd_sc_hd__clkbuf_4_179/A
+ sky130_fd_sc_hd__clkbuf_4_180/A sky130_fd_sc_hd__clkbuf_4_181/A sky130_fd_sc_hd__clkbuf_4_182/A
+ sky130_fd_sc_hd__clkbuf_4_183/A sky130_fd_sc_hd__clkbuf_4_184/A sky130_fd_sc_hd__clkbuf_4_185/A
+ sky130_fd_sc_hd__clkbuf_4_186/A sky130_fd_sc_hd__clkbuf_4_187/A sky130_fd_sc_hd__clkbuf_4_188/A
+ sky130_fd_sc_hd__clkbuf_1_529/A sky130_fd_sc_hd__clkbuf_4_190/A sky130_fd_sc_hd__clkbuf_4_191/A
+ sky130_fd_sc_hd__clkbuf_4_192/A VDD VSS sky130_sram_2kbyte_1rw1r_32x512_8
Xsky130_fd_sc_hd__dfxtp_1_1205 VDD VSS sky130_fd_sc_hd__fa_2_1254/A sky130_fd_sc_hd__clkinv_8_75/Y
+ sky130_fd_sc_hd__mux2_2_184/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1216 VDD VSS sky130_fd_sc_hd__fa_2_1228/A sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__mux2_2_207/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1227 VDD VSS sky130_fd_sc_hd__fa_2_1239/A sky130_fd_sc_hd__clkinv_8_116/Y
+ sky130_fd_sc_hd__mux2_2_179/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1238 VDD VSS sky130_fd_sc_hd__fa_2_1267/A sky130_fd_sc_hd__clkinv_8_65/Y
+ sky130_fd_sc_hd__mux2_2_208/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_810 VDD VSS sky130_fd_sc_hd__fa_2_1062/A sky130_fd_sc_hd__clkinv_4_26/Y
+ sky130_fd_sc_hd__mux2_2_53/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1249 VDD VSS sky130_fd_sc_hd__nor2_4_18/B sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__nor2b_1_121/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_821 VDD VSS sky130_fd_sc_hd__fa_2_1095/A sky130_fd_sc_hd__clkinv_8_59/Y
+ sky130_fd_sc_hd__and2_0_297/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_832 VDD VSS sky130_fd_sc_hd__fa_2_1106/A sky130_fd_sc_hd__clkinv_4_26/Y
+ sky130_fd_sc_hd__mux2_2_68/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_843 VDD VSS sky130_fd_sc_hd__mux2_2_69/A0 sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__o21ai_1_160/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_854 VDD VSS sky130_fd_sc_hd__mux2_2_45/A1 sky130_fd_sc_hd__clkinv_4_25/Y
+ sky130_fd_sc_hd__o21ai_1_171/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_865 VDD VSS sky130_fd_sc_hd__mux2_2_62/A1 sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__o21ai_1_179/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_876 VDD VSS sky130_fd_sc_hd__mux2_2_39/A1 sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__o21ai_1_190/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_887 VDD VSS sky130_fd_sc_hd__fa_2_855/A sky130_fd_sc_hd__dfxtp_1_904/CLK
+ sky130_fd_sc_hd__dfxtp_1_887/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_898 VDD VSS sky130_fd_sc_hd__fa_2_933/B sky130_fd_sc_hd__dfxtp_1_904/CLK
+ sky130_fd_sc_hd__dfxtp_1_898/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_430 VSS VDD sky130_fd_sc_hd__clkbuf_1_430/X sky130_fd_sc_hd__clkbuf_1_430/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_441 VSS VDD sky130_fd_sc_hd__a22oi_2_29/A2 sky130_fd_sc_hd__clkbuf_1_441/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_452 VSS VDD sky130_fd_sc_hd__a22oi_2_16/A2 sky130_fd_sc_hd__clkbuf_1_539/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_463 VSS VDD sky130_fd_sc_hd__clkbuf_1_463/X sky130_fd_sc_hd__clkbuf_1_463/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_474 VSS VDD sky130_fd_sc_hd__nand4_1_63/D sky130_fd_sc_hd__a22oi_1_254/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_485 VSS VDD sky130_fd_sc_hd__clkbuf_1_485/X sky130_fd_sc_hd__nand3_2_7/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_704 sky130_fd_sc_hd__fa_2_703/CIN sky130_fd_sc_hd__fa_2_704/SUM
+ sky130_fd_sc_hd__fa_2_704/A sky130_fd_sc_hd__fa_2_704/B sky130_fd_sc_hd__fa_2_704/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_496 VSS VDD sky130_fd_sc_hd__a22oi_2_27/B2 sky130_fd_sc_hd__clkbuf_1_496/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_715 sky130_fd_sc_hd__fa_2_714/CIN sky130_fd_sc_hd__fa_2_715/SUM
+ sky130_fd_sc_hd__fa_2_715/A sky130_fd_sc_hd__fa_2_715/B sky130_fd_sc_hd__fa_2_715/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_726 sky130_fd_sc_hd__maj3_1_153/B sky130_fd_sc_hd__maj3_1_154/A
+ sky130_fd_sc_hd__fa_2_726/A sky130_fd_sc_hd__fa_2_726/B sky130_fd_sc_hd__fa_2_727/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_737 sky130_fd_sc_hd__fa_2_739/B sky130_fd_sc_hd__fa_2_735/A
+ sky130_fd_sc_hd__fa_2_817/B sky130_fd_sc_hd__ha_2_140/B sky130_fd_sc_hd__fa_2_834/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_748 sky130_fd_sc_hd__maj3_1_146/B sky130_fd_sc_hd__maj3_1_147/A
+ sky130_fd_sc_hd__fa_2_748/A sky130_fd_sc_hd__fa_2_748/B sky130_fd_sc_hd__fa_2_749/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_759 sky130_fd_sc_hd__fa_2_761/CIN sky130_fd_sc_hd__fa_2_756/A
+ sky130_fd_sc_hd__fa_2_826/A sky130_fd_sc_hd__fa_2_759/B sky130_fd_sc_hd__fa_2_759/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor2b_1_101 sky130_fd_sc_hd__nor2b_1_97/Y sky130_fd_sc_hd__nor2b_1_101/Y
+ sky130_fd_sc_hd__buf_2_262/X VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_112 sky130_fd_sc_hd__nor2b_2_3/A sky130_fd_sc_hd__nor2b_1_112/Y
+ sky130_fd_sc_hd__o32ai_1_5/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_123 sky130_fd_sc_hd__o32ai_1_8/Y sky130_fd_sc_hd__nor2b_1_123/Y
+ sky130_fd_sc_hd__buf_2_262/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_134 sky130_fd_sc_hd__a21oi_1_481/Y sky130_fd_sc_hd__nor2b_1_134/Y
+ sky130_fd_sc_hd__nor4_1_13/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__buf_6_2 VDD VSS sky130_fd_sc_hd__buf_6_2/X sky130_fd_sc_hd__buf_6_2/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__bufbuf_8_5 sky130_fd_sc_hd__a22o_1_19/X sky130_fd_sc_hd__bufbuf_8_5/X
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufbuf_8
Xsky130_fd_sc_hd__buf_6_18 VDD VSS sky130_fd_sc_hd__buf_6_18/X sky130_fd_sc_hd__buf_6_18/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_29 VDD VSS sky130_fd_sc_hd__buf_6_29/X sky130_fd_sc_hd__buf_6_29/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__o22ai_1_202 sky130_fd_sc_hd__nor2_1_137/A sky130_fd_sc_hd__o22ai_1_204/B1
+ sky130_fd_sc_hd__o22ai_1_202/Y sky130_fd_sc_hd__o22ai_1_206/B1 sky130_fd_sc_hd__nor2_1_138/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__sdlclkp_4_0 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__clkinv_8_118/Y
+ sky130_fd_sc_hd__dfxtp_1_61/CLK sky130_fd_sc_hd__clkbuf_1_0/X VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__o22ai_1_213 sky130_fd_sc_hd__nand2_1_358/Y sky130_fd_sc_hd__nand2_1_357/Y
+ sky130_fd_sc_hd__o22ai_1_213/Y sky130_fd_sc_hd__o22ai_1_226/A1 sky130_fd_sc_hd__a21o_2_7/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_224 sky130_fd_sc_hd__nand2_1_360/Y sky130_fd_sc_hd__nand2_1_359/Y
+ sky130_fd_sc_hd__o22ai_1_224/Y sky130_fd_sc_hd__o22ai_1_224/A1 sky130_fd_sc_hd__a21o_2_6/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_235 sky130_fd_sc_hd__nand2_1_360/Y sky130_fd_sc_hd__nand2_1_359/Y
+ sky130_fd_sc_hd__o22ai_1_235/Y sky130_fd_sc_hd__o22ai_1_235/A1 sky130_fd_sc_hd__o21ai_1_283/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_246 sky130_fd_sc_hd__o22ai_1_265/A2 sky130_fd_sc_hd__o22ai_1_247/A1
+ sky130_fd_sc_hd__o22ai_1_246/Y sky130_fd_sc_hd__nor2_1_146/B sky130_fd_sc_hd__o32ai_1_2/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_257 sky130_fd_sc_hd__o22ai_1_265/A2 sky130_fd_sc_hd__o22ai_1_265/B1
+ sky130_fd_sc_hd__o22ai_1_257/Y sky130_fd_sc_hd__o21a_1_29/A2 sky130_fd_sc_hd__o22ai_1_261/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_1_3 sky130_fd_sc_hd__inv_2_2/Y sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__nor2_4_2/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_1_909 sky130_fd_sc_hd__nor2_1_218/A sky130_fd_sc_hd__fa_2_1188/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_909/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_268 sky130_fd_sc_hd__nand2_1_410/Y sky130_fd_sc_hd__nand2_1_409/Y
+ sky130_fd_sc_hd__o22ai_1_268/Y sky130_fd_sc_hd__o22ai_1_281/A1 sky130_fd_sc_hd__a21o_2_12/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_279 sky130_fd_sc_hd__nand2_1_410/Y sky130_fd_sc_hd__nand2_1_409/Y
+ sky130_fd_sc_hd__o22ai_1_279/Y sky130_fd_sc_hd__o22ai_1_292/A1 sky130_fd_sc_hd__o21ai_1_337/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__bufinv_8_5 sky130_fd_sc_hd__bufinv_8_6/A sky130_fd_sc_hd__buf_6_46/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufinv_8
Xsky130_fd_sc_hd__dfxtp_1_106 VDD VSS sky130_fd_sc_hd__nor4_1_4/C sky130_fd_sc_hd__dfxtp_1_111/CLK
+ sky130_fd_sc_hd__and2_0_2/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_117 VDD VSS sky130_fd_sc_hd__nor2_1_9/A sky130_fd_sc_hd__dfxtp_1_117/CLK
+ sky130_fd_sc_hd__xor2_1_0/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_128 VDD VSS sky130_fd_sc_hd__buf_2_32/A sky130_fd_sc_hd__clkinv_2_2/Y
+ sky130_fd_sc_hd__and2_0_14/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_139 VDD VSS sky130_fd_sc_hd__ha_2_23/A sky130_fd_sc_hd__dfxtp_1_140/CLK
+ sky130_fd_sc_hd__nor2b_1_10/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_440 VSS VDD sky130_fd_sc_hd__nand2_1_524/B sky130_fd_sc_hd__nor2_1_294/Y
+ sky130_fd_sc_hd__nor2_1_293/B sky130_fd_sc_hd__o21ai_1_440/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_451 VSS VDD sky130_fd_sc_hd__a222oi_1_36/Y sky130_fd_sc_hd__nor2_1_309/A
+ sky130_fd_sc_hd__nand2_1_529/Y sky130_fd_sc_hd__xor2_1_301/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_462 VSS VDD sky130_fd_sc_hd__o22ai_1_436/A2 sky130_fd_sc_hd__nor2_1_303/A
+ sky130_fd_sc_hd__a22oi_1_398/Y sky130_fd_sc_hd__o21ai_1_462/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_473 VSS VDD sky130_fd_sc_hd__o21ai_1_473/A2 sky130_fd_sc_hd__nor2_1_309/A
+ sky130_fd_sc_hd__nand2_1_538/Y sky130_fd_sc_hd__xor2_1_281/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_484 VSS VDD sky130_fd_sc_hd__o22ai_1_432/A2 sky130_fd_sc_hd__nor2_1_308/A
+ sky130_fd_sc_hd__a21oi_1_472/Y sky130_fd_sc_hd__o21ai_1_484/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_495 VSS VDD sky130_fd_sc_hd__nand2_1_556/A sky130_fd_sc_hd__o21ai_1_507/A1
+ sky130_fd_sc_hd__nand2_1_556/Y sky130_fd_sc_hd__and2_0_345/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_1205 sky130_fd_sc_hd__fa_2_1206/CIN sky130_fd_sc_hd__mux2_2_132/A0
+ sky130_fd_sc_hd__fa_2_1205/A sky130_fd_sc_hd__fa_2_1205/B sky130_fd_sc_hd__fa_2_1205/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1216 sky130_fd_sc_hd__fa_2_1217/CIN sky130_fd_sc_hd__mux2_2_160/A1
+ sky130_fd_sc_hd__fa_2_1216/A sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__fa_2_1216/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1227 sky130_fd_sc_hd__fa_2_1228/CIN sky130_fd_sc_hd__mux2_2_210/A1
+ sky130_fd_sc_hd__fa_2_1227/A sky130_fd_sc_hd__fa_2_1227/B sky130_fd_sc_hd__fa_2_1227/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1238 sky130_fd_sc_hd__fa_2_1239/CIN sky130_fd_sc_hd__mux2_2_181/A0
+ sky130_fd_sc_hd__fa_2_1238/A sky130_fd_sc_hd__fa_2_1238/B sky130_fd_sc_hd__fa_2_1238/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1249 sky130_fd_sc_hd__fa_2_1250/CIN sky130_fd_sc_hd__mux2_2_197/A1
+ sky130_fd_sc_hd__fa_2_1249/A sky130_fd_sc_hd__fa_2_1249/B sky130_fd_sc_hd__fa_2_1249/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1002 VDD VSS sky130_fd_sc_hd__mux2_2_116/A0 sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__nor2_1_159/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_11 VSS VDD sky130_fd_sc_hd__o31ai_1_1/Y sky130_fd_sc_hd__or4_1_1/D
+ sky130_fd_sc_hd__o31ai_1_0/Y sky130_fd_sc_hd__o21ai_1_11/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1013 VDD VSS sky130_fd_sc_hd__mux2_2_86/A1 sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__o22ai_1_226/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_22 VSS VDD sky130_fd_sc_hd__a21oi_2_0/Y sky130_fd_sc_hd__nor2_1_11/B
+ sky130_fd_sc_hd__nand2_1_41/Y sky130_fd_sc_hd__o21ai_1_22/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1024 VDD VSS sky130_fd_sc_hd__fa_2_845/A sky130_fd_sc_hd__dfxtp_1_1026/CLK
+ sky130_fd_sc_hd__a21oi_1_313/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_33 VSS VDD sky130_fd_sc_hd__xnor2_1_28/B sky130_fd_sc_hd__nor4_1_7/B
+ sky130_fd_sc_hd__nor4_1_7/A sky130_fd_sc_hd__o31ai_1_3/B1 VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1035 VDD VSS sky130_fd_sc_hd__fa_2_902/CIN sky130_fd_sc_hd__dfxtp_1_1047/CLK
+ sky130_fd_sc_hd__o32ai_1_3/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_44 VSS VDD sky130_fd_sc_hd__o21ai_1_53/A2 sky130_fd_sc_hd__xnor2_1_42/Y
+ sky130_fd_sc_hd__a21oi_1_32/Y sky130_fd_sc_hd__o21ai_1_44/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1046 VDD VSS sky130_fd_sc_hd__fa_2_912/B sky130_fd_sc_hd__dfxtp_1_1050/CLK
+ sky130_fd_sc_hd__a21oi_1_302/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_55 VSS VDD sky130_fd_sc_hd__nand2_2_3/Y sky130_fd_sc_hd__o21ai_1_72/A2
+ sky130_fd_sc_hd__o21ai_1_56/B1 sky130_fd_sc_hd__o21ai_1_55/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1057 VDD VSS sky130_fd_sc_hd__fa_2_1196/A sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__mux2_2_155/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_66 VSS VDD sky130_fd_sc_hd__nand2_2_3/Y sky130_fd_sc_hd__xnor2_1_52/Y
+ sky130_fd_sc_hd__a21oi_1_52/Y sky130_fd_sc_hd__o21ai_1_66/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1068 VDD VSS sky130_fd_sc_hd__fa_2_1207/A sky130_fd_sc_hd__clkinv_8_70/Y
+ sky130_fd_sc_hd__mux2_2_128/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_640 VDD VSS sky130_fd_sc_hd__fa_2_1004/A sky130_fd_sc_hd__clkinv_8_44/Y
+ sky130_fd_sc_hd__mux2_2_24/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_77 VSS VDD sky130_fd_sc_hd__xnor2_1_48/A sky130_fd_sc_hd__o21ai_1_77/A1
+ sky130_fd_sc_hd__o21ai_1_77/B1 sky130_fd_sc_hd__xnor2_1_50/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1079 VDD VSS sky130_fd_sc_hd__fa_2_1181/A sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__mux2_2_147/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_88 VSS VDD sky130_fd_sc_hd__nand4_1_85/Y sky130_fd_sc_hd__fa_2_974/A
+ sky130_fd_sc_hd__fa_2_975/A sky130_fd_sc_hd__o21ai_1_88/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_651 VDD VSS sky130_fd_sc_hd__fa_2_1015/A sky130_fd_sc_hd__clkinv_8_44/Y
+ sky130_fd_sc_hd__mux2_2_1/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_99 VSS VDD sky130_fd_sc_hd__nor2_1_80/Y sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__a21oi_1_86/Y sky130_fd_sc_hd__xor2_1_69/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_662 VDD VSS sky130_fd_sc_hd__fa_2_979/A sky130_fd_sc_hd__clkinv_8_41/Y
+ sky130_fd_sc_hd__mux2_2_31/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_673 VDD VSS sky130_fd_sc_hd__fa_2_990/A sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__mux2_2_7/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_684 VDD VSS sky130_fd_sc_hd__fa_2_1023/A sky130_fd_sc_hd__clkinv_8_59/Y
+ sky130_fd_sc_hd__and2_0_280/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_695 VDD VSS sky130_fd_sc_hd__buf_2_253/A sky130_fd_sc_hd__clkinv_8_41/Y
+ sky130_fd_sc_hd__nor2b_1_94/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_260 VSS VDD sky130_fd_sc_hd__clkbuf_1_260/X sky130_fd_sc_hd__clkbuf_1_260/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_271 VSS VDD sky130_fd_sc_hd__clkbuf_1_271/X sky130_fd_sc_hd__clkbuf_1_271/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_282 VSS VDD sky130_fd_sc_hd__clkbuf_1_282/X sky130_fd_sc_hd__clkbuf_1_282/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_293 VSS VDD sky130_fd_sc_hd__clkbuf_1_293/X sky130_fd_sc_hd__clkbuf_1_293/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_501 sky130_fd_sc_hd__fa_2_499/B sky130_fd_sc_hd__fa_2_495/B
+ sky130_fd_sc_hd__fa_2_551/A sky130_fd_sc_hd__fa_2_543/A sky130_fd_sc_hd__ha_2_121/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_512 sky130_fd_sc_hd__fa_2_514/CIN sky130_fd_sc_hd__fa_2_508/A
+ sky130_fd_sc_hd__fa_2_512/A sky130_fd_sc_hd__fa_2_512/B sky130_fd_sc_hd__fa_2_512/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_523 sky130_fd_sc_hd__fa_2_525/CIN sky130_fd_sc_hd__fa_2_519/A
+ sky130_fd_sc_hd__fa_2_523/A sky130_fd_sc_hd__fa_2_523/B sky130_fd_sc_hd__fa_2_523/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o2bb2ai_1_19 sky130_fd_sc_hd__dfxtp_1_558/D sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__dfxtp_1_558/Q sky130_fd_sc_hd__nor4_1_5/C sky130_fd_sc_hd__nand3_1_45/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_534 sky130_fd_sc_hd__fa_2_538/B sky130_fd_sc_hd__fa_2_534/SUM
+ sky130_fd_sc_hd__fa_2_534/A sky130_fd_sc_hd__fa_2_534/B sky130_fd_sc_hd__fa_2_534/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_545 sky130_fd_sc_hd__fa_2_548/B sky130_fd_sc_hd__fa_2_545/SUM
+ sky130_fd_sc_hd__fa_2_545/A sky130_fd_sc_hd__fa_2_545/B sky130_fd_sc_hd__fa_2_545/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_556 sky130_fd_sc_hd__maj3_1_82/B sky130_fd_sc_hd__maj3_1_83/A
+ sky130_fd_sc_hd__fa_2_556/A sky130_fd_sc_hd__fa_2_556/B sky130_fd_sc_hd__fa_2_557/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_567 sky130_fd_sc_hd__fa_2_565/A sky130_fd_sc_hd__fa_2_567/SUM
+ sky130_fd_sc_hd__fa_2_567/A sky130_fd_sc_hd__fa_2_567/B sky130_fd_sc_hd__fa_2_546/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_578 sky130_fd_sc_hd__fa_2_577/CIN sky130_fd_sc_hd__and2_0_96/A
+ sky130_fd_sc_hd__fa_2_578/A sky130_fd_sc_hd__fa_2_578/B sky130_fd_sc_hd__fa_2_578/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_589 sky130_fd_sc_hd__fa_2_590/B sky130_fd_sc_hd__fa_2_589/SUM
+ sky130_fd_sc_hd__fa_2_683/B sky130_fd_sc_hd__ha_2_126/A sky130_fd_sc_hd__ha_2_132/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_280 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_280/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__and2_0_280/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_291 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_291/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__and2_0_291/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_506 sky130_fd_sc_hd__buf_12_506/A sky130_fd_sc_hd__buf_12_506/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_517 sky130_fd_sc_hd__buf_12_517/A sky130_fd_sc_hd__buf_12_517/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__nand2_1_107 sky130_fd_sc_hd__nand2_1_107/Y sky130_fd_sc_hd__buf_2_270/X
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_706 sky130_fd_sc_hd__clkinv_1_706/Y sky130_fd_sc_hd__nor2_1_130/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_706/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_118 sky130_fd_sc_hd__nand2_1_118/Y sky130_fd_sc_hd__fa_2_702/SUM
+ sky130_fd_sc_hd__and2_0_235/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_717 sky130_fd_sc_hd__nand4_1_86/A sky130_fd_sc_hd__fa_2_1049/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_717/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_129 sky130_fd_sc_hd__nand2_1_129/Y sky130_fd_sc_hd__nand2_1_130/Y
+ sky130_fd_sc_hd__buf_2_264/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_728 sky130_fd_sc_hd__clkinv_1_728/Y sky130_fd_sc_hd__a21oi_1_238/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_728/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_739 sky130_fd_sc_hd__nor2_1_137/A sky130_fd_sc_hd__fa_2_1087/A
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_270 VSS VDD sky130_fd_sc_hd__o21ai_1_270/A2 sky130_fd_sc_hd__o22ai_1_206/A1
+ sky130_fd_sc_hd__a22oi_1_366/Y sky130_fd_sc_hd__a21o_2_4/B1 VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_281 VSS VDD sky130_fd_sc_hd__nand2_1_371/B sky130_fd_sc_hd__nor2_1_170/Y
+ sky130_fd_sc_hd__a21o_2_9/A2 sky130_fd_sc_hd__o21ai_1_281/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkinv_8_9 sky130_fd_sc_hd__clkinv_8_9/Y sky130_fd_sc_hd__clkinv_8_9/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_9/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__o21ai_1_292 VSS VDD sky130_fd_sc_hd__nor2_1_175/B sky130_fd_sc_hd__nor2_1_182/A
+ sky130_fd_sc_hd__a21oi_1_263/Y sky130_fd_sc_hd__xor2_1_169/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor3_1_17 sky130_fd_sc_hd__nor3_1_17/C sky130_fd_sc_hd__nor3_1_17/Y
+ sky130_fd_sc_hd__nor3_2_5/A sky130_fd_sc_hd__nor3_2_6/A VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_28 sky130_fd_sc_hd__xor2_1_17/X sky130_fd_sc_hd__nor3_1_28/Y
+ sky130_fd_sc_hd__nor3_1_28/A sky130_fd_sc_hd__nor3_1_28/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_39 sky130_fd_sc_hd__nor3_1_39/C sky130_fd_sc_hd__nor3_1_39/Y
+ sky130_fd_sc_hd__nor3_1_39/A sky130_fd_sc_hd__nor3_1_39/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__fa_2_1002 sky130_fd_sc_hd__fa_2_1003/CIN sky130_fd_sc_hd__mux2_2_29/A1
+ sky130_fd_sc_hd__fa_2_1002/A sky130_fd_sc_hd__xor2_1_74/X sky130_fd_sc_hd__fa_2_1002/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1013 sky130_fd_sc_hd__fa_2_1014/CIN sky130_fd_sc_hd__mux2_2_6/A0
+ sky130_fd_sc_hd__fa_2_1013/A sky130_fd_sc_hd__xor2_1_63/X sky130_fd_sc_hd__fa_2_1013/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1024 sky130_fd_sc_hd__fa_2_1025/CIN sky130_fd_sc_hd__and2_0_281/A
+ sky130_fd_sc_hd__fa_2_1024/A sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_1024/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1035 sky130_fd_sc_hd__fa_2_1036/CIN sky130_fd_sc_hd__fa_2_1035/SUM
+ sky130_fd_sc_hd__fa_2_1035/A sky130_fd_sc_hd__nor2_1_53/A sky130_fd_sc_hd__fa_2_1035/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1046 sky130_fd_sc_hd__fa_2_1047/CIN sky130_fd_sc_hd__and2_0_301/A
+ sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1046/B sky130_fd_sc_hd__xor2_1_111/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1057 sky130_fd_sc_hd__fa_2_1058/CIN sky130_fd_sc_hd__mux2_2_63/A0
+ sky130_fd_sc_hd__fa_2_1057/A sky130_fd_sc_hd__fa_2_1057/B sky130_fd_sc_hd__fa_2_1057/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1068 sky130_fd_sc_hd__xor2_1_86/B sky130_fd_sc_hd__mux2_2_41/A0
+ sky130_fd_sc_hd__fa_2_1068/A sky130_fd_sc_hd__xor2_1_89/X sky130_fd_sc_hd__fa_2_1068/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1079 sky130_fd_sc_hd__fa_2_1080/CIN sky130_fd_sc_hd__mux2_2_64/A0
+ sky130_fd_sc_hd__fa_2_1079/A sky130_fd_sc_hd__fa_2_1079/B sky130_fd_sc_hd__fa_2_1079/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_11 sky130_fd_sc_hd__inv_2_11/A sky130_fd_sc_hd__inv_2_11/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_22 sky130_fd_sc_hd__inv_2_22/A sky130_fd_sc_hd__inv_2_22/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_33 sky130_fd_sc_hd__inv_2_33/A sky130_fd_sc_hd__buf_8_3/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_44 sky130_fd_sc_hd__inv_2_44/A sky130_fd_sc_hd__inv_2_44/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_55 sky130_fd_sc_hd__inv_2_55/A sky130_fd_sc_hd__inv_2_55/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_66 sky130_fd_sc_hd__inv_2_66/A sky130_fd_sc_hd__inv_2_66/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_470 VDD VSS sky130_fd_sc_hd__buf_2_2/A sky130_fd_sc_hd__dfxtp_1_472/CLK
+ sky130_fd_sc_hd__and2_0_121/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_77 sky130_fd_sc_hd__inv_2_77/A sky130_fd_sc_hd__inv_2_77/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_481 VDD VSS sky130_fd_sc_hd__nor2_1_40/B sky130_fd_sc_hd__dfxtp_1_483/CLK
+ sky130_fd_sc_hd__nor2b_1_68/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_2_1 sky130_fd_sc_hd__nand2_2_1/Y sky130_fd_sc_hd__nor2_1_6/Y
+ sky130_fd_sc_hd__or2_1_2/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__inv_2_88 sky130_fd_sc_hd__inv_2_88/A sky130_fd_sc_hd__inv_2_88/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_492 VDD VSS sky130_fd_sc_hd__o21ai_1_39/A1 sky130_fd_sc_hd__dfxtp_1_496/CLK
+ sky130_fd_sc_hd__nor2b_1_59/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_99 sky130_fd_sc_hd__inv_2_99/A sky130_fd_sc_hd__inv_2_99/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__fa_2_320 sky130_fd_sc_hd__fa_2_317/B sky130_fd_sc_hd__fa_2_321/CIN
+ sky130_fd_sc_hd__fa_2_320/A sky130_fd_sc_hd__fa_2_320/B sky130_fd_sc_hd__fa_2_320/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_331 sky130_fd_sc_hd__maj3_1_75/B sky130_fd_sc_hd__maj3_1_76/A
+ sky130_fd_sc_hd__fa_2_331/A sky130_fd_sc_hd__fa_2_331/B sky130_fd_sc_hd__fa_2_332/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_342 sky130_fd_sc_hd__fa_2_344/CIN sky130_fd_sc_hd__fa_2_340/A
+ sky130_fd_sc_hd__ha_2_115/B sky130_fd_sc_hd__fa_2_395/A sky130_fd_sc_hd__fa_2_342/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_353 sky130_fd_sc_hd__fa_2_356/B sky130_fd_sc_hd__fa_2_353/SUM
+ sky130_fd_sc_hd__fa_2_353/A sky130_fd_sc_hd__fa_2_353/B sky130_fd_sc_hd__fa_2_353/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_364 sky130_fd_sc_hd__fa_2_365/B sky130_fd_sc_hd__fa_2_357/A
+ sky130_fd_sc_hd__ha_2_109/B sky130_fd_sc_hd__ha_2_113/B sky130_fd_sc_hd__fa_2_413/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_375 sky130_fd_sc_hd__fa_2_376/B sky130_fd_sc_hd__fa_2_367/A
+ sky130_fd_sc_hd__fa_2_404/A sky130_fd_sc_hd__ha_2_114/A sky130_fd_sc_hd__fa_2_360/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_16 sky130_fd_sc_hd__conb_1_10/LO sky130_fd_sc_hd__clkinv_4_63/Y
+ sky130_fd_sc_hd__dfxtp_1_155/CLK sky130_fd_sc_hd__nand2b_1_1/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_386 sky130_fd_sc_hd__fa_2_388/CIN sky130_fd_sc_hd__fa_2_382/A
+ sky130_fd_sc_hd__fa_2_386/A sky130_fd_sc_hd__fa_2_386/B sky130_fd_sc_hd__fa_2_386/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_27 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_96/A
+ sky130_fd_sc_hd__dfxtp_1_463/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__and2_1_2 VDD VSS sky130_fd_sc_hd__inv_2_96/A sky130_fd_sc_hd__ha_2_52/A
+ sky130_fd_sc_hd__nor2_4_2/Y VDD VSS sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__fa_2_397 sky130_fd_sc_hd__fa_2_402/B sky130_fd_sc_hd__fa_2_397/SUM
+ sky130_fd_sc_hd__fa_2_397/A sky130_fd_sc_hd__fa_2_397/B sky130_fd_sc_hd__fa_2_397/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22oi_2_8 sky130_fd_sc_hd__nor2_4_5/Y sky130_fd_sc_hd__a22oi_2_8/A2
+ sky130_fd_sc_hd__a22oi_2_9/B1 sky130_fd_sc_hd__a22oi_2_8/B2 sky130_fd_sc_hd__a22oi_2_8/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__diode_2_203 sky130_fd_sc_hd__buf_2_267/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__sdlclkp_4_38 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_100/Y
+ sky130_fd_sc_hd__dfxtp_1_325/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__diode_2_214 amplitude_adc_done VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__sdlclkp_4_49 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_4_53/Y
+ sky130_fd_sc_hd__dfxtp_1_448/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__diode_2_225 sig_amplitude[0] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkinv_8_80 sky130_fd_sc_hd__clkinv_8_80/Y sky130_fd_sc_hd__clkinv_8_80/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_80/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_91 sky130_fd_sc_hd__clkinv_8_97/A sky130_fd_sc_hd__clkinv_8_91/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_91/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__nor2_1_107 sky130_fd_sc_hd__nor2_1_107/B sky130_fd_sc_hd__nor2_1_107/Y
+ sky130_fd_sc_hd__fa_2_1110/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_118 sky130_fd_sc_hd__nor2_1_118/B sky130_fd_sc_hd__nor2_1_118/Y
+ sky130_fd_sc_hd__o21a_1_14/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_129 sky130_fd_sc_hd__nor2_1_129/B sky130_fd_sc_hd__nor2_1_129/Y
+ sky130_fd_sc_hd__nor2_1_129/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_16 sky130_fd_sc_hd__nor2_2_0/Y sky130_fd_sc_hd__clkinv_1_4/Y
+ sky130_fd_sc_hd__nand4_1_23/Y sky130_fd_sc_hd__nand4_1_7/Y sky130_fd_sc_hd__a22oi_1_16/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_27 sky130_fd_sc_hd__nor2_2_0/Y sky130_fd_sc_hd__clkinv_1_4/Y
+ sky130_fd_sc_hd__nand4_1_16/Y sky130_fd_sc_hd__nand4_1_0/Y sky130_fd_sc_hd__a22oi_1_27/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_38 sky130_fd_sc_hd__a22oi_2_9/B1 sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__clkbuf_4_39/X sky130_fd_sc_hd__a22oi_1_38/A2 sky130_fd_sc_hd__a22oi_1_38/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_49 sky130_fd_sc_hd__clkbuf_4_8/X sky130_fd_sc_hd__clkbuf_4_9/X
+ sky130_fd_sc_hd__clkbuf_1_28/X sky130_fd_sc_hd__a22oi_1_49/A2 sky130_fd_sc_hd__a22oi_1_49/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_303 sky130_fd_sc_hd__buf_8_150/X sky130_fd_sc_hd__buf_12_303/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_314 sky130_fd_sc_hd__buf_4_84/X sky130_fd_sc_hd__buf_12_314/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_325 sky130_fd_sc_hd__buf_4_79/X sky130_fd_sc_hd__buf_12_325/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_336 sky130_fd_sc_hd__buf_4_75/X sky130_fd_sc_hd__buf_12_336/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_347 sky130_fd_sc_hd__buf_4_97/X sky130_fd_sc_hd__buf_12_369/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_206 sky130_fd_sc_hd__clkbuf_1_264/X sky130_fd_sc_hd__nor2_2_3/Y
+ sky130_fd_sc_hd__a22oi_1_206/B2 sky130_fd_sc_hd__clkbuf_4_123/X sky130_fd_sc_hd__nand4_1_46/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_358 sky130_fd_sc_hd__buf_12_358/A sky130_fd_sc_hd__buf_12_358/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_217 sky130_fd_sc_hd__buf_2_166/X sky130_fd_sc_hd__buf_2_167/X
+ sky130_fd_sc_hd__clkbuf_1_436/X sky130_fd_sc_hd__buf_2_181/X sky130_fd_sc_hd__nand4_1_50/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_369 sky130_fd_sc_hd__buf_12_369/A sky130_fd_sc_hd__buf_12_369/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_228 sky130_fd_sc_hd__nor3_1_19/Y sky130_fd_sc_hd__nor3_1_20/Y
+ sky130_fd_sc_hd__clkbuf_1_434/X sky130_fd_sc_hd__buf_2_177/X sky130_fd_sc_hd__nand4_1_54/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_239 sky130_fd_sc_hd__buf_2_166/X sky130_fd_sc_hd__buf_2_167/X
+ sky130_fd_sc_hd__clkbuf_1_499/X sky130_fd_sc_hd__buf_2_173/X sky130_fd_sc_hd__nand4_1_58/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_503 sky130_fd_sc_hd__o21ai_1_79/A1 sky130_fd_sc_hd__o21ai_1_86/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_503/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_514 sky130_fd_sc_hd__nor2_1_55/B sky130_fd_sc_hd__fa_2_1031/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_514/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_525 sky130_fd_sc_hd__nor2_1_61/B sky130_fd_sc_hd__fa_2_1042/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_525/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_536 sky130_fd_sc_hd__nand2_1_262/A sky130_fd_sc_hd__a222oi_1_0/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_536/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_547 sky130_fd_sc_hd__o22ai_1_110/B1 sky130_fd_sc_hd__fa_2_986/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_547/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_558 sky130_fd_sc_hd__nor2_1_68/B sky130_fd_sc_hd__fa_2_980/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_558/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_569 sky130_fd_sc_hd__clkinv_1_569/Y sky130_fd_sc_hd__nor2_1_73/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_569/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_50 sky130_fd_sc_hd__nor2_1_50/B sky130_fd_sc_hd__nor2_1_50/Y
+ sky130_fd_sc_hd__nor2_1_50/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_61 sky130_fd_sc_hd__nor2_1_61/B sky130_fd_sc_hd__nor2_1_61/Y
+ sky130_fd_sc_hd__nor2_1_61/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_16 sky130_fd_sc_hd__clkinv_4_16/A sky130_fd_sc_hd__inv_16_6/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_16/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_72 sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_1_72/Y
+ sky130_fd_sc_hd__nor2_2_9/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_27 sky130_fd_sc_hd__clkinv_4_27/A sky130_fd_sc_hd__clkinv_4_27/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_27/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_83 sky130_fd_sc_hd__nor2_1_83/B sky130_fd_sc_hd__nor2_1_83/Y
+ sky130_fd_sc_hd__nor2_1_83/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_38 sky130_fd_sc_hd__clkinv_4_38/A sky130_fd_sc_hd__buf_6_55/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_38/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_94 sky130_fd_sc_hd__nor2_1_94/B sky130_fd_sc_hd__nor2_1_94/Y
+ sky130_fd_sc_hd__nor2_1_94/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_49 sky130_fd_sc_hd__clkinv_4_49/A sky130_fd_sc_hd__clkinv_4_50/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_49/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_sram_2kbyte_1rw1r_32x512_8_2 sky130_fd_sc_hd__buf_6_1/X sky130_fd_sc_hd__clkbuf_4_0/X
+ sky130_fd_sc_hd__buf_4_2/X sky130_fd_sc_hd__buf_4_3/X sky130_fd_sc_hd__buf_4_5/X
+ sky130_fd_sc_hd__buf_6_4/X sky130_fd_sc_hd__buf_4_7/X sky130_fd_sc_hd__buf_6_6/X
+ sky130_fd_sc_hd__clkbuf_4_1/X sky130_fd_sc_hd__buf_4_8/X sky130_fd_sc_hd__buf_4_9/X
+ sky130_fd_sc_hd__clkbuf_4_5/X sky130_fd_sc_hd__clkbuf_4_6/X sky130_fd_sc_hd__buf_4_11/X
+ sky130_fd_sc_hd__buf_12_0/X sky130_fd_sc_hd__buf_6_9/X sky130_fd_sc_hd__buf_6_1/X
+ sky130_fd_sc_hd__clkbuf_4_0/X sky130_fd_sc_hd__buf_4_2/X sky130_fd_sc_hd__buf_4_3/X
+ sky130_fd_sc_hd__buf_4_5/X sky130_fd_sc_hd__buf_6_4/X sky130_fd_sc_hd__buf_4_7/X
+ sky130_fd_sc_hd__buf_6_6/X sky130_fd_sc_hd__clkbuf_4_1/X sky130_fd_sc_hd__buf_4_8/X
+ sky130_fd_sc_hd__buf_4_9/X sky130_fd_sc_hd__clkbuf_4_5/X sky130_fd_sc_hd__clkbuf_4_6/X
+ sky130_fd_sc_hd__buf_4_11/X sky130_fd_sc_hd__buf_12_0/X sky130_fd_sc_hd__buf_6_9/X
+ sky130_fd_sc_hd__buf_12_39/X sky130_fd_sc_hd__buf_8_61/X sky130_fd_sc_hd__buf_12_92/X
+ sky130_fd_sc_hd__buf_12_90/X sky130_fd_sc_hd__buf_12_119/X sky130_fd_sc_hd__buf_12_91/X
+ sky130_fd_sc_hd__buf_12_55/X sky130_fd_sc_hd__buf_12_28/X sky130_fd_sc_hd__buf_12_27/X
+ sky130_fd_sc_hd__buf_12_5/X sky130_fd_sc_hd__buf_12_23/X sky130_fd_sc_hd__buf_12_120/X
+ sky130_fd_sc_hd__buf_12_118/X sky130_fd_sc_hd__buf_12_117/X sky130_fd_sc_hd__buf_12_60/X
+ sky130_fd_sc_hd__buf_12_38/X sky130_fd_sc_hd__buf_12_98/X sky130_fd_sc_hd__buf_12_96/X
+ sky130_fd_sc_hd__clkbuf_1_71/X sky130_fd_sc_hd__clkbuf_1_89/X sky130_fd_sc_hd__clkbuf_1_71/X
+ sky130_fd_sc_hd__clkinv_8_1/Y sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__buf_12_101/X
+ sky130_fd_sc_hd__buf_8_62/X sky130_fd_sc_hd__buf_12_88/X sky130_fd_sc_hd__buf_12_34/X
+ sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[0] sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[1]
+ sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[2] sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[3]
+ sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[4] sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[5]
+ sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[6] sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[7]
+ sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[8] sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[9]
+ sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[10] sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[11]
+ sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[12] sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[13]
+ sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[14] sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[15]
+ sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[16] sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[17]
+ sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[18] sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[19]
+ sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[20] sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[21]
+ sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[22] sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[23]
+ sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[24] sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[25]
+ sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[26] sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[27]
+ sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[28] sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[29]
+ sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[30] sky130_sram_2kbyte_1rw1r_32x512_8_2/dout0[31]
+ sky130_fd_sc_hd__clkbuf_4_10/A sky130_fd_sc_hd__clkbuf_4_11/A sky130_fd_sc_hd__clkbuf_4_12/A
+ sky130_fd_sc_hd__clkbuf_4_13/A sky130_fd_sc_hd__clkbuf_4_14/A sky130_fd_sc_hd__clkbuf_4_15/A
+ sky130_fd_sc_hd__clkbuf_4_16/A sky130_fd_sc_hd__clkbuf_4_17/A sky130_fd_sc_hd__clkbuf_4_18/A
+ sky130_fd_sc_hd__clkbuf_4_19/A sky130_fd_sc_hd__clkbuf_4_20/A sky130_fd_sc_hd__clkbuf_4_21/A
+ sky130_fd_sc_hd__clkbuf_4_22/A sky130_fd_sc_hd__clkbuf_4_23/A sky130_fd_sc_hd__clkbuf_4_24/A
+ sky130_fd_sc_hd__clkbuf_4_25/A sky130_fd_sc_hd__clkbuf_4_26/A sky130_fd_sc_hd__clkbuf_4_27/A
+ sky130_fd_sc_hd__clkbuf_4_28/A sky130_fd_sc_hd__clkbuf_4_29/A sky130_fd_sc_hd__clkbuf_4_30/A
+ sky130_fd_sc_hd__clkbuf_4_31/A sky130_fd_sc_hd__clkbuf_4_32/A sky130_fd_sc_hd__clkbuf_4_33/A
+ sky130_fd_sc_hd__clkbuf_4_34/A sky130_fd_sc_hd__clkbuf_4_35/A sky130_fd_sc_hd__clkbuf_4_36/A
+ sky130_fd_sc_hd__clkbuf_4_37/A sky130_fd_sc_hd__clkbuf_4_38/A sky130_fd_sc_hd__clkbuf_4_39/A
+ sky130_fd_sc_hd__clkbuf_4_40/A sky130_fd_sc_hd__clkbuf_4_41/A VDD VSS sky130_sram_2kbyte_1rw1r_32x512_8
Xsky130_fd_sc_hd__a21oi_1_400 sky130_fd_sc_hd__fa_2_1234/A sky130_fd_sc_hd__o22ai_1_366/Y
+ sky130_fd_sc_hd__a21oi_1_400/Y sky130_fd_sc_hd__nor2_2_17/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_411 sky130_fd_sc_hd__or2_0_11/B sky130_fd_sc_hd__o21ai_1_429/Y
+ sky130_fd_sc_hd__a21oi_1_411/Y sky130_fd_sc_hd__o21ai_1_430/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_422 sky130_fd_sc_hd__o21a_1_58/B1 sky130_fd_sc_hd__o21a_1_57/A1
+ sky130_fd_sc_hd__a21oi_1_422/Y sky130_fd_sc_hd__nor2_1_270/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_433 sky130_fd_sc_hd__nor2_1_281/A sky130_fd_sc_hd__o21a_1_66/A1
+ sky130_fd_sc_hd__a21oi_1_433/Y sky130_fd_sc_hd__nor2_1_281/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_444 sky130_fd_sc_hd__a21oi_1_447/A1 sky130_fd_sc_hd__a21oi_1_444/B1
+ sky130_fd_sc_hd__a21oi_1_444/Y sky130_fd_sc_hd__nand2_1_543/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_455 sky130_fd_sc_hd__fa_2_1283/A sky130_fd_sc_hd__o22ai_1_417/Y
+ sky130_fd_sc_hd__a21oi_1_455/Y sky130_fd_sc_hd__nor2_2_18/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_466 sky130_fd_sc_hd__o21ai_1_484/Y sky130_fd_sc_hd__o21ai_1_479/Y
+ sky130_fd_sc_hd__a21oi_1_466/Y sky130_fd_sc_hd__nor2b_1_126/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_477 sky130_fd_sc_hd__a22oi_1_400/B1 sky130_fd_sc_hd__o22ai_1_434/Y
+ sky130_fd_sc_hd__a21oi_1_477/Y sky130_fd_sc_hd__fa_2_1308/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_488 sky130_fd_sc_hd__nor2_1_319/Y sky130_fd_sc_hd__or2_0_0/B
+ sky130_fd_sc_hd__nand2_1_556/A sky130_fd_sc_hd__nor2_1_322/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_8_102 sky130_fd_sc_hd__clkinv_8_102/Y sky130_fd_sc_hd__clkinv_8_63/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_102/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__a21oi_1_499 sky130_fd_sc_hd__nor2_1_318/Y sky130_fd_sc_hd__or2_0_0/B
+ sky130_fd_sc_hd__nand2_1_567/A sky130_fd_sc_hd__or2_0_13/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_8_113 sky130_fd_sc_hd__dfxtp_1_83/CLK sky130_fd_sc_hd__clkinv_8_15/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_113/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_124 sky130_fd_sc_hd__clkinv_8_124/Y sky130_fd_sc_hd__clkinv_8_6/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_135 sky130_fd_sc_hd__clkinv_8_136/A sky130_fd_sc_hd__clkinv_8_135/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__o21a_1_4 sky130_fd_sc_hd__o21a_1_4/X sky130_fd_sc_hd__o21a_1_4/A1
+ sky130_fd_sc_hd__o21a_1_4/B1 sky130_fd_sc_hd__fa_2_984/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__nand2_1_460 sky130_fd_sc_hd__o32ai_1_8/B1 sky130_fd_sc_hd__o32ai_1_8/A3
+ sky130_fd_sc_hd__o21bai_1_4/A2 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_471 sky130_fd_sc_hd__o31ai_1_9/A1 sky130_fd_sc_hd__nand2_1_471/B
+ sky130_fd_sc_hd__nor2_1_251/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_482 sky130_fd_sc_hd__nand2_1_482/Y sky130_fd_sc_hd__nand2_1_491/B
+ sky130_fd_sc_hd__o21ai_1_402/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_493 sky130_fd_sc_hd__nand2_1_493/Y sky130_fd_sc_hd__nor2b_1_119/Y
+ sky130_fd_sc_hd__o21ai_1_431/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_40 sky130_fd_sc_hd__ha_2_80/SUM sky130_fd_sc_hd__nor2b_1_40/Y
+ sky130_fd_sc_hd__or2_0_3/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_51 sky130_fd_sc_hd__nor2_1_22/A sky130_fd_sc_hd__nor2b_1_51/Y
+ sky130_fd_sc_hd__o21ai_1_9/A2 VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_62 sky130_fd_sc_hd__nor2_1_36/B sky130_fd_sc_hd__nor2b_1_62/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_73 sky130_fd_sc_hd__nor4_1_12/B sky130_fd_sc_hd__nor2b_1_73/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1040 sky130_fd_sc_hd__o32ai_1_9/A2 sky130_fd_sc_hd__fa_2_1275/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1040/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_84 sky130_fd_sc_hd__nor2b_1_85/A sky130_fd_sc_hd__nor2b_1_84/Y
+ sky130_fd_sc_hd__fa_2_953/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1051 sky130_fd_sc_hd__o22ai_1_397/A1 sky130_fd_sc_hd__fa_2_7/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1051/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1062 sky130_fd_sc_hd__nor2_1_275/B sky130_fd_sc_hd__fa_2_1279/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1062/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_95 sky130_fd_sc_hd__o22ai_1_90/Y sky130_fd_sc_hd__nor2b_1_95/Y
+ sky130_fd_sc_hd__buf_2_262/X VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__xnor2_1_3 VSS VDD sky130_fd_sc_hd__xnor2_1_3/B sky130_fd_sc_hd__xnor2_1_3/Y
+ sky130_fd_sc_hd__xnor2_1_3/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_1073 sky130_fd_sc_hd__o22ai_1_415/A1 sky130_fd_sc_hd__o21ai_1_460/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1073/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1084 sky130_fd_sc_hd__nor2_1_274/B sky130_fd_sc_hd__fa_2_1281/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1084/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1095 sky130_fd_sc_hd__o22ai_1_430/B1 sky130_fd_sc_hd__fa_2_1310/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1095/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_150 sky130_fd_sc_hd__fa_2_143/CIN sky130_fd_sc_hd__nor2_1_254/A
+ sky130_fd_sc_hd__fa_2_150/A sky130_fd_sc_hd__fa_2_150/B sky130_fd_sc_hd__fa_2_150/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_161 sky130_fd_sc_hd__fa_2_158/CIN sky130_fd_sc_hd__nor2_1_255/A
+ sky130_fd_sc_hd__fa_2_161/A sky130_fd_sc_hd__fa_2_161/B sky130_fd_sc_hd__fa_2_161/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_18 VDD VSS sky130_fd_sc_hd__fa_2_360/B sky130_fd_sc_hd__dfxtp_1_26/CLK
+ sky130_fd_sc_hd__nand4_1_36/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_172 sky130_fd_sc_hd__maj3_1_55/B sky130_fd_sc_hd__fa_2_172/SUM
+ sky130_fd_sc_hd__fa_2_67/B sky130_fd_sc_hd__ha_2_93/A sky130_fd_sc_hd__ha_2_99/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_29 VDD VSS sky130_fd_sc_hd__ha_2_108/B sky130_fd_sc_hd__dfxtp_1_29/CLK
+ sky130_fd_sc_hd__nand4_1_47/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_183 sky130_fd_sc_hd__maj3_1_48/B sky130_fd_sc_hd__maj3_1_49/A
+ sky130_fd_sc_hd__fa_2_183/A sky130_fd_sc_hd__fa_2_183/B sky130_fd_sc_hd__fa_2_184/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_194 sky130_fd_sc_hd__fa_2_197/CIN sky130_fd_sc_hd__fa_2_192/B
+ sky130_fd_sc_hd__fa_2_15/B sky130_fd_sc_hd__fa_2_194/B sky130_fd_sc_hd__fa_2_194/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o22ai_1_60 sky130_fd_sc_hd__o22ai_1_60/A2 sky130_fd_sc_hd__fa_2_965/A
+ sky130_fd_sc_hd__o22ai_1_60/Y sky130_fd_sc_hd__fa_2_966/A sky130_fd_sc_hd__o22ai_1_60/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_71 sky130_fd_sc_hd__o22ai_1_88/B1 sky130_fd_sc_hd__nand2_2_3/Y
+ sky130_fd_sc_hd__o22ai_1_71/Y sky130_fd_sc_hd__xnor2_1_53/Y sky130_fd_sc_hd__o22ai_1_85/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkbuf_4_108 sky130_fd_sc_hd__clkbuf_4_108/X sky130_fd_sc_hd__dfxtp_1_1450/Q
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o22ai_1_82 sky130_fd_sc_hd__o22ai_1_89/A1 sky130_fd_sc_hd__o22ai_1_88/B1
+ sky130_fd_sc_hd__o22ai_1_82/Y sky130_fd_sc_hd__xnor2_1_47/Y sky130_fd_sc_hd__o22ai_1_82/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkbuf_4_119 sky130_fd_sc_hd__clkbuf_4_119/X sky130_fd_sc_hd__clkbuf_4_119/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o22ai_1_93 sky130_fd_sc_hd__nor2_2_9/B sky130_fd_sc_hd__nor2_1_76/A
+ sky130_fd_sc_hd__o22ai_1_93/Y sky130_fd_sc_hd__o22ai_1_99/A2 sky130_fd_sc_hd__nor2_1_84/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_4_40 VDD VSS sky130_fd_sc_hd__buf_4_40/X sky130_fd_sc_hd__buf_4_40/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_51 VDD VSS sky130_fd_sc_hd__buf_4_51/X sky130_fd_sc_hd__buf_4_51/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_62 VDD VSS sky130_fd_sc_hd__buf_4_62/X sky130_fd_sc_hd__buf_4_62/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_73 VDD VSS sky130_fd_sc_hd__buf_4_73/X sky130_fd_sc_hd__buf_4_73/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_84 VDD VSS sky130_fd_sc_hd__buf_4_84/X sky130_fd_sc_hd__buf_4_84/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_95 VDD VSS sky130_fd_sc_hd__buf_4_95/X sky130_fd_sc_hd__buf_4_95/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_12_100 sky130_fd_sc_hd__buf_12_42/X sky130_fd_sc_hd__buf_12_100/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_111 sky130_fd_sc_hd__buf_12_111/A sky130_fd_sc_hd__buf_12_111/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_122 sky130_fd_sc_hd__buf_2_37/X sky130_fd_sc_hd__buf_12_122/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_133 sky130_fd_sc_hd__buf_12_133/A sky130_fd_sc_hd__buf_12_240/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_144 sky130_fd_sc_hd__buf_12_144/A sky130_fd_sc_hd__buf_12_250/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_155 sky130_fd_sc_hd__buf_4_43/A sky130_fd_sc_hd__buf_12_201/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_166 sky130_fd_sc_hd__buf_8_85/X sky130_fd_sc_hd__buf_12_166/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_4_3 sky130_fd_sc_hd__clkbuf_4_3/X sky130_fd_sc_hd__buf_2_7/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_12_177 sky130_fd_sc_hd__buf_8_93/X sky130_fd_sc_hd__buf_12_177/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_188 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__buf_12_188/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_199 sky130_fd_sc_hd__buf_4_42/X sky130_fd_sc_hd__buf_12_244/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_300 sky130_fd_sc_hd__fa_2_250/A sky130_fd_sc_hd__fa_2_242/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_300/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_311 sky130_fd_sc_hd__fa_2_424/B sky130_fd_sc_hd__fa_2_404/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_311/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_322 sky130_fd_sc_hd__fa_2_416/B sky130_fd_sc_hd__ha_2_110/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_322/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_333 sky130_fd_sc_hd__fa_2_537/A sky130_fd_sc_hd__ha_2_123/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_333/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_344 sky130_fd_sc_hd__fa_2_692/A sky130_fd_sc_hd__fa_2_700/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_344/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_355 sky130_fd_sc_hd__fa_2_817/B sky130_fd_sc_hd__fa_2_793/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_355/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_366 sky130_fd_sc_hd__ha_2_142/A sky130_fd_sc_hd__fa_2_820/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_366/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_377 sky130_fd_sc_hd__fa_2_871/B sky130_fd_sc_hd__dfxtp_1_271/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_377/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_388 sky130_fd_sc_hd__fa_2_884/B sky130_fd_sc_hd__nand2_1_36/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_388/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_399 sky130_fd_sc_hd__nand2_1_204/B sky130_fd_sc_hd__nand2_1_36/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_399/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21a_1_18 sky130_fd_sc_hd__o21a_1_18/X sky130_fd_sc_hd__o21a_1_18/A1
+ sky130_fd_sc_hd__o21a_1_18/B1 sky130_fd_sc_hd__fa_2_1136/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_29 sky130_fd_sc_hd__o21a_1_29/X sky130_fd_sc_hd__o21a_1_29/A1
+ sky130_fd_sc_hd__o21a_1_29/B1 sky130_fd_sc_hd__o21a_1_29/A2 VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__a21oi_1_230 sky130_fd_sc_hd__a21o_2_5/A2 sky130_fd_sc_hd__o21ai_1_265/Y
+ sky130_fd_sc_hd__a21oi_1_230/Y sky130_fd_sc_hd__fa_2_1074/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_241 sky130_fd_sc_hd__o21a_1_18/B1 sky130_fd_sc_hd__o21a_1_17/A1
+ sky130_fd_sc_hd__dfxtp_1_907/D sky130_fd_sc_hd__nor2_1_176/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_252 sky130_fd_sc_hd__o21a_1_27/B1 sky130_fd_sc_hd__o21a_1_26/A1
+ sky130_fd_sc_hd__dfxtp_1_885/D sky130_fd_sc_hd__nor2_1_153/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_263 sky130_fd_sc_hd__o21ai_1_298/Y sky130_fd_sc_hd__clkinv_1_818/Y
+ sky130_fd_sc_hd__a21oi_1_263/Y sky130_fd_sc_hd__nor2b_1_104/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_274 sky130_fd_sc_hd__fa_2_1136/A sky130_fd_sc_hd__o22ai_1_245/Y
+ sky130_fd_sc_hd__a21oi_1_274/Y sky130_fd_sc_hd__nor3_1_38/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_285 sky130_fd_sc_hd__fa_2_1154/A sky130_fd_sc_hd__o22ai_1_254/Y
+ sky130_fd_sc_hd__a21oi_1_285/Y sky130_fd_sc_hd__clkinv_1_779/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_4_3 sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__buf_12_23/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_3/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__a21oi_1_296 sky130_fd_sc_hd__fa_2_1146/A sky130_fd_sc_hd__o22ai_1_261/Y
+ sky130_fd_sc_hd__a21oi_1_296/Y sky130_fd_sc_hd__nor3_1_38/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_204 sky130_fd_sc_hd__buf_8_204/A sky130_fd_sc_hd__buf_8_204/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_215 sky130_fd_sc_hd__inv_2_133/Y sky130_fd_sc_hd__buf_8_215/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__xor2_1_107 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1050/B
+ sky130_fd_sc_hd__xor2_1_107/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_290 sky130_fd_sc_hd__xnor2_1_77/B sky130_fd_sc_hd__nand2_1_290/B
+ sky130_fd_sc_hd__nand2_1_297/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_118 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1088/B
+ sky130_fd_sc_hd__xor2_1_118/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_129 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1077/B
+ sky130_fd_sc_hd__xor2_1_129/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_1409 VDD VSS sky130_fd_sc_hd__mux2_2_223/A1 sky130_fd_sc_hd__clkinv_8_75/Y
+ sky130_fd_sc_hd__o31ai_1_12/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_109 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_109/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_850/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_17 sky130_fd_sc_hd__nand3_2_0/C sky130_fd_sc_hd__xor2_1_2/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_17/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_28 sky130_fd_sc_hd__inv_2_17/A sky130_fd_sc_hd__ha_2_26/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_28/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_39 sky130_fd_sc_hd__inv_2_28/A sky130_fd_sc_hd__buf_2_12/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_39/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_4 sky130_fd_sc_hd__fa_2_3/CIN sky130_fd_sc_hd__fa_2_4/SUM sky130_fd_sc_hd__fa_2_4/A
+ sky130_fd_sc_hd__fa_2_4/B sky130_fd_sc_hd__fa_2_4/CIN VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_908 sky130_fd_sc_hd__fa_2_894/A sky130_fd_sc_hd__fa_2_895/B
+ sky130_fd_sc_hd__fa_2_908/A sky130_fd_sc_hd__fa_2_908/B sky130_fd_sc_hd__fa_2_908/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_919 sky130_fd_sc_hd__fa_2_918/CIN sky130_fd_sc_hd__fa_2_919/SUM
+ sky130_fd_sc_hd__fa_2_919/A sky130_fd_sc_hd__fa_2_919/B sky130_fd_sc_hd__fa_2_919/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a211o_1_10 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_105/A sky130_fd_sc_hd__a211o_1_9/A2
+ sky130_fd_sc_hd__nor2_1_123/Y sky130_fd_sc_hd__nand2_1_331/B sky130_fd_sc_hd__o22ai_1_166/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__a211o_1_21 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_227/A sky130_fd_sc_hd__nor2b_1_112/Y
+ sky130_fd_sc_hd__o22ai_1_297/Y sky130_fd_sc_hd__o21ai_1_348/Y sky130_fd_sc_hd__o22ai_1_296/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__mux2_2_208 VSS VDD sky130_fd_sc_hd__mux2_2_208/A1 sky130_fd_sc_hd__mux2_2_208/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_208/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_219 VSS VDD sky130_fd_sc_hd__mux2_2_219/A1 sky130_fd_sc_hd__mux2_2_219/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_219/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__clkinv_1_130 sky130_fd_sc_hd__clkinv_2_8/A sky130_fd_sc_hd__clkinv_1_130/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_130/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_141 sky130_fd_sc_hd__buf_12_267/A sky130_fd_sc_hd__clkinv_1_141/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_141/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_152 sky130_fd_sc_hd__clkinv_1_153/A sky130_fd_sc_hd__and2_1_7/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_152/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_163 sky130_fd_sc_hd__inv_2_94/A sky130_fd_sc_hd__inv_2_77/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_163/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_174 sky130_fd_sc_hd__inv_2_103/A sky130_fd_sc_hd__clkinv_1_174/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_174/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_6 sky130_fd_sc_hd__buf_8_6/A sky130_fd_sc_hd__buf_8_6/X VSS
+ VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__a22o_1_8 sky130_fd_sc_hd__a22o_1_8/A1 sky130_fd_sc_hd__nor2_1_1/Y
+ sky130_fd_sc_hd__a22o_1_8/X sky130_fd_sc_hd__a22o_1_8/B2 sky130_fd_sc_hd__nor2_1_0/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_10 sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__ha_2_61/A
+ sky130_fd_sc_hd__a22o_1_10/X sky130_fd_sc_hd__dfxtp_1_10/Q sky130_fd_sc_hd__a22o_2_3/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_185 sky130_fd_sc_hd__nor2b_1_38/B_N sky130_fd_sc_hd__ha_2_89/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_185/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_196 sky130_fd_sc_hd__clkinv_2_20/A sky130_fd_sc_hd__a22o_2_7/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_196/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_21 sky130_fd_sc_hd__nor2_4_4/Y sky130_fd_sc_hd__ha_2_79/A
+ sky130_fd_sc_hd__inv_2_116/A sky130_fd_sc_hd__a22o_1_21/B2 sky130_fd_sc_hd__a22o_2_6/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_32 sky130_fd_sc_hd__or2_1_1/B sky130_fd_sc_hd__ha_2_89/B
+ sky130_fd_sc_hd__a22o_1_32/X sky130_fd_sc_hd__a22o_1_32/B2 sky130_fd_sc_hd__a22o_4_0/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_43 sky130_fd_sc_hd__a22o_1_43/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_43/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__fa_2_949/SUM
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_54 sky130_fd_sc_hd__a22o_1_54/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_54/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__nor4_1_10/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_65 sky130_fd_sc_hd__a22o_1_65/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_65/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__nor4_1_12/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__nand4_1_4 sky130_fd_sc_hd__nand4_1_4/C sky130_fd_sc_hd__nand4_1_4/B
+ sky130_fd_sc_hd__nand4_1_4/Y sky130_fd_sc_hd__nand4_1_4/D sky130_fd_sc_hd__nand4_1_4/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__clkinv_2_0 sky130_fd_sc_hd__inv_2_4/A sky130_fd_sc_hd__ha_2_19/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_0/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__nor2_1_290 sky130_fd_sc_hd__nor2_1_290/B sky130_fd_sc_hd__nor2_1_290/Y
+ sky130_fd_sc_hd__nor2_1_290/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__maj3_1_16 sky130_fd_sc_hd__maj3_1_17/X sky130_fd_sc_hd__maj3_1_16/X
+ sky130_fd_sc_hd__maj3_1_16/B sky130_fd_sc_hd__maj3_1_16/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_27 sky130_fd_sc_hd__maj3_1_28/X sky130_fd_sc_hd__maj3_1_27/X
+ sky130_fd_sc_hd__o22ai_1_2/Y sky130_fd_sc_hd__maj3_1_27/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_406 sky130_fd_sc_hd__nand2_1_516/Y sky130_fd_sc_hd__nand2_1_515/Y
+ sky130_fd_sc_hd__o22ai_1_406/Y sky130_fd_sc_hd__o22ai_1_406/A1 sky130_fd_sc_hd__o21ai_1_445/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_38 sky130_fd_sc_hd__maj3_1_39/X sky130_fd_sc_hd__maj3_1_38/X
+ sky130_fd_sc_hd__maj3_1_38/B sky130_fd_sc_hd__maj3_1_38/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_417 sky130_fd_sc_hd__o22ai_1_436/A2 sky130_fd_sc_hd__o22ai_1_418/A1
+ sky130_fd_sc_hd__o22ai_1_417/Y sky130_fd_sc_hd__nor2_1_273/B sky130_fd_sc_hd__o32ai_1_11/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_49 sky130_fd_sc_hd__maj3_1_50/X sky130_fd_sc_hd__maj3_1_49/X
+ sky130_fd_sc_hd__maj3_1_49/B sky130_fd_sc_hd__maj3_1_49/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_428 sky130_fd_sc_hd__o22ai_1_436/A2 sky130_fd_sc_hd__o22ai_1_436/B1
+ sky130_fd_sc_hd__o22ai_1_428/Y sky130_fd_sc_hd__o21a_1_68/A2 sky130_fd_sc_hd__o22ai_1_432/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_11 sky130_fd_sc_hd__nand3_1_11/C sky130_fd_sc_hd__nand4_1_68/Y
+ sky130_fd_sc_hd__nand2_1_9/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_22 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor3_2_2/B
+ sky130_fd_sc_hd__nor3_2_3/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_33 sky130_fd_sc_hd__nand2_1_33/Y sky130_fd_sc_hd__nor2b_1_50/Y
+ sky130_fd_sc_hd__nand2_1_33/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_44 sky130_fd_sc_hd__nand2_1_44/Y sky130_fd_sc_hd__nand2_1_44/B
+ sky130_fd_sc_hd__a21oi_2_0/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_55 sky130_fd_sc_hd__nand2_1_55/Y sky130_fd_sc_hd__nand2_1_2/B
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_66 sky130_fd_sc_hd__nand2_1_66/Y sky130_fd_sc_hd__nand2_1_67/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_77 sky130_fd_sc_hd__nand2_1_77/Y sky130_fd_sc_hd__nand4_1_66/Y
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_88 sky130_fd_sc_hd__nand2_1_88/Y sky130_fd_sc_hd__nand2_1_89/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_99 sky130_fd_sc_hd__nand2_1_99/Y sky130_fd_sc_hd__buf_2_267/X
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__fa_2_18 sky130_fd_sc_hd__fa_2_8/A sky130_fd_sc_hd__fa_2_16/A sky130_fd_sc_hd__fa_2_86/A
+ sky130_fd_sc_hd__fa_2_18/B sky130_fd_sc_hd__fa_2_18/CIN VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_29 sky130_fd_sc_hd__fa_2_27/CIN sky130_fd_sc_hd__or3_1_5/C
+ sky130_fd_sc_hd__fa_2_29/A sky130_fd_sc_hd__fa_2_29/B sky130_fd_sc_hd__fa_2_29/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_sram_2kbyte_1rw1r_32x512_8_14 sky130_fd_sc_hd__clkbuf_4_160/X sky130_fd_sc_hd__clkbuf_4_161/X
+ sky130_fd_sc_hd__buf_4_120/X sky130_fd_sc_hd__clkbuf_4_162/X sky130_fd_sc_hd__buf_4_98/X
+ sky130_fd_sc_hd__clkbuf_4_210/A sky130_fd_sc_hd__clkbuf_4_163/X sky130_fd_sc_hd__clkbuf_4_164/X
+ sky130_fd_sc_hd__buf_4_99/X sky130_fd_sc_hd__buf_4_100/X sky130_fd_sc_hd__buf_6_54/X
+ sky130_fd_sc_hd__buf_4_101/X sky130_fd_sc_hd__buf_4_102/X sky130_fd_sc_hd__buf_4_103/X
+ sky130_fd_sc_hd__buf_4_104/X sky130_fd_sc_hd__buf_4_105/X sky130_fd_sc_hd__clkbuf_4_160/X
+ sky130_fd_sc_hd__clkbuf_4_161/X sky130_fd_sc_hd__buf_4_120/A sky130_fd_sc_hd__clkbuf_4_162/X
+ sky130_fd_sc_hd__buf_4_98/X sky130_fd_sc_hd__clkbuf_4_210/A sky130_fd_sc_hd__clkbuf_4_163/X
+ sky130_fd_sc_hd__clkbuf_4_164/X sky130_fd_sc_hd__buf_4_99/X sky130_fd_sc_hd__buf_4_100/X
+ sky130_fd_sc_hd__buf_6_54/X sky130_fd_sc_hd__buf_4_101/X sky130_fd_sc_hd__buf_4_102/X
+ sky130_fd_sc_hd__buf_4_103/X sky130_fd_sc_hd__buf_4_104/X sky130_fd_sc_hd__buf_4_105/X
+ sky130_fd_sc_hd__buf_12_469/X sky130_fd_sc_hd__buf_12_507/X sky130_fd_sc_hd__buf_12_478/X
+ sky130_fd_sc_hd__buf_12_505/X sky130_fd_sc_hd__buf_12_461/X sky130_fd_sc_hd__buf_12_404/X
+ sky130_fd_sc_hd__buf_12_479/X sky130_fd_sc_hd__buf_12_474/X sky130_fd_sc_hd__buf_12_455/X
+ sky130_fd_sc_hd__buf_12_503/X sky130_fd_sc_hd__buf_12_496/X sky130_fd_sc_hd__buf_12_500/X
+ sky130_fd_sc_hd__buf_12_425/X sky130_fd_sc_hd__buf_12_482/X sky130_fd_sc_hd__buf_12_396/X
+ sky130_fd_sc_hd__buf_12_424/X sky130_fd_sc_hd__buf_12_446/X sky130_fd_sc_hd__buf_12_506/X
+ sky130_fd_sc_hd__clkbuf_1_484/X sky130_fd_sc_hd__clkbuf_1_374/X sky130_fd_sc_hd__clkbuf_1_485/X
+ sky130_fd_sc_hd__clkinv_8_36/Y sky130_fd_sc_hd__clkinv_8_19/Y sky130_fd_sc_hd__buf_12_470/X
+ sky130_fd_sc_hd__buf_12_447/X sky130_fd_sc_hd__bufbuf_8_9/A sky130_fd_sc_hd__buf_12_519/X
+ sky130_fd_sc_hd__buf_2_249/A sky130_fd_sc_hd__buf_2_169/A sky130_fd_sc_hd__buf_2_170/A
+ sky130_fd_sc_hd__buf_2_171/A sky130_fd_sc_hd__clkbuf_1_531/A sky130_fd_sc_hd__buf_2_173/A
+ sky130_fd_sc_hd__buf_2_174/A sky130_fd_sc_hd__buf_2_175/A sky130_fd_sc_hd__buf_2_176/A
+ sky130_fd_sc_hd__buf_2_177/A sky130_fd_sc_hd__buf_2_178/A sky130_fd_sc_hd__buf_2_179/A
+ sky130_fd_sc_hd__buf_2_180/A sky130_fd_sc_hd__clkbuf_1_528/A sky130_fd_sc_hd__buf_2_182/A
+ sky130_fd_sc_hd__buf_2_183/A sky130_fd_sc_hd__clkbuf_1_414/A sky130_fd_sc_hd__buf_2_184/A
+ sky130_fd_sc_hd__clkbuf_1_415/A sky130_fd_sc_hd__clkbuf_1_416/A sky130_fd_sc_hd__clkbuf_1_417/A
+ sky130_fd_sc_hd__buf_2_251/A sky130_fd_sc_hd__clkbuf_1_419/A sky130_fd_sc_hd__clkbuf_1_420/A
+ sky130_fd_sc_hd__clkbuf_1_421/A sky130_fd_sc_hd__clkbuf_1_527/A sky130_fd_sc_hd__buf_2_185/A
+ sky130_fd_sc_hd__buf_2_186/A sky130_fd_sc_hd__clkbuf_1_423/A sky130_fd_sc_hd__clkbuf_1_536/A
+ sky130_fd_sc_hd__clkbuf_1_425/A sky130_fd_sc_hd__clkbuf_1_426/A sky130_fd_sc_hd__buf_2_187/A
+ sky130_fd_sc_hd__buf_2_188/A sky130_fd_sc_hd__buf_2_189/A sky130_fd_sc_hd__buf_2_190/A
+ sky130_fd_sc_hd__buf_2_191/A sky130_fd_sc_hd__buf_2_192/A sky130_fd_sc_hd__buf_2_193/A
+ sky130_fd_sc_hd__buf_2_194/A sky130_fd_sc_hd__buf_2_195/A sky130_fd_sc_hd__buf_2_196/A
+ sky130_fd_sc_hd__buf_2_197/A sky130_fd_sc_hd__buf_2_198/A sky130_fd_sc_hd__buf_2_199/A
+ sky130_fd_sc_hd__buf_2_200/A sky130_fd_sc_hd__buf_2_201/A sky130_fd_sc_hd__buf_2_202/A
+ sky130_fd_sc_hd__buf_2_203/A sky130_fd_sc_hd__buf_2_204/A sky130_fd_sc_hd__clkbuf_1_427/A
+ sky130_fd_sc_hd__buf_2_205/A sky130_fd_sc_hd__buf_2_206/A sky130_fd_sc_hd__buf_2_207/A
+ sky130_fd_sc_hd__buf_2_208/A sky130_fd_sc_hd__buf_2_209/A sky130_fd_sc_hd__buf_2_210/A
+ sky130_fd_sc_hd__clkbuf_1_530/A sky130_fd_sc_hd__buf_2_212/A sky130_fd_sc_hd__buf_2_213/A
+ sky130_fd_sc_hd__buf_2_214/A sky130_fd_sc_hd__buf_2_247/A sky130_fd_sc_hd__buf_2_216/A
+ sky130_fd_sc_hd__buf_2_217/A VDD VSS sky130_sram_2kbyte_1rw1r_32x512_8
Xsky130_fd_sc_hd__dfxtp_1_1206 VDD VSS sky130_fd_sc_hd__fa_2_1255/A sky130_fd_sc_hd__clkinv_8_116/Y
+ sky130_fd_sc_hd__mux2_2_182/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1217 VDD VSS sky130_fd_sc_hd__fa_2_1229/A sky130_fd_sc_hd__clkinv_8_78/Y
+ sky130_fd_sc_hd__mux2_2_204/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1228 VDD VSS sky130_fd_sc_hd__fa_2_1240/A sky130_fd_sc_hd__clkinv_8_116/Y
+ sky130_fd_sc_hd__mux2_2_177/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_800 VDD VSS sky130_fd_sc_hd__fa_2_1052/A sky130_fd_sc_hd__clkinv_8_55/Y
+ sky130_fd_sc_hd__mux2_2_75/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1239 VDD VSS sky130_fd_sc_hd__fa_2_1268/A sky130_fd_sc_hd__clkinv_8_65/Y
+ sky130_fd_sc_hd__mux2_2_205/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_811 VDD VSS sky130_fd_sc_hd__fa_2_1063/A sky130_fd_sc_hd__clkinv_4_26/Y
+ sky130_fd_sc_hd__mux2_2_51/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_822 VDD VSS sky130_fd_sc_hd__fa_2_1096/A sky130_fd_sc_hd__clkinv_8_59/Y
+ sky130_fd_sc_hd__and2_0_298/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_833 VDD VSS sky130_fd_sc_hd__xor2_1_139/A sky130_fd_sc_hd__clkinv_4_26/Y
+ sky130_fd_sc_hd__mux2_2_66/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_844 VDD VSS sky130_fd_sc_hd__mux2_2_65/A1 sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__o21ai_1_161/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_855 VDD VSS sky130_fd_sc_hd__mux2_2_43/A1 sky130_fd_sc_hd__clkinv_4_25/Y
+ sky130_fd_sc_hd__o21ai_1_172/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_866 VDD VSS sky130_fd_sc_hd__mux2_2_60/A1 sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__o21ai_1_180/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_877 VDD VSS sky130_fd_sc_hd__mux2_2_38/A1 sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__o21ai_1_191/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_888 VDD VSS sky130_fd_sc_hd__fa_2_854/A sky130_fd_sc_hd__dfxtp_1_904/CLK
+ sky130_fd_sc_hd__o21a_1_25/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_899 VDD VSS sky130_fd_sc_hd__fa_2_934/B sky130_fd_sc_hd__dfxtp_1_899/CLK
+ sky130_fd_sc_hd__dfxtp_1_899/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_420 VSS VDD sky130_fd_sc_hd__clkbuf_1_420/X sky130_fd_sc_hd__clkbuf_1_420/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_431 VSS VDD sky130_fd_sc_hd__clkbuf_1_431/X sky130_fd_sc_hd__clkbuf_1_431/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_442 VSS VDD sky130_fd_sc_hd__a22oi_2_28/A2 sky130_fd_sc_hd__clkbuf_1_442/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_453 VSS VDD sky130_fd_sc_hd__clkbuf_1_453/X sky130_fd_sc_hd__clkbuf_1_453/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_464 VSS VDD sky130_fd_sc_hd__clkbuf_1_464/X sky130_fd_sc_hd__clkbuf_1_464/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_475 VSS VDD sky130_fd_sc_hd__nand4_1_61/D sky130_fd_sc_hd__a22oi_1_247/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_486 VSS VDD sky130_fd_sc_hd__buf_8_196/A sky130_fd_sc_hd__inv_2_112/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_497 VSS VDD sky130_fd_sc_hd__clkbuf_1_497/X sky130_fd_sc_hd__clkbuf_1_497/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_705 sky130_fd_sc_hd__fa_2_704/CIN sky130_fd_sc_hd__fa_2_705/SUM
+ sky130_fd_sc_hd__fa_2_705/A sky130_fd_sc_hd__fa_2_705/B sky130_fd_sc_hd__fa_2_705/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_716 sky130_fd_sc_hd__fa_2_715/CIN sky130_fd_sc_hd__fa_2_716/SUM
+ sky130_fd_sc_hd__fa_2_716/A sky130_fd_sc_hd__fa_2_716/B sky130_fd_sc_hd__maj3_1_135/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_727 sky130_fd_sc_hd__fa_2_729/B sky130_fd_sc_hd__fa_2_727/SUM
+ sky130_fd_sc_hd__ha_2_142/A sky130_fd_sc_hd__fa_2_758/B sky130_fd_sc_hd__fa_2_736/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_738 sky130_fd_sc_hd__maj3_1_149/B sky130_fd_sc_hd__maj3_1_150/A
+ sky130_fd_sc_hd__fa_2_738/A sky130_fd_sc_hd__fa_2_738/B sky130_fd_sc_hd__fa_2_739/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_749 sky130_fd_sc_hd__fa_2_752/B sky130_fd_sc_hd__fa_2_749/SUM
+ sky130_fd_sc_hd__fa_2_749/A sky130_fd_sc_hd__fa_2_749/B sky130_fd_sc_hd__o22ai_1_50/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor2b_1_102 sky130_fd_sc_hd__o22ai_1_164/Y sky130_fd_sc_hd__nor2b_1_102/Y
+ sky130_fd_sc_hd__buf_2_262/X VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_113 sky130_fd_sc_hd__or2_0_10/X sky130_fd_sc_hd__nor2b_1_113/Y
+ sky130_fd_sc_hd__buf_2_262/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_124 sky130_fd_sc_hd__and2_0_333/X sky130_fd_sc_hd__nor2b_1_124/Y
+ sky130_fd_sc_hd__buf_2_262/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_135 sky130_fd_sc_hd__nand2b_1_17/Y sky130_fd_sc_hd__nor2b_1_135/Y
+ sky130_fd_sc_hd__nor4_1_13/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__buf_6_3 VDD VSS sky130_fd_sc_hd__buf_6_3/X sky130_fd_sc_hd__buf_6_3/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__bufbuf_8_6 sky130_fd_sc_hd__a22o_1_25/X sky130_fd_sc_hd__buf_6_70/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufbuf_8
Xsky130_fd_sc_hd__buf_6_19 VDD VSS sky130_fd_sc_hd__buf_6_19/X sky130_fd_sc_hd__buf_6_19/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__o22ai_1_203 sky130_fd_sc_hd__nor2_1_126/A sky130_fd_sc_hd__nor2_2_13/B
+ sky130_fd_sc_hd__o22ai_1_203/Y sky130_fd_sc_hd__a21oi_1_238/Y sky130_fd_sc_hd__a211oi_1_9/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__sdlclkp_4_1 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__clkinv_8_118/Y
+ sky130_fd_sc_hd__dfxtp_1_60/CLK sky130_fd_sc_hd__clkbuf_1_0/X VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__o22ai_1_214 sky130_fd_sc_hd__nand2_1_358/Y sky130_fd_sc_hd__nand2_1_357/Y
+ sky130_fd_sc_hd__o22ai_1_214/Y sky130_fd_sc_hd__nand2_1_369/B sky130_fd_sc_hd__o21ai_1_279/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_225 sky130_fd_sc_hd__nand2_1_360/Y sky130_fd_sc_hd__nand2_1_359/Y
+ sky130_fd_sc_hd__o22ai_1_225/Y sky130_fd_sc_hd__nand2_1_368/B sky130_fd_sc_hd__o21ai_1_278/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_236 sky130_fd_sc_hd__nor2_1_183/A sky130_fd_sc_hd__nor2_1_180/A
+ sky130_fd_sc_hd__o22ai_1_236/Y sky130_fd_sc_hd__a21boi_1_2/Y sky130_fd_sc_hd__nor2_1_164/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_247 sky130_fd_sc_hd__o22ai_1_265/A2 sky130_fd_sc_hd__nor2_1_143/B
+ sky130_fd_sc_hd__o22ai_1_247/Y sky130_fd_sc_hd__o22ai_1_247/A1 sky130_fd_sc_hd__o32ai_1_2/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_258 sky130_fd_sc_hd__o22ai_1_265/A2 sky130_fd_sc_hd__o22ai_1_258/B1
+ sky130_fd_sc_hd__o22ai_1_258/Y sky130_fd_sc_hd__nor2_1_154/B sky130_fd_sc_hd__o32ai_1_2/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_1_4 sky130_fd_sc_hd__nor2_4_6/B sky130_fd_sc_hd__nor2_1_4/Y
+ sky130_fd_sc_hd__nor3_2_4/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__o22ai_1_269 sky130_fd_sc_hd__nand2_1_410/Y sky130_fd_sc_hd__nand2_1_409/Y
+ sky130_fd_sc_hd__o22ai_1_269/Y sky130_fd_sc_hd__nand2_1_420/B sky130_fd_sc_hd__o21ai_1_332/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__bufinv_8_6 sky130_fd_sc_hd__bufinv_8_6/A sky130_fd_sc_hd__bufinv_8_6/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufinv_8
Xsky130_fd_sc_hd__dfxtp_1_107 VDD VSS sky130_fd_sc_hd__xor2_1_9/A sky130_fd_sc_hd__dfxtp_1_111/CLK
+ sky130_fd_sc_hd__ha_2_9/SUM VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_118 VDD VSS sky130_fd_sc_hd__o21ai_1_1/A2 sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__and2_0_0/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_129 VDD VSS sky130_fd_sc_hd__ha_2_11/A sky130_fd_sc_hd__dfxtp_1_129/CLK
+ sky130_fd_sc_hd__and2_0_23/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_430 VSS VDD sky130_fd_sc_hd__o22ai_1_375/A2 sky130_fd_sc_hd__nor2_1_266/A
+ sky130_fd_sc_hd__a21oi_1_412/Y sky130_fd_sc_hd__o21ai_1_430/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_441 VSS VDD sky130_fd_sc_hd__nand2_1_525/B sky130_fd_sc_hd__nor2_1_295/Y
+ sky130_fd_sc_hd__nor2_1_294/B sky130_fd_sc_hd__o21ai_1_441/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_452 VSS VDD sky130_fd_sc_hd__nor2_1_299/B sky130_fd_sc_hd__nor2_1_309/A
+ sky130_fd_sc_hd__nand2_1_529/Y sky130_fd_sc_hd__xor2_1_302/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_463 VSS VDD sky130_fd_sc_hd__nor2_1_270/B sky130_fd_sc_hd__o21a_1_68/A1
+ sky130_fd_sc_hd__a21oi_1_454/Y sky130_fd_sc_hd__o21ai_1_463/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_474 VSS VDD sky130_fd_sc_hd__a211oi_1_37/Y sky130_fd_sc_hd__nor2_1_309/A
+ sky130_fd_sc_hd__nand2_1_538/Y sky130_fd_sc_hd__xor2_1_282/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_485 VSS VDD sky130_fd_sc_hd__nor2_1_278/B sky130_fd_sc_hd__o21a_1_68/A1
+ sky130_fd_sc_hd__a21oi_1_473/Y sky130_fd_sc_hd__o21ai_1_485/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_496 VSS VDD sky130_fd_sc_hd__nand2_1_557/A sky130_fd_sc_hd__o21ai_1_507/A1
+ sky130_fd_sc_hd__nand2_1_557/Y sky130_fd_sc_hd__and2_0_341/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_1206 sky130_fd_sc_hd__fa_2_1207/CIN sky130_fd_sc_hd__mux2_2_130/A0
+ sky130_fd_sc_hd__fa_2_1206/A sky130_fd_sc_hd__fa_2_1206/B sky130_fd_sc_hd__fa_2_1206/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1217 sky130_fd_sc_hd__fa_2_1218/CIN sky130_fd_sc_hd__mux2_2_157/A1
+ sky130_fd_sc_hd__fa_2_1217/A sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__fa_2_1217/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1228 sky130_fd_sc_hd__fa_2_1229/CIN sky130_fd_sc_hd__mux2_2_207/A1
+ sky130_fd_sc_hd__fa_2_1228/A sky130_fd_sc_hd__fa_2_1228/B sky130_fd_sc_hd__fa_2_1228/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1239 sky130_fd_sc_hd__fa_2_1240/CIN sky130_fd_sc_hd__mux2_2_179/A0
+ sky130_fd_sc_hd__fa_2_1239/A sky130_fd_sc_hd__fa_2_1239/B sky130_fd_sc_hd__fa_2_1239/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1003 VDD VSS sky130_fd_sc_hd__mux2_2_113/A0 sky130_fd_sc_hd__clkinv_8_55/Y
+ sky130_fd_sc_hd__a21oi_1_259/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_12 VSS VDD sky130_fd_sc_hd__o21ai_1_13/Y sky130_fd_sc_hd__or4_1_1/B
+ sky130_fd_sc_hd__a21oi_1_9/Y sky130_fd_sc_hd__nor4_1_1/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1014 VDD VSS sky130_fd_sc_hd__mux2_2_84/A1 sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__o22ai_1_225/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_23 VSS VDD sky130_fd_sc_hd__a21oi_2_0/Y sky130_fd_sc_hd__nor2_1_12/B
+ sky130_fd_sc_hd__nand2_1_42/Y sky130_fd_sc_hd__o21ai_1_23/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1025 VDD VSS sky130_fd_sc_hd__fa_2_844/A sky130_fd_sc_hd__dfxtp_1_1038/CLK
+ sky130_fd_sc_hd__o21a_1_40/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_34 VSS VDD sky130_fd_sc_hd__nor2b_1_84/Y sky130_fd_sc_hd__nor3_1_35/Y
+ sky130_fd_sc_hd__nand4_1_84/C sky130_fd_sc_hd__o21ai_1_34/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1036 VDD VSS sky130_fd_sc_hd__fa_2_901/A sky130_fd_sc_hd__dfxtp_1_1038/CLK
+ sky130_fd_sc_hd__a21oi_1_308/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_45 VSS VDD sky130_fd_sc_hd__o21ai_1_53/A2 sky130_fd_sc_hd__xnor2_1_44/Y
+ sky130_fd_sc_hd__a21oi_1_33/Y sky130_fd_sc_hd__o21ai_1_45/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1047 VDD VSS sky130_fd_sc_hd__fa_2_913/B sky130_fd_sc_hd__dfxtp_1_1047/CLK
+ sky130_fd_sc_hd__o21a_1_31/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_56 VSS VDD sky130_fd_sc_hd__nand2_2_3/Y sky130_fd_sc_hd__o21ai_1_73/A2
+ sky130_fd_sc_hd__o21ai_1_56/B1 sky130_fd_sc_hd__o21ai_1_56/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1058 VDD VSS sky130_fd_sc_hd__fa_2_1197/A sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__mux2_2_152/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_67 VSS VDD sky130_fd_sc_hd__nand2_2_3/Y sky130_fd_sc_hd__xnor2_1_54/Y
+ sky130_fd_sc_hd__a21oi_1_53/Y sky130_fd_sc_hd__o21ai_1_67/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_290 sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1281/B
+ sky130_fd_sc_hd__xor2_1_290/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_630 VDD VSS sky130_fd_sc_hd__fa_2_994/A sky130_fd_sc_hd__clkinv_8_41/Y
+ sky130_fd_sc_hd__and2_0_279/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1069 VDD VSS sky130_fd_sc_hd__fa_2_1208/A sky130_fd_sc_hd__clkinv_8_70/Y
+ sky130_fd_sc_hd__mux2_2_126/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_641 VDD VSS sky130_fd_sc_hd__fa_2_1005/A sky130_fd_sc_hd__clkinv_8_44/Y
+ sky130_fd_sc_hd__mux2_2_22/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_78 VSS VDD sky130_fd_sc_hd__xnor2_1_44/A sky130_fd_sc_hd__o21ai_1_78/A1
+ sky130_fd_sc_hd__o21ai_1_78/B1 sky130_fd_sc_hd__xnor2_1_46/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_652 VDD VSS sky130_fd_sc_hd__nor2_4_9/B sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__mux2_2_0/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_89 VSS VDD sky130_fd_sc_hd__nor2_1_77/A sky130_fd_sc_hd__o22ai_1_90/A2
+ sky130_fd_sc_hd__o21ai_1_89/B1 sky130_fd_sc_hd__o21ai_1_89/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_663 VDD VSS sky130_fd_sc_hd__fa_2_980/A sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__mux2_2_27/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_674 VDD VSS sky130_fd_sc_hd__fa_2_991/A sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__mux2_2_5/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_685 VDD VSS sky130_fd_sc_hd__fa_2_1024/A sky130_fd_sc_hd__clkinv_8_59/Y
+ sky130_fd_sc_hd__and2_0_281/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_696 VDD VSS sky130_fd_sc_hd__nor2_1_89/A sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__o21bai_1_0/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_250 VSS VDD sky130_fd_sc_hd__clkbuf_1_250/X sky130_fd_sc_hd__clkbuf_1_251/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_261 VSS VDD sky130_fd_sc_hd__nand2_2_0/B sky130_fd_sc_hd__nor2b_1_1/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_272 VSS VDD sky130_fd_sc_hd__clkbuf_1_272/X sky130_fd_sc_hd__clkbuf_1_272/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_283 VSS VDD sky130_fd_sc_hd__clkbuf_1_283/X sky130_fd_sc_hd__clkbuf_1_283/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_294 VSS VDD sky130_fd_sc_hd__clkbuf_1_294/X sky130_fd_sc_hd__clkbuf_1_294/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_502 sky130_fd_sc_hd__fa_2_503/B sky130_fd_sc_hd__fa_2_495/A
+ sky130_fd_sc_hd__ha_2_124/A sky130_fd_sc_hd__fa_2_502/B sky130_fd_sc_hd__fa_2_554/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_513 sky130_fd_sc_hd__maj3_1_91/B sky130_fd_sc_hd__maj3_1_92/A
+ sky130_fd_sc_hd__fa_2_513/A sky130_fd_sc_hd__fa_2_513/B sky130_fd_sc_hd__fa_2_514/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_524 sky130_fd_sc_hd__maj3_1_89/B sky130_fd_sc_hd__maj3_1_90/A
+ sky130_fd_sc_hd__fa_2_524/A sky130_fd_sc_hd__fa_2_524/B sky130_fd_sc_hd__fa_2_525/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_535 sky130_fd_sc_hd__fa_2_532/B sky130_fd_sc_hd__fa_2_528/B
+ sky130_fd_sc_hd__fa_2_535/A sky130_fd_sc_hd__ha_2_124/B sky130_fd_sc_hd__fa_2_567/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_546 sky130_fd_sc_hd__fa_2_545/A sky130_fd_sc_hd__fa_2_539/B
+ sky130_fd_sc_hd__fa_2_546/A sky130_fd_sc_hd__fa_2_546/B sky130_fd_sc_hd__fa_2_558/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_557 sky130_fd_sc_hd__fa_2_560/B sky130_fd_sc_hd__fa_2_557/SUM
+ sky130_fd_sc_hd__fa_2_557/A sky130_fd_sc_hd__fa_2_557/B sky130_fd_sc_hd__fa_2_557/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_568 sky130_fd_sc_hd__xnor2_1_4/B sky130_fd_sc_hd__and2_0_86/A
+ sky130_fd_sc_hd__fa_2_698/A sky130_fd_sc_hd__fa_2_568/B sky130_fd_sc_hd__fa_2_568/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_579 sky130_fd_sc_hd__fa_2_578/CIN sky130_fd_sc_hd__and2_0_97/A
+ sky130_fd_sc_hd__fa_2_579/A sky130_fd_sc_hd__fa_2_579/B sky130_fd_sc_hd__fa_2_579/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_4_0 VDD VSS sky130_fd_sc_hd__buf_4_0/X sky130_fd_sc_hd__buf_4_0/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__and2_0_270 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_270/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__and2_0_270/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_281 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_281/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__and2_0_281/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_292 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_292/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__and2_0_292/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_507 sky130_fd_sc_hd__buf_12_507/A sky130_fd_sc_hd__buf_12_507/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_518 sky130_fd_sc_hd__buf_12_518/A sky130_fd_sc_hd__buf_12_518/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__inv_4_0 sky130_fd_sc_hd__inv_4_0/Y sky130_fd_sc_hd__inv_4_0/A VDD
+ VSS VDD VSS sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__nand2_1_108 sky130_fd_sc_hd__nand2_1_108/Y sky130_fd_sc_hd__nand2_1_109/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_707 sky130_fd_sc_hd__nor2_1_114/B sky130_fd_sc_hd__fa_2_1063/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_707/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_119 sky130_fd_sc_hd__nand2_1_119/Y sky130_fd_sc_hd__nand2_1_120/Y
+ sky130_fd_sc_hd__buf_2_264/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_718 sky130_fd_sc_hd__nand4_1_86/D sky130_fd_sc_hd__fa_2_1046/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_718/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_729 sky130_fd_sc_hd__clkinv_1_729/Y sky130_fd_sc_hd__a211oi_1_10/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_729/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_260 VSS VDD sky130_fd_sc_hd__a21oi_1_231/Y sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__a21oi_1_225/Y sky130_fd_sc_hd__xor2_1_104/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_271 VSS VDD sky130_fd_sc_hd__o21ai_1_271/A2 sky130_fd_sc_hd__o22ai_1_206/A1
+ sky130_fd_sc_hd__a22oi_1_367/Y sky130_fd_sc_hd__o21ai_1_271/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_282 VSS VDD sky130_fd_sc_hd__nand2_1_372/B sky130_fd_sc_hd__nor2_1_171/Y
+ sky130_fd_sc_hd__nor2_1_170/B sky130_fd_sc_hd__o21ai_1_282/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_293 VSS VDD sky130_fd_sc_hd__a222oi_1_6/Y sky130_fd_sc_hd__nor2_1_180/A
+ sky130_fd_sc_hd__a21oi_1_264/Y sky130_fd_sc_hd__xor2_1_170/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor3_1_18 sky130_fd_sc_hd__nor3_2_10/B sky130_fd_sc_hd__nor3_1_18/Y
+ sky130_fd_sc_hd__nor2_2_5/A sky130_fd_sc_hd__nor3_2_10/A VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_29 sky130_fd_sc_hd__xor2_1_9/A sky130_fd_sc_hd__xor2_1_22/B
+ sky130_fd_sc_hd__nor4_1_4/B sky130_fd_sc_hd__nor4_1_4/C VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor2b_2_0 sky130_fd_sc_hd__ha_2_44/SUM sky130_fd_sc_hd__or2_1_0/B
+ sky130_fd_sc_hd__nor2b_2_0/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_2
Xsky130_fd_sc_hd__fa_2_1003 sky130_fd_sc_hd__fa_2_1004/CIN sky130_fd_sc_hd__mux2_2_26/A0
+ sky130_fd_sc_hd__fa_2_1003/A sky130_fd_sc_hd__xor2_1_73/X sky130_fd_sc_hd__fa_2_1003/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1014 sky130_fd_sc_hd__fa_2_1015/CIN sky130_fd_sc_hd__mux2_2_4/A0
+ sky130_fd_sc_hd__fa_2_1014/A sky130_fd_sc_hd__xor2_1_62/X sky130_fd_sc_hd__fa_2_1014/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1025 sky130_fd_sc_hd__fa_2_1026/CIN sky130_fd_sc_hd__and2_0_285/A
+ sky130_fd_sc_hd__fa_2_1025/A sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_1025/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1036 sky130_fd_sc_hd__fa_2_1037/CIN sky130_fd_sc_hd__fa_2_1036/SUM
+ sky130_fd_sc_hd__nor2_1_58/A sky130_fd_sc_hd__fa_2_1036/B sky130_fd_sc_hd__fa_2_1036/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1047 sky130_fd_sc_hd__fa_2_1048/CIN sky130_fd_sc_hd__and2_0_303/A
+ sky130_fd_sc_hd__fa_2_1047/A sky130_fd_sc_hd__fa_2_1047/B sky130_fd_sc_hd__fa_2_1047/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1058 sky130_fd_sc_hd__fa_2_1059/CIN sky130_fd_sc_hd__mux2_2_61/A0
+ sky130_fd_sc_hd__fa_2_1058/A sky130_fd_sc_hd__xor2_1_99/X sky130_fd_sc_hd__fa_2_1058/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1069 sky130_fd_sc_hd__fa_2_1070/CIN sky130_fd_sc_hd__and2_0_302/A
+ sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1069/B sky130_fd_sc_hd__xor2_1_137/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_12 sky130_fd_sc_hd__inv_2_12/A sky130_fd_sc_hd__inv_2_12/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_23 sky130_fd_sc_hd__inv_2_23/A sky130_fd_sc_hd__inv_2_23/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_34 sky130_fd_sc_hd__inv_2_34/A sky130_fd_sc_hd__inv_2_34/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_45 sky130_fd_sc_hd__inv_2_45/A sky130_fd_sc_hd__inv_2_45/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_56 sky130_fd_sc_hd__ha_2_49/A sky130_fd_sc_hd__inv_2_56/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_460 VDD VSS sky130_fd_sc_hd__buf_2_10/A sky130_fd_sc_hd__dfxtp_1_463/CLK
+ sky130_fd_sc_hd__and2_0_238/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_67 sky130_fd_sc_hd__inv_2_67/A sky130_fd_sc_hd__inv_2_67/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_471 VDD VSS sky130_fd_sc_hd__clkbuf_1_3/A sky130_fd_sc_hd__dfxtp_1_473/CLK
+ sky130_fd_sc_hd__and2_0_116/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_78 sky130_fd_sc_hd__inv_2_78/A sky130_fd_sc_hd__inv_2_78/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_482 VDD VSS sky130_fd_sc_hd__nand2_1_223/A sky130_fd_sc_hd__dfxtp_1_483/CLK
+ sky130_fd_sc_hd__nor2b_1_63/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_2_2 sky130_fd_sc_hd__nand2_2_2/Y sky130_fd_sc_hd__nor2_1_16/Y
+ sky130_fd_sc_hd__nor3_1_26/C VDD VSS VSS VDD sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__inv_2_89 sky130_fd_sc_hd__inv_2_89/A sky130_fd_sc_hd__inv_2_89/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_493 VDD VSS sky130_fd_sc_hd__dfxtp_1_493/Q sky130_fd_sc_hd__dfxtp_1_496/CLK
+ sky130_fd_sc_hd__nor2b_1_60/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_310 sky130_fd_sc_hd__fa_2_306/CIN sky130_fd_sc_hd__nor2_1_213/A
+ sky130_fd_sc_hd__fa_2_310/A sky130_fd_sc_hd__fa_2_310/B sky130_fd_sc_hd__fa_2_310/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_321 sky130_fd_sc_hd__fa_2_314/A sky130_fd_sc_hd__fa_2_318/B
+ sky130_fd_sc_hd__fa_2_321/A sky130_fd_sc_hd__fa_2_321/B sky130_fd_sc_hd__fa_2_321/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_332 sky130_fd_sc_hd__fa_2_334/B sky130_fd_sc_hd__fa_2_332/SUM
+ sky130_fd_sc_hd__ha_2_110/B sky130_fd_sc_hd__fa_2_422/B sky130_fd_sc_hd__fa_2_332/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_343 sky130_fd_sc_hd__maj3_1_71/B sky130_fd_sc_hd__maj3_1_72/A
+ sky130_fd_sc_hd__fa_2_343/A sky130_fd_sc_hd__fa_2_343/B sky130_fd_sc_hd__fa_2_344/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_354 sky130_fd_sc_hd__fa_2_355/CIN sky130_fd_sc_hd__fa_2_348/A
+ sky130_fd_sc_hd__ha_2_110/A sky130_fd_sc_hd__fa_2_412/A sky130_fd_sc_hd__fa_2_413/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_365 sky130_fd_sc_hd__fa_2_367/CIN sky130_fd_sc_hd__fa_2_362/A
+ sky130_fd_sc_hd__fa_2_365/A sky130_fd_sc_hd__fa_2_365/B sky130_fd_sc_hd__fa_2_373/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_376 sky130_fd_sc_hd__fa_2_378/CIN sky130_fd_sc_hd__fa_2_371/A
+ sky130_fd_sc_hd__fa_2_376/A sky130_fd_sc_hd__fa_2_376/B sky130_fd_sc_hd__fa_2_376/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_17 sky130_fd_sc_hd__conb_1_11/LO sky130_fd_sc_hd__clkinv_8_131/A
+ sky130_fd_sc_hd__dfxtp_1_170/CLK sky130_fd_sc_hd__or2_1_0/X VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_387 sky130_fd_sc_hd__maj3_1_62/B sky130_fd_sc_hd__maj3_1_63/A
+ sky130_fd_sc_hd__fa_2_387/A sky130_fd_sc_hd__fa_2_387/B sky130_fd_sc_hd__fa_2_388/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_28 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_61/Y
+ sky130_fd_sc_hd__dfxtp_1_258/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__and2_1_3 VDD VSS sky130_fd_sc_hd__and2_1_3/X sky130_fd_sc_hd__ha_2_53/A
+ sky130_fd_sc_hd__nor2_4_2/Y VDD VSS sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__fa_2_398 sky130_fd_sc_hd__fa_2_395/B sky130_fd_sc_hd__fa_2_398/SUM
+ sky130_fd_sc_hd__ha_2_116/A sky130_fd_sc_hd__ha_2_116/B sky130_fd_sc_hd__ha_2_115/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22oi_2_9 sky130_fd_sc_hd__nor2_4_5/Y sky130_fd_sc_hd__a22oi_2_9/A2
+ sky130_fd_sc_hd__a22oi_2_9/B1 sky130_fd_sc_hd__a22oi_2_9/B2 sky130_fd_sc_hd__a22oi_2_9/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__diode_2_204 sky130_fd_sc_hd__inv_2_141/Y VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__sdlclkp_4_39 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_100/Y
+ sky130_fd_sc_hd__dfxtp_1_361/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__diode_2_215 amplitude_adc_done VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_226 sig_amplitude[0] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkinv_8_70 sky130_fd_sc_hd__clkinv_8_70/Y sky130_fd_sc_hd__clkinv_8_70/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_70/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_81 sky130_fd_sc_hd__clkinv_8_82/A sky130_fd_sc_hd__clkinv_8_81/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_81/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_92 sky130_fd_sc_hd__clkinv_8_93/A sky130_fd_sc_hd__clkinv_8_97/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_92/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_90 sky130_fd_sc_hd__buf_12_90/A sky130_fd_sc_hd__buf_12_90/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__nor2_1_108 sky130_fd_sc_hd__nor2_1_108/B sky130_fd_sc_hd__nor2_1_108/Y
+ sky130_fd_sc_hd__fa_2_1112/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_119 sky130_fd_sc_hd__nor2_1_119/B sky130_fd_sc_hd__o21a_1_14/A1
+ sky130_fd_sc_hd__o21a_1_15/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_17 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__a22oi_1_9/A1
+ sky130_fd_sc_hd__nand4_1_39/Y sky130_fd_sc_hd__buf_2_291/X sky130_fd_sc_hd__nand3_1_8/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_28 sky130_fd_sc_hd__clkbuf_4_8/X sky130_fd_sc_hd__clkbuf_4_9/X
+ sky130_fd_sc_hd__clkbuf_1_34/X sky130_fd_sc_hd__a22oi_1_28/A2 sky130_fd_sc_hd__a22oi_1_28/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_39 sky130_fd_sc_hd__clkbuf_4_8/X sky130_fd_sc_hd__clkbuf_4_9/X
+ sky130_fd_sc_hd__clkbuf_1_31/X sky130_fd_sc_hd__a22oi_1_39/A2 sky130_fd_sc_hd__a22oi_1_39/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_304 sky130_fd_sc_hd__buf_8_136/X sky130_fd_sc_hd__buf_8_177/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_315 sky130_fd_sc_hd__buf_4_76/X sky130_fd_sc_hd__buf_12_315/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_326 sky130_fd_sc_hd__buf_4_72/X sky130_fd_sc_hd__buf_12_326/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_337 sky130_fd_sc_hd__buf_4_80/X sky130_fd_sc_hd__buf_12_337/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_348 sky130_fd_sc_hd__buf_6_47/X sky130_fd_sc_hd__buf_12_348/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_207 sky130_fd_sc_hd__clkbuf_1_265/X sky130_fd_sc_hd__clkbuf_1_266/X
+ sky130_fd_sc_hd__clkbuf_1_267/X sky130_fd_sc_hd__a22oi_1_207/A2 sky130_fd_sc_hd__a22oi_1_207/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_359 sky130_fd_sc_hd__buf_12_359/A sky130_fd_sc_hd__buf_12_359/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_218 sky130_fd_sc_hd__buf_2_164/X sky130_fd_sc_hd__nor2_4_8/Y
+ sky130_fd_sc_hd__clkbuf_1_424/X sky130_fd_sc_hd__buf_2_233/X sky130_fd_sc_hd__nand4_1_50/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_229 sky130_fd_sc_hd__nor2_4_7/Y sky130_fd_sc_hd__buf_2_165/X
+ sky130_fd_sc_hd__a22oi_1_229/B2 sky130_fd_sc_hd__clkbuf_1_448/X sky130_fd_sc_hd__a22oi_1_229/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_504 sky130_fd_sc_hd__a21oi_1_63/A1 sky130_fd_sc_hd__nor2_1_53/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_504/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_515 sky130_fd_sc_hd__nor2_1_56/B sky130_fd_sc_hd__fa_2_1032/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_515/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_526 sky130_fd_sc_hd__nor2_1_49/B sky130_fd_sc_hd__fa_2_1043/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_526/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_537 sky130_fd_sc_hd__a21oi_1_88/A2 sky130_fd_sc_hd__a21oi_1_97/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_537/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_548 sky130_fd_sc_hd__nand4_1_85/B sky130_fd_sc_hd__fa_2_972/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_548/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_559 sky130_fd_sc_hd__o22ai_1_120/B1 sky130_fd_sc_hd__fa_2_977/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_559/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_40 sky130_fd_sc_hd__nor2_1_40/B sky130_fd_sc_hd__nor3_1_37/C
+ sky130_fd_sc_hd__nor2_1_40/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_51 sky130_fd_sc_hd__nor2_1_51/B sky130_fd_sc_hd__nor2_1_51/Y
+ sky130_fd_sc_hd__nor2_1_51/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_62 sky130_fd_sc_hd__nor2_1_62/B sky130_fd_sc_hd__nor2_1_62/Y
+ sky130_fd_sc_hd__nor2_1_62/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_17 sky130_fd_sc_hd__clkinv_8_87/A sky130_fd_sc_hd__clkinv_8_20/A
+ VSS VDD VDD VSS VSS sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_73 sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__nor2_1_73/Y
+ sky130_fd_sc_hd__nor2_1_76/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_28 sky130_fd_sc_hd__clkinv_4_53/Y sky130_fd_sc_hd__clkinv_8_65/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_28/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_84 sky130_fd_sc_hd__nor2_1_84/B sky130_fd_sc_hd__nor2_1_84/Y
+ sky130_fd_sc_hd__nor2_1_84/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_39 sky130_fd_sc_hd__clkinv_4_39/A sky130_fd_sc_hd__dfxtp_1_87/D
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_39/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_95 sky130_fd_sc_hd__nor2_1_95/B sky130_fd_sc_hd__nor2_1_95/Y
+ sky130_fd_sc_hd__nor2_1_95/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_sram_2kbyte_1rw1r_32x512_8_3 sky130_fd_sc_hd__buf_6_1/A sky130_fd_sc_hd__buf_4_0/X
+ sky130_fd_sc_hd__buf_4_1/X sky130_fd_sc_hd__buf_6_2/X sky130_fd_sc_hd__buf_4_4/X
+ sky130_fd_sc_hd__buf_6_3/X sky130_fd_sc_hd__buf_4_6/X sky130_fd_sc_hd__buf_6_5/X
+ sky130_fd_sc_hd__buf_6_7/X sky130_fd_sc_hd__clkbuf_4_2/X sky130_fd_sc_hd__clkbuf_4_3/X
+ sky130_fd_sc_hd__clkbuf_1_127/X sky130_fd_sc_hd__buf_4_10/X sky130_fd_sc_hd__clkbuf_4_7/X
+ sky130_fd_sc_hd__buf_6_8/X sky130_fd_sc_hd__buf_4_12/X sky130_fd_sc_hd__buf_6_1/A
+ sky130_fd_sc_hd__buf_4_0/X sky130_fd_sc_hd__buf_4_1/X sky130_fd_sc_hd__buf_6_2/X
+ sky130_fd_sc_hd__buf_4_4/X sky130_fd_sc_hd__buf_6_3/X sky130_fd_sc_hd__buf_4_6/X
+ sky130_fd_sc_hd__buf_6_5/X sky130_fd_sc_hd__buf_6_7/X sky130_fd_sc_hd__clkbuf_4_2/X
+ sky130_fd_sc_hd__clkbuf_4_3/X sky130_fd_sc_hd__clkbuf_4_4/X sky130_fd_sc_hd__buf_4_10/X
+ sky130_fd_sc_hd__clkbuf_4_7/X sky130_fd_sc_hd__buf_6_8/X sky130_fd_sc_hd__buf_4_12/X
+ sky130_fd_sc_hd__buf_12_29/X sky130_fd_sc_hd__buf_12_31/X sky130_fd_sc_hd__buf_12_56/X
+ sky130_fd_sc_hd__buf_12_37/X sky130_fd_sc_hd__buf_12_14/X sky130_fd_sc_hd__buf_12_65/X
+ sky130_fd_sc_hd__buf_12_71/X sky130_fd_sc_hd__buf_12_17/X sky130_fd_sc_hd__buf_12_18/X
+ sky130_fd_sc_hd__buf_12_87/X sky130_fd_sc_hd__buf_12_22/X sky130_fd_sc_hd__buf_12_111/X
+ sky130_fd_sc_hd__buf_12_61/X sky130_fd_sc_hd__buf_12_104/X sky130_fd_sc_hd__buf_12_47/X
+ sky130_fd_sc_hd__buf_12_97/X sky130_fd_sc_hd__buf_12_107/X sky130_fd_sc_hd__buf_12_99/X
+ sky130_fd_sc_hd__buf_2_22/X sky130_fd_sc_hd__clkbuf_1_88/X sky130_fd_sc_hd__buf_2_22/X
+ sky130_fd_sc_hd__clkinv_8_0/Y sky130_fd_sc_hd__clkinv_8_5/Y sky130_fd_sc_hd__buf_12_83/X
+ sky130_fd_sc_hd__buf_12_82/X sky130_fd_sc_hd__buf_12_102/X sky130_fd_sc_hd__buf_12_85/X
+ sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[0] sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[1]
+ sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[2] sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[3]
+ sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[4] sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[5]
+ sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[6] sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[7]
+ sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[8] sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[9]
+ sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[10] sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[11]
+ sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[12] sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[13]
+ sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[14] sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[15]
+ sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[16] sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[17]
+ sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[18] sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[19]
+ sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[20] sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[21]
+ sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[22] sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[23]
+ sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[24] sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[25]
+ sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[26] sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[27]
+ sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[28] sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[29]
+ sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[30] sky130_sram_2kbyte_1rw1r_32x512_8_3/dout0[31]
+ sky130_fd_sc_hd__clkbuf_1_19/A sky130_fd_sc_hd__clkbuf_1_20/A sky130_fd_sc_hd__clkbuf_1_21/A
+ sky130_fd_sc_hd__clkbuf_1_22/A sky130_fd_sc_hd__clkbuf_1_23/A sky130_fd_sc_hd__clkbuf_1_24/A
+ sky130_fd_sc_hd__clkbuf_1_25/A sky130_fd_sc_hd__clkbuf_1_26/A sky130_fd_sc_hd__clkbuf_1_125/A
+ sky130_fd_sc_hd__clkbuf_1_28/A sky130_fd_sc_hd__clkbuf_1_29/A sky130_fd_sc_hd__clkbuf_1_30/A
+ sky130_fd_sc_hd__clkbuf_1_31/A sky130_fd_sc_hd__clkbuf_1_32/A sky130_fd_sc_hd__clkbuf_1_33/A
+ sky130_fd_sc_hd__clkbuf_1_34/A sky130_fd_sc_hd__a22oi_1_80/A2 sky130_fd_sc_hd__a22oi_1_76/A2
+ sky130_fd_sc_hd__a22oi_1_72/A2 sky130_fd_sc_hd__a22oi_1_68/A2 sky130_fd_sc_hd__a22oi_1_64/A2
+ sky130_fd_sc_hd__a22oi_1_61/A2 sky130_fd_sc_hd__a22oi_1_58/A2 sky130_fd_sc_hd__a22oi_1_55/A2
+ sky130_fd_sc_hd__a22oi_1_52/A2 sky130_fd_sc_hd__a22oi_1_49/A2 sky130_fd_sc_hd__a22oi_1_46/A2
+ sky130_fd_sc_hd__a22oi_1_43/A2 sky130_fd_sc_hd__a22oi_1_39/A2 sky130_fd_sc_hd__a22oi_1_35/A2
+ sky130_fd_sc_hd__a22oi_1_31/A2 sky130_fd_sc_hd__a22oi_1_28/A2 VDD VSS sky130_sram_2kbyte_1rw1r_32x512_8
Xsky130_fd_sc_hd__a21oi_1_401 sky130_fd_sc_hd__a21oi_1_404/A1 sky130_fd_sc_hd__a21oi_1_401/B1
+ sky130_fd_sc_hd__a21oi_1_401/Y sky130_fd_sc_hd__nand2_1_491/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_412 sky130_fd_sc_hd__nor3_1_40/A sky130_fd_sc_hd__o22ai_1_370/Y
+ sky130_fd_sc_hd__a21oi_1_412/Y sky130_fd_sc_hd__fa_2_1257/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_423 sky130_fd_sc_hd__o21a_1_59/B1 sky130_fd_sc_hd__o21a_1_58/A1
+ sky130_fd_sc_hd__a21oi_1_423/Y sky130_fd_sc_hd__nor2_1_271/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_434 sky130_fd_sc_hd__o21a_1_67/B1 sky130_fd_sc_hd__nor2_1_282/Y
+ sky130_fd_sc_hd__a21oi_1_434/Y sky130_fd_sc_hd__nor2_1_282/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_445 sky130_fd_sc_hd__o21ai_1_460/Y sky130_fd_sc_hd__nor2_1_300/Y
+ sky130_fd_sc_hd__a21oi_1_445/Y sky130_fd_sc_hd__nor2b_1_126/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_456 sky130_fd_sc_hd__nor2_2_18/Y sky130_fd_sc_hd__o21ai_1_466/Y
+ sky130_fd_sc_hd__nor2_1_301/B sky130_fd_sc_hd__fa_2_1290/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_467 sky130_fd_sc_hd__nor2b_2_5/Y sky130_fd_sc_hd__o21ai_1_481/Y
+ sky130_fd_sc_hd__a21oi_1_467/Y sky130_fd_sc_hd__o21ai_1_488/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_478 sky130_fd_sc_hd__nor3_1_41/A sky130_fd_sc_hd__o22ai_1_435/Y
+ sky130_fd_sc_hd__a21oi_1_478/Y sky130_fd_sc_hd__fa_2_1298/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_489 sky130_fd_sc_hd__nand2_1_569/A sky130_fd_sc_hd__or2_0_0/B
+ sky130_fd_sc_hd__nand2_1_557/A sky130_fd_sc_hd__nor2_1_317/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_8_103 sky130_fd_sc_hd__clkinv_8_104/A sky130_fd_sc_hd__clkinv_4_54/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_103/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_114 sky130_fd_sc_hd__clkinv_8_115/A sky130_fd_sc_hd__clkinv_8_114/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_114/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_125 sky130_fd_sc_hd__clkinv_4_64/A sky130_fd_sc_hd__clkinv_8_87/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_136 sky130_fd_sc_hd__clkinv_8_137/A sky130_fd_sc_hd__clkinv_8_136/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__o21a_1_5 sky130_fd_sc_hd__o21a_1_5/X sky130_fd_sc_hd__o21a_1_5/A1
+ sky130_fd_sc_hd__o21a_1_5/B1 sky130_fd_sc_hd__fa_2_982/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__nand2_1_450 sky130_fd_sc_hd__o21a_1_47/B1 sky130_fd_sc_hd__fa_2_1232/A
+ sky130_fd_sc_hd__o21a_1_47/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_461 sky130_fd_sc_hd__nand2_1_461/Y sky130_fd_sc_hd__xnor2_1_99/Y
+ sky130_fd_sc_hd__xor2_1_230/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_472 sky130_fd_sc_hd__nor2_1_251/B sky130_fd_sc_hd__nand2_1_472/B
+ sky130_fd_sc_hd__nor2_1_252/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_483 sky130_fd_sc_hd__nand2_1_483/Y sky130_fd_sc_hd__nor2b_2_4/Y
+ sky130_fd_sc_hd__o21ai_1_409/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_494 sky130_fd_sc_hd__o21a_1_55/A1 sky130_fd_sc_hd__nor2_2_17/B
+ sky130_fd_sc_hd__nor2_4_18/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_30 sky130_fd_sc_hd__ha_2_60/SUM sky130_fd_sc_hd__nor2b_1_30/Y
+ sky130_fd_sc_hd__or2_0_2/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_41 sky130_fd_sc_hd__ha_2_81/SUM sky130_fd_sc_hd__nor2b_1_41/Y
+ sky130_fd_sc_hd__or2_0_3/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_52 sky130_fd_sc_hd__nor2_1_23/A sky130_fd_sc_hd__nor2b_1_52/Y
+ sky130_fd_sc_hd__nor2b_1_52/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_63 sky130_fd_sc_hd__dfxtp_1_483/Q sky130_fd_sc_hd__nor2b_1_63/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1030 sky130_fd_sc_hd__nor2_4_20/B sky130_fd_sc_hd__nor2_8_2/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1030/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_74 sky130_fd_sc_hd__nor2_1_39/A sky130_fd_sc_hd__nor2b_1_74/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1041 sky130_fd_sc_hd__nor2_1_273/A sky130_fd_sc_hd__nor2_1_274/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1041/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_85 sky130_fd_sc_hd__fa_2_953/A sky130_fd_sc_hd__nor3_1_35/C
+ sky130_fd_sc_hd__nor2b_1_85/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1052 sky130_fd_sc_hd__o22ai_1_399/A1 sky130_fd_sc_hd__fa_2_0/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1052/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_96 sky130_fd_sc_hd__o21ai_1_89/Y sky130_fd_sc_hd__nor2b_1_96/Y
+ sky130_fd_sc_hd__buf_2_262/X VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1063 sky130_fd_sc_hd__nor2_1_290/B sky130_fd_sc_hd__xor2_1_275/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1063/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_4 VSS VDD sky130_fd_sc_hd__xnor2_1_4/B sky130_fd_sc_hd__xnor2_1_4/Y
+ sky130_fd_sc_hd__fa_2_699/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_1074 sky130_fd_sc_hd__nor2_1_300/A sky130_fd_sc_hd__xor2_1_299/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1074/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1085 sky130_fd_sc_hd__o21ai_1_468/A1 sky130_fd_sc_hd__o21ai_1_470/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1085/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1096 sky130_fd_sc_hd__nor2_1_277/B sky130_fd_sc_hd__fa_2_1308/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1096/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_290 VDD VSS sky130_fd_sc_hd__a22o_1_57/A1 sky130_fd_sc_hd__clkinv_4_31/Y
+ sky130_fd_sc_hd__nand2_1_129/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_140 sky130_fd_sc_hd__fa_2_23/CIN sky130_fd_sc_hd__fa_2_136/A
+ sky130_fd_sc_hd__ha_2_97/A sky130_fd_sc_hd__ha_2_99/A sky130_fd_sc_hd__fa_2_76/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_151 sky130_fd_sc_hd__fa_2_142/A sky130_fd_sc_hd__fa_2_143/B
+ sky130_fd_sc_hd__fa_2_238/B sky130_fd_sc_hd__fa_2_151/B sky130_fd_sc_hd__fa_2_154/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_162 sky130_fd_sc_hd__fa_2_158/B sky130_fd_sc_hd__fa_2_161/B
+ sky130_fd_sc_hd__fa_2_162/A sky130_fd_sc_hd__fa_2_162/B sky130_fd_sc_hd__fa_2_162/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_19 VDD VSS sky130_fd_sc_hd__ha_2_113/B sky130_fd_sc_hd__dfxtp_1_26/CLK
+ sky130_fd_sc_hd__nand4_1_37/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_173 sky130_fd_sc_hd__maj3_1_54/B sky130_fd_sc_hd__maj3_1_55/A
+ sky130_fd_sc_hd__fa_2_31/A sky130_fd_sc_hd__ha_2_99/B sky130_fd_sc_hd__fa_2_67/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_184 sky130_fd_sc_hd__fa_2_186/B sky130_fd_sc_hd__fa_2_184/SUM
+ sky130_fd_sc_hd__fa_2_242/B sky130_fd_sc_hd__fa_2_280/B sky130_fd_sc_hd__fa_2_184/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_195 sky130_fd_sc_hd__fa_2_194/CIN sky130_fd_sc_hd__fa_2_195/SUM
+ sky130_fd_sc_hd__fa_2_5/B sky130_fd_sc_hd__ha_2_91/A sky130_fd_sc_hd__fa_2_280/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o22ai_1_50 sky130_fd_sc_hd__fa_2_807/B sky130_fd_sc_hd__ha_2_142/B
+ sky130_fd_sc_hd__o22ai_1_50/Y sky130_fd_sc_hd__fa_2_806/A sky130_fd_sc_hd__ha_2_140/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_61 sky130_fd_sc_hd__o22ai_1_88/B1 sky130_fd_sc_hd__nand2_2_3/Y
+ sky130_fd_sc_hd__o22ai_1_61/Y sky130_fd_sc_hd__xnor2_1_33/Y sky130_fd_sc_hd__o22ai_1_75/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_72 sky130_fd_sc_hd__o22ai_1_88/B1 sky130_fd_sc_hd__nand2_2_3/Y
+ sky130_fd_sc_hd__o22ai_1_72/Y sky130_fd_sc_hd__xnor2_1_55/Y sky130_fd_sc_hd__o22ai_1_86/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_190 VDD VSS sky130_fd_sc_hd__buf_2_190/X sky130_fd_sc_hd__buf_2_190/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__clkbuf_4_109 sky130_fd_sc_hd__clkbuf_4_109/X sky130_fd_sc_hd__nand2_1_568/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o22ai_1_83 sky130_fd_sc_hd__o22ai_1_89/A1 sky130_fd_sc_hd__o22ai_1_88/B1
+ sky130_fd_sc_hd__o22ai_1_83/Y sky130_fd_sc_hd__xnor2_1_49/Y sky130_fd_sc_hd__o22ai_1_83/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_94 sky130_fd_sc_hd__nor2_2_9/B sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__o22ai_1_94/Y sky130_fd_sc_hd__a21oi_1_95/Y sky130_fd_sc_hd__nor2_1_83/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_4_30 VDD VSS sky130_fd_sc_hd__buf_4_30/X sky130_fd_sc_hd__inv_2_44/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_41 VDD VSS sky130_fd_sc_hd__buf_4_41/X sky130_fd_sc_hd__buf_4_41/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_52 VDD VSS sky130_fd_sc_hd__buf_4_52/X sky130_fd_sc_hd__buf_8_80/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_63 VDD VSS sky130_fd_sc_hd__buf_4_63/X sky130_fd_sc_hd__buf_4_63/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_74 VDD VSS sky130_fd_sc_hd__buf_4_74/X sky130_fd_sc_hd__buf_4_74/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_85 VDD VSS sky130_fd_sc_hd__buf_4_85/X sky130_fd_sc_hd__buf_4_85/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_96 VDD VSS sky130_fd_sc_hd__buf_4_96/X sky130_fd_sc_hd__buf_4_96/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_12_101 sky130_fd_sc_hd__buf_12_79/X sky130_fd_sc_hd__buf_12_101/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_112 sky130_fd_sc_hd__buf_12_112/A sky130_fd_sc_hd__buf_12_119/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_123 sky130_fd_sc_hd__buf_12_133/A sky130_fd_sc_hd__buf_12_248/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_134 sky130_fd_sc_hd__buf_12_134/A sky130_fd_sc_hd__buf_12_251/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_145 sky130_fd_sc_hd__buf_12_145/A sky130_fd_sc_hd__buf_12_235/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_156 sky130_fd_sc_hd__buf_4_44/A sky130_fd_sc_hd__buf_12_246/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_167 sky130_fd_sc_hd__buf_12_167/A sky130_fd_sc_hd__buf_12_242/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_90 VSS VDD sky130_fd_sc_hd__clkbuf_1_91/A sky130_fd_sc_hd__nand3_1_20/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_4_4 sky130_fd_sc_hd__clkbuf_4_4/X sky130_fd_sc_hd__buf_2_8/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_12_178 sky130_fd_sc_hd__buf_8_103/X sky130_fd_sc_hd__buf_12_178/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_189 sky130_fd_sc_hd__bufinv_8_3/Y sky130_fd_sc_hd__buf_12_189/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_301 sky130_fd_sc_hd__fa_2_283/A sky130_fd_sc_hd__fa_2_32/A
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_312 sky130_fd_sc_hd__fa_2_425/B sky130_fd_sc_hd__ha_2_116/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_312/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_323 sky130_fd_sc_hd__fa_2_546/B sky130_fd_sc_hd__ha_2_122/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_323/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_334 sky130_fd_sc_hd__fa_2_564/B sky130_fd_sc_hd__ha_2_121/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_334/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_345 sky130_fd_sc_hd__ha_2_132/B sky130_fd_sc_hd__fa_2_672/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_345/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_356 sky130_fd_sc_hd__ha_2_139/B sky130_fd_sc_hd__ha_2_144/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_356/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_367 sky130_fd_sc_hd__ha_2_138/A sky130_fd_sc_hd__ha_2_143/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_367/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_378 sky130_fd_sc_hd__fa_2_870/B sky130_fd_sc_hd__dfxtp_1_270/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_378/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_389 sky130_fd_sc_hd__fa_2_883/B sky130_fd_sc_hd__nor2_1_23/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_389/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21a_1_19 sky130_fd_sc_hd__o21a_1_19/X sky130_fd_sc_hd__o21a_1_19/A1
+ sky130_fd_sc_hd__o21a_1_19/B1 sky130_fd_sc_hd__fa_2_1134/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__a21oi_1_220 sky130_fd_sc_hd__a21o_2_5/A2 sky130_fd_sc_hd__o21ai_1_255/Y
+ sky130_fd_sc_hd__a21oi_1_220/Y sky130_fd_sc_hd__fa_2_1089/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_231 sky130_fd_sc_hd__a21o_2_5/A2 sky130_fd_sc_hd__o21ai_1_267/Y
+ sky130_fd_sc_hd__a21oi_1_231/Y sky130_fd_sc_hd__fa_2_1078/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_242 sky130_fd_sc_hd__o21a_1_19/B1 sky130_fd_sc_hd__o21a_1_18/A1
+ sky130_fd_sc_hd__dfxtp_1_905/D sky130_fd_sc_hd__nor2_1_143/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_253 sky130_fd_sc_hd__nor2_1_154/A sky130_fd_sc_hd__o21a_1_27/A1
+ sky130_fd_sc_hd__dfxtp_1_883/D sky130_fd_sc_hd__nor2_1_154/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_264 sky130_fd_sc_hd__clkinv_1_819/Y sky130_fd_sc_hd__clkinv_1_818/Y
+ sky130_fd_sc_hd__a21oi_1_264/Y sky130_fd_sc_hd__nand2_1_387/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_275 sky130_fd_sc_hd__fa_2_1130/A sky130_fd_sc_hd__o22ai_1_246/Y
+ sky130_fd_sc_hd__a21oi_1_275/Y sky130_fd_sc_hd__nor2_2_15/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_286 sky130_fd_sc_hd__o21ai_1_322/Y sky130_fd_sc_hd__o21ai_1_317/Y
+ sky130_fd_sc_hd__a21oi_1_286/Y sky130_fd_sc_hd__nor2b_1_105/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_4_4 sky130_fd_sc_hd__clkinv_8_7/Y sky130_fd_sc_hd__clkinv_4_7/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_4/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__a21oi_1_297 sky130_fd_sc_hd__clkinv_1_779/Y sky130_fd_sc_hd__o22ai_1_263/Y
+ sky130_fd_sc_hd__a21oi_1_297/Y sky130_fd_sc_hd__fa_2_1155/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_205 sky130_fd_sc_hd__buf_8_205/A sky130_fd_sc_hd__buf_8_205/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_216 sky130_fd_sc_hd__buf_8_216/A sky130_fd_sc_hd__buf_8_216/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nand2_1_280 sky130_fd_sc_hd__o21a_1_8/A2 sky130_fd_sc_hd__nor2_2_8/B
+ sky130_fd_sc_hd__nor2_2_7/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_108 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1049/B
+ sky130_fd_sc_hd__xor2_1_108/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_291 sky130_fd_sc_hd__xnor2_1_81/B sky130_fd_sc_hd__nand2_1_291/B
+ sky130_fd_sc_hd__nand2_1_296/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_890 sky130_fd_sc_hd__nor2_1_198/B sky130_fd_sc_hd__fa_2_1195/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_890/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor2_1_119 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1087/B
+ sky130_fd_sc_hd__xor2_1_119/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkinv_1_18 sky130_fd_sc_hd__nand3_2_0/B sky130_fd_sc_hd__ha_2_20/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_18/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_29 sky130_fd_sc_hd__inv_2_18/A sky130_fd_sc_hd__inv_2_9/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_29/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_5 sky130_fd_sc_hd__fa_2_3/B sky130_fd_sc_hd__fa_2_4/B sky130_fd_sc_hd__fa_2_5/A
+ sky130_fd_sc_hd__fa_2_5/B sky130_fd_sc_hd__fa_2_2/B VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_909 sky130_fd_sc_hd__fa_2_893/A sky130_fd_sc_hd__fa_2_894/B
+ sky130_fd_sc_hd__fa_2_909/A sky130_fd_sc_hd__fa_2_909/B sky130_fd_sc_hd__fa_2_909/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a211o_1_11 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_133/A sky130_fd_sc_hd__o21ai_1_239/Y
+ sky130_fd_sc_hd__nor2_1_124/Y sky130_fd_sc_hd__nand2_1_331/B sky130_fd_sc_hd__o22ai_1_167/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__a211o_1_22 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_223/A sky130_fd_sc_hd__o21ai_1_348/Y
+ sky130_fd_sc_hd__nor2_1_207/Y sky130_fd_sc_hd__nor2b_2_3/Y sky130_fd_sc_hd__o22ai_1_298/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__mux2_2_209 VSS VDD sky130_fd_sc_hd__mux2_2_209/A1 sky130_fd_sc_hd__mux2_2_209/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_209/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__clkinv_1_120 sky130_fd_sc_hd__a22o_2_3/B1 sky130_fd_sc_hd__nor2_1_3/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_120/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_131 sky130_fd_sc_hd__clkinv_2_9/A sky130_fd_sc_hd__clkinv_1_131/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_131/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_142 sky130_fd_sc_hd__inv_2_77/A sky130_fd_sc_hd__a22o_2_0/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_142/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_153 sky130_fd_sc_hd__clkinv_1_155/A sky130_fd_sc_hd__clkinv_1_153/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_153/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_164 sky130_fd_sc_hd__inv_2_95/A sky130_fd_sc_hd__inv_2_74/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_164/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_175 sky130_fd_sc_hd__bufinv_8_4/A sky130_fd_sc_hd__buf_8_155/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_175/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_7 sky130_fd_sc_hd__inv_2_8/Y sky130_fd_sc_hd__buf_8_7/X VSS
+ VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__a22o_1_9 sky130_fd_sc_hd__a22o_1_9/A1 sky130_fd_sc_hd__nor2_1_1/Y
+ sky130_fd_sc_hd__a22o_1_9/X sky130_fd_sc_hd__a22o_1_9/B2 sky130_fd_sc_hd__nor2_1_0/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_186 sky130_fd_sc_hd__nor2_1_6/B sky130_fd_sc_hd__nor2_1_7/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_186/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_11 sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__ha_2_62/A
+ sky130_fd_sc_hd__buf_8_140/A sky130_fd_sc_hd__dfxtp_1_9/Q sky130_fd_sc_hd__a22o_2_3/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_197 sky130_fd_sc_hd__inv_2_105/A sky130_fd_sc_hd__a22o_2_7/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_197/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_22 sky130_fd_sc_hd__nor2_4_4/Y sky130_fd_sc_hd__ha_2_79/B
+ sky130_fd_sc_hd__a22o_1_22/X sky130_fd_sc_hd__a22o_1_22/B2 sky130_fd_sc_hd__a22o_2_6/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_33 sky130_fd_sc_hd__nor4_1_5/Y sky130_fd_sc_hd__nor4_1_9/Y
+ sky130_fd_sc_hd__a22o_1_33/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__a22o_1_33/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_44 sky130_fd_sc_hd__a22o_1_44/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_44/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__fa_2_950/SUM
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_55 sky130_fd_sc_hd__a22o_1_55/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_55/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__nor4_1_10/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_66 sky130_fd_sc_hd__a22o_1_68/A1 sky130_fd_sc_hd__a22o_1_68/B2
+ sky130_fd_sc_hd__a22o_1_66/X sky130_fd_sc_hd__ha_2_185/SUM sky130_fd_sc_hd__a22o_1_68/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__nand4_1_5 sky130_fd_sc_hd__nand4_1_5/C sky130_fd_sc_hd__nand4_1_5/B
+ sky130_fd_sc_hd__nand4_1_5/Y sky130_fd_sc_hd__nand4_1_5/D sky130_fd_sc_hd__nand4_1_5/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__clkinv_2_1 sky130_fd_sc_hd__clkinv_8_1/A sky130_fd_sc_hd__clkinv_8_9/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_1/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__nor2_1_280 sky130_fd_sc_hd__nor2_1_280/B sky130_fd_sc_hd__o21a_1_65/A1
+ sky130_fd_sc_hd__o21a_1_66/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_291 sky130_fd_sc_hd__nor2_1_291/B sky130_fd_sc_hd__nor2_1_291/Y
+ sky130_fd_sc_hd__nor2_1_309/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__maj3_1_17 sky130_fd_sc_hd__maj3_1_18/X sky130_fd_sc_hd__maj3_1_17/X
+ sky130_fd_sc_hd__maj3_1_17/B sky130_fd_sc_hd__maj3_1_17/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_28 sky130_fd_sc_hd__maj3_1_29/X sky130_fd_sc_hd__maj3_1_28/X
+ sky130_fd_sc_hd__maj3_1_28/B sky130_fd_sc_hd__maj3_1_28/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_407 sky130_fd_sc_hd__nor2_1_310/A sky130_fd_sc_hd__nor2_1_307/A
+ sky130_fd_sc_hd__o22ai_1_407/Y sky130_fd_sc_hd__a21boi_1_8/Y sky130_fd_sc_hd__nor2_1_291/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__maj3_1_39 sky130_fd_sc_hd__maj3_1_40/X sky130_fd_sc_hd__maj3_1_39/X
+ sky130_fd_sc_hd__maj3_1_39/B sky130_fd_sc_hd__maj3_1_39/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_418 sky130_fd_sc_hd__o22ai_1_436/A2 sky130_fd_sc_hd__nor2_1_270/B
+ sky130_fd_sc_hd__o22ai_1_418/Y sky130_fd_sc_hd__o22ai_1_418/A1 sky130_fd_sc_hd__o32ai_1_11/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_429 sky130_fd_sc_hd__o22ai_1_436/A2 sky130_fd_sc_hd__o22ai_1_429/B1
+ sky130_fd_sc_hd__o22ai_1_429/Y sky130_fd_sc_hd__nor2_1_281/B sky130_fd_sc_hd__o32ai_1_11/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__a22oi_1_390 sky130_fd_sc_hd__nor3_1_40/B sky130_fd_sc_hd__fa_2_1241/A
+ sky130_fd_sc_hd__xor2_1_254/A sky130_fd_sc_hd__clkinv_1_946/Y sky130_fd_sc_hd__a22oi_1_390/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nand2_1_12 sky130_fd_sc_hd__nand3_1_12/C sky130_fd_sc_hd__nand4_1_67/Y
+ sky130_fd_sc_hd__nand2_1_9/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_23 sky130_fd_sc_hd__nor2_4_6/B sky130_fd_sc_hd__nor3_2_4/B
+ sky130_fd_sc_hd__nor3_1_9/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_34 sky130_fd_sc_hd__xor2_1_11/A sky130_fd_sc_hd__nor2b_1_51/Y
+ sky130_fd_sc_hd__nand2_1_34/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_45 sky130_fd_sc_hd__nand2_1_45/Y sky130_fd_sc_hd__nand2_1_45/B
+ sky130_fd_sc_hd__a21oi_2_0/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_56 sky130_fd_sc_hd__nand2_1_56/Y sky130_fd_sc_hd__nand2_1_57/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_67 sky130_fd_sc_hd__nand2_1_67/Y sky130_fd_sc_hd__nand2_1_8/B
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_78 sky130_fd_sc_hd__nand2_1_78/Y sky130_fd_sc_hd__nand2_1_79/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_89 sky130_fd_sc_hd__nand2_1_89/Y sky130_fd_sc_hd__nand2_1_89/B
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__fa_2_19 sky130_fd_sc_hd__fa_2_16/CIN sky130_fd_sc_hd__fa_2_19/SUM
+ sky130_fd_sc_hd__fa_2_19/A sky130_fd_sc_hd__fa_2_19/B sky130_fd_sc_hd__fa_2_19/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_sram_2kbyte_1rw1r_32x512_8_15 sky130_fd_sc_hd__clkbuf_4_160/X sky130_fd_sc_hd__clkbuf_4_161/X
+ sky130_fd_sc_hd__buf_4_120/A sky130_fd_sc_hd__clkbuf_4_162/X sky130_fd_sc_hd__buf_4_98/X
+ sky130_fd_sc_hd__clkbuf_4_210/A sky130_fd_sc_hd__clkbuf_4_163/X sky130_fd_sc_hd__clkbuf_4_164/X
+ sky130_fd_sc_hd__buf_4_99/X sky130_fd_sc_hd__buf_4_100/X sky130_fd_sc_hd__buf_6_54/X
+ sky130_fd_sc_hd__buf_4_101/X sky130_fd_sc_hd__buf_4_102/X sky130_fd_sc_hd__buf_4_103/X
+ sky130_fd_sc_hd__buf_4_104/X sky130_fd_sc_hd__buf_4_105/X sky130_fd_sc_hd__clkbuf_4_160/X
+ sky130_fd_sc_hd__clkbuf_4_161/X sky130_fd_sc_hd__buf_4_120/A sky130_fd_sc_hd__clkbuf_4_162/X
+ sky130_fd_sc_hd__buf_4_98/X sky130_fd_sc_hd__clkbuf_4_210/X sky130_fd_sc_hd__clkbuf_4_163/X
+ sky130_fd_sc_hd__clkbuf_4_164/X sky130_fd_sc_hd__buf_4_99/X sky130_fd_sc_hd__buf_4_100/X
+ sky130_fd_sc_hd__buf_6_54/X sky130_fd_sc_hd__buf_4_101/X sky130_fd_sc_hd__buf_4_102/X
+ sky130_fd_sc_hd__buf_4_103/X sky130_fd_sc_hd__buf_4_104/X sky130_fd_sc_hd__buf_4_105/X
+ sky130_fd_sc_hd__buf_12_490/X sky130_fd_sc_hd__buf_12_516/X sky130_fd_sc_hd__buf_12_495/X
+ sky130_fd_sc_hd__buf_12_399/X sky130_fd_sc_hd__buf_12_413/X sky130_fd_sc_hd__buf_12_390/X
+ sky130_fd_sc_hd__buf_12_475/X sky130_fd_sc_hd__buf_12_480/X sky130_fd_sc_hd__buf_12_465/X
+ sky130_fd_sc_hd__buf_12_412/X sky130_fd_sc_hd__buf_12_439/X sky130_fd_sc_hd__buf_12_491/X
+ sky130_fd_sc_hd__buf_12_514/X sky130_fd_sc_hd__buf_12_388/X sky130_fd_sc_hd__buf_12_494/X
+ sky130_fd_sc_hd__buf_12_484/X sky130_fd_sc_hd__buf_12_435/X sky130_fd_sc_hd__buf_12_428/X
+ sky130_fd_sc_hd__clkinv_1_225/Y sky130_fd_sc_hd__buf_2_163/X sky130_fd_sc_hd__buf_2_242/X
+ sky130_fd_sc_hd__clkinv_8_36/Y sky130_fd_sc_hd__clkinv_8_32/Y sky130_fd_sc_hd__buf_12_416/X
+ sky130_fd_sc_hd__buf_12_411/X sky130_fd_sc_hd__buf_12_487/X sky130_fd_sc_hd__buf_12_466/X
+ sky130_fd_sc_hd__clkbuf_1_541/A sky130_fd_sc_hd__clkbuf_1_383/A sky130_fd_sc_hd__clkbuf_1_384/A
+ sky130_fd_sc_hd__inv_2_136/A sky130_fd_sc_hd__clkbuf_1_386/A sky130_fd_sc_hd__clkbuf_1_387/A
+ sky130_fd_sc_hd__clkbuf_1_388/A sky130_fd_sc_hd__clkbuf_1_389/A sky130_fd_sc_hd__clkbuf_1_390/A
+ sky130_fd_sc_hd__clkbuf_1_391/A sky130_fd_sc_hd__clkbuf_1_392/A sky130_fd_sc_hd__clkbuf_1_393/A
+ sky130_fd_sc_hd__clkbuf_1_394/A sky130_fd_sc_hd__clkbuf_1_395/A sky130_fd_sc_hd__clkbuf_1_396/A
+ sky130_fd_sc_hd__clkbuf_1_397/A sky130_fd_sc_hd__a22oi_1_254/A2 sky130_fd_sc_hd__a22oi_1_250/A2
+ sky130_fd_sc_hd__a22oi_1_247/A2 sky130_fd_sc_hd__a22oi_1_244/A2 sky130_fd_sc_hd__a22oi_1_241/A2
+ sky130_fd_sc_hd__a22oi_2_25/A2 sky130_fd_sc_hd__a22oi_2_24/A2 sky130_fd_sc_hd__a22oi_2_22/A2
+ sky130_fd_sc_hd__a22oi_1_231/A2 sky130_fd_sc_hd__a22oi_2_20/A2 sky130_fd_sc_hd__a22oi_1_224/A2
+ sky130_fd_sc_hd__a22oi_2_19/A2 sky130_fd_sc_hd__a22oi_2_17/A2 sky130_fd_sc_hd__a22oi_2_15/A2
+ sky130_fd_sc_hd__a22oi_2_14/A2 sky130_fd_sc_hd__a22oi_2_13/A2 sky130_fd_sc_hd__clkbuf_1_398/A
+ sky130_fd_sc_hd__clkbuf_1_399/A sky130_fd_sc_hd__clkbuf_1_400/A sky130_fd_sc_hd__clkbuf_1_401/A
+ sky130_fd_sc_hd__clkbuf_1_402/A sky130_fd_sc_hd__clkbuf_1_403/A sky130_fd_sc_hd__clkbuf_1_404/A
+ sky130_fd_sc_hd__clkbuf_1_405/A sky130_fd_sc_hd__clkbuf_1_406/A sky130_fd_sc_hd__clkbuf_1_407/A
+ sky130_fd_sc_hd__clkbuf_1_408/A sky130_fd_sc_hd__clkbuf_1_409/A sky130_fd_sc_hd__clkbuf_1_410/A
+ sky130_fd_sc_hd__clkbuf_1_524/A sky130_fd_sc_hd__clkbuf_1_412/A sky130_fd_sc_hd__clkbuf_1_413/A
+ sky130_fd_sc_hd__a22oi_1_317/A2 sky130_fd_sc_hd__a22oi_1_313/A2 sky130_fd_sc_hd__a22oi_1_309/A2
+ sky130_fd_sc_hd__a22oi_1_305/A2 sky130_fd_sc_hd__a22oi_1_301/A2 sky130_fd_sc_hd__a22oi_1_297/A2
+ sky130_fd_sc_hd__a22oi_1_293/A2 sky130_fd_sc_hd__a22oi_1_289/A2 sky130_fd_sc_hd__a22oi_1_285/A2
+ sky130_fd_sc_hd__a22oi_1_281/A2 sky130_fd_sc_hd__clkbuf_1_532/A sky130_fd_sc_hd__a22oi_1_273/A2
+ sky130_fd_sc_hd__a22oi_1_269/A2 sky130_fd_sc_hd__a22oi_1_265/A2 sky130_fd_sc_hd__a22oi_1_261/A2
+ sky130_fd_sc_hd__a22oi_1_257/A2 VDD VSS sky130_sram_2kbyte_1rw1r_32x512_8
Xsky130_fd_sc_hd__dfxtp_1_1207 VDD VSS sky130_fd_sc_hd__fa_2_1256/A sky130_fd_sc_hd__clkinv_8_116/Y
+ sky130_fd_sc_hd__mux2_2_180/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1218 VDD VSS sky130_fd_sc_hd__fa_2_1230/A sky130_fd_sc_hd__clkinv_8_78/Y
+ sky130_fd_sc_hd__mux2_2_201/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1229 VDD VSS sky130_fd_sc_hd__fa_2_1241/A sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__mux2_2_175/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_801 VDD VSS sky130_fd_sc_hd__fa_2_1053/A sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__mux2_2_73/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_812 VDD VSS sky130_fd_sc_hd__fa_2_1064/A sky130_fd_sc_hd__clkinv_4_26/Y
+ sky130_fd_sc_hd__mux2_2_49/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_823 VDD VSS sky130_fd_sc_hd__fa_2_1097/A sky130_fd_sc_hd__clkinv_8_59/Y
+ sky130_fd_sc_hd__and2_0_299/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_834 VDD VSS sky130_fd_sc_hd__nand2_1_339/A sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__nor2b_1_102/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_845 VDD VSS sky130_fd_sc_hd__mux2_2_63/A1 sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__o21ai_1_162/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_856 VDD VSS sky130_fd_sc_hd__mux2_2_41/A1 sky130_fd_sc_hd__clkinv_4_25/Y
+ sky130_fd_sc_hd__o21ai_1_173/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_867 VDD VSS sky130_fd_sc_hd__mux2_2_58/A1 sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__o21ai_1_181/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_878 VDD VSS sky130_fd_sc_hd__ha_2_147/A sky130_fd_sc_hd__dfxtp_1_899/CLK
+ sky130_fd_sc_hd__o32ai_1_1/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_889 VDD VSS sky130_fd_sc_hd__fa_2_853/A sky130_fd_sc_hd__clkinv_4_22/Y
+ sky130_fd_sc_hd__dfxtp_1_889/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_410 VSS VDD sky130_fd_sc_hd__clkbuf_1_410/X sky130_fd_sc_hd__clkbuf_1_410/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_421 VSS VDD sky130_fd_sc_hd__clkbuf_1_421/X sky130_fd_sc_hd__clkbuf_1_421/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_432 VSS VDD sky130_fd_sc_hd__clkbuf_1_432/X sky130_fd_sc_hd__clkbuf_1_432/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_443 VSS VDD sky130_fd_sc_hd__a22oi_2_27/A2 sky130_fd_sc_hd__clkbuf_1_443/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_454 VSS VDD sky130_fd_sc_hd__clkbuf_1_454/X sky130_fd_sc_hd__clkbuf_1_454/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_465 VSS VDD sky130_fd_sc_hd__clkbuf_1_465/X sky130_fd_sc_hd__clkbuf_1_465/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_476 VSS VDD sky130_fd_sc_hd__nand4_1_60/D sky130_fd_sc_hd__a22oi_1_244/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_487 VSS VDD sky130_fd_sc_hd__buf_8_207/A sky130_fd_sc_hd__inv_2_112/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_706 sky130_fd_sc_hd__fa_2_705/CIN sky130_fd_sc_hd__fa_2_706/SUM
+ sky130_fd_sc_hd__fa_2_706/A sky130_fd_sc_hd__fa_2_706/B sky130_fd_sc_hd__fa_2_706/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_498 VSS VDD sky130_fd_sc_hd__a22oi_2_26/B2 sky130_fd_sc_hd__clkbuf_1_498/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_717 sky130_fd_sc_hd__maj3_1_159/B sky130_fd_sc_hd__maj3_1_160/A
+ sky130_fd_sc_hd__ha_2_143/A sky130_fd_sc_hd__ha_2_141/B sky130_fd_sc_hd__fa_2_758/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_728 sky130_fd_sc_hd__fa_2_730/CIN sky130_fd_sc_hd__fa_2_726/A
+ sky130_fd_sc_hd__ha_2_145/B sky130_fd_sc_hd__ha_2_142/B sky130_fd_sc_hd__ha_2_139/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_739 sky130_fd_sc_hd__fa_2_741/B sky130_fd_sc_hd__fa_2_739/SUM
+ sky130_fd_sc_hd__fa_2_739/A sky130_fd_sc_hd__fa_2_739/B sky130_fd_sc_hd__fa_2_743/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor2b_1_103 sky130_fd_sc_hd__o21ai_1_207/Y sky130_fd_sc_hd__nor2b_1_103/Y
+ sky130_fd_sc_hd__buf_2_262/X VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_114 sky130_fd_sc_hd__nor3_1_39/Y sky130_fd_sc_hd__nor2b_1_114/Y
+ sky130_fd_sc_hd__buf_2_262/X VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_125 sky130_fd_sc_hd__o22ai_1_323/Y sky130_fd_sc_hd__nor2b_1_125/Y
+ sky130_fd_sc_hd__buf_2_262/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_136 sky130_fd_sc_hd__o2bb2ai_1_33/Y sky130_fd_sc_hd__nor2b_1_136/Y
+ sky130_fd_sc_hd__nor4_1_13/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__buf_6_4 VDD VSS sky130_fd_sc_hd__buf_6_4/X sky130_fd_sc_hd__buf_6_4/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__bufbuf_8_7 sky130_fd_sc_hd__buf_2_240/X sky130_fd_sc_hd__bufbuf_8_7/X
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufbuf_8
Xsky130_fd_sc_hd__o22ai_1_204 sky130_fd_sc_hd__nor2_1_138/A sky130_fd_sc_hd__o22ai_1_204/B1
+ sky130_fd_sc_hd__o22ai_1_204/Y sky130_fd_sc_hd__o22ai_1_206/B1 sky130_fd_sc_hd__o22ai_1_206/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__sdlclkp_4_2 sky130_fd_sc_hd__conb_1_1/LO sky130_fd_sc_hd__clkinv_8_47/A
+ sky130_fd_sc_hd__clkinv_4_79/A sky130_fd_sc_hd__nor3_2_1/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__o22ai_1_215 sky130_fd_sc_hd__nand2_1_358/Y sky130_fd_sc_hd__nand2_1_357/Y
+ sky130_fd_sc_hd__o22ai_1_215/Y sky130_fd_sc_hd__o22ai_1_228/A1 sky130_fd_sc_hd__a21o_2_8/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_226 sky130_fd_sc_hd__nand2_1_360/Y sky130_fd_sc_hd__nand2_1_359/Y
+ sky130_fd_sc_hd__o22ai_1_226/Y sky130_fd_sc_hd__o22ai_1_226/A1 sky130_fd_sc_hd__a21o_2_7/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_237 sky130_fd_sc_hd__o32ai_1_1/B2 sky130_fd_sc_hd__nor2_1_182/A
+ sky130_fd_sc_hd__o22ai_1_237/Y sky130_fd_sc_hd__o22ai_1_262/A1 sky130_fd_sc_hd__a222oi_1_4/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_248 sky130_fd_sc_hd__o22ai_1_261/A2 sky130_fd_sc_hd__nor2_1_145/B
+ sky130_fd_sc_hd__o22ai_1_248/Y sky130_fd_sc_hd__nor2_1_146/B sky130_fd_sc_hd__o32ai_1_2/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_259 sky130_fd_sc_hd__o22ai_1_261/A2 sky130_fd_sc_hd__o22ai_1_259/B1
+ sky130_fd_sc_hd__o22ai_1_259/Y sky130_fd_sc_hd__nor2_1_150/B sky130_fd_sc_hd__o32ai_1_2/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_1_5 sky130_fd_sc_hd__nor2_2_3/B sky130_fd_sc_hd__nor2_1_5/Y
+ sky130_fd_sc_hd__nor3_2_6/C VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__bufinv_8_7 sky130_fd_sc_hd__bufinv_8_7/A sky130_fd_sc_hd__bufinv_8_7/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufinv_8
Xsky130_fd_sc_hd__dfxtp_1_108 VDD VSS sky130_fd_sc_hd__nor4_1_4/B sky130_fd_sc_hd__dfxtp_1_111/CLK
+ sky130_fd_sc_hd__ha_2_8/SUM VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_119 VDD VSS sky130_fd_sc_hd__or2_0_0/A sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__and2_0_1/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_420 VSS VDD sky130_fd_sc_hd__a211oi_1_30/Y sky130_fd_sc_hd__nor2_1_267/A
+ sky130_fd_sc_hd__nand2_1_486/Y sky130_fd_sc_hd__xor2_1_237/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_431 VSS VDD sky130_fd_sc_hd__nor2_1_236/B sky130_fd_sc_hd__o21a_1_55/A1
+ sky130_fd_sc_hd__a21oi_1_413/Y sky130_fd_sc_hd__o21ai_1_431/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_442 VSS VDD sky130_fd_sc_hd__nand2_1_526/B sky130_fd_sc_hd__nor2_1_296/Y
+ sky130_fd_sc_hd__nor2_1_295/B sky130_fd_sc_hd__o21ai_1_442/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_453 VSS VDD sky130_fd_sc_hd__nor2_1_301/B sky130_fd_sc_hd__nor2_1_309/A
+ sky130_fd_sc_hd__nand2_1_529/Y sky130_fd_sc_hd__xor2_1_303/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_464 VSS VDD sky130_fd_sc_hd__nor2_1_307/A sky130_fd_sc_hd__a21oi_1_458/Y
+ sky130_fd_sc_hd__a211oi_1_33/Y sky130_fd_sc_hd__xor2_1_315/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_475 VSS VDD sky130_fd_sc_hd__a222oi_1_40/Y sky130_fd_sc_hd__nor2_1_307/A
+ sky130_fd_sc_hd__a21oi_1_461/Y sky130_fd_sc_hd__xor2_1_284/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_486 VSS VDD sky130_fd_sc_hd__nor2_1_307/A sky130_fd_sc_hd__a21oi_1_476/Y
+ sky130_fd_sc_hd__a211oi_1_36/Y sky130_fd_sc_hd__xor2_1_294/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_497 VSS VDD sky130_fd_sc_hd__nand2_1_558/A sky130_fd_sc_hd__o21ai_1_507/A1
+ sky130_fd_sc_hd__nand2_1_558/Y sky130_fd_sc_hd__and2_0_342/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_1207 sky130_fd_sc_hd__fa_2_1208/CIN sky130_fd_sc_hd__mux2_2_128/A0
+ sky130_fd_sc_hd__fa_2_1207/A sky130_fd_sc_hd__fa_2_1207/B sky130_fd_sc_hd__fa_2_1207/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1218 sky130_fd_sc_hd__fa_2_1219/CIN sky130_fd_sc_hd__mux2_2_154/A1
+ sky130_fd_sc_hd__fa_2_1218/A sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__fa_2_1218/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1229 sky130_fd_sc_hd__fa_2_1230/CIN sky130_fd_sc_hd__mux2_2_204/A1
+ sky130_fd_sc_hd__fa_2_1229/A sky130_fd_sc_hd__fa_2_1229/B sky130_fd_sc_hd__fa_2_1229/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1004 VDD VSS sky130_fd_sc_hd__mux2_2_110/A0 sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__o22ai_1_235/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_13 VSS VDD sky130_fd_sc_hd__nor2b_1_53/Y sky130_fd_sc_hd__nand2_1_36/A
+ sky130_fd_sc_hd__nor2b_1_52/A sky130_fd_sc_hd__o21ai_1_13/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1015 VDD VSS sky130_fd_sc_hd__mux2_2_82/A1 sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__o22ai_1_224/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_24 VSS VDD sky130_fd_sc_hd__a21oi_2_0/Y sky130_fd_sc_hd__o21ai_1_29/B1
+ sky130_fd_sc_hd__nand2_1_43/Y sky130_fd_sc_hd__o21ai_1_24/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1026 VDD VSS sky130_fd_sc_hd__fa_2_843/A sky130_fd_sc_hd__dfxtp_1_1026/CLK
+ sky130_fd_sc_hd__a21oi_1_312/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_35 VSS VDD sky130_fd_sc_hd__o21ai_1_35/A2 sky130_fd_sc_hd__o21ai_1_35/A1
+ sky130_fd_sc_hd__o21ai_1_35/B1 sky130_fd_sc_hd__o21ai_1_35/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1037 VDD VSS sky130_fd_sc_hd__fa_2_903/B sky130_fd_sc_hd__dfxtp_1_1047/CLK
+ sky130_fd_sc_hd__a21oi_1_307/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_46 VSS VDD sky130_fd_sc_hd__o21ai_1_53/A2 sky130_fd_sc_hd__xnor2_1_46/Y
+ sky130_fd_sc_hd__a21oi_1_34/Y sky130_fd_sc_hd__o21ai_1_46/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1048 VDD VSS sky130_fd_sc_hd__fa_2_914/B sky130_fd_sc_hd__dfxtp_1_1050/CLK
+ sky130_fd_sc_hd__a21oi_1_301/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_620 VDD VSS sky130_fd_sc_hd__ha_2_144/A sky130_fd_sc_hd__dfxtp_1_626/CLK
+ sky130_fd_sc_hd__o21a_1_4/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_280 sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1291/B
+ sky130_fd_sc_hd__xor2_1_280/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o21ai_1_57 VSS VDD sky130_fd_sc_hd__nand2_2_3/Y sky130_fd_sc_hd__xnor2_1_34/Y
+ sky130_fd_sc_hd__a21oi_1_43/Y sky130_fd_sc_hd__o21ai_1_57/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1059 VDD VSS sky130_fd_sc_hd__fa_2_1198/A sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__mux2_2_149/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_291 sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1280/B
+ sky130_fd_sc_hd__xor2_1_291/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_631 VDD VSS sky130_fd_sc_hd__fa_2_995/A sky130_fd_sc_hd__clkinv_8_41/Y
+ sky130_fd_sc_hd__and2_0_283/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_68 VSS VDD sky130_fd_sc_hd__nand2_2_3/Y sky130_fd_sc_hd__xnor2_1_56/Y
+ sky130_fd_sc_hd__a21oi_1_54/Y sky130_fd_sc_hd__o21ai_1_68/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_642 VDD VSS sky130_fd_sc_hd__fa_2_1006/A sky130_fd_sc_hd__clkinv_8_44/Y
+ sky130_fd_sc_hd__mux2_2_20/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_79 VSS VDD sky130_fd_sc_hd__xnor2_1_40/A sky130_fd_sc_hd__o21ai_1_79/A1
+ sky130_fd_sc_hd__o21ai_1_79/B1 sky130_fd_sc_hd__xnor2_1_42/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_653 VDD VSS sky130_fd_sc_hd__fa_2_970/B sky130_fd_sc_hd__clkinv_8_41/Y
+ sky130_fd_sc_hd__and2_0_276/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_664 VDD VSS sky130_fd_sc_hd__fa_2_981/A sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__mux2_2_25/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_675 VDD VSS sky130_fd_sc_hd__fa_2_992/A sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__mux2_2_3/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_686 VDD VSS sky130_fd_sc_hd__fa_2_1025/A sky130_fd_sc_hd__clkinv_8_54/Y
+ sky130_fd_sc_hd__and2_0_285/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_697 VDD VSS sky130_fd_sc_hd__nand2_1_282/B sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__nor2b_1_96/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_240 VSS VDD sky130_fd_sc_hd__buf_4_47/A sky130_fd_sc_hd__buf_8_78/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_251 VSS VDD sky130_fd_sc_hd__clkbuf_1_251/X sky130_fd_sc_hd__clkbuf_1_251/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_262 VSS VDD sky130_fd_sc_hd__nand2_2_0/A sky130_fd_sc_hd__buf_6_86/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_273 VSS VDD sky130_fd_sc_hd__clkbuf_1_273/X sky130_fd_sc_hd__clkbuf_1_273/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_284 VSS VDD sky130_fd_sc_hd__clkbuf_1_284/X sky130_fd_sc_hd__clkbuf_1_284/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_295 VSS VDD sky130_fd_sc_hd__clkbuf_1_295/X sky130_fd_sc_hd__clkbuf_1_295/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_503 sky130_fd_sc_hd__fa_2_505/CIN sky130_fd_sc_hd__fa_2_498/A
+ sky130_fd_sc_hd__fa_2_503/A sky130_fd_sc_hd__fa_2_503/B sky130_fd_sc_hd__fa_2_510/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_514 sky130_fd_sc_hd__fa_2_519/B sky130_fd_sc_hd__fa_2_514/SUM
+ sky130_fd_sc_hd__fa_2_514/A sky130_fd_sc_hd__fa_2_514/B sky130_fd_sc_hd__fa_2_514/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_525 sky130_fd_sc_hd__fa_2_529/B sky130_fd_sc_hd__fa_2_525/SUM
+ sky130_fd_sc_hd__fa_2_525/A sky130_fd_sc_hd__fa_2_525/B sky130_fd_sc_hd__fa_2_525/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_536 sky130_fd_sc_hd__fa_2_537/CIN sky130_fd_sc_hd__fa_2_530/A
+ sky130_fd_sc_hd__ha_2_123/B sky130_fd_sc_hd__fa_2_546/B sky130_fd_sc_hd__fa_2_564/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_547 sky130_fd_sc_hd__fa_2_549/B sky130_fd_sc_hd__fa_2_544/A
+ sky130_fd_sc_hd__fa_2_555/A sky130_fd_sc_hd__fa_2_547/B sky130_fd_sc_hd__ha_2_125/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_558 sky130_fd_sc_hd__fa_2_557/A sky130_fd_sc_hd__fa_2_553/A
+ sky130_fd_sc_hd__fa_2_566/A sky130_fd_sc_hd__fa_2_558/B sky130_fd_sc_hd__fa_2_564/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_569 sky130_fd_sc_hd__fa_2_568/CIN sky130_fd_sc_hd__and2_0_87/A
+ sky130_fd_sc_hd__fa_2_569/A sky130_fd_sc_hd__fa_2_569/B sky130_fd_sc_hd__fa_2_569/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_4_1 VDD VSS sky130_fd_sc_hd__buf_4_1/X sky130_fd_sc_hd__buf_4_1/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__and2_0_260 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_260/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__fa_2_961/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_271 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_271/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__and2_0_271/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_282 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_282/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__fa_2_972/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_293 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_293/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__fa_2_998/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_508 sky130_fd_sc_hd__buf_12_508/A sky130_fd_sc_hd__buf_12_518/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_519 sky130_fd_sc_hd__bufbuf_8_9/X sky130_fd_sc_hd__buf_12_519/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__inv_4_1 sky130_fd_sc_hd__inv_4_1/Y sky130_fd_sc_hd__inv_4_1/A VDD
+ VSS VDD VSS sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__nand2_1_109 sky130_fd_sc_hd__nand2_1_109/Y sky130_fd_sc_hd__buf_2_271/X
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_708 sky130_fd_sc_hd__o22ai_1_184/B1 sky130_fd_sc_hd__fa_2_1062/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_708/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_719 sky130_fd_sc_hd__nor2_1_117/B sky130_fd_sc_hd__fa_2_1057/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_719/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_250 VSS VDD sky130_fd_sc_hd__o21a_1_16/X sky130_fd_sc_hd__nor2_1_126/A
+ sky130_fd_sc_hd__nand2b_1_16/Y sky130_fd_sc_hd__o21ai_1_250/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_261 VSS VDD sky130_fd_sc_hd__o21a_1_16/A2 sky130_fd_sc_hd__o21ai_1_261/A1
+ sky130_fd_sc_hd__a22oi_1_361/Y sky130_fd_sc_hd__o21ai_1_261/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_272 VSS VDD sky130_fd_sc_hd__nor2_1_126/A sky130_fd_sc_hd__a21oi_1_240/Y
+ sky130_fd_sc_hd__a21oi_1_236/Y sky130_fd_sc_hd__xor2_1_111/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_90 sky130_fd_sc_hd__nand4_1_25/A sky130_fd_sc_hd__clkbuf_4_90/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_283 VSS VDD sky130_fd_sc_hd__o22ai_1_235/A1 sky130_fd_sc_hd__nor2_1_162/Y
+ sky130_fd_sc_hd__or3_1_2/X sky130_fd_sc_hd__o21ai_1_283/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_294 VSS VDD sky130_fd_sc_hd__o22ai_1_247/A1 sky130_fd_sc_hd__o21a_1_29/A1
+ sky130_fd_sc_hd__a21oi_1_266/Y sky130_fd_sc_hd__o21ai_1_294/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor3_1_19 sky130_fd_sc_hd__nor3_2_8/C sky130_fd_sc_hd__nor3_1_19/Y
+ sky130_fd_sc_hd__nor3_2_9/B sky130_fd_sc_hd__nor3_2_9/C VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor2b_2_1 sky130_fd_sc_hd__ha_2_43/SUM sky130_fd_sc_hd__or2_1_0/B
+ sky130_fd_sc_hd__nor2b_2_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_2
Xsky130_fd_sc_hd__fa_2_1004 sky130_fd_sc_hd__fa_2_1005/CIN sky130_fd_sc_hd__mux2_2_24/A0
+ sky130_fd_sc_hd__fa_2_1004/A sky130_fd_sc_hd__xor2_1_72/X sky130_fd_sc_hd__fa_2_1004/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1015 sky130_fd_sc_hd__xor2_1_58/B sky130_fd_sc_hd__mux2_2_1/A0
+ sky130_fd_sc_hd__fa_2_1015/A sky130_fd_sc_hd__xor2_1_61/X sky130_fd_sc_hd__fa_2_1015/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1026 sky130_fd_sc_hd__fa_2_1027/CIN sky130_fd_sc_hd__and2_0_290/A
+ sky130_fd_sc_hd__fa_2_1026/A sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_1026/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1037 sky130_fd_sc_hd__fa_2_1038/CIN sky130_fd_sc_hd__fa_2_1037/SUM
+ sky130_fd_sc_hd__fa_2_1037/A sky130_fd_sc_hd__nor2_1_52/A sky130_fd_sc_hd__fa_2_1037/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1048 sky130_fd_sc_hd__fa_2_1049/CIN sky130_fd_sc_hd__and2_0_307/A
+ sky130_fd_sc_hd__fa_2_1048/A sky130_fd_sc_hd__fa_2_1048/B sky130_fd_sc_hd__fa_2_1048/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1059 sky130_fd_sc_hd__fa_2_1060/CIN sky130_fd_sc_hd__mux2_2_59/A0
+ sky130_fd_sc_hd__fa_2_1059/A sky130_fd_sc_hd__xor2_1_98/X sky130_fd_sc_hd__fa_2_1059/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_13 sky130_fd_sc_hd__inv_2_13/A sky130_fd_sc_hd__inv_2_13/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_24 sky130_fd_sc_hd__inv_2_24/A sky130_fd_sc_hd__inv_2_24/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_35 sky130_fd_sc_hd__inv_2_35/A sky130_fd_sc_hd__inv_2_35/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_46 sky130_fd_sc_hd__inv_2_46/A sky130_fd_sc_hd__inv_2_46/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_450 VDD VSS sky130_fd_sc_hd__dfxtp_1_996/D sky130_fd_sc_hd__dfxtp_1_454/CLK
+ sky130_fd_sc_hd__nand2_1_64/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_57 sky130_fd_sc_hd__inv_2_57/A sky130_fd_sc_hd__inv_2_57/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_461 VDD VSS sky130_fd_sc_hd__buf_2_9/A sky130_fd_sc_hd__dfxtp_1_463/CLK
+ sky130_fd_sc_hd__and2_0_237/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_68 sky130_fd_sc_hd__inv_2_68/A sky130_fd_sc_hd__inv_2_68/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_472 VDD VSS sky130_fd_sc_hd__clkbuf_1_2/A sky130_fd_sc_hd__dfxtp_1_472/CLK
+ sky130_fd_sc_hd__and2_0_111/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_79 sky130_fd_sc_hd__inv_2_79/A sky130_fd_sc_hd__inv_2_81/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_483 VDD VSS sky130_fd_sc_hd__dfxtp_1_483/Q sky130_fd_sc_hd__dfxtp_1_483/CLK
+ sky130_fd_sc_hd__nor2b_1_75/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_2_3 sky130_fd_sc_hd__nand2_2_3/Y sky130_fd_sc_hd__nor2_2_6/A
+ sky130_fd_sc_hd__nor2_1_41/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__dfxtp_1_494 VDD VSS sky130_fd_sc_hd__dfxtp_1_494/Q sky130_fd_sc_hd__dfxtp_1_502/CLK
+ sky130_fd_sc_hd__nor2b_1_57/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_300 sky130_fd_sc_hd__fa_2_293/CIN sky130_fd_sc_hd__fa_2_300/SUM
+ sky130_fd_sc_hd__fa_2_300/A sky130_fd_sc_hd__fa_2_300/B sky130_fd_sc_hd__fa_2_300/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_311 sky130_fd_sc_hd__fa_2_307/CIN sky130_fd_sc_hd__fa_2_313/A
+ sky130_fd_sc_hd__ha_2_116/A sky130_fd_sc_hd__ha_2_112/B sky130_fd_sc_hd__fa_2_409/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_322 sky130_fd_sc_hd__fa_2_318/CIN sky130_fd_sc_hd__or3_1_3/B
+ sky130_fd_sc_hd__fa_2_322/A sky130_fd_sc_hd__fa_2_322/B sky130_fd_sc_hd__maj3_1_56/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_333 sky130_fd_sc_hd__fa_2_335/CIN sky130_fd_sc_hd__fa_2_331/B
+ sky130_fd_sc_hd__ha_2_115/B sky130_fd_sc_hd__fa_2_393/A sky130_fd_sc_hd__fa_2_417/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_344 sky130_fd_sc_hd__fa_2_347/A sky130_fd_sc_hd__fa_2_344/SUM
+ sky130_fd_sc_hd__fa_2_344/A sky130_fd_sc_hd__fa_2_344/B sky130_fd_sc_hd__fa_2_344/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_355 sky130_fd_sc_hd__fa_2_357/CIN sky130_fd_sc_hd__fa_2_352/A
+ sky130_fd_sc_hd__fa_2_355/A sky130_fd_sc_hd__fa_2_355/B sky130_fd_sc_hd__fa_2_355/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_366 sky130_fd_sc_hd__maj3_1_66/B sky130_fd_sc_hd__maj3_1_67/A
+ sky130_fd_sc_hd__fa_2_366/A sky130_fd_sc_hd__fa_2_366/B sky130_fd_sc_hd__fa_2_367/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_377 sky130_fd_sc_hd__maj3_1_64/B sky130_fd_sc_hd__maj3_1_65/A
+ sky130_fd_sc_hd__fa_2_377/A sky130_fd_sc_hd__fa_2_377/B sky130_fd_sc_hd__fa_2_378/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_18 sky130_fd_sc_hd__conb_1_11/LO sky130_fd_sc_hd__clkinv_8_131/A
+ sky130_fd_sc_hd__clkinv_4_10/A sky130_fd_sc_hd__or2_1_0/X VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_388 sky130_fd_sc_hd__fa_2_391/B sky130_fd_sc_hd__fa_2_388/SUM
+ sky130_fd_sc_hd__fa_2_388/A sky130_fd_sc_hd__fa_2_388/B sky130_fd_sc_hd__fa_2_388/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_29 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_61/Y
+ sky130_fd_sc_hd__dfxtp_1_262/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__and2_1_4 VDD VSS sky130_fd_sc_hd__and2_1_4/X sky130_fd_sc_hd__ha_2_55/A
+ sky130_fd_sc_hd__nor2_4_2/Y VDD VSS sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__fa_2_399 sky130_fd_sc_hd__fa_2_401/CIN sky130_fd_sc_hd__fa_2_392/B
+ sky130_fd_sc_hd__ha_2_108/B sky130_fd_sc_hd__ha_2_110/B sky130_fd_sc_hd__fa_2_286/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__diode_2_205 sky130_fd_sc_hd__buf_2_282/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_216 amplitude_adc_done VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_227 sig_amplitude[0] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkinv_8_60 sky130_fd_sc_hd__clkinv_8_62/A sky130_fd_sc_hd__clkinv_8_94/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_60/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_71 sky130_fd_sc_hd__clkinv_8_72/A sky130_fd_sc_hd__clkinv_8_71/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_82 sky130_fd_sc_hd__clkinv_8_83/A sky130_fd_sc_hd__clkinv_8_82/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_82/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_93 sky130_fd_sc_hd__clkinv_8_94/A sky130_fd_sc_hd__clkinv_8_93/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_80 sky130_fd_sc_hd__buf_6_12/X sky130_fd_sc_hd__buf_12_80/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_91 sky130_fd_sc_hd__buf_12_91/A sky130_fd_sc_hd__buf_12_91/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__dfxtp_1_1390 VDD VSS sky130_fd_sc_hd__nor2_4_19/B sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__nor2b_1_128/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nor2_1_109 sky130_fd_sc_hd__nor2_1_109/B sky130_fd_sc_hd__nor2_1_109/Y
+ sky130_fd_sc_hd__fa_2_1114/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_18 sky130_fd_sc_hd__nor2_2_0/Y sky130_fd_sc_hd__clkinv_1_4/Y
+ sky130_fd_sc_hd__nand4_1_22/Y sky130_fd_sc_hd__nand4_1_6/Y sky130_fd_sc_hd__a22oi_1_18/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_29 sky130_fd_sc_hd__a22oi_1_81/B1 sky130_fd_sc_hd__clkbuf_1_99/X
+ sky130_fd_sc_hd__clkbuf_1_50/X sky130_fd_sc_hd__clkbuf_4_25/X sky130_fd_sc_hd__nand4_1_0/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_305 sky130_fd_sc_hd__buf_8_130/X sky130_fd_sc_hd__buf_12_305/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_316 sky130_fd_sc_hd__buf_4_82/X sky130_fd_sc_hd__buf_12_316/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_327 sky130_fd_sc_hd__buf_4_81/X sky130_fd_sc_hd__buf_12_327/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_338 sky130_fd_sc_hd__buf_6_35/X sky130_fd_sc_hd__buf_12_338/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_349 sky130_fd_sc_hd__buf_6_46/X sky130_fd_sc_hd__buf_12_349/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_208 sky130_fd_sc_hd__clkbuf_1_351/X sky130_fd_sc_hd__clkbuf_1_353/X
+ sky130_fd_sc_hd__clkbuf_4_113/X sky130_fd_sc_hd__a22oi_1_208/A2 sky130_fd_sc_hd__nand4_1_47/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_219 sky130_fd_sc_hd__buf_2_166/X sky130_fd_sc_hd__buf_2_167/X
+ sky130_fd_sc_hd__clkbuf_1_435/X sky130_fd_sc_hd__buf_2_180/X sky130_fd_sc_hd__nand4_1_51/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor3_2_0 sky130_fd_sc_hd__nor4_1_0/B sky130_fd_sc_hd__nor3_2_0/Y
+ sky130_fd_sc_hd__nor3_2_0/A sky130_fd_sc_hd__nor4_1_0/A VDD VSS VSS VDD sky130_fd_sc_hd__nor3_2
Xsky130_fd_sc_hd__clkinv_1_505 sky130_fd_sc_hd__o21ai_1_78/A1 sky130_fd_sc_hd__o21ai_1_85/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_505/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_516 sky130_fd_sc_hd__nor2_1_54/B sky130_fd_sc_hd__fa_2_1033/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_516/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_527 sky130_fd_sc_hd__nor2_1_62/B sky130_fd_sc_hd__fa_2_1044/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_527/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_538 sky130_fd_sc_hd__o211ai_1_6/A1 sky130_fd_sc_hd__fa_2_990/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_538/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_549 sky130_fd_sc_hd__nor2_1_69/B sky130_fd_sc_hd__fa_2_978/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_549/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_30 sky130_fd_sc_hd__nor2_1_30/B sky130_fd_sc_hd__nor2_1_30/Y
+ sky130_fd_sc_hd__nor4_1_7/C VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_41 sky130_fd_sc_hd__nor2_1_41/B sky130_fd_sc_hd__nor2_1_41/Y
+ sky130_fd_sc_hd__nor2_2_6/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_52 sky130_fd_sc_hd__nor2_1_52/B sky130_fd_sc_hd__nor2_1_52/Y
+ sky130_fd_sc_hd__nor2_1_52/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_63 sky130_fd_sc_hd__nor2_1_63/B sky130_fd_sc_hd__o21a_1_1/A1
+ sky130_fd_sc_hd__o21a_1_2/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_18 sky130_fd_sc_hd__clkinv_8_33/Y sky130_fd_sc_hd__clkinv_8_34/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_18/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_74 sky130_fd_sc_hd__nor2_1_85/Y sky130_fd_sc_hd__nor2_1_74/Y
+ sky130_fd_sc_hd__nor2_1_74/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_29 sky130_fd_sc_hd__clkinv_4_29/A sky130_fd_sc_hd__clkinv_8_76/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_29/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_85 sky130_fd_sc_hd__nor2_1_85/B sky130_fd_sc_hd__nor2_1_85/Y
+ sky130_fd_sc_hd__nor2_1_85/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_96 sky130_fd_sc_hd__nor2_1_96/B sky130_fd_sc_hd__nor2_1_96/Y
+ sky130_fd_sc_hd__nor2_1_96/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_sram_2kbyte_1rw1r_32x512_8_4 sky130_fd_sc_hd__buf_6_19/X sky130_fd_sc_hd__buf_4_33/X
+ sky130_fd_sc_hd__clkbuf_4_60/X sky130_fd_sc_hd__buf_12_121/X sky130_fd_sc_hd__clkbuf_4_61/X
+ sky130_fd_sc_hd__clkbuf_4_64/X sky130_fd_sc_hd__buf_4_35/X sky130_fd_sc_hd__buf_12_122/X
+ sky130_fd_sc_hd__buf_4_37/X sky130_fd_sc_hd__buf_4_38/X sky130_fd_sc_hd__buf_4_39/X
+ sky130_fd_sc_hd__clkbuf_8_0/X sky130_fd_sc_hd__buf_4_40/X sky130_fd_sc_hd__clkbuf_4_67/X
+ sky130_fd_sc_hd__clkbuf_4_69/X sky130_fd_sc_hd__clkbuf_4_71/X sky130_fd_sc_hd__buf_6_19/X
+ sky130_fd_sc_hd__buf_4_33/X sky130_fd_sc_hd__clkbuf_4_60/X sky130_fd_sc_hd__buf_12_121/X
+ sky130_fd_sc_hd__clkbuf_4_61/X sky130_fd_sc_hd__clkbuf_4_64/X sky130_fd_sc_hd__buf_4_35/X
+ sky130_fd_sc_hd__buf_12_122/X sky130_fd_sc_hd__buf_4_37/X sky130_fd_sc_hd__buf_4_38/X
+ sky130_fd_sc_hd__buf_4_39/X sky130_fd_sc_hd__clkbuf_8_0/X sky130_fd_sc_hd__buf_4_40/X
+ sky130_fd_sc_hd__clkbuf_4_67/X sky130_fd_sc_hd__clkbuf_4_69/X sky130_fd_sc_hd__clkbuf_4_71/X
+ sky130_fd_sc_hd__buf_12_234/X sky130_fd_sc_hd__buf_12_200/X sky130_fd_sc_hd__buf_12_231/X
+ sky130_fd_sc_hd__buf_12_230/X sky130_fd_sc_hd__buf_12_213/X sky130_fd_sc_hd__buf_12_229/X
+ sky130_fd_sc_hd__buf_12_212/X sky130_fd_sc_hd__buf_12_259/X sky130_fd_sc_hd__buf_12_260/X
+ sky130_fd_sc_hd__buf_12_257/X sky130_fd_sc_hd__buf_12_236/X sky130_fd_sc_hd__buf_12_211/X
+ sky130_fd_sc_hd__buf_12_216/X sky130_fd_sc_hd__buf_12_235/X sky130_fd_sc_hd__buf_12_223/X
+ sky130_fd_sc_hd__buf_12_249/X sky130_fd_sc_hd__buf_12_177/X sky130_fd_sc_hd__buf_12_126/X
+ sky130_fd_sc_hd__buf_2_99/X sky130_fd_sc_hd__clkbuf_1_242/X sky130_fd_sc_hd__buf_2_99/X
+ sky130_fd_sc_hd__clkinv_8_132/Y sky130_fd_sc_hd__clkinv_8_12/Y sky130_fd_sc_hd__buf_12_189/X
+ sky130_fd_sc_hd__buf_12_183/X sky130_fd_sc_hd__buf_12_157/X sky130_fd_sc_hd__buf_12_158/X
+ sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[0] sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[1]
+ sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[2] sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[3]
+ sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[4] sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[5]
+ sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[6] sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[7]
+ sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[8] sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[9]
+ sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[10] sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[11]
+ sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[12] sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[13]
+ sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[14] sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[15]
+ sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[16] sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[17]
+ sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[18] sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[19]
+ sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[20] sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[21]
+ sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[22] sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[23]
+ sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[24] sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[25]
+ sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[26] sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[27]
+ sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[28] sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[29]
+ sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[30] sky130_sram_2kbyte_1rw1r_32x512_8_4/dout0[31]
+ sky130_fd_sc_hd__buf_2_66/A sky130_fd_sc_hd__buf_2_67/A sky130_fd_sc_hd__buf_2_68/A
+ sky130_fd_sc_hd__clkbuf_1_254/A sky130_fd_sc_hd__buf_2_70/A sky130_fd_sc_hd__buf_2_71/A
+ sky130_fd_sc_hd__buf_2_72/A sky130_fd_sc_hd__buf_2_73/A sky130_fd_sc_hd__buf_2_74/A
+ sky130_fd_sc_hd__buf_2_75/A sky130_fd_sc_hd__buf_2_76/A sky130_fd_sc_hd__buf_2_77/A
+ sky130_fd_sc_hd__buf_2_78/A sky130_fd_sc_hd__buf_2_79/A sky130_fd_sc_hd__buf_2_80/A
+ sky130_fd_sc_hd__buf_2_81/A sky130_fd_sc_hd__buf_2_82/A sky130_fd_sc_hd__buf_2_83/A
+ sky130_fd_sc_hd__buf_2_84/A sky130_fd_sc_hd__buf_2_85/A sky130_fd_sc_hd__buf_2_86/A
+ sky130_fd_sc_hd__buf_2_87/A sky130_fd_sc_hd__buf_2_88/A sky130_fd_sc_hd__buf_2_89/A
+ sky130_fd_sc_hd__buf_2_90/A sky130_fd_sc_hd__buf_2_91/A sky130_fd_sc_hd__buf_2_92/A
+ sky130_fd_sc_hd__buf_2_93/A sky130_fd_sc_hd__buf_2_94/A sky130_fd_sc_hd__buf_2_95/A
+ sky130_fd_sc_hd__buf_2_96/A sky130_fd_sc_hd__buf_2_97/A VDD VSS sky130_sram_2kbyte_1rw1r_32x512_8
Xsky130_fd_sc_hd__a21oi_1_402 sky130_fd_sc_hd__nor2b_2_4/Y sky130_fd_sc_hd__o21ai_1_423/Y
+ sky130_fd_sc_hd__a21oi_1_402/Y sky130_fd_sc_hd__o21ai_1_436/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_413 sky130_fd_sc_hd__fa_2_1256/A sky130_fd_sc_hd__o22ai_1_371/Y
+ sky130_fd_sc_hd__a21oi_1_413/Y sky130_fd_sc_hd__nor3_1_40/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_424 sky130_fd_sc_hd__o21a_1_60/B1 sky130_fd_sc_hd__o21a_1_59/A1
+ sky130_fd_sc_hd__a21oi_1_424/Y sky130_fd_sc_hd__nor2_1_272/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_435 sky130_fd_sc_hd__nor2_1_283/A sky130_fd_sc_hd__o21a_1_67/A1
+ sky130_fd_sc_hd__a21oi_1_435/Y sky130_fd_sc_hd__nor2_1_283/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_446 sky130_fd_sc_hd__fa_2_1283/A sky130_fd_sc_hd__o22ai_1_413/Y
+ sky130_fd_sc_hd__a21oi_1_446/Y sky130_fd_sc_hd__nor3_1_41/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_457 sky130_fd_sc_hd__fa_2_1286/A sky130_fd_sc_hd__o22ai_1_418/Y
+ sky130_fd_sc_hd__a21oi_1_457/Y sky130_fd_sc_hd__nor2_2_18/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_468 sky130_fd_sc_hd__nor2_1_309/Y sky130_fd_sc_hd__nor2_1_304/Y
+ sky130_fd_sc_hd__a21oi_1_468/Y sky130_fd_sc_hd__fa_2_1301/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_479 sky130_fd_sc_hd__fa_2_1303/A sky130_fd_sc_hd__o22ai_1_436/Y
+ sky130_fd_sc_hd__o21a_1_68/B1 sky130_fd_sc_hd__nor2_2_18/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_8_104 sky130_fd_sc_hd__clkinv_8_67/A sky130_fd_sc_hd__clkinv_8_104/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_104/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_115 sky130_fd_sc_hd__clkinv_8_71/A sky130_fd_sc_hd__clkinv_8_115/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_115/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_126 sky130_fd_sc_hd__clkinv_8_127/A sky130_fd_sc_hd__clkinv_4_64/Y
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_137 sky130_fd_sc_hd__clkinv_8_18/A sky130_fd_sc_hd__clkinv_8_137/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__o21a_1_6 sky130_fd_sc_hd__o21a_1_6/X sky130_fd_sc_hd__o21a_1_6/A1
+ sky130_fd_sc_hd__o21a_1_6/B1 sky130_fd_sc_hd__fa_2_979/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__maj3_1_160 sky130_fd_sc_hd__maj3_1_161/X sky130_fd_sc_hd__maj3_1_160/X
+ sky130_fd_sc_hd__maj3_1_160/B sky130_fd_sc_hd__maj3_1_160/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_440 sky130_fd_sc_hd__nand2_1_440/Y sky130_fd_sc_hd__nor2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_377/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_451 sky130_fd_sc_hd__o21a_1_48/B1 sky130_fd_sc_hd__fa_2_1229/A
+ sky130_fd_sc_hd__o21a_1_48/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_462 sky130_fd_sc_hd__nand2_1_462/Y sky130_fd_sc_hd__nor2_1_246/B
+ sky130_fd_sc_hd__xnor2_1_99/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_473 sky130_fd_sc_hd__nor2_1_252/B sky130_fd_sc_hd__nand2_1_473/B
+ sky130_fd_sc_hd__nor2_1_253/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_484 sky130_fd_sc_hd__nand2_1_484/Y sky130_fd_sc_hd__fa_2_1241/A
+ sky130_fd_sc_hd__nor3_1_40/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_495 sky130_fd_sc_hd__nor2_1_268/A sky130_fd_sc_hd__nor2b_2_4/A
+ sky130_fd_sc_hd__o32ai_1_8/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_20 sky130_fd_sc_hd__ha_2_42/SUM sky130_fd_sc_hd__nor2b_1_20/Y
+ sky130_fd_sc_hd__or2_1_0/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_31 sky130_fd_sc_hd__ha_2_65/SUM sky130_fd_sc_hd__nor2b_1_31/Y
+ sky130_fd_sc_hd__or2_0_2/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_42 sky130_fd_sc_hd__ha_2_89/SUM sky130_fd_sc_hd__nor2b_1_42/Y
+ sky130_fd_sc_hd__or2_0_3/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_53 sky130_fd_sc_hd__nor4_1_4/A sky130_fd_sc_hd__nor2b_1_53/Y
+ sky130_fd_sc_hd__o31ai_1_1/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1020 sky130_fd_sc_hd__nor2_1_239/B sky130_fd_sc_hd__fa_2_1249/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1020/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_64 sky130_fd_sc_hd__o21ai_1_36/A1 sky130_fd_sc_hd__nor2b_1_64/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1031 sky130_fd_sc_hd__a22oi_1_400/B1 sky130_fd_sc_hd__o21a_1_68/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1031/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_75 sky130_fd_sc_hd__nor2b_1_88/A sky130_fd_sc_hd__nor2b_1_75/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1042 sky130_fd_sc_hd__nor2_1_275/A sky130_fd_sc_hd__nor2_1_276/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1042/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_86 sky130_fd_sc_hd__fa_2_951/A sky130_fd_sc_hd__nor2b_1_86/Y
+ sky130_fd_sc_hd__nor2b_1_86/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1053 sky130_fd_sc_hd__o22ai_1_401/A1 sky130_fd_sc_hd__fa_2_8/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1053/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1064 sky130_fd_sc_hd__o31ai_1_12/A3 sky130_fd_sc_hd__xnor2_1_0/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1064/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_97 sky130_fd_sc_hd__buf_2_263/A sky130_fd_sc_hd__nor2b_1_97/Y
+ sky130_fd_sc_hd__a32o_1_1/A3 VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__xnor2_1_5 VSS VDD sky130_fd_sc_hd__xnor2_1_5/B sky130_fd_sc_hd__xnor2_1_5/Y
+ sky130_fd_sc_hd__fa_2_833/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_1075 sky130_fd_sc_hd__a21oi_1_452/A2 sky130_fd_sc_hd__nor2_1_299/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1075/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1086 sky130_fd_sc_hd__o22ai_1_423/B1 sky130_fd_sc_hd__fa_2_1287/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1086/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1097 sky130_fd_sc_hd__nor2_1_284/B sky130_fd_sc_hd__fa_2_1296/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1097/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_280 VDD VSS sky130_fd_sc_hd__buf_2_263/A sky130_fd_sc_hd__dfxtp_1_282/CLK
+ sky130_fd_sc_hd__or2_0_4/B VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_291 VDD VSS sky130_fd_sc_hd__a22o_1_56/A1 sky130_fd_sc_hd__clkinv_4_31/Y
+ sky130_fd_sc_hd__nand2_1_127/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o22ai_1_0 sky130_fd_sc_hd__o22ai_1_0/A2 sky130_fd_sc_hd__xnor2_1_19/Y
+ sky130_fd_sc_hd__o22ai_1_0/Y sky130_fd_sc_hd__xnor2_1_12/B sky130_fd_sc_hd__o22ai_1_0/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_130 sky130_fd_sc_hd__fa_2_129/B sky130_fd_sc_hd__fa_2_130/SUM
+ sky130_fd_sc_hd__fa_2_130/A sky130_fd_sc_hd__fa_2_130/B sky130_fd_sc_hd__fa_2_135/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_141 sky130_fd_sc_hd__fa_2_25/B sky130_fd_sc_hd__fa_2_141/SUM
+ sky130_fd_sc_hd__fa_2_49/B sky130_fd_sc_hd__fa_2_141/B sky130_fd_sc_hd__fa_2_141/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_152 sky130_fd_sc_hd__fa_2_143/A sky130_fd_sc_hd__fa_2_150/B
+ sky130_fd_sc_hd__fa_2_280/A sky130_fd_sc_hd__fa_2_152/B sky130_fd_sc_hd__fa_2_155/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_163 sky130_fd_sc_hd__fa_2_160/B sky130_fd_sc_hd__fa_2_162/B
+ sky130_fd_sc_hd__fa_2_15/B sky130_fd_sc_hd__fa_2_31/A sky130_fd_sc_hd__fa_2_281/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_174 sky130_fd_sc_hd__fa_2_175/CIN sky130_fd_sc_hd__maj3_1_54/A
+ sky130_fd_sc_hd__fa_2_32/A sky130_fd_sc_hd__ha_2_99/A sky130_fd_sc_hd__fa_2_31/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_185 sky130_fd_sc_hd__fa_2_187/CIN sky130_fd_sc_hd__fa_2_183/A
+ sky130_fd_sc_hd__fa_2_15/B sky130_fd_sc_hd__ha_2_104/B sky130_fd_sc_hd__fa_2_273/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_196 sky130_fd_sc_hd__maj3_1_44/B sky130_fd_sc_hd__maj3_1_45/A
+ sky130_fd_sc_hd__fa_2_196/A sky130_fd_sc_hd__fa_2_196/B sky130_fd_sc_hd__fa_2_197/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o22ai_1_40 sky130_fd_sc_hd__fa_2_531/B sky130_fd_sc_hd__fa_2_558/B
+ sky130_fd_sc_hd__fa_2_561/A sky130_fd_sc_hd__ha_2_119/A sky130_fd_sc_hd__ha_2_124/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_51 sky130_fd_sc_hd__fa_2_811/A sky130_fd_sc_hd__ha_2_141/B
+ sky130_fd_sc_hd__o22ai_1_51/Y sky130_fd_sc_hd__fa_2_812/B sky130_fd_sc_hd__ha_2_136/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_62 sky130_fd_sc_hd__o22ai_1_88/B1 sky130_fd_sc_hd__nand2_2_3/Y
+ sky130_fd_sc_hd__o22ai_1_62/Y sky130_fd_sc_hd__xnor2_1_35/Y sky130_fd_sc_hd__o22ai_1_76/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_180 VDD VSS sky130_fd_sc_hd__buf_2_180/X sky130_fd_sc_hd__buf_2_180/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_73 sky130_fd_sc_hd__o22ai_1_88/B1 sky130_fd_sc_hd__nand2_2_3/Y
+ sky130_fd_sc_hd__o22ai_1_73/Y sky130_fd_sc_hd__xnor2_1_57/Y sky130_fd_sc_hd__o22ai_1_87/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_191 VDD VSS sky130_fd_sc_hd__buf_2_191/X sky130_fd_sc_hd__buf_2_191/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_84 sky130_fd_sc_hd__o22ai_1_89/A1 sky130_fd_sc_hd__o22ai_1_88/B1
+ sky130_fd_sc_hd__o22ai_1_84/Y sky130_fd_sc_hd__xnor2_1_51/Y sky130_fd_sc_hd__o22ai_1_84/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_95 sky130_fd_sc_hd__nor2_2_9/B sky130_fd_sc_hd__nor2_1_77/A
+ sky130_fd_sc_hd__o22ai_1_95/Y sky130_fd_sc_hd__a21oi_1_92/Y sky130_fd_sc_hd__nor2_1_81/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_4_20 VDD VSS sky130_fd_sc_hd__buf_4_20/X sky130_fd_sc_hd__buf_8_23/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_31 VDD VSS sky130_fd_sc_hd__buf_4_31/X sky130_fd_sc_hd__buf_8_41/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_42 VDD VSS sky130_fd_sc_hd__buf_4_42/X sky130_fd_sc_hd__buf_8_84/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_53 VDD VSS sky130_fd_sc_hd__buf_4_53/X sky130_fd_sc_hd__buf_8_66/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_64 VDD VSS sky130_fd_sc_hd__buf_4_64/X sky130_fd_sc_hd__buf_4_64/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_75 VDD VSS sky130_fd_sc_hd__buf_4_75/X sky130_fd_sc_hd__buf_4_75/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_86 VDD VSS sky130_fd_sc_hd__buf_4_86/X sky130_fd_sc_hd__buf_4_86/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_97 VDD VSS sky130_fd_sc_hd__buf_4_97/X sky130_fd_sc_hd__buf_4_97/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_12_102 sky130_fd_sc_hd__buf_12_20/X sky130_fd_sc_hd__buf_12_102/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_113 sky130_fd_sc_hd__buf_12_113/A sky130_fd_sc_hd__buf_12_116/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_124 sky130_fd_sc_hd__inv_2_58/Y sky130_fd_sc_hd__buf_12_124/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_135 sky130_fd_sc_hd__buf_12_135/A sky130_fd_sc_hd__buf_12_257/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_146 sky130_fd_sc_hd__buf_8_69/X sky130_fd_sc_hd__buf_12_146/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_157 sky130_fd_sc_hd__buf_8_105/X sky130_fd_sc_hd__buf_12_157/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_80 VSS VDD sky130_fd_sc_hd__nand4_1_7/A sky130_fd_sc_hd__a22oi_2_8/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_91 VSS VDD sky130_fd_sc_hd__clkbuf_1_91/X sky130_fd_sc_hd__clkbuf_1_91/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_168 sky130_fd_sc_hd__buf_8_64/X sky130_fd_sc_hd__buf_12_227/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_4_5 sky130_fd_sc_hd__clkbuf_4_5/X sky130_fd_sc_hd__clkbuf_4_5/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_12_179 sky130_fd_sc_hd__buf_8_109/X sky130_fd_sc_hd__buf_12_220/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_1_302 sky130_fd_sc_hd__fa_2_280/B sky130_fd_sc_hd__fa_2_209/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_302/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_313 sky130_fd_sc_hd__fa_2_409/A sky130_fd_sc_hd__ha_2_110/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_313/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_324 sky130_fd_sc_hd__fa_2_554/A sky130_fd_sc_hd__ha_2_117/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_324/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_335 sky130_fd_sc_hd__fa_2_567/A sky130_fd_sc_hd__ha_2_118/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_335/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_346 sky130_fd_sc_hd__ha_2_130/A sky130_fd_sc_hd__fa_2_673/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_346/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_357 sky130_fd_sc_hd__fa_2_823/B sky130_fd_sc_hd__ha_2_144/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_357/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_368 sky130_fd_sc_hd__ha_2_141/A sky130_fd_sc_hd__ha_2_143/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_368/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_379 sky130_fd_sc_hd__fa_2_869/B sky130_fd_sc_hd__dfxtp_1_269/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_379/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_210 sky130_fd_sc_hd__fa_2_1058/A sky130_fd_sc_hd__o22ai_1_186/Y
+ sky130_fd_sc_hd__a21oi_1_210/Y sky130_fd_sc_hd__nor2_2_12/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_221 sky130_fd_sc_hd__a21o_2_5/A2 sky130_fd_sc_hd__o21ai_1_256/Y
+ sky130_fd_sc_hd__nor2_1_123/B sky130_fd_sc_hd__fa_2_1085/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_232 sky130_fd_sc_hd__a21o_2_4/X sky130_fd_sc_hd__o22ai_1_207/Y
+ sky130_fd_sc_hd__a21oi_1_232/Y sky130_fd_sc_hd__nand2_1_331/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_243 sky130_fd_sc_hd__o21a_1_20/B1 sky130_fd_sc_hd__o21a_1_19/A1
+ sky130_fd_sc_hd__dfxtp_1_903/D sky130_fd_sc_hd__nor2_1_144/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_254 sky130_fd_sc_hd__o21a_1_28/B1 sky130_fd_sc_hd__nor2_1_155/Y
+ sky130_fd_sc_hd__dfxtp_1_882/D sky130_fd_sc_hd__nor2_1_155/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_265 sky130_fd_sc_hd__o21ai_1_298/Y sky130_fd_sc_hd__nor2_1_173/Y
+ sky130_fd_sc_hd__a21oi_1_265/Y sky130_fd_sc_hd__nor2b_1_105/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_276 sky130_fd_sc_hd__nor2_2_15/Y sky130_fd_sc_hd__o21ai_1_304/Y
+ sky130_fd_sc_hd__nor2_1_174/B sky130_fd_sc_hd__fa_2_1137/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_287 sky130_fd_sc_hd__nor2b_1_104/Y sky130_fd_sc_hd__o21ai_1_319/Y
+ sky130_fd_sc_hd__a21oi_1_287/Y sky130_fd_sc_hd__o21ai_1_326/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_4_5 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_4_5/Y
+ VSS VDD VDD VSS VSS sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__a21oi_1_298 sky130_fd_sc_hd__nor3_1_38/A sky130_fd_sc_hd__o22ai_1_264/Y
+ sky130_fd_sc_hd__a21oi_1_298/Y sky130_fd_sc_hd__fa_2_1145/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_206 sky130_fd_sc_hd__inv_2_111/Y sky130_fd_sc_hd__buf_6_61/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_217 sky130_fd_sc_hd__buf_8_217/A sky130_fd_sc_hd__buf_6_69/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__o2111ai_1_0 sky130_fd_sc_hd__o21ai_1_8/Y sky130_fd_sc_hd__nand2_1_31/Y
+ sky130_fd_sc_hd__or4_1_0/D sky130_fd_sc_hd__o21ai_1_14/Y sky130_fd_sc_hd__nor4_1_1/Y
+ sky130_fd_sc_hd__a21oi_1_4/B1 VDD VSS VSS VDD sky130_fd_sc_hd__o2111ai_1
Xsky130_fd_sc_hd__nand2_1_270 sky130_fd_sc_hd__o211ai_1_8/B1 sky130_fd_sc_hd__a211o_1_8/A2
+ sky130_fd_sc_hd__o21ai_1_117/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_281 sky130_fd_sc_hd__a22o_1_68/B1 sky130_fd_sc_hd__nand2_2_3/Y
+ sky130_fd_sc_hd__o22ai_1_89/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_880 sky130_fd_sc_hd__o22ai_1_281/A1 sky130_fd_sc_hd__nor2_1_208/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_880/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_292 sky130_fd_sc_hd__xnor2_1_85/B sky130_fd_sc_hd__nand2_1_292/B
+ sky130_fd_sc_hd__nand2_1_295/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_109 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1048/B
+ sky130_fd_sc_hd__a211o_1_9/X VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkinv_1_891 sky130_fd_sc_hd__o32ai_1_3/B2 sky130_fd_sc_hd__fa_2_1175/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_891/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_19 sky130_fd_sc_hd__inv_2_5/A sky130_fd_sc_hd__ha_2_23/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_19/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_6 sky130_fd_sc_hd__fa_2_7/CIN sky130_fd_sc_hd__fa_2_6/SUM sky130_fd_sc_hd__fa_2_6/A
+ sky130_fd_sc_hd__fa_2_6/B sky130_fd_sc_hd__fa_2_6/CIN VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a211o_1_12 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_132/A sky130_fd_sc_hd__o21ai_1_236/Y
+ sky130_fd_sc_hd__nor2_1_125/Y sky130_fd_sc_hd__nand2_1_331/B sky130_fd_sc_hd__o22ai_1_168/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__a211o_1_23 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_251/A sky130_fd_sc_hd__nor2b_1_119/Y
+ sky130_fd_sc_hd__o22ai_1_351/Y sky130_fd_sc_hd__o21ai_1_424/Y sky130_fd_sc_hd__o22ai_1_350/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__clkinv_1_110 sky130_fd_sc_hd__inv_2_72/A sky130_fd_sc_hd__ha_2_43/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_110/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_121 sky130_fd_sc_hd__nor2b_1_26/B_N sky130_fd_sc_hd__ha_2_69/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_121/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_132 sky130_fd_sc_hd__clkinv_2_10/A sky130_fd_sc_hd__clkinv_1_132/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_132/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_143 sky130_fd_sc_hd__inv_2_80/A sky130_fd_sc_hd__inv_2_79/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_143/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_154 sky130_fd_sc_hd__buf_12_269/A sky130_fd_sc_hd__inv_2_85/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_154/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_165 sky130_fd_sc_hd__clkinv_1_166/A sky130_fd_sc_hd__inv_2_90/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_165/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_176 sky130_fd_sc_hd__bufinv_8_6/A sky130_fd_sc_hd__buf_8_128/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_176/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_8 sky130_fd_sc_hd__ha_2_19/A sky130_fd_sc_hd__buf_8_8/X VSS
+ VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__a22o_1_12 sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__ha_2_63/A
+ sky130_fd_sc_hd__a22o_1_12/X sky130_fd_sc_hd__dfxtp_1_8/Q sky130_fd_sc_hd__a22o_2_3/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_187 sky130_fd_sc_hd__nor3_2_8/C sky130_fd_sc_hd__nor3_2_9/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_187/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_23 sky130_fd_sc_hd__nor2_4_4/Y sky130_fd_sc_hd__ha_2_74/A
+ sky130_fd_sc_hd__a22o_1_23/X sky130_fd_sc_hd__a22o_1_23/B2 sky130_fd_sc_hd__a22o_2_6/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_198 sky130_fd_sc_hd__inv_2_106/A sky130_fd_sc_hd__a22o_1_30/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_198/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_34 sky130_fd_sc_hd__nor3_1_30/Y sky130_fd_sc_hd__nor2_1_29/Y
+ sky130_fd_sc_hd__a22o_1_34/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__a22o_1_34/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_45 sky130_fd_sc_hd__a22o_1_45/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_45/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__fa_2_951/SUM
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_56 sky130_fd_sc_hd__a22o_1_56/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_56/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__nor4_1_10/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_67 sky130_fd_sc_hd__nor2_1_41/Y sky130_fd_sc_hd__a22o_1_67/A2
+ sky130_fd_sc_hd__a22o_1_67/X sky130_fd_sc_hd__o21ai_1_74/Y sky130_fd_sc_hd__nor2_2_6/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__nand4_1_6 sky130_fd_sc_hd__nand4_1_6/C sky130_fd_sc_hd__nand4_1_6/B
+ sky130_fd_sc_hd__nand4_1_6/Y sky130_fd_sc_hd__nand4_1_6/D sky130_fd_sc_hd__nand4_1_6/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__clkinv_2_2 sky130_fd_sc_hd__clkinv_2_2/Y sky130_fd_sc_hd__clkinv_8_8/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_2/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__nor2_1_270 sky130_fd_sc_hd__nor2_1_270/B sky130_fd_sc_hd__o21a_1_57/A1
+ sky130_fd_sc_hd__o21a_1_58/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_281 sky130_fd_sc_hd__nor2_1_281/B sky130_fd_sc_hd__o21a_1_66/A1
+ sky130_fd_sc_hd__nor2_1_281/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_292 sky130_fd_sc_hd__nor2_1_292/B sky130_fd_sc_hd__nor2_1_292/Y
+ sky130_fd_sc_hd__nor2_1_309/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__maj3_1_18 sky130_fd_sc_hd__maj3_1_19/X sky130_fd_sc_hd__maj3_1_18/X
+ sky130_fd_sc_hd__maj3_1_18/B sky130_fd_sc_hd__maj3_1_18/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_29 sky130_fd_sc_hd__maj3_1_29/C sky130_fd_sc_hd__maj3_1_29/X
+ sky130_fd_sc_hd__maj3_1_29/B sky130_fd_sc_hd__maj3_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_408 sky130_fd_sc_hd__o32ai_1_10/B2 sky130_fd_sc_hd__nor2_1_309/A
+ sky130_fd_sc_hd__o22ai_1_408/Y sky130_fd_sc_hd__o22ai_1_433/A1 sky130_fd_sc_hd__a222oi_1_34/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_419 sky130_fd_sc_hd__o22ai_1_432/A2 sky130_fd_sc_hd__nor2_1_272/B
+ sky130_fd_sc_hd__o22ai_1_419/Y sky130_fd_sc_hd__nor2_1_273/B sky130_fd_sc_hd__o32ai_1_11/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__a22oi_1_380 sky130_fd_sc_hd__clkinv_1_861/Y sky130_fd_sc_hd__nor3_1_39/B
+ sky130_fd_sc_hd__fa_2_1179/A sky130_fd_sc_hd__fa_2_1180/A sky130_fd_sc_hd__a22oi_1_380/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_391 sky130_fd_sc_hd__fa_2_1232/A sky130_fd_sc_hd__nor2_1_267/Y
+ sky130_fd_sc_hd__nor2_1_265/Y sky130_fd_sc_hd__fa_2_1228/A sky130_fd_sc_hd__a22oi_1_391/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nand2_1_13 sky130_fd_sc_hd__nand3_1_13/C sky130_fd_sc_hd__nand4_1_66/Y
+ sky130_fd_sc_hd__nand2_1_9/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_24 sky130_fd_sc_hd__or2_0_2/B sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__nor2_1_3/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_35 sky130_fd_sc_hd__o21ai_1_9/A2 sky130_fd_sc_hd__nor2b_1_52/Y
+ sky130_fd_sc_hd__nand2_1_35/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_46 sky130_fd_sc_hd__nand2_1_46/Y sky130_fd_sc_hd__nand2_1_46/B
+ sky130_fd_sc_hd__a21oi_2_0/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_57 sky130_fd_sc_hd__nand2_1_57/Y sky130_fd_sc_hd__nand2_1_3/B
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_68 sky130_fd_sc_hd__nand2_1_68/Y sky130_fd_sc_hd__nand2_1_69/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_79 sky130_fd_sc_hd__nand2_1_79/Y sky130_fd_sc_hd__nand4_1_65/Y
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_1208 VDD VSS sky130_fd_sc_hd__fa_2_1257/A sky130_fd_sc_hd__clkinv_8_116/Y
+ sky130_fd_sc_hd__mux2_2_178/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1219 VDD VSS sky130_fd_sc_hd__fa_2_1231/A sky130_fd_sc_hd__clkinv_8_78/Y
+ sky130_fd_sc_hd__mux2_2_198/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_802 VDD VSS sky130_fd_sc_hd__fa_2_1054/A sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__mux2_2_71/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_813 VDD VSS sky130_fd_sc_hd__fa_2_1065/A sky130_fd_sc_hd__clkinv_4_25/Y
+ sky130_fd_sc_hd__mux2_2_47/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_824 VDD VSS sky130_fd_sc_hd__fa_2_1098/A sky130_fd_sc_hd__clkinv_8_59/Y
+ sky130_fd_sc_hd__and2_0_300/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_835 VDD VSS sky130_fd_sc_hd__nor2_4_13/A sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__nor2b_1_100/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_846 VDD VSS sky130_fd_sc_hd__mux2_2_61/A1 sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__o21ai_1_163/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_857 VDD VSS sky130_fd_sc_hd__mux2_2_40/A1 sky130_fd_sc_hd__clkinv_4_25/Y
+ sky130_fd_sc_hd__o21ai_1_174/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_868 VDD VSS sky130_fd_sc_hd__mux2_2_56/A1 sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__o21ai_1_182/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_879 VDD VSS sky130_fd_sc_hd__fa_2_863/A sky130_fd_sc_hd__dfxtp_1_899/CLK
+ sky130_fd_sc_hd__dfxtp_1_879/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_400 VSS VDD sky130_fd_sc_hd__clkbuf_1_400/X sky130_fd_sc_hd__clkbuf_1_400/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_411 VSS VDD sky130_fd_sc_hd__clkbuf_1_411/X sky130_fd_sc_hd__clkbuf_1_524/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_422 VSS VDD sky130_fd_sc_hd__clkbuf_1_422/X sky130_fd_sc_hd__clkbuf_1_526/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_433 VSS VDD sky130_fd_sc_hd__clkbuf_1_433/X sky130_fd_sc_hd__clkbuf_1_433/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_444 VSS VDD sky130_fd_sc_hd__a22oi_2_26/A2 sky130_fd_sc_hd__clkbuf_1_444/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_455 VSS VDD sky130_fd_sc_hd__clkbuf_1_455/X sky130_fd_sc_hd__clkbuf_1_455/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_466 VSS VDD sky130_fd_sc_hd__clkbuf_1_466/X sky130_fd_sc_hd__clkbuf_1_466/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_477 VSS VDD sky130_fd_sc_hd__nand4_1_59/D sky130_fd_sc_hd__a22oi_1_241/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_488 VSS VDD sky130_fd_sc_hd__buf_4_107/A sky130_fd_sc_hd__inv_2_132/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_499 VSS VDD sky130_fd_sc_hd__clkbuf_1_499/X sky130_fd_sc_hd__clkbuf_1_499/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_707 sky130_fd_sc_hd__fa_2_706/CIN sky130_fd_sc_hd__fa_2_707/SUM
+ sky130_fd_sc_hd__fa_2_707/A sky130_fd_sc_hd__fa_2_707/B sky130_fd_sc_hd__fa_2_707/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_718 sky130_fd_sc_hd__maj3_1_158/B sky130_fd_sc_hd__maj3_1_159/A
+ sky130_fd_sc_hd__ha_2_142/A sky130_fd_sc_hd__ha_2_142/B sky130_fd_sc_hd__ha_2_137/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_729 sky130_fd_sc_hd__maj3_1_152/B sky130_fd_sc_hd__maj3_1_153/A
+ sky130_fd_sc_hd__fa_2_729/A sky130_fd_sc_hd__fa_2_729/B sky130_fd_sc_hd__fa_2_730/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor2b_1_104 sky130_fd_sc_hd__o32ai_1_2/A1 sky130_fd_sc_hd__nor2b_1_104/Y
+ sky130_fd_sc_hd__nor2b_1_104/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_115 sky130_fd_sc_hd__nor2_1_200/Y sky130_fd_sc_hd__nor2b_1_115/Y
+ sky130_fd_sc_hd__buf_2_262/X VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_126 sky130_fd_sc_hd__nor2b_2_5/A sky130_fd_sc_hd__nor2b_1_126/Y
+ sky130_fd_sc_hd__o32ai_1_11/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_137 sky130_fd_sc_hd__nor2_1_322/Y sky130_fd_sc_hd__nor2_1_316/A
+ sky130_fd_sc_hd__nor2_1_321/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__buf_6_5 VDD VSS sky130_fd_sc_hd__buf_6_5/X sky130_fd_sc_hd__buf_6_5/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__bufbuf_8_8 sky130_fd_sc_hd__inv_2_132/Y sky130_fd_sc_hd__buf_6_68/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufbuf_8
Xsky130_fd_sc_hd__clkinv_2_40 sky130_fd_sc_hd__clkinv_4_32/A sky130_fd_sc_hd__clkinv_2_40/A
+ VSS VDD VDD VSS VSS sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__or2_1_0 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__or2_1_0/X sky130_fd_sc_hd__or2_1_0/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__or2_1
Xsky130_fd_sc_hd__o22ai_1_205 sky130_fd_sc_hd__nand2_2_6/Y sky130_fd_sc_hd__nor2_2_13/B
+ sky130_fd_sc_hd__o22ai_1_205/Y sky130_fd_sc_hd__a21oi_1_230/Y sky130_fd_sc_hd__a211oi_1_10/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__sdlclkp_4_3 sky130_fd_sc_hd__conb_1_1/LO sky130_fd_sc_hd__clkinv_8_47/A
+ sky130_fd_sc_hd__dfxtp_1_39/CLK sky130_fd_sc_hd__nor3_2_1/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__o22ai_1_216 sky130_fd_sc_hd__nand2_1_358/Y sky130_fd_sc_hd__nand2_1_357/Y
+ sky130_fd_sc_hd__o22ai_1_216/Y sky130_fd_sc_hd__nand2_1_370/B sky130_fd_sc_hd__o21ai_1_280/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_227 sky130_fd_sc_hd__nand2_1_360/Y sky130_fd_sc_hd__nand2_1_359/Y
+ sky130_fd_sc_hd__o22ai_1_227/Y sky130_fd_sc_hd__nand2_1_369/B sky130_fd_sc_hd__o21ai_1_279/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_238 sky130_fd_sc_hd__nor2_1_172/A sky130_fd_sc_hd__nor2_1_183/A
+ sky130_fd_sc_hd__o22ai_1_238/Y sky130_fd_sc_hd__a21boi_1_2/Y sky130_fd_sc_hd__a222oi_1_10/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_249 sky130_fd_sc_hd__nor2_1_149/B sky130_fd_sc_hd__nor2_1_182/A
+ sky130_fd_sc_hd__o22ai_1_249/Y sky130_fd_sc_hd__o22ai_1_262/A1 sky130_fd_sc_hd__a222oi_1_9/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_1_6 sky130_fd_sc_hd__nor2_1_6/B sky130_fd_sc_hd__nor2_1_6/Y
+ sky130_fd_sc_hd__nor2_1_7/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__bufinv_8_8 sky130_fd_sc_hd__bufinv_8_8/A sky130_fd_sc_hd__bufinv_8_8/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufinv_8
Xsky130_fd_sc_hd__dfxtp_1_109 VDD VSS sky130_fd_sc_hd__nor4_1_4/A sky130_fd_sc_hd__dfxtp_1_111/CLK
+ sky130_fd_sc_hd__ha_2_7/SUM VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_410 VSS VDD sky130_fd_sc_hd__nor2_1_265/A sky130_fd_sc_hd__a21oi_1_398/Y
+ sky130_fd_sc_hd__a211oi_1_26/Y sky130_fd_sc_hd__xor2_1_270/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_421 VSS VDD sky130_fd_sc_hd__a222oi_1_30/Y sky130_fd_sc_hd__nor2_1_265/A
+ sky130_fd_sc_hd__a21oi_1_401/Y sky130_fd_sc_hd__xor2_1_239/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_432 VSS VDD sky130_fd_sc_hd__nor2_1_265/A sky130_fd_sc_hd__a21oi_1_416/Y
+ sky130_fd_sc_hd__a211oi_1_29/Y sky130_fd_sc_hd__xor2_1_249/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_443 VSS VDD sky130_fd_sc_hd__nand2_1_527/B sky130_fd_sc_hd__nor2_1_297/Y
+ sky130_fd_sc_hd__nor2_1_296/B sky130_fd_sc_hd__o21ai_1_443/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_454 VSS VDD sky130_fd_sc_hd__nor2_1_302/B sky130_fd_sc_hd__nor2_1_309/A
+ sky130_fd_sc_hd__a21oi_1_443/Y sky130_fd_sc_hd__xor2_1_304/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_465 VSS VDD sky130_fd_sc_hd__a222oi_1_38/Y sky130_fd_sc_hd__nor2_1_309/A
+ sky130_fd_sc_hd__a22oi_1_399/Y sky130_fd_sc_hd__o21ai_1_465/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_476 VSS VDD sky130_fd_sc_hd__o21a_1_68/X sky130_fd_sc_hd__nor2_1_309/A
+ sky130_fd_sc_hd__a21oi_1_462/Y sky130_fd_sc_hd__xor2_1_287/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_487 VSS VDD sky130_fd_sc_hd__a211oi_1_37/Y sky130_fd_sc_hd__nor2_1_310/A
+ sky130_fd_sc_hd__a22oi_1_402/Y sky130_fd_sc_hd__o21ai_1_487/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_498 VSS VDD sky130_fd_sc_hd__nand2_1_559/A sky130_fd_sc_hd__o21ai_1_507/A1
+ sky130_fd_sc_hd__nand2_1_559/Y sky130_fd_sc_hd__and2_0_346/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_1208 sky130_fd_sc_hd__xor2_1_207/B sky130_fd_sc_hd__mux2_2_126/A0
+ sky130_fd_sc_hd__fa_2_1208/A sky130_fd_sc_hd__fa_2_1208/B sky130_fd_sc_hd__fa_2_1208/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1219 sky130_fd_sc_hd__fa_2_1220/CIN sky130_fd_sc_hd__mux2_2_151/A1
+ sky130_fd_sc_hd__fa_2_1219/A sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__fa_2_1219/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1005 VDD VSS sky130_fd_sc_hd__mux2_2_107/A0 sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__o22ai_1_234/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_14 VSS VDD sky130_fd_sc_hd__nor2b_1_52/Y sky130_fd_sc_hd__nand2_1_35/A
+ sky130_fd_sc_hd__o21ai_1_9/A2 sky130_fd_sc_hd__o21ai_1_14/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1016 VDD VSS sky130_fd_sc_hd__mux2_2_80/A1 sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__o22ai_1_223/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_25 VSS VDD sky130_fd_sc_hd__a21oi_2_0/Y sky130_fd_sc_hd__maj3_1_2/B
+ sky130_fd_sc_hd__nand2_1_44/Y sky130_fd_sc_hd__o21ai_1_25/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1027 VDD VSS sky130_fd_sc_hd__fa_2_842/A sky130_fd_sc_hd__dfxtp_1_1047/CLK
+ sky130_fd_sc_hd__o21a_1_39/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_36 VSS VDD sky130_fd_sc_hd__o21ai_1_36/A2 sky130_fd_sc_hd__o21ai_1_36/A1
+ sky130_fd_sc_hd__o21ai_1_36/B1 sky130_fd_sc_hd__o21ai_1_36/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1038 VDD VSS sky130_fd_sc_hd__fa_2_904/B sky130_fd_sc_hd__dfxtp_1_1038/CLK
+ sky130_fd_sc_hd__o21a_1_35/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_47 VSS VDD sky130_fd_sc_hd__o21ai_1_53/A2 sky130_fd_sc_hd__xnor2_1_48/Y
+ sky130_fd_sc_hd__a21oi_1_35/Y sky130_fd_sc_hd__o21ai_1_47/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_610 VDD VSS sky130_fd_sc_hd__and2_0_224/A sky130_fd_sc_hd__dfxtp_1_611/CLK
+ sky130_fd_sc_hd__fa_2_1030/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_270 sky130_fd_sc_hd__fa_2_1242/A sky130_fd_sc_hd__fa_2_1244/B
+ sky130_fd_sc_hd__xor2_1_270/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_1049 VDD VSS sky130_fd_sc_hd__fa_2_915/B sky130_fd_sc_hd__dfxtp_1_1050/CLK
+ sky130_fd_sc_hd__o21a_1_30/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_58 VSS VDD sky130_fd_sc_hd__nand2_2_3/Y sky130_fd_sc_hd__xnor2_1_36/Y
+ sky130_fd_sc_hd__a21oi_1_44/Y sky130_fd_sc_hd__o21ai_1_58/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_621 VDD VSS sky130_fd_sc_hd__fa_2_793/A sky130_fd_sc_hd__dfxtp_1_626/CLK
+ sky130_fd_sc_hd__a21oi_1_75/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_281 sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1290/B
+ sky130_fd_sc_hd__xor2_1_281/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o21ai_1_69 VSS VDD sky130_fd_sc_hd__nand2_2_3/Y sky130_fd_sc_hd__xnor2_1_58/Y
+ sky130_fd_sc_hd__a21oi_1_55/Y sky130_fd_sc_hd__o21ai_1_69/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_632 VDD VSS sky130_fd_sc_hd__fa_2_996/A sky130_fd_sc_hd__clkinv_8_41/Y
+ sky130_fd_sc_hd__and2_0_286/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_292 sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1279/B
+ sky130_fd_sc_hd__xor2_1_292/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_643 VDD VSS sky130_fd_sc_hd__fa_2_1007/A sky130_fd_sc_hd__clkinv_8_44/Y
+ sky130_fd_sc_hd__mux2_2_18/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_654 VDD VSS sky130_fd_sc_hd__fa_2_971/A sky130_fd_sc_hd__clkinv_8_41/Y
+ sky130_fd_sc_hd__and2_0_278/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_665 VDD VSS sky130_fd_sc_hd__fa_2_982/A sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__mux2_2_23/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_676 VDD VSS sky130_fd_sc_hd__xor2_1_60/A sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__mux2_2_2/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_687 VDD VSS sky130_fd_sc_hd__fa_2_1026/A sky130_fd_sc_hd__clkinv_8_54/Y
+ sky130_fd_sc_hd__and2_0_290/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_698 VDD VSS sky130_fd_sc_hd__nor2_4_10/B sky130_fd_sc_hd__clkinv_8_41/Y
+ sky130_fd_sc_hd__nor2b_1_92/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_230 VSS VDD sky130_fd_sc_hd__clkbuf_1_230/X sky130_fd_sc_hd__clkbuf_1_230/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_241 VSS VDD sky130_fd_sc_hd__buf_12_136/A sky130_fd_sc_hd__buf_8_66/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_252 VSS VDD sky130_fd_sc_hd__buf_2_123/A sky130_fd_sc_hd__clkbuf_1_252/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_263 VSS VDD sky130_fd_sc_hd__clkbuf_1_263/X sky130_fd_sc_hd__nand3_1_34/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_274 VSS VDD sky130_fd_sc_hd__clkbuf_1_274/X sky130_fd_sc_hd__clkbuf_1_274/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_285 VSS VDD sky130_fd_sc_hd__clkbuf_1_285/X sky130_fd_sc_hd__clkbuf_1_285/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_296 VSS VDD sky130_fd_sc_hd__clkbuf_1_296/X sky130_fd_sc_hd__clkbuf_1_296/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_504 sky130_fd_sc_hd__maj3_1_93/B sky130_fd_sc_hd__maj3_1_94/A
+ sky130_fd_sc_hd__fa_2_504/A sky130_fd_sc_hd__fa_2_504/B sky130_fd_sc_hd__fa_2_505/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_515 sky130_fd_sc_hd__fa_2_512/B sky130_fd_sc_hd__fa_2_515/SUM
+ sky130_fd_sc_hd__ha_2_123/A sky130_fd_sc_hd__fa_2_554/A sky130_fd_sc_hd__fa_2_566/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_526 sky130_fd_sc_hd__fa_2_528/CIN sky130_fd_sc_hd__fa_2_520/B
+ sky130_fd_sc_hd__fa_2_566/B sky130_fd_sc_hd__fa_2_559/B sky130_fd_sc_hd__fa_2_526/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_537 sky130_fd_sc_hd__fa_2_539/CIN sky130_fd_sc_hd__fa_2_533/A
+ sky130_fd_sc_hd__fa_2_537/A sky130_fd_sc_hd__fa_2_537/B sky130_fd_sc_hd__fa_2_537/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_548 sky130_fd_sc_hd__maj3_1_84/B sky130_fd_sc_hd__maj3_1_85/A
+ sky130_fd_sc_hd__fa_2_548/A sky130_fd_sc_hd__fa_2_548/B sky130_fd_sc_hd__fa_2_549/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_559 sky130_fd_sc_hd__fa_2_560/A sky130_fd_sc_hd__fa_2_556/A
+ sky130_fd_sc_hd__fa_2_559/A sky130_fd_sc_hd__fa_2_559/B sky130_fd_sc_hd__fa_2_559/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_4_2 VDD VSS sky130_fd_sc_hd__buf_4_2/X sky130_fd_sc_hd__buf_4_2/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__and2_0_250 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_250/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__and2_0_250/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_261 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_261/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__fa_2_962/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_272 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_272/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__and2_0_272/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_283 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_283/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__fa_2_995/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_294 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_294/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_294/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_509 sky130_fd_sc_hd__buf_12_509/A sky130_fd_sc_hd__buf_12_509/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__sdlclkp_2_0 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__clkinv_4_53/Y
+ sky130_fd_sc_hd__dfxtp_1_99/CLK sky130_fd_sc_hd__or2_0_0/X VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__clkinv_1_709 sky130_fd_sc_hd__nand4_1_86/B sky130_fd_sc_hd__fa_2_1048/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_709/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_240 VSS VDD sky130_fd_sc_hd__o22ai_1_196/B1 sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__nand2_1_330/Y sky130_fd_sc_hd__xor2_1_89/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_251 VSS VDD sky130_fd_sc_hd__o21ai_1_251/A2 sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__a21oi_1_218/Y sky130_fd_sc_hd__xor2_1_100/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_262 VSS VDD sky130_fd_sc_hd__nor2_1_127/A sky130_fd_sc_hd__a21oi_1_235/Y
+ sky130_fd_sc_hd__a21oi_1_227/Y sky130_fd_sc_hd__xor2_1_106/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_80 sky130_fd_sc_hd__clkbuf_4_80/X sky130_fd_sc_hd__clkbuf_4_80/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_273 VSS VDD sky130_fd_sc_hd__o21a_1_16/A2 sky130_fd_sc_hd__o21ai_1_273/A1
+ sky130_fd_sc_hd__a22oi_1_368/Y sky130_fd_sc_hd__o21ai_1_273/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_91 sky130_fd_sc_hd__nand4_1_24/A sky130_fd_sc_hd__clkbuf_4_91/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_284 VSS VDD sky130_fd_sc_hd__nor2_1_163/Y sky130_fd_sc_hd__or3_1_2/C
+ sky130_fd_sc_hd__o31ai_1_6/A1 sky130_fd_sc_hd__o21ai_1_284/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_295 VSS VDD sky130_fd_sc_hd__nor2_1_182/A sky130_fd_sc_hd__a21oi_1_278/Y
+ sky130_fd_sc_hd__a21oi_1_269/Y sky130_fd_sc_hd__xor2_1_176/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2b_2_2 sky130_fd_sc_hd__or2_1_1/A sky130_fd_sc_hd__or2_1_1/B
+ sky130_fd_sc_hd__nor2b_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_2
Xsky130_fd_sc_hd__fa_2_1005 sky130_fd_sc_hd__fa_2_1006/CIN sky130_fd_sc_hd__mux2_2_22/A0
+ sky130_fd_sc_hd__fa_2_1005/A sky130_fd_sc_hd__xor2_1_71/X sky130_fd_sc_hd__fa_2_1005/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1016 sky130_fd_sc_hd__fa_2_1017/CIN sky130_fd_sc_hd__and2_0_269/A
+ sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_1016/B sky130_fd_sc_hd__fa_2_970/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1027 sky130_fd_sc_hd__fa_2_1028/CIN sky130_fd_sc_hd__and2_0_291/A
+ sky130_fd_sc_hd__fa_2_1027/A sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_1027/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1038 sky130_fd_sc_hd__fa_2_1039/CIN sky130_fd_sc_hd__fa_2_1038/SUM
+ sky130_fd_sc_hd__nor2_1_59/A sky130_fd_sc_hd__fa_2_1038/B sky130_fd_sc_hd__fa_2_1038/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1049 sky130_fd_sc_hd__fa_2_1050/CIN sky130_fd_sc_hd__and2_0_309/A
+ sky130_fd_sc_hd__fa_2_1049/A sky130_fd_sc_hd__fa_2_1049/B sky130_fd_sc_hd__fa_2_1049/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_14 sky130_fd_sc_hd__inv_2_14/A sky130_fd_sc_hd__inv_2_14/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_25 sky130_fd_sc_hd__inv_2_25/A sky130_fd_sc_hd__inv_2_25/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_36 sky130_fd_sc_hd__inv_2_36/A sky130_fd_sc_hd__inv_2_36/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_440 VDD VSS sky130_fd_sc_hd__xor2_1_275/A sky130_fd_sc_hd__dfxtp_1_454/CLK
+ sky130_fd_sc_hd__nand2_1_84/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_47 sky130_fd_sc_hd__inv_2_47/A sky130_fd_sc_hd__inv_2_47/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_451 VDD VSS sky130_fd_sc_hd__dfxtp_1_997/D sky130_fd_sc_hd__dfxtp_1_454/CLK
+ sky130_fd_sc_hd__nand2_1_62/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_58 sky130_fd_sc_hd__inv_2_58/A sky130_fd_sc_hd__inv_2_58/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_462 VDD VSS sky130_fd_sc_hd__buf_2_8/A sky130_fd_sc_hd__dfxtp_1_462/CLK
+ sky130_fd_sc_hd__and2_0_239/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_69 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__inv_2_69/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_473 VDD VSS sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__dfxtp_1_473/CLK
+ sky130_fd_sc_hd__and2_0_107/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_484 VDD VSS sky130_fd_sc_hd__nor2b_1_88/A sky130_fd_sc_hd__dfxtp_1_488/CLK
+ sky130_fd_sc_hd__nor2b_1_74/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_2_4 sky130_fd_sc_hd__nor2_1_74/A sky130_fd_sc_hd__nand2_2_4/A
+ sky130_fd_sc_hd__nand2_2_4/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__dfxtp_1_495 VDD VSS sky130_fd_sc_hd__nor2b_1_85/A sky130_fd_sc_hd__dfxtp_1_502/CLK
+ sky130_fd_sc_hd__nor2b_1_58/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2b_1_10 sky130_fd_sc_hd__fa_2_969/CIN sky130_fd_sc_hd__xor2_1_30/A
+ sky130_fd_sc_hd__xor2_1_30/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__fa_2_301 sky130_fd_sc_hd__fa_2_295/B sky130_fd_sc_hd__fa_2_302/CIN
+ sky130_fd_sc_hd__fa_2_404/A sky130_fd_sc_hd__ha_2_114/A sky130_fd_sc_hd__fa_2_409/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_312 sky130_fd_sc_hd__fa_2_309/B sky130_fd_sc_hd__fa_2_313/CIN
+ sky130_fd_sc_hd__fa_2_395/A sky130_fd_sc_hd__fa_2_312/B sky130_fd_sc_hd__fa_2_312/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_323 sky130_fd_sc_hd__maj3_1_81/B sky130_fd_sc_hd__fa_2_323/SUM
+ sky130_fd_sc_hd__fa_2_360/B sky130_fd_sc_hd__ha_2_112/A sky130_fd_sc_hd__ha_2_112/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_334 sky130_fd_sc_hd__maj3_1_74/B sky130_fd_sc_hd__maj3_1_75/A
+ sky130_fd_sc_hd__fa_2_334/A sky130_fd_sc_hd__fa_2_334/B sky130_fd_sc_hd__fa_2_335/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_345 sky130_fd_sc_hd__fa_2_348/CIN sky130_fd_sc_hd__fa_2_343/B
+ sky130_fd_sc_hd__ha_2_116/B sky130_fd_sc_hd__fa_2_345/B sky130_fd_sc_hd__fa_2_345/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_356 sky130_fd_sc_hd__maj3_1_68/B sky130_fd_sc_hd__maj3_1_69/A
+ sky130_fd_sc_hd__fa_2_356/A sky130_fd_sc_hd__fa_2_356/B sky130_fd_sc_hd__fa_2_357/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_367 sky130_fd_sc_hd__fa_2_371/B sky130_fd_sc_hd__fa_2_367/SUM
+ sky130_fd_sc_hd__fa_2_367/A sky130_fd_sc_hd__fa_2_367/B sky130_fd_sc_hd__fa_2_367/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_378 sky130_fd_sc_hd__fa_2_382/B sky130_fd_sc_hd__fa_2_378/SUM
+ sky130_fd_sc_hd__fa_2_378/A sky130_fd_sc_hd__fa_2_378/B sky130_fd_sc_hd__fa_2_378/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_19 sky130_fd_sc_hd__conb_1_12/LO sky130_fd_sc_hd__clkinv_2_7/Y
+ sky130_fd_sc_hd__dfxtp_1_182/CLK sky130_fd_sc_hd__nand3b_1_0/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__fa_2_389 sky130_fd_sc_hd__fa_2_388/B sky130_fd_sc_hd__fa_2_383/B
+ sky130_fd_sc_hd__fa_2_417/A sky130_fd_sc_hd__fa_2_389/B sky130_fd_sc_hd__fa_2_389/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_1_5 VDD VSS sky130_fd_sc_hd__and2_1_5/X sky130_fd_sc_hd__ha_2_57/A
+ sky130_fd_sc_hd__nor2_4_2/Y VDD VSS sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__diode_2_206 sig_frequency[7] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_217 amplitude_adc_done VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_228 sig_amplitude[0] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkinv_8_50 sky130_fd_sc_hd__clkinv_8_50/Y sky130_fd_sc_hd__clkinv_8_70/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_50/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_61 sky130_fd_sc_hd__clkinv_8_61/Y sky130_fd_sc_hd__clkinv_8_62/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_61/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_72 sky130_fd_sc_hd__clkinv_8_74/A sky130_fd_sc_hd__clkinv_8_72/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_72/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_83 sky130_fd_sc_hd__clkinv_8_84/A sky130_fd_sc_hd__clkinv_8_83/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_83/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_94 sky130_fd_sc_hd__clkinv_8_95/A sky130_fd_sc_hd__clkinv_8_94/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_70 sky130_fd_sc_hd__buf_4_15/X sky130_fd_sc_hd__buf_12_93/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_81 sky130_fd_sc_hd__buf_8_57/X sky130_fd_sc_hd__buf_12_82/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_92 sky130_fd_sc_hd__buf_12_92/A sky130_fd_sc_hd__buf_12_92/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__dfxtp_1_1380 VDD VSS sky130_fd_sc_hd__fa_2_1319/A sky130_fd_sc_hd__clkinv_8_65/Y
+ sky130_fd_sc_hd__mux2_2_253/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1391 VDD VSS sky130_fd_sc_hd__nor2_8_2/A sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__nor2b_1_131/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a22oi_1_19 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__nor3_2_0/A
+ sky130_fd_sc_hd__nand4_1_38/Y sig_frequency[6] sky130_fd_sc_hd__a22oi_1_19/Y VDD
+ VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_306 sky130_fd_sc_hd__buf_8_149/X sky130_fd_sc_hd__buf_12_306/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_317 sky130_fd_sc_hd__buf_4_91/X sky130_fd_sc_hd__buf_12_361/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_328 sky130_fd_sc_hd__buf_4_70/X sky130_fd_sc_hd__buf_12_328/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_339 sky130_fd_sc_hd__buf_6_41/X sky130_fd_sc_hd__buf_8_175/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_209 sky130_fd_sc_hd__clkbuf_4_111/X sky130_fd_sc_hd__clkbuf_4_112/X
+ sky130_fd_sc_hd__a22oi_1_209/B2 sky130_fd_sc_hd__clkbuf_1_282/X sky130_fd_sc_hd__a22oi_1_209/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__fa_2_890 sky130_fd_sc_hd__fa_2_889/CIN sky130_fd_sc_hd__fa_2_890/SUM
+ sky130_fd_sc_hd__fa_2_890/A sky130_fd_sc_hd__fa_2_890/B sky130_fd_sc_hd__fa_2_890/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor3_2_1 sky130_fd_sc_hd__or2_0_0/B sky130_fd_sc_hd__nor3_2_1/Y
+ sky130_fd_sc_hd__nor3_2_1/A sky130_fd_sc_hd__nor3_2_1/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_2
Xsky130_fd_sc_hd__clkinv_1_506 sky130_fd_sc_hd__a21oi_1_62/A1 sky130_fd_sc_hd__nor2_1_52/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_506/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_517 sky130_fd_sc_hd__nor2_1_57/B sky130_fd_sc_hd__fa_2_1034/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_517/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_528 sky130_fd_sc_hd__o21ai_1_73/A2 sky130_fd_sc_hd__nor2_1_91/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_528/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_539 sky130_fd_sc_hd__a21oi_1_91/A1 sky130_fd_sc_hd__nor2_1_81/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_539/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_20 sky130_fd_sc_hd__nor2_1_20/B sky130_fd_sc_hd__nor3_1_28/B
+ sky130_fd_sc_hd__nor2_1_9/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_31 sky130_fd_sc_hd__nor2_1_31/B sky130_fd_sc_hd__nor2_1_31/Y
+ sky130_fd_sc_hd__nor4_1_6/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_42 sky130_fd_sc_hd__nor2_1_42/B sky130_fd_sc_hd__nor2_1_42/Y
+ sky130_fd_sc_hd__nor2_1_55/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_53 sky130_fd_sc_hd__nor2_1_53/B sky130_fd_sc_hd__nor2_1_53/Y
+ sky130_fd_sc_hd__nor2_1_53/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_64 sky130_fd_sc_hd__nor2_1_64/B sky130_fd_sc_hd__o21a_1_2/A1
+ sky130_fd_sc_hd__o21a_1_3/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_4_19 sky130_fd_sc_hd__clkinv_8_34/A sky130_fd_sc_hd__clkinv_8_37/A
+ VSS VDD VDD VSS VSS sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nor2_1_75 sky130_fd_sc_hd__nor2_1_82/Y sky130_fd_sc_hd__nor2_1_75/Y
+ sky130_fd_sc_hd__nor2_1_76/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_86 sky130_fd_sc_hd__o21a_1_8/A2 sky130_fd_sc_hd__nor2_1_86/Y
+ sky130_fd_sc_hd__nor2_1_86/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_190 VSS VDD sky130_fd_sc_hd__mux2_2_190/A1 sky130_fd_sc_hd__mux2_2_190/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_190/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_97 sky130_fd_sc_hd__nor2_1_97/B sky130_fd_sc_hd__nor2_1_97/Y
+ sky130_fd_sc_hd__nor2_1_97/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_sram_2kbyte_1rw1r_32x512_8_5 sky130_fd_sc_hd__buf_6_19/X sky130_fd_sc_hd__buf_4_33/X
+ sky130_fd_sc_hd__clkbuf_4_60/X sky130_fd_sc_hd__buf_12_121/X sky130_fd_sc_hd__clkbuf_4_61/X
+ sky130_fd_sc_hd__clkbuf_4_64/X sky130_fd_sc_hd__buf_4_35/X sky130_fd_sc_hd__buf_12_122/X
+ sky130_fd_sc_hd__buf_4_37/X sky130_fd_sc_hd__buf_4_38/X sky130_fd_sc_hd__buf_4_39/X
+ sky130_fd_sc_hd__clkbuf_8_0/X sky130_fd_sc_hd__buf_4_40/X sky130_fd_sc_hd__clkbuf_4_67/X
+ sky130_fd_sc_hd__clkbuf_4_69/X sky130_fd_sc_hd__clkbuf_4_71/X sky130_fd_sc_hd__buf_6_19/X
+ sky130_fd_sc_hd__buf_4_33/X sky130_fd_sc_hd__clkbuf_4_60/X sky130_fd_sc_hd__buf_12_121/X
+ sky130_fd_sc_hd__clkbuf_4_61/X sky130_fd_sc_hd__clkbuf_4_64/X sky130_fd_sc_hd__buf_4_35/X
+ sky130_fd_sc_hd__buf_12_122/X sky130_fd_sc_hd__buf_4_37/X sky130_fd_sc_hd__buf_4_38/X
+ sky130_fd_sc_hd__buf_4_39/X sky130_fd_sc_hd__clkbuf_8_0/X sky130_fd_sc_hd__buf_4_40/X
+ sky130_fd_sc_hd__clkbuf_4_67/X sky130_fd_sc_hd__clkbuf_4_69/X sky130_fd_sc_hd__clkbuf_4_71/X
+ sky130_fd_sc_hd__buf_12_140/X sky130_fd_sc_hd__buf_12_198/X sky130_fd_sc_hd__buf_12_142/X
+ sky130_fd_sc_hd__buf_12_139/X sky130_fd_sc_hd__buf_12_176/X sky130_fd_sc_hd__buf_12_265/X
+ sky130_fd_sc_hd__buf_12_197/X sky130_fd_sc_hd__buf_12_190/X sky130_fd_sc_hd__buf_12_261/X
+ sky130_fd_sc_hd__buf_12_124/X sky130_fd_sc_hd__buf_12_256/X sky130_fd_sc_hd__buf_12_263/X
+ sky130_fd_sc_hd__buf_12_217/X sky130_fd_sc_hd__buf_12_244/X sky130_fd_sc_hd__buf_12_245/X
+ sky130_fd_sc_hd__buf_12_172/X sky130_fd_sc_hd__buf_12_251/X sky130_fd_sc_hd__buf_12_262/X
+ sky130_fd_sc_hd__clkbuf_1_174/X sky130_fd_sc_hd__clkbuf_1_192/X sky130_fd_sc_hd__clkbuf_1_174/X
+ sky130_fd_sc_hd__clkinv_8_132/Y sky130_fd_sc_hd__clkinv_8_129/Y sky130_fd_sc_hd__buf_12_196/X
+ sky130_fd_sc_hd__buf_12_201/X sky130_fd_sc_hd__buf_12_233/X sky130_fd_sc_hd__buf_12_166/X
+ sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[0] sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[1]
+ sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[2] sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[3]
+ sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[4] sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[5]
+ sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[6] sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[7]
+ sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[8] sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[9]
+ sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[10] sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[11]
+ sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[12] sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[13]
+ sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[14] sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[15]
+ sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[16] sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[17]
+ sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[18] sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[19]
+ sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[20] sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[21]
+ sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[22] sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[23]
+ sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[24] sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[25]
+ sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[26] sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[27]
+ sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[28] sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[29]
+ sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[30] sky130_sram_2kbyte_1rw1r_32x512_8_5/dout0[31]
+ sky130_fd_sc_hd__buf_2_52/A sky130_fd_sc_hd__clkbuf_1_155/A sky130_fd_sc_hd__clkbuf_1_200/A
+ sky130_fd_sc_hd__buf_2_53/A sky130_fd_sc_hd__buf_2_54/A sky130_fd_sc_hd__buf_2_55/A
+ sky130_fd_sc_hd__buf_2_56/A sky130_fd_sc_hd__buf_2_57/A sky130_fd_sc_hd__buf_2_58/A
+ sky130_fd_sc_hd__buf_2_59/A sky130_fd_sc_hd__buf_2_60/A sky130_fd_sc_hd__buf_2_61/A
+ sky130_fd_sc_hd__buf_2_62/A sky130_fd_sc_hd__buf_2_63/A sky130_fd_sc_hd__buf_2_64/A
+ sky130_fd_sc_hd__buf_2_65/A sky130_fd_sc_hd__clkbuf_1_157/A sky130_fd_sc_hd__clkbuf_1_158/A
+ sky130_fd_sc_hd__clkbuf_1_159/A sky130_fd_sc_hd__clkbuf_1_160/A sky130_fd_sc_hd__clkbuf_1_161/A
+ sky130_fd_sc_hd__clkbuf_1_162/A sky130_fd_sc_hd__clkbuf_1_163/A sky130_fd_sc_hd__clkbuf_1_249/A
+ sky130_fd_sc_hd__clkbuf_1_165/A sky130_fd_sc_hd__clkbuf_1_166/A sky130_fd_sc_hd__clkbuf_1_247/A
+ sky130_fd_sc_hd__clkbuf_1_252/A sky130_fd_sc_hd__clkbuf_1_169/A sky130_fd_sc_hd__clkbuf_1_170/A
+ sky130_fd_sc_hd__clkbuf_1_171/A sky130_fd_sc_hd__clkbuf_1_172/A VDD VSS sky130_sram_2kbyte_1rw1r_32x512_8
Xsky130_fd_sc_hd__a21oi_1_403 sky130_fd_sc_hd__fa_2_1250/A sky130_fd_sc_hd__o22ai_1_367/Y
+ sky130_fd_sc_hd__a21oi_1_403/Y sky130_fd_sc_hd__nor3_1_40/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_414 sky130_fd_sc_hd__fa_2_1250/A sky130_fd_sc_hd__o22ai_1_372/Y
+ sky130_fd_sc_hd__a21oi_1_414/Y sky130_fd_sc_hd__nor2_2_17/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_425 sky130_fd_sc_hd__nor2_1_273/A sky130_fd_sc_hd__o21a_1_60/A1
+ sky130_fd_sc_hd__a21oi_1_425/Y sky130_fd_sc_hd__nor2_1_273/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_436 sky130_fd_sc_hd__nor2_1_284/A sky130_fd_sc_hd__nor2_1_284/Y
+ sky130_fd_sc_hd__a21oi_1_436/Y sky130_fd_sc_hd__nor2_1_284/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_447 sky130_fd_sc_hd__a21oi_1_447/A1 sky130_fd_sc_hd__nor2_1_300/Y
+ sky130_fd_sc_hd__a21oi_1_447/Y sky130_fd_sc_hd__nor2b_2_5/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_458 sky130_fd_sc_hd__fa_2_1281/A sky130_fd_sc_hd__o22ai_1_419/Y
+ sky130_fd_sc_hd__a21oi_1_458/Y sky130_fd_sc_hd__nor3_1_41/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_469 sky130_fd_sc_hd__nand2_1_543/B sky130_fd_sc_hd__o22ai_1_426/Y
+ sky130_fd_sc_hd__a21oi_1_469/Y sky130_fd_sc_hd__o21ai_1_491/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_8_105 sky130_fd_sc_hd__clkinv_8_105/Y sky130_fd_sc_hd__clkinv_8_67/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_105/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_116 sky130_fd_sc_hd__clkinv_8_116/Y sky130_fd_sc_hd__clkinv_8_75/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_116/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_127 sky130_fd_sc_hd__clkinv_8_128/A sky130_fd_sc_hd__clkinv_8_127/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_127/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_138 sky130_fd_sc_hd__clkinv_8_17/A sky130_fd_sc_hd__clkinv_4_75/Y
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__o21a_1_7 sky130_fd_sc_hd__o21a_1_7/X sky130_fd_sc_hd__o21a_1_7/A1
+ sky130_fd_sc_hd__o21a_1_7/B1 sky130_fd_sc_hd__fa_2_977/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__maj3_1_150 sky130_fd_sc_hd__maj3_1_151/X sky130_fd_sc_hd__maj3_1_150/X
+ sky130_fd_sc_hd__maj3_1_150/B sky130_fd_sc_hd__maj3_1_150/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_161 sky130_fd_sc_hd__fa_2_758/B sky130_fd_sc_hd__maj3_1_161/X
+ sky130_fd_sc_hd__ha_2_142/B sky130_fd_sc_hd__maj3_1_161/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_430 sky130_fd_sc_hd__nand2_1_430/Y sky130_fd_sc_hd__nand2_1_439/B
+ sky130_fd_sc_hd__o21ai_1_348/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_441 sky130_fd_sc_hd__nand2_1_441/Y sky130_fd_sc_hd__nor2b_1_112/Y
+ sky130_fd_sc_hd__o21ai_1_377/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_452 sky130_fd_sc_hd__nor2_1_234/A sky130_fd_sc_hd__fa_2_1226/A
+ sky130_fd_sc_hd__fa_2_1225/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_463 sky130_fd_sc_hd__nand2_1_463/Y sky130_fd_sc_hd__xor2_1_275/B
+ sky130_fd_sc_hd__nor2_1_245/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_474 sky130_fd_sc_hd__nor2_1_253/B sky130_fd_sc_hd__nand2_1_474/B
+ sky130_fd_sc_hd__nor2_1_254/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_485 sky130_fd_sc_hd__nand2_1_485/Y sky130_fd_sc_hd__nor2b_1_119/Y
+ sky130_fd_sc_hd__o21ai_1_409/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_496 sky130_fd_sc_hd__o32ai_1_11/A3 sky130_fd_sc_hd__nor2_4_19/B
+ sky130_fd_sc_hd__nor2_4_19/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_10 sky130_fd_sc_hd__ha_2_23/SUM sky130_fd_sc_hd__nor2b_1_10/Y
+ sky130_fd_sc_hd__or2_0_1/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_21 sky130_fd_sc_hd__ha_2_45/SUM sky130_fd_sc_hd__nor2b_1_21/Y
+ sky130_fd_sc_hd__or2_1_0/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_32 sky130_fd_sc_hd__ha_2_68/SUM sky130_fd_sc_hd__nor2b_1_32/Y
+ sky130_fd_sc_hd__or2_0_2/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_43 sky130_fd_sc_hd__ha_2_88/SUM sky130_fd_sc_hd__nor2b_1_43/Y
+ sky130_fd_sc_hd__or2_0_3/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1010 sky130_fd_sc_hd__o22ai_1_373/B1 sky130_fd_sc_hd__fa_2_1259/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1010/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1021 sky130_fd_sc_hd__o22ai_1_378/A1 sky130_fd_sc_hd__fa_2_1250/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1021/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_54 sky130_fd_sc_hd__a21oi_2_0/Y sky130_fd_sc_hd__nor2b_1_54/Y
+ sky130_fd_sc_hd__o31ai_1_0/A3 VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_65 sky130_fd_sc_hd__nor2b_1_89/A sky130_fd_sc_hd__nor2b_1_65/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1032 sky130_fd_sc_hd__o22ai_1_432/A2 sky130_fd_sc_hd__nor2_2_18/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1032/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_76 sky130_fd_sc_hd__dfxtp_1_490/Q sky130_fd_sc_hd__nor2b_1_76/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1043 sky130_fd_sc_hd__o32ai_1_10/A3 sky130_fd_sc_hd__fa_2_1294/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1043/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_87 sky130_fd_sc_hd__fa_2_949/A sky130_fd_sc_hd__or3_1_0/A
+ sky130_fd_sc_hd__nor2b_1_87/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1054 sky130_fd_sc_hd__o22ai_1_403/A1 sky130_fd_sc_hd__fa_2_19/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1054/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_98 sky130_fd_sc_hd__or2_0_8/X sky130_fd_sc_hd__nor2b_1_98/Y
+ sky130_fd_sc_hd__buf_2_262/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1065 sky130_fd_sc_hd__nand2_1_523/B sky130_fd_sc_hd__fa_2_2/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1065/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_6 VSS VDD sky130_fd_sc_hd__xnor2_1_6/B sky130_fd_sc_hd__xnor2_1_6/Y
+ sky130_fd_sc_hd__xnor2_1_7/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_1076 sky130_fd_sc_hd__o21ai_1_466/A2 sky130_fd_sc_hd__fa_2_1289/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1076/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1087 sky130_fd_sc_hd__nor2_1_272/B sky130_fd_sc_hd__fa_2_1284/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1087/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1098 sky130_fd_sc_hd__o22ai_1_433/A1 sky130_fd_sc_hd__nor2_1_309/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1098/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_270 VDD VSS sky130_fd_sc_hd__dfxtp_1_270/Q sky130_fd_sc_hd__dfxtp_1_277/CLK
+ sky130_fd_sc_hd__and2_0_214/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_281 VDD VSS sky130_fd_sc_hd__buf_2_284/A sky130_fd_sc_hd__dfxtp_1_282/CLK
+ sky130_fd_sc_hd__o21ai_1_30/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_292 VDD VSS sky130_fd_sc_hd__a22o_1_55/A1 sky130_fd_sc_hd__clkinv_4_31/Y
+ sky130_fd_sc_hd__nand2_1_125/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o22ai_1_1 sky130_fd_sc_hd__fa_2_80/B sky130_fd_sc_hd__fa_2_2/B sky130_fd_sc_hd__xnor2_1_0/B
+ sky130_fd_sc_hd__ha_2_97/A sky130_fd_sc_hd__fa_2_5/A VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_120 sky130_fd_sc_hd__fa_2_122/CIN sky130_fd_sc_hd__fa_2_117/A
+ sky130_fd_sc_hd__fa_2_139/B sky130_fd_sc_hd__fa_2_120/B sky130_fd_sc_hd__fa_2_120/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_131 sky130_fd_sc_hd__fa_2_130/A sky130_fd_sc_hd__fa_2_131/SUM
+ sky130_fd_sc_hd__fa_2_87/B sky130_fd_sc_hd__fa_2_86/A sky130_fd_sc_hd__fa_2_45/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_142 sky130_fd_sc_hd__fa_2_148/CIN sky130_fd_sc_hd__nor2_1_253/A
+ sky130_fd_sc_hd__fa_2_142/A sky130_fd_sc_hd__fa_2_142/B sky130_fd_sc_hd__fa_2_142/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_153 sky130_fd_sc_hd__fa_2_148/A sky130_fd_sc_hd__fa_2_142/B
+ sky130_fd_sc_hd__fa_2_280/A sky130_fd_sc_hd__fa_2_153/B sky130_fd_sc_hd__fa_2_241/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_164 sky130_fd_sc_hd__fa_2_161/CIN sky130_fd_sc_hd__fa_2_164/SUM
+ sky130_fd_sc_hd__fa_2_164/A sky130_fd_sc_hd__fa_2_164/B sky130_fd_sc_hd__fa_2_164/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_175 sky130_fd_sc_hd__maj3_1_52/B sky130_fd_sc_hd__maj3_1_53/A
+ sky130_fd_sc_hd__fa_2_67/B sky130_fd_sc_hd__fa_2_265/B sky130_fd_sc_hd__fa_2_175/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_186 sky130_fd_sc_hd__maj3_1_47/B sky130_fd_sc_hd__maj3_1_48/A
+ sky130_fd_sc_hd__fa_2_186/A sky130_fd_sc_hd__fa_2_186/B sky130_fd_sc_hd__fa_2_187/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_197 sky130_fd_sc_hd__fa_2_201/B sky130_fd_sc_hd__fa_2_197/SUM
+ sky130_fd_sc_hd__fa_2_197/A sky130_fd_sc_hd__fa_2_197/B sky130_fd_sc_hd__fa_2_197/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o22ai_1_30 sky130_fd_sc_hd__fa_2_389/B sky130_fd_sc_hd__fa_2_416/B
+ sky130_fd_sc_hd__fa_2_419/A sky130_fd_sc_hd__ha_2_110/A sky130_fd_sc_hd__ha_2_115/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_41 sky130_fd_sc_hd__fa_2_695/A sky130_fd_sc_hd__ha_2_130/A
+ sky130_fd_sc_hd__fa_2_607/A sky130_fd_sc_hd__fa_2_673/B sky130_fd_sc_hd__ha_2_135/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_52 sky130_fd_sc_hd__fa_2_793/A sky130_fd_sc_hd__ha_2_138/A
+ sky130_fd_sc_hd__fa_2_772/A sky130_fd_sc_hd__ha_2_143/B sky130_fd_sc_hd__fa_2_817/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_170 VDD VSS sky130_fd_sc_hd__buf_2_170/X sky130_fd_sc_hd__buf_2_170/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_63 sky130_fd_sc_hd__o22ai_1_88/B1 sky130_fd_sc_hd__nand2_2_3/Y
+ sky130_fd_sc_hd__o22ai_1_63/Y sky130_fd_sc_hd__xnor2_1_37/Y sky130_fd_sc_hd__o22ai_1_77/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_181 VDD VSS sky130_fd_sc_hd__buf_2_181/X sky130_fd_sc_hd__buf_2_248/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_74 sky130_fd_sc_hd__o22ai_1_88/B1 sky130_fd_sc_hd__nand2_2_3/Y
+ sky130_fd_sc_hd__o22ai_1_74/Y sky130_fd_sc_hd__xnor2_1_59/Y sky130_fd_sc_hd__o22ai_1_88/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_192 VDD VSS sky130_fd_sc_hd__buf_2_192/X sky130_fd_sc_hd__buf_2_192/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_85 sky130_fd_sc_hd__o22ai_1_89/A1 sky130_fd_sc_hd__o22ai_1_88/B1
+ sky130_fd_sc_hd__o22ai_1_85/Y sky130_fd_sc_hd__xnor2_1_53/Y sky130_fd_sc_hd__o22ai_1_85/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_96 sky130_fd_sc_hd__a21oi_1_90/Y sky130_fd_sc_hd__a21oi_1_99/Y
+ sky130_fd_sc_hd__o22ai_1_96/Y sky130_fd_sc_hd__nor2_2_9/B sky130_fd_sc_hd__nor2_1_76/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_4_10 VDD VSS sky130_fd_sc_hd__buf_4_10/X sky130_fd_sc_hd__buf_2_9/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_21 VDD VSS sky130_fd_sc_hd__buf_4_21/X sky130_fd_sc_hd__buf_8_2/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_32 VDD VSS sky130_fd_sc_hd__buf_4_32/X sky130_fd_sc_hd__buf_4_32/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_43 VDD VSS sky130_fd_sc_hd__buf_4_43/X sky130_fd_sc_hd__buf_4_43/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_54 VDD VSS sky130_fd_sc_hd__buf_4_54/X sky130_fd_sc_hd__buf_8_88/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_65 VDD VSS sky130_fd_sc_hd__buf_4_65/X sky130_fd_sc_hd__buf_6_85/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_76 VDD VSS sky130_fd_sc_hd__buf_4_76/X sky130_fd_sc_hd__buf_4_76/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_87 VDD VSS sky130_fd_sc_hd__buf_4_87/X sky130_fd_sc_hd__buf_4_87/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_98 VDD VSS sky130_fd_sc_hd__buf_4_98/X sky130_fd_sc_hd__buf_4_98/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_12_103 sky130_fd_sc_hd__buf_12_2/X sky130_fd_sc_hd__buf_12_103/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_114 sky130_fd_sc_hd__buf_12_114/A sky130_fd_sc_hd__buf_12_114/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_125 sky130_fd_sc_hd__inv_2_65/Y sky130_fd_sc_hd__buf_12_125/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_136 sky130_fd_sc_hd__buf_12_136/A sky130_fd_sc_hd__buf_12_247/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_147 sky130_fd_sc_hd__buf_8_73/X sky130_fd_sc_hd__buf_12_241/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_70 VSS VDD sky130_fd_sc_hd__clkbuf_1_70/X sky130_fd_sc_hd__clkbuf_1_70/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_158 sky130_fd_sc_hd__buf_8_105/X sky130_fd_sc_hd__buf_12_158/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_81 VSS VDD sky130_fd_sc_hd__nand4_1_6/A sky130_fd_sc_hd__a22oi_2_7/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_169 sky130_fd_sc_hd__buf_8_102/X sky130_fd_sc_hd__buf_12_169/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_92 VSS VDD sky130_fd_sc_hd__buf_6_11/A sky130_fd_sc_hd__ha_2_17/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_4_6 sky130_fd_sc_hd__clkbuf_4_6/X sky130_fd_sc_hd__clkbuf_4_6/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_1_303 sky130_fd_sc_hd__fa_2_277/B sky130_fd_sc_hd__ha_2_99/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_303/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_314 sky130_fd_sc_hd__fa_2_413/A sky130_fd_sc_hd__ha_2_114/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_314/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_325 sky130_fd_sc_hd__fa_2_427/B sky130_fd_sc_hd__ha_2_125/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_325/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_336 sky130_fd_sc_hd__fa_2_559/A sky130_fd_sc_hd__fa_2_502/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_336/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_347 sky130_fd_sc_hd__ha_2_131/B sky130_fd_sc_hd__fa_2_678/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_347/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_358 sky130_fd_sc_hd__fa_2_832/A sky130_fd_sc_hd__fa_2_833/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_358/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_369 sky130_fd_sc_hd__ha_2_140/B sky130_fd_sc_hd__ha_2_145/B
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_200 sky130_fd_sc_hd__fa_2_1068/A sky130_fd_sc_hd__nor2_1_128/Y
+ sky130_fd_sc_hd__a21oi_1_200/Y sky130_fd_sc_hd__nor2_4_12/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_211 sky130_fd_sc_hd__a21o_2_5/A2 sky130_fd_sc_hd__o22ai_1_187/Y
+ sky130_fd_sc_hd__a21oi_1_211/Y sky130_fd_sc_hd__fa_2_1049/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_222 sky130_fd_sc_hd__nor2_2_12/Y sky130_fd_sc_hd__o22ai_1_197/Y
+ sky130_fd_sc_hd__a21oi_1_222/Y sky130_fd_sc_hd__fa_2_1082/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_233 sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__a22o_1_74/X
+ sky130_fd_sc_hd__a21oi_1_233/Y sky130_fd_sc_hd__fa_2_1070/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_244 sky130_fd_sc_hd__o21a_1_21/B1 sky130_fd_sc_hd__o21a_1_20/A1
+ sky130_fd_sc_hd__dfxtp_1_901/D sky130_fd_sc_hd__nor2_1_145/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_255 sky130_fd_sc_hd__nor2_1_156/A sky130_fd_sc_hd__o21a_1_28/A1
+ sky130_fd_sc_hd__dfxtp_1_880/D sky130_fd_sc_hd__nor2_1_156/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_266 sky130_fd_sc_hd__fa_2_1130/A sky130_fd_sc_hd__o22ai_1_242/Y
+ sky130_fd_sc_hd__a21oi_1_266/Y sky130_fd_sc_hd__nor3_1_38/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_277 sky130_fd_sc_hd__fa_2_1133/A sky130_fd_sc_hd__o22ai_1_247/Y
+ sky130_fd_sc_hd__a21oi_1_277/Y sky130_fd_sc_hd__nor2_2_15/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_288 sky130_fd_sc_hd__nor2_1_182/Y sky130_fd_sc_hd__nor2_1_177/Y
+ sky130_fd_sc_hd__a21oi_1_288/Y sky130_fd_sc_hd__fa_2_1148/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_4_6 sky130_fd_sc_hd__clkinv_4_6/A sky130_fd_sc_hd__clkinv_8_8/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_6/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__a21oi_1_299 sky130_fd_sc_hd__fa_2_1150/A sky130_fd_sc_hd__o22ai_1_265/Y
+ sky130_fd_sc_hd__o21a_1_29/B1 sky130_fd_sc_hd__nor2_2_15/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_207 sky130_fd_sc_hd__buf_8_207/A sky130_fd_sc_hd__buf_8_207/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_218 sky130_fd_sc_hd__buf_8_218/A sky130_fd_sc_hd__buf_8_218/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__o2111ai_1_1 sky130_fd_sc_hd__nor4_1_11/Y sky130_fd_sc_hd__nor4_1_12/Y
+ sky130_fd_sc_hd__o21ai_1_35/Y sky130_fd_sc_hd__a21oi_1_21/Y sky130_fd_sc_hd__o22a_1_0/X
+ sky130_fd_sc_hd__o2111ai_1_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__o2111ai_1
Xsky130_fd_sc_hd__nand2_1_260 sky130_fd_sc_hd__o21ai_1_96/B1 sky130_fd_sc_hd__xor2_1_60/A
+ sky130_fd_sc_hd__nor2_1_74/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_271 sky130_fd_sc_hd__o211ai_1_9/B1 sky130_fd_sc_hd__a211o_1_8/A2
+ sky130_fd_sc_hd__o21ai_1_119/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_870 sky130_fd_sc_hd__o32ai_1_3/A2 sky130_fd_sc_hd__fa_2_1173/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_870/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_282 sky130_fd_sc_hd__nor2_2_9/B sky130_fd_sc_hd__nand2_1_282/B
+ sky130_fd_sc_hd__o22ai_1_90/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_881 sky130_fd_sc_hd__o22ai_1_283/A1 sky130_fd_sc_hd__nor2_1_209/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_881/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_293 sky130_fd_sc_hd__xnor2_1_89/B sky130_fd_sc_hd__nand2_1_293/B
+ sky130_fd_sc_hd__nand2_1_294/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_892 sky130_fd_sc_hd__nor2_1_190/B sky130_fd_sc_hd__fa_2_1177/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_892/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__fa_2_7 sky130_fd_sc_hd__fa_2_4/CIN sky130_fd_sc_hd__fa_2_7/SUM sky130_fd_sc_hd__fa_2_7/A
+ sky130_fd_sc_hd__fa_2_7/B sky130_fd_sc_hd__fa_2_7/CIN VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a211o_1_13 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_131/A sky130_fd_sc_hd__o21ai_1_234/Y
+ sky130_fd_sc_hd__nor2_1_126/Y sky130_fd_sc_hd__nand2_1_333/B sky130_fd_sc_hd__o22ai_1_169/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__a211o_1_24 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_247/A sky130_fd_sc_hd__o21ai_1_424/Y
+ sky130_fd_sc_hd__nor2_1_249/Y sky130_fd_sc_hd__nor2b_2_4/Y sky130_fd_sc_hd__o22ai_1_352/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__clkinv_1_100 sky130_fd_sc_hd__inv_2_64/A sky130_fd_sc_hd__ha_2_35/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_100/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_111 sky130_fd_sc_hd__clkbuf_4_97/A sky130_fd_sc_hd__buf_12_148/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_111/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_122 sky130_fd_sc_hd__nor3_2_6/C sky130_fd_sc_hd__nor3_2_5/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_122/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_133 sky130_fd_sc_hd__clkinv_2_11/A sky130_fd_sc_hd__clkinv_1_133/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_133/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_144 sky130_fd_sc_hd__inv_2_82/A sky130_fd_sc_hd__buf_8_119/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_144/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_155 sky130_fd_sc_hd__inv_2_86/A sky130_fd_sc_hd__clkinv_1_155/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_155/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_166 sky130_fd_sc_hd__buf_8_122/A sky130_fd_sc_hd__clkinv_1_166/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_166/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_177 sky130_fd_sc_hd__buf_8_152/A sky130_fd_sc_hd__bufinv_8_6/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_177/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_9 sky130_fd_sc_hd__buf_8_9/A sky130_fd_sc_hd__buf_8_9/X VSS
+ VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__a22o_1_13 sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__ha_2_65/A
+ sky130_fd_sc_hd__a22o_1_13/X sky130_fd_sc_hd__dfxtp_1_6/Q sky130_fd_sc_hd__a22o_2_3/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_188 sky130_fd_sc_hd__nor3_2_9/C sky130_fd_sc_hd__nor3_2_8/A
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_199 sky130_fd_sc_hd__clkinv_1_201/A sky130_fd_sc_hd__buf_2_243/X
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_24 sky130_fd_sc_hd__nor2_4_4/Y sky130_fd_sc_hd__ha_2_75/A
+ sky130_fd_sc_hd__a22o_1_24/X sky130_fd_sc_hd__a22o_1_24/B2 sky130_fd_sc_hd__a22o_2_6/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_35 sky130_fd_sc_hd__nor2_1_26/Y sky130_fd_sc_hd__nor2_1_29/Y
+ sky130_fd_sc_hd__a22o_1_35/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__a22o_1_35/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__o21ai_1_0 VSS VDD sky130_fd_sc_hd__nor3_1_4/B sky130_fd_sc_hd__o21ai_1_0/A1
+ sky130_fd_sc_hd__nor3_1_2/C sky130_fd_sc_hd__o21ai_1_0/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a22o_1_46 sky130_fd_sc_hd__a22o_1_46/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_46/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__fa_2_952/SUM
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_57 sky130_fd_sc_hd__a22o_1_57/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_57/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__nor4_1_9/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_68 sky130_fd_sc_hd__a22o_1_68/A1 sky130_fd_sc_hd__ha_2_185/SUM
+ sky130_fd_sc_hd__a22o_1_68/X sky130_fd_sc_hd__a22o_1_68/B2 sky130_fd_sc_hd__a22o_1_68/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__nand4_1_7 sky130_fd_sc_hd__nand4_1_7/C sky130_fd_sc_hd__nand4_1_7/B
+ sky130_fd_sc_hd__nand4_1_7/Y sky130_fd_sc_hd__nand4_1_7/D sky130_fd_sc_hd__nand4_1_7/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__clkinv_2_3 sky130_fd_sc_hd__clkinv_8_9/A sky130_fd_sc_hd__clkinv_4_5/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_3/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__nor2_1_260 sky130_fd_sc_hd__nor2_1_260/B sky130_fd_sc_hd__nor2_1_260/Y
+ sky130_fd_sc_hd__nor2_1_268/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_271 sky130_fd_sc_hd__nor2_1_271/B sky130_fd_sc_hd__o21a_1_58/A1
+ sky130_fd_sc_hd__o21a_1_59/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_282 sky130_fd_sc_hd__nor2_1_282/B sky130_fd_sc_hd__nor2_1_282/Y
+ sky130_fd_sc_hd__o21a_1_67/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_293 sky130_fd_sc_hd__nor2_1_293/B sky130_fd_sc_hd__nor2_1_293/Y
+ sky130_fd_sc_hd__fa_2_3/SUM VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__maj3_1_19 sky130_fd_sc_hd__maj3_1_20/X sky130_fd_sc_hd__maj3_1_19/X
+ sky130_fd_sc_hd__maj3_1_19/B sky130_fd_sc_hd__maj3_1_19/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_409 sky130_fd_sc_hd__nor2_1_299/A sky130_fd_sc_hd__nor2_1_310/A
+ sky130_fd_sc_hd__o22ai_1_409/Y sky130_fd_sc_hd__a21boi_1_8/Y sky130_fd_sc_hd__a222oi_1_40/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__a22oi_1_370 sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__nor2_4_13/Y
+ sky130_fd_sc_hd__fa_2_1077/A sky130_fd_sc_hd__fa_2_1078/A sky130_fd_sc_hd__a22oi_1_370/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_381 sky130_fd_sc_hd__nor2_1_222/Y sky130_fd_sc_hd__nor2_1_224/Y
+ sky130_fd_sc_hd__fa_2_1182/A sky130_fd_sc_hd__fa_2_1178/A sky130_fd_sc_hd__a22oi_1_381/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_392 sky130_fd_sc_hd__clkinv_1_946/Y sky130_fd_sc_hd__nor3_1_40/B
+ sky130_fd_sc_hd__fa_2_1240/A sky130_fd_sc_hd__fa_2_1241/A sky130_fd_sc_hd__a22oi_1_392/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nand2_1_14 sky130_fd_sc_hd__nand3_1_14/C sky130_fd_sc_hd__nand4_1_65/Y
+ sky130_fd_sc_hd__nand2_1_9/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_25 sky130_fd_sc_hd__nor2_2_3/B sky130_fd_sc_hd__nor3_2_6/B
+ sky130_fd_sc_hd__nor3_2_6/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_36 sky130_fd_sc_hd__nor2b_1_52/A sky130_fd_sc_hd__nor2b_1_53/Y
+ sky130_fd_sc_hd__nand2_1_36/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_47 sky130_fd_sc_hd__nand2_1_47/Y sky130_fd_sc_hd__nand2_1_47/B
+ sky130_fd_sc_hd__a21oi_2_0/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_58 sky130_fd_sc_hd__nand2_1_58/Y sky130_fd_sc_hd__nand2_1_59/Y
+ sky130_fd_sc_hd__nand2_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_69 sky130_fd_sc_hd__nand2_1_69/Y sky130_fd_sc_hd__nand2_1_9/B
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2_8_0 sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__nor2_8_0/A
+ sky130_fd_sc_hd__nor2_8_0/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_8
Xsky130_fd_sc_hd__dfxtp_1_1209 VDD VSS sky130_fd_sc_hd__fa_2_1258/A sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__mux2_2_176/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_803 VDD VSS sky130_fd_sc_hd__fa_2_1055/A sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__mux2_2_69/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_814 VDD VSS sky130_fd_sc_hd__o21a_1_9/A2 sky130_fd_sc_hd__clkinv_4_26/Y
+ sky130_fd_sc_hd__mux2_2_45/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_825 VDD VSS sky130_fd_sc_hd__fa_2_1099/A sky130_fd_sc_hd__clkinv_8_59/Y
+ sky130_fd_sc_hd__and2_0_305/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_836 VDD VSS sky130_fd_sc_hd__buf_2_254/A sky130_fd_sc_hd__clkinv_8_55/Y
+ sky130_fd_sc_hd__nor2b_1_101/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_847 VDD VSS sky130_fd_sc_hd__mux2_2_59/A1 sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__o21ai_1_164/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_858 VDD VSS sky130_fd_sc_hd__mux2_2_68/A1 sky130_fd_sc_hd__clkinv_4_26/Y
+ sky130_fd_sc_hd__a22o_1_73/A1 VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_869 VDD VSS sky130_fd_sc_hd__mux2_2_54/A1 sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__o21ai_1_183/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_401 VSS VDD sky130_fd_sc_hd__clkbuf_1_401/X sky130_fd_sc_hd__clkbuf_1_401/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_412 VSS VDD sky130_fd_sc_hd__clkbuf_1_412/X sky130_fd_sc_hd__clkbuf_1_412/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_423 VSS VDD sky130_fd_sc_hd__clkbuf_1_423/X sky130_fd_sc_hd__clkbuf_1_423/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_434 VSS VDD sky130_fd_sc_hd__clkbuf_1_434/X sky130_fd_sc_hd__clkbuf_1_434/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_445 VSS VDD sky130_fd_sc_hd__clkbuf_1_445/X sky130_fd_sc_hd__clkbuf_1_445/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_456 VSS VDD sky130_fd_sc_hd__clkbuf_1_456/X sky130_fd_sc_hd__clkbuf_1_456/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_467 VSS VDD sky130_fd_sc_hd__clkbuf_1_467/X sky130_fd_sc_hd__clkbuf_1_467/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_478 VSS VDD sky130_fd_sc_hd__nand4_1_54/B sky130_fd_sc_hd__a22oi_1_229/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_489 VSS VDD sky130_fd_sc_hd__clkbuf_1_489/X sky130_fd_sc_hd__clkbuf_1_540/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_708 sky130_fd_sc_hd__fa_2_707/CIN sky130_fd_sc_hd__fa_2_708/SUM
+ sky130_fd_sc_hd__fa_2_708/A sky130_fd_sc_hd__fa_2_708/B sky130_fd_sc_hd__fa_2_708/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_719 sky130_fd_sc_hd__maj3_1_157/B sky130_fd_sc_hd__maj3_1_158/A
+ sky130_fd_sc_hd__ha_2_136/A sky130_fd_sc_hd__fa_2_719/B sky130_fd_sc_hd__ha_2_138/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor2b_1_105 sky130_fd_sc_hd__nor2b_1_104/A sky130_fd_sc_hd__nor2b_1_105/Y
+ sky130_fd_sc_hd__o32ai_1_2/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_116 sky130_fd_sc_hd__o32ai_1_5/Y sky130_fd_sc_hd__nor2b_1_116/Y
+ sky130_fd_sc_hd__buf_2_262/X VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_127 sky130_fd_sc_hd__or2_0_12/X sky130_fd_sc_hd__nor2b_1_127/Y
+ sky130_fd_sc_hd__buf_2_262/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_138 sky130_fd_sc_hd__nor2_1_316/A sky130_fd_sc_hd__nor2b_1_138/Y
+ sky130_fd_sc_hd__nor2b_1_142/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__buf_6_6 VDD VSS sky130_fd_sc_hd__buf_6_6/X sky130_fd_sc_hd__buf_6_6/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__bufbuf_8_9 sky130_fd_sc_hd__bufbuf_8_9/A sky130_fd_sc_hd__bufbuf_8_9/X
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufbuf_8
Xsky130_fd_sc_hd__clkinv_2_30 sky130_fd_sc_hd__buf_8_186/A sky130_fd_sc_hd__clkinv_2_30/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_30/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_41 sky130_fd_sc_hd__clkinv_2_41/Y sky130_fd_sc_hd__clkinv_4_78/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_41/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__or2_1_1 sky130_fd_sc_hd__or2_1_1/A sky130_fd_sc_hd__or2_1_1/X sky130_fd_sc_hd__or2_1_1/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__or2_1
Xsky130_fd_sc_hd__o22ai_1_206 sky130_fd_sc_hd__nor2_1_137/A sky130_fd_sc_hd__o22ai_1_206/B1
+ sky130_fd_sc_hd__o22ai_1_206/Y sky130_fd_sc_hd__o22ai_1_206/A1 sky130_fd_sc_hd__o22ai_1_206/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__sdlclkp_4_4 sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__clkinv_8_69/A
+ sky130_fd_sc_hd__dfxtp_1_77/CLK sky130_fd_sc_hd__nor3_1_3/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__o22ai_1_217 sky130_fd_sc_hd__nand2_1_358/Y sky130_fd_sc_hd__nand2_1_357/Y
+ sky130_fd_sc_hd__o22ai_1_217/Y sky130_fd_sc_hd__o22ai_1_230/A1 sky130_fd_sc_hd__a21o_2_9/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_228 sky130_fd_sc_hd__nand2_1_360/Y sky130_fd_sc_hd__nand2_1_359/Y
+ sky130_fd_sc_hd__o22ai_1_228/Y sky130_fd_sc_hd__o22ai_1_228/A1 sky130_fd_sc_hd__a21o_2_8/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_239 sky130_fd_sc_hd__nor2_1_183/A sky130_fd_sc_hd__nor2_1_180/A
+ sky130_fd_sc_hd__o22ai_1_239/Y sky130_fd_sc_hd__a21boi_1_1/Y sky130_fd_sc_hd__nor2_1_165/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_1_7 sky130_fd_sc_hd__nor2_1_7/B sky130_fd_sc_hd__nor2_1_7/Y
+ sky130_fd_sc_hd__nor2_1_7/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__o21ai_1_400 VSS VDD sky130_fd_sc_hd__nor2_1_260/B sky130_fd_sc_hd__nor2_1_267/A
+ sky130_fd_sc_hd__a21oi_1_383/Y sky130_fd_sc_hd__xor2_1_259/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_411 VSS VDD sky130_fd_sc_hd__a222oi_1_28/Y sky130_fd_sc_hd__nor2_1_267/A
+ sky130_fd_sc_hd__a22oi_1_391/Y sky130_fd_sc_hd__o21ai_1_411/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_422 VSS VDD sky130_fd_sc_hd__o21a_1_55/X sky130_fd_sc_hd__nor2_1_267/A
+ sky130_fd_sc_hd__a21oi_1_402/Y sky130_fd_sc_hd__xor2_1_242/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_433 VSS VDD sky130_fd_sc_hd__a211oi_1_30/Y sky130_fd_sc_hd__nor2_1_268/A
+ sky130_fd_sc_hd__a22oi_1_394/Y sky130_fd_sc_hd__o21ai_1_433/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_444 VSS VDD sky130_fd_sc_hd__nand2_1_528/B sky130_fd_sc_hd__nor2_1_298/Y
+ sky130_fd_sc_hd__nor2_1_297/B sky130_fd_sc_hd__o21ai_1_444/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_455 VSS VDD sky130_fd_sc_hd__a222oi_1_36/Y sky130_fd_sc_hd__nor2_1_307/A
+ sky130_fd_sc_hd__a21oi_1_444/Y sky130_fd_sc_hd__xor2_1_305/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_466 VSS VDD sky130_fd_sc_hd__o21ai_1_466/A2 sky130_fd_sc_hd__o22ai_1_436/A2
+ sky130_fd_sc_hd__a22oi_1_400/Y sky130_fd_sc_hd__o21ai_1_466/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_477 VSS VDD sky130_fd_sc_hd__a21oi_1_470/Y sky130_fd_sc_hd__nor2_1_299/A
+ sky130_fd_sc_hd__o21ai_1_479/B1 sky130_fd_sc_hd__o21ai_1_477/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_488 VSS VDD sky130_fd_sc_hd__o22ai_1_432/A2 sky130_fd_sc_hd__o21a_1_68/A2
+ sky130_fd_sc_hd__a21oi_1_475/Y sky130_fd_sc_hd__o21ai_1_488/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_499 VSS VDD sky130_fd_sc_hd__nand2_1_560/A sky130_fd_sc_hd__o21ai_1_507/A1
+ sky130_fd_sc_hd__nand2_1_560/Y sky130_fd_sc_hd__and2_0_351/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_4_20 sky130_fd_sc_hd__nor2_4_20/Y sky130_fd_sc_hd__nor2_8_2/A
+ sky130_fd_sc_hd__nor2_4_20/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__fa_2_1209 sky130_fd_sc_hd__fa_2_1210/CIN sky130_fd_sc_hd__mux2_2_171/A1
+ sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__fa_2_1209/B sky130_fd_sc_hd__nor2_8_0/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1006 VDD VSS sky130_fd_sc_hd__mux2_2_104/A0 sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__o22ai_1_233/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_15 VSS VDD sky130_fd_sc_hd__nor2b_1_51/Y sky130_fd_sc_hd__nand2_1_34/A
+ sky130_fd_sc_hd__xor2_1_11/A sky130_fd_sc_hd__o21ai_1_7/A2 VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1017 VDD VSS sky130_fd_sc_hd__mux2_2_78/A1 sky130_fd_sc_hd__clkinv_8_46/Y
+ sky130_fd_sc_hd__o31ai_1_5/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_26 VSS VDD sky130_fd_sc_hd__a21oi_2_0/Y sky130_fd_sc_hd__maj3_1_3/C
+ sky130_fd_sc_hd__nand2_1_45/Y sky130_fd_sc_hd__o21ai_1_26/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1028 VDD VSS sky130_fd_sc_hd__fa_2_841/A sky130_fd_sc_hd__dfxtp_1_1038/CLK
+ sky130_fd_sc_hd__a21oi_1_311/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_37 VSS VDD sky130_fd_sc_hd__nand3_1_48/A sky130_fd_sc_hd__nand3_1_48/C
+ sky130_fd_sc_hd__nand3_1_48/B sky130_fd_sc_hd__o21ai_1_37/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_600 VDD VSS sky130_fd_sc_hd__and2_0_210/A sky130_fd_sc_hd__dfxtp_1_601/CLK
+ sky130_fd_sc_hd__fa_2_1020/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_260 sky130_fd_sc_hd__xor2_1_267/B sky130_fd_sc_hd__fa_2_1254/B
+ sky130_fd_sc_hd__xor2_1_260/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_1039 VDD VSS sky130_fd_sc_hd__fa_2_905/B sky130_fd_sc_hd__dfxtp_1_1050/CLK
+ sky130_fd_sc_hd__a21oi_1_306/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_611 VDD VSS sky130_fd_sc_hd__and2_0_227/A sky130_fd_sc_hd__dfxtp_1_611/CLK
+ sky130_fd_sc_hd__xor2_1_85/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_48 VSS VDD sky130_fd_sc_hd__o21ai_1_53/A2 sky130_fd_sc_hd__xnor2_1_50/Y
+ sky130_fd_sc_hd__a21oi_1_36/Y sky130_fd_sc_hd__o21ai_1_48/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_271 sky130_fd_sc_hd__fa_2_1242/A sky130_fd_sc_hd__fa_2_1243/B
+ sky130_fd_sc_hd__xor2_1_271/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_622 VDD VSS sky130_fd_sc_hd__ha_2_144/B sky130_fd_sc_hd__dfxtp_1_626/CLK
+ sky130_fd_sc_hd__o21a_1_3/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_282 sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1289/B
+ sky130_fd_sc_hd__xor2_1_282/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o21ai_1_59 VSS VDD sky130_fd_sc_hd__nand2_2_3/Y sky130_fd_sc_hd__xnor2_1_38/Y
+ sky130_fd_sc_hd__a21oi_1_45/Y sky130_fd_sc_hd__o21ai_1_59/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_633 VDD VSS sky130_fd_sc_hd__fa_2_997/A sky130_fd_sc_hd__clkinv_8_41/Y
+ sky130_fd_sc_hd__and2_0_287/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_293 sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1278/B
+ sky130_fd_sc_hd__xor2_1_293/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_644 VDD VSS sky130_fd_sc_hd__fa_2_1008/A sky130_fd_sc_hd__clkinv_8_44/Y
+ sky130_fd_sc_hd__mux2_2_16/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_655 VDD VSS sky130_fd_sc_hd__fa_2_972/A sky130_fd_sc_hd__clkinv_8_41/Y
+ sky130_fd_sc_hd__and2_0_282/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_666 VDD VSS sky130_fd_sc_hd__fa_2_983/A sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__mux2_2_21/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_677 VDD VSS sky130_fd_sc_hd__fa_2_1016/B sky130_fd_sc_hd__clkinv_8_59/Y
+ sky130_fd_sc_hd__and2_0_269/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_688 VDD VSS sky130_fd_sc_hd__fa_2_1027/A sky130_fd_sc_hd__clkinv_8_59/Y
+ sky130_fd_sc_hd__and2_0_291/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_699 VDD VSS sky130_fd_sc_hd__mux2_2_37/A0 sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__a22o_1_66/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_220 VSS VDD sky130_fd_sc_hd__buf_8_95/A sky130_fd_sc_hd__clkbuf_1_232/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_231 VSS VDD sky130_fd_sc_hd__clkbuf_1_232/A sky130_fd_sc_hd__buf_8_82/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_242 VSS VDD sky130_fd_sc_hd__clkbuf_1_242/X sky130_fd_sc_hd__clkinv_1_92/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_253 VSS VDD sky130_fd_sc_hd__buf_2_69/A sky130_fd_sc_hd__clkbuf_1_254/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_264 VSS VDD sky130_fd_sc_hd__clkbuf_1_264/X sky130_fd_sc_hd__nor3_1_17/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_275 VSS VDD sky130_fd_sc_hd__clkbuf_1_275/X sky130_fd_sc_hd__clkbuf_1_275/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_286 VSS VDD sky130_fd_sc_hd__clkbuf_1_286/X sky130_fd_sc_hd__clkbuf_1_286/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_297 VSS VDD sky130_fd_sc_hd__clkbuf_1_297/X sky130_fd_sc_hd__clkbuf_1_297/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_505 sky130_fd_sc_hd__fa_2_508/B sky130_fd_sc_hd__fa_2_505/SUM
+ sky130_fd_sc_hd__fa_2_505/A sky130_fd_sc_hd__fa_2_505/B sky130_fd_sc_hd__fa_2_505/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_516 sky130_fd_sc_hd__fa_2_518/CIN sky130_fd_sc_hd__fa_2_509/B
+ sky130_fd_sc_hd__fa_2_535/A sky130_fd_sc_hd__fa_2_566/A sky130_fd_sc_hd__fa_2_559/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_527 sky130_fd_sc_hd__fa_2_528/A sky130_fd_sc_hd__fa_2_520/A
+ sky130_fd_sc_hd__ha_2_119/B sky130_fd_sc_hd__fa_2_564/B sky130_fd_sc_hd__fa_2_427/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_538 sky130_fd_sc_hd__maj3_1_86/B sky130_fd_sc_hd__maj3_1_87/A
+ sky130_fd_sc_hd__fa_2_538/A sky130_fd_sc_hd__fa_2_538/B sky130_fd_sc_hd__fa_2_539/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_549 sky130_fd_sc_hd__fa_2_552/B sky130_fd_sc_hd__fa_2_549/SUM
+ sky130_fd_sc_hd__fa_2_549/A sky130_fd_sc_hd__fa_2_549/B sky130_fd_sc_hd__o22ai_1_37/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_4_3 VDD VSS sky130_fd_sc_hd__buf_4_3/X sky130_fd_sc_hd__buf_4_3/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__and2_0_240 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_240/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__o211ai_1_1/Y sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_251 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_251/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__xnor2_1_26/Y sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_262 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_262/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__fa_2_963/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_273 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_273/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__and2_0_273/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_284 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_284/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__fa_2_973/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_295 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_295/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_295/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__sdlclkp_2_1 sky130_fd_sc_hd__conb_1_7/LO sky130_fd_sc_hd__clkinv_8_100/Y
+ sky130_fd_sc_hd__dfxtp_1_111/CLK sky130_fd_sc_hd__a21oi_1_0/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__o21ai_1_230 VSS VDD sky130_fd_sc_hd__o21a_1_16/A2 sky130_fd_sc_hd__o21ai_1_230/A1
+ sky130_fd_sc_hd__a22oi_1_351/Y sky130_fd_sc_hd__o21ai_1_230/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_241 VSS VDD sky130_fd_sc_hd__a222oi_1_3/Y sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__nand2_1_330/Y sky130_fd_sc_hd__xor2_1_90/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_252 VSS VDD sky130_fd_sc_hd__a21oi_1_226/Y sky130_fd_sc_hd__nor2_1_126/A
+ sky130_fd_sc_hd__nand2b_1_16/Y sky130_fd_sc_hd__o21ai_1_252/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_70 sky130_fd_sc_hd__buf_2_42/A sky130_fd_sc_hd__dfxtp_1_262/Q
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_263 VSS VDD sky130_fd_sc_hd__nor2_1_127/A sky130_fd_sc_hd__a21oi_1_240/Y
+ sky130_fd_sc_hd__a21oi_1_228/Y sky130_fd_sc_hd__xor2_1_107/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_81 sky130_fd_sc_hd__clkbuf_4_81/X sky130_fd_sc_hd__clkbuf_4_81/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_274 VSS VDD sky130_fd_sc_hd__o21ai_1_274/A2 sky130_fd_sc_hd__o22ai_1_206/A1
+ sky130_fd_sc_hd__a22oi_1_369/Y sky130_fd_sc_hd__o21ai_1_274/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_92 sky130_fd_sc_hd__nand4_1_23/A sky130_fd_sc_hd__clkbuf_4_92/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_285 VSS VDD sky130_fd_sc_hd__nor2_1_156/B sky130_fd_sc_hd__o22ai_1_265/A2
+ sky130_fd_sc_hd__a22oi_1_371/Y sky130_fd_sc_hd__o21ai_1_285/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_296 VSS VDD sky130_fd_sc_hd__nor2_1_174/B sky130_fd_sc_hd__nor2_1_172/A
+ sky130_fd_sc_hd__a21oi_1_270/Y sky130_fd_sc_hd__o21ai_1_296/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2b_2_3 sky130_fd_sc_hd__o32ai_1_5/A1 sky130_fd_sc_hd__nor2b_2_3/A
+ sky130_fd_sc_hd__nor2b_2_3/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_2
Xsky130_fd_sc_hd__fa_2_1006 sky130_fd_sc_hd__fa_2_1007/CIN sky130_fd_sc_hd__mux2_2_20/A0
+ sky130_fd_sc_hd__fa_2_1006/A sky130_fd_sc_hd__xor2_1_70/X sky130_fd_sc_hd__fa_2_1006/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1017 sky130_fd_sc_hd__fa_2_1018/CIN sky130_fd_sc_hd__and2_0_270/A
+ sky130_fd_sc_hd__fa_2_1017/A sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_1017/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1028 sky130_fd_sc_hd__fa_2_1029/CIN sky130_fd_sc_hd__and2_0_292/A
+ sky130_fd_sc_hd__fa_2_1028/A sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_1028/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1039 sky130_fd_sc_hd__fa_2_1040/CIN sky130_fd_sc_hd__fa_2_1039/SUM
+ sky130_fd_sc_hd__fa_2_1039/A sky130_fd_sc_hd__nor2_1_51/A sky130_fd_sc_hd__fa_2_1039/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_15 sky130_fd_sc_hd__inv_2_15/A sky130_fd_sc_hd__inv_2_15/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_26 sky130_fd_sc_hd__inv_2_26/A sky130_fd_sc_hd__inv_2_26/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_430 VDD VSS sky130_fd_sc_hd__dfxtp_1_430/Q sky130_fd_sc_hd__dfxtp_1_433/CLK
+ sky130_fd_sc_hd__nand2_1_104/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_37 sky130_fd_sc_hd__inv_2_37/A sky130_fd_sc_hd__inv_2_37/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_441 VDD VSS sky130_fd_sc_hd__xor2_1_275/B sky130_fd_sc_hd__dfxtp_1_454/CLK
+ sky130_fd_sc_hd__nand2_1_82/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_48 sky130_fd_sc_hd__inv_2_48/A sky130_fd_sc_hd__inv_2_48/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_452 VDD VSS sky130_fd_sc_hd__dfxtp_1_998/D sky130_fd_sc_hd__dfxtp_1_452/CLK
+ sky130_fd_sc_hd__nand2_1_60/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_59 sky130_fd_sc_hd__inv_2_59/A sky130_fd_sc_hd__inv_2_59/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_463 VDD VSS sky130_fd_sc_hd__buf_2_7/A sky130_fd_sc_hd__dfxtp_1_463/CLK
+ sky130_fd_sc_hd__and2_0_156/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_474 VDD VSS sky130_fd_sc_hd__nor3_1_26/A sky130_fd_sc_hd__dfxtp_1_476/CLK
+ sky130_fd_sc_hd__and2_0_241/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_485 VDD VSS sky130_fd_sc_hd__nor2_1_39/A sky130_fd_sc_hd__dfxtp_1_488/CLK
+ sky130_fd_sc_hd__nor2b_1_56/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_2_5 sky130_fd_sc_hd__nand2_2_5/Y sky130_fd_sc_hd__nor2_2_11/A
+ sky130_fd_sc_hd__nor2_2_10/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__dfxtp_1_496 VDD VSS sky130_fd_sc_hd__nand2b_1_7/B sky130_fd_sc_hd__dfxtp_1_496/CLK
+ sky130_fd_sc_hd__nor2b_1_69/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2b_1_11 sky130_fd_sc_hd__xnor2_1_34/B sky130_fd_sc_hd__ha_2_185/B
+ sky130_fd_sc_hd__ha_2_185/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__fa_2_302 sky130_fd_sc_hd__fa_2_293/A sky130_fd_sc_hd__fa_2_300/A
+ sky130_fd_sc_hd__fa_2_425/B sky130_fd_sc_hd__fa_2_302/B sky130_fd_sc_hd__fa_2_302/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_313 sky130_fd_sc_hd__fa_2_306/A sky130_fd_sc_hd__fa_2_310/B
+ sky130_fd_sc_hd__fa_2_313/A sky130_fd_sc_hd__fa_2_313/B sky130_fd_sc_hd__fa_2_313/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_324 sky130_fd_sc_hd__maj3_1_80/B sky130_fd_sc_hd__maj3_1_81/A
+ sky130_fd_sc_hd__ha_2_113/B sky130_fd_sc_hd__ha_2_109/B sky130_fd_sc_hd__fa_2_360/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_335 sky130_fd_sc_hd__fa_2_337/B sky130_fd_sc_hd__fa_2_335/SUM
+ sky130_fd_sc_hd__ha_2_115/B sky130_fd_sc_hd__fa_2_417/A sky130_fd_sc_hd__fa_2_335/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_346 sky130_fd_sc_hd__fa_2_345/CIN sky130_fd_sc_hd__fa_2_346/SUM
+ sky130_fd_sc_hd__fa_2_404/A sky130_fd_sc_hd__ha_2_110/A sky130_fd_sc_hd__fa_2_417/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_357 sky130_fd_sc_hd__fa_2_362/B sky130_fd_sc_hd__fa_2_357/SUM
+ sky130_fd_sc_hd__fa_2_357/A sky130_fd_sc_hd__fa_2_357/B sky130_fd_sc_hd__fa_2_357/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_368 sky130_fd_sc_hd__fa_2_365/A sky130_fd_sc_hd__fa_2_368/SUM
+ sky130_fd_sc_hd__ha_2_115/B sky130_fd_sc_hd__ha_2_116/A sky130_fd_sc_hd__fa_2_360/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_379 sky130_fd_sc_hd__fa_2_381/CIN sky130_fd_sc_hd__fa_2_372/B
+ sky130_fd_sc_hd__fa_2_425/B sky130_fd_sc_hd__fa_2_424/B sky130_fd_sc_hd__fa_2_416/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_1_6 VDD VSS sky130_fd_sc_hd__and2_1_6/X sky130_fd_sc_hd__ha_2_58/A
+ sky130_fd_sc_hd__nor2_4_2/Y VDD VSS sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__diode_2_207 sig_frequency[7] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_218 sig_amplitude[3] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkinv_8_40 sky130_fd_sc_hd__clkinv_8_43/A sky130_fd_sc_hd__clkinv_8_40/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_40/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__diode_2_229 sig_amplitude[0] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkinv_8_51 sky130_fd_sc_hd__clkinv_8_51/Y sky130_fd_sc_hd__clkinv_8_70/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_51/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_62 sky130_fd_sc_hd__clkinv_8_62/Y sky130_fd_sc_hd__clkinv_8_62/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_62/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_73 sky130_fd_sc_hd__clkinv_8_73/Y sky130_fd_sc_hd__clkinv_8_74/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_73/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_84 sky130_fd_sc_hd__clkinv_8_84/Y sky130_fd_sc_hd__clkinv_8_84/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_84/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_95 sky130_fd_sc_hd__clkinv_8_96/A sky130_fd_sc_hd__clkinv_8_95/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_60 sky130_fd_sc_hd__buf_4_16/X sky130_fd_sc_hd__buf_12_60/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_71 sky130_fd_sc_hd__buf_4_27/X sky130_fd_sc_hd__buf_12_71/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_82 sky130_fd_sc_hd__buf_12_82/A sky130_fd_sc_hd__buf_12_82/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_93 sky130_fd_sc_hd__buf_12_93/A sky130_fd_sc_hd__buf_12_93/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_2_0 VDD VSS sky130_fd_sc_hd__buf_6_0/A sky130_fd_sc_hd__buf_2_0/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1370 VDD VSS sky130_fd_sc_hd__fa_2_1292/A sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__mux2_2_223/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1381 VDD VSS sky130_fd_sc_hd__fa_2_1320/A sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__mux2_2_250/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1392 VDD VSS sky130_fd_sc_hd__nor3_1_41/C sky130_fd_sc_hd__clkinv_8_78/Y
+ sky130_fd_sc_hd__o21bai_1_5/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_12_307 sky130_fd_sc_hd__buf_8_152/X sky130_fd_sc_hd__buf_12_360/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_318 sky130_fd_sc_hd__buf_4_89/X sky130_fd_sc_hd__buf_12_318/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_329 sky130_fd_sc_hd__buf_4_78/X sky130_fd_sc_hd__buf_12_329/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__fa_2_880 sky130_fd_sc_hd__fa_2_879/CIN sky130_fd_sc_hd__nand2_1_40/B
+ sky130_fd_sc_hd__ha_2_151/A sky130_fd_sc_hd__fa_2_880/B sky130_fd_sc_hd__fa_2_880/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_891 sky130_fd_sc_hd__fa_2_890/CIN sky130_fd_sc_hd__fa_2_891/SUM
+ sky130_fd_sc_hd__fa_2_891/A sky130_fd_sc_hd__fa_2_891/B sky130_fd_sc_hd__fa_2_891/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_0 load_en sky130_fd_sc_hd__inv_2_0/Y VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__nor3_2_2 sky130_fd_sc_hd__nor3_2_2/C sky130_fd_sc_hd__nor3_2_2/Y
+ sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__nor3_2_2/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_2
Xsky130_fd_sc_hd__clkinv_1_507 sky130_fd_sc_hd__o21ai_1_77/A1 sky130_fd_sc_hd__o21ai_1_84/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_507/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_518 sky130_fd_sc_hd__nor2_1_53/B sky130_fd_sc_hd__fa_2_1035/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_518/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_529 sky130_fd_sc_hd__nor2_1_67/A sky130_fd_sc_hd__nor2_1_68/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_529/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_10 sky130_fd_sc_hd__nor2_1_10/B sky130_fd_sc_hd__nor2_1_10/Y
+ sky130_fd_sc_hd__nor2_1_10/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_21 sky130_fd_sc_hd__nor2_1_21/B sky130_fd_sc_hd__nor2_1_21/Y
+ sky130_fd_sc_hd__nor2_1_21/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_32 sky130_fd_sc_hd__or4_1_2/D sky130_fd_sc_hd__xor2_1_28/B
+ sky130_fd_sc_hd__or4_1_2/C VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_43 sky130_fd_sc_hd__nor2_1_43/B sky130_fd_sc_hd__nor2_1_43/Y
+ sky130_fd_sc_hd__nor2_1_54/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_54 sky130_fd_sc_hd__nor2_1_54/B sky130_fd_sc_hd__nor2_1_54/Y
+ sky130_fd_sc_hd__nor2_1_54/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_65 sky130_fd_sc_hd__nor2_1_65/B sky130_fd_sc_hd__o21a_1_3/A1
+ sky130_fd_sc_hd__o21a_1_4/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_76 sky130_fd_sc_hd__nor2_1_80/Y sky130_fd_sc_hd__nor2_1_76/Y
+ sky130_fd_sc_hd__nor2_1_76/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_180 VSS VDD sky130_fd_sc_hd__mux2_2_180/A1 sky130_fd_sc_hd__mux2_2_180/A0
+ sky130_fd_sc_hd__nor2_8_1/A sky130_fd_sc_hd__mux2_2_180/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_87 sky130_fd_sc_hd__o21a_1_8/A2 sky130_fd_sc_hd__nor2_1_87/Y
+ sky130_fd_sc_hd__nor2_1_87/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_191 VSS VDD sky130_fd_sc_hd__mux2_2_191/A1 sky130_fd_sc_hd__mux2_2_191/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_191/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_98 sky130_fd_sc_hd__nor2_1_98/B sky130_fd_sc_hd__nor2_1_98/Y
+ sky130_fd_sc_hd__nor2_1_99/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_sram_2kbyte_1rw1r_32x512_8_6 sky130_fd_sc_hd__buf_4_32/X sky130_fd_sc_hd__buf_8_63/X
+ sky130_fd_sc_hd__buf_2_35/A sky130_fd_sc_hd__buf_4_34/X sky130_fd_sc_hd__inv_12_0/Y
+ sky130_fd_sc_hd__clkbuf_4_63/X sky130_fd_sc_hd__buf_2_36/A sky130_fd_sc_hd__buf_4_36/X
+ sky130_fd_sc_hd__clkbuf_1_198/X sky130_fd_sc_hd__clkbuf_1_201/X sky130_fd_sc_hd__buf_2_38/A
+ sky130_fd_sc_hd__buf_2_39/A sky130_fd_sc_hd__clkbuf_4_95/X sky130_fd_sc_hd__buf_2_40/A
+ sky130_fd_sc_hd__buf_2_41/A sky130_fd_sc_hd__buf_2_42/A sky130_fd_sc_hd__buf_4_32/X
+ sky130_fd_sc_hd__buf_8_63/X sky130_fd_sc_hd__buf_2_35/A sky130_fd_sc_hd__buf_4_34/X
+ sky130_fd_sc_hd__inv_12_0/Y sky130_fd_sc_hd__clkbuf_4_63/X sky130_fd_sc_hd__buf_2_36/A
+ sky130_fd_sc_hd__buf_4_36/X sky130_fd_sc_hd__buf_2_116/X sky130_fd_sc_hd__buf_2_117/X
+ sky130_fd_sc_hd__buf_2_38/A sky130_fd_sc_hd__buf_2_39/A sky130_fd_sc_hd__clkbuf_4_95/X
+ sky130_fd_sc_hd__buf_2_40/A sky130_fd_sc_hd__buf_2_41/A sky130_fd_sc_hd__buf_2_42/A
+ sky130_fd_sc_hd__buf_12_129/X sky130_fd_sc_hd__buf_12_238/X sky130_fd_sc_hd__buf_12_205/X
+ sky130_fd_sc_hd__buf_12_202/X sky130_fd_sc_hd__buf_12_187/X sky130_fd_sc_hd__buf_12_228/X
+ sky130_fd_sc_hd__buf_12_188/X sky130_fd_sc_hd__buf_12_169/X sky130_fd_sc_hd__buf_12_224/X
+ sky130_fd_sc_hd__buf_12_146/X sky130_fd_sc_hd__buf_12_148/X sky130_fd_sc_hd__buf_12_242/X
+ sky130_fd_sc_hd__buf_12_209/X sky130_fd_sc_hd__buf_12_252/X sky130_fd_sc_hd__buf_12_250/X
+ sky130_fd_sc_hd__buf_12_153/X sky130_fd_sc_hd__buf_12_239/X sky130_fd_sc_hd__buf_12_247/X
+ sky130_fd_sc_hd__clkbuf_1_173/X sky130_fd_sc_hd__clkbuf_1_190/X sky130_fd_sc_hd__clkbuf_1_173/X
+ sky130_fd_sc_hd__clkinv_8_124/Y sky130_fd_sc_hd__clkinv_8_13/Y sky130_fd_sc_hd__buf_12_191/X
+ sky130_fd_sc_hd__buf_12_208/X sky130_fd_sc_hd__buf_12_181/X sky130_fd_sc_hd__buf_12_182/X
+ sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[0] sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[1]
+ sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[2] sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[3]
+ sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[4] sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[5]
+ sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[6] sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[7]
+ sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[8] sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[9]
+ sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[10] sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[11]
+ sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[12] sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[13]
+ sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[14] sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[15]
+ sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[16] sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[17]
+ sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[18] sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[19]
+ sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[20] sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[21]
+ sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[22] sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[23]
+ sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[24] sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[25]
+ sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[26] sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[27]
+ sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[28] sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[29]
+ sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[30] sky130_sram_2kbyte_1rw1r_32x512_8_6/dout0[31]
+ sky130_fd_sc_hd__clkbuf_1_258/A sky130_fd_sc_hd__clkbuf_4_75/A sky130_fd_sc_hd__clkbuf_4_76/A
+ sky130_fd_sc_hd__clkbuf_4_77/A sky130_fd_sc_hd__clkbuf_4_78/A sky130_fd_sc_hd__clkbuf_4_79/A
+ sky130_fd_sc_hd__clkbuf_4_80/A sky130_fd_sc_hd__clkbuf_4_81/A sky130_fd_sc_hd__clkbuf_4_82/A
+ sky130_fd_sc_hd__clkbuf_4_83/A sky130_fd_sc_hd__clkbuf_4_84/A sky130_fd_sc_hd__clkbuf_4_85/A
+ sky130_fd_sc_hd__clkbuf_4_86/A sky130_fd_sc_hd__clkbuf_4_87/A sky130_fd_sc_hd__clkbuf_4_88/A
+ sky130_fd_sc_hd__clkbuf_4_89/A sky130_fd_sc_hd__a22oi_1_146/B2 sky130_fd_sc_hd__a22oi_1_142/B2
+ sky130_fd_sc_hd__a22oi_1_138/B2 sky130_fd_sc_hd__a22oi_1_134/B2 sky130_fd_sc_hd__a22oi_1_130/B2
+ sky130_fd_sc_hd__a22oi_1_127/B2 sky130_fd_sc_hd__a22oi_1_123/B2 sky130_fd_sc_hd__a22oi_1_119/B2
+ sky130_fd_sc_hd__a22oi_1_115/B2 sky130_fd_sc_hd__a22oi_1_111/B2 sky130_fd_sc_hd__a22oi_1_107/B2
+ sky130_fd_sc_hd__clkbuf_1_260/A sky130_fd_sc_hd__a22oi_1_99/B2 sky130_fd_sc_hd__a22oi_1_95/B2
+ sky130_fd_sc_hd__a22oi_1_91/B2 sky130_fd_sc_hd__a22oi_1_87/B2 VDD VSS sky130_sram_2kbyte_1rw1r_32x512_8
Xsky130_fd_sc_hd__a21oi_1_404 sky130_fd_sc_hd__a21oi_1_404/A1 sky130_fd_sc_hd__nor2_1_262/Y
+ sky130_fd_sc_hd__a21oi_1_404/Y sky130_fd_sc_hd__nor2b_2_4/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_415 sky130_fd_sc_hd__nor3_1_40/A sky130_fd_sc_hd__o22ai_1_374/Y
+ sky130_fd_sc_hd__a21oi_1_415/Y sky130_fd_sc_hd__fa_2_1252/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_426 sky130_fd_sc_hd__o21a_1_61/B1 sky130_fd_sc_hd__nor2_1_274/Y
+ sky130_fd_sc_hd__a21oi_1_426/Y sky130_fd_sc_hd__nor2_1_274/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_437 sky130_fd_sc_hd__nor3_1_41/B sky130_fd_sc_hd__nor2b_1_126/Y
+ sky130_fd_sc_hd__a21oi_1_437/Y sky130_fd_sc_hd__nor2b_2_5/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_448 sky130_fd_sc_hd__fa_2_1289/A sky130_fd_sc_hd__o22ai_1_414/Y
+ sky130_fd_sc_hd__a21oi_1_448/Y sky130_fd_sc_hd__a22oi_1_400/B1 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_459 sky130_fd_sc_hd__nor3_1_41/A sky130_fd_sc_hd__o22ai_1_422/Y
+ sky130_fd_sc_hd__a21oi_1_459/Y sky130_fd_sc_hd__fa_2_1280/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_8_106 sky130_fd_sc_hd__clkinv_8_107/A sky130_fd_sc_hd__clkinv_8_91/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_106/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_117 sky130_fd_sc_hd__clkinv_4_60/A sky130_fd_sc_hd__clkinv_8_71/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_117/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_128 sky130_fd_sc_hd__clkinv_4_70/A sky130_fd_sc_hd__clkinv_8_128/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_139 sky130_fd_sc_hd__clkinv_4_78/A sky130_fd_sc_hd__clkinv_4_76/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_139/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__o21a_1_8 sky130_fd_sc_hd__o21a_1_8/X sky130_fd_sc_hd__o21a_1_8/A1
+ sky130_fd_sc_hd__o21a_1_8/B1 sky130_fd_sc_hd__o21a_1_8/A2 VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__maj3_1_140 sky130_fd_sc_hd__maj3_1_141/X sky130_fd_sc_hd__maj3_1_140/X
+ sky130_fd_sc_hd__maj3_1_140/B sky130_fd_sc_hd__maj3_1_140/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_420 sky130_fd_sc_hd__nor2_1_208/B sky130_fd_sc_hd__nand2_1_420/B
+ sky130_fd_sc_hd__nor2_1_209/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_151 sky130_fd_sc_hd__maj3_1_152/X sky130_fd_sc_hd__maj3_1_151/X
+ sky130_fd_sc_hd__maj3_1_151/B sky130_fd_sc_hd__maj3_1_151/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_431 sky130_fd_sc_hd__nand2_1_431/Y sky130_fd_sc_hd__nor2b_2_3/Y
+ sky130_fd_sc_hd__o21ai_1_355/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_442 sky130_fd_sc_hd__o21a_1_42/A1 sky130_fd_sc_hd__nor2_2_16/B
+ sky130_fd_sc_hd__nor2_4_16/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_453 sky130_fd_sc_hd__xnor2_1_98/B sky130_fd_sc_hd__fa_2_1258/A
+ sky130_fd_sc_hd__o21a_1_49/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_464 sky130_fd_sc_hd__nand2_1_464/Y sky130_fd_sc_hd__nor2_1_248/B
+ sky130_fd_sc_hd__nor2_1_245/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_475 sky130_fd_sc_hd__nor2_1_254/B sky130_fd_sc_hd__nand2_1_475/B
+ sky130_fd_sc_hd__nor2_1_255/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_486 sky130_fd_sc_hd__nand2_1_486/Y sky130_fd_sc_hd__xor2_1_253/A
+ sky130_fd_sc_hd__nor2_1_267/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_497 sky130_fd_sc_hd__nor2_1_309/A sky130_fd_sc_hd__nand2_1_497/B
+ sky130_fd_sc_hd__o32ai_1_11/B2 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_11 sky130_fd_sc_hd__ha_2_20/SUM sky130_fd_sc_hd__nor2b_1_11/Y
+ sky130_fd_sc_hd__or2_0_1/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_22 sky130_fd_sc_hd__ha_2_41/SUM sky130_fd_sc_hd__nor2b_1_22/Y
+ sky130_fd_sc_hd__or2_1_0/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_33 sky130_fd_sc_hd__ha_2_64/SUM sky130_fd_sc_hd__nor2b_1_33/Y
+ sky130_fd_sc_hd__or2_0_2/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1000 sky130_fd_sc_hd__o21ai_1_414/A1 sky130_fd_sc_hd__o21ai_1_416/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1000/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_44 sky130_fd_sc_hd__ha_2_87/SUM sky130_fd_sc_hd__nor2b_1_44/Y
+ sky130_fd_sc_hd__or2_0_3/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1011 sky130_fd_sc_hd__nor2_1_235/B sky130_fd_sc_hd__fa_2_1257/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1011/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_55 sky130_fd_sc_hd__xnor2_1_12/B sky130_fd_sc_hd__nor2_1_10/A
+ sky130_fd_sc_hd__ha_2_151/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1022 sky130_fd_sc_hd__nor2_1_240/B sky130_fd_sc_hd__fa_2_1248/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1022/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_66 sky130_fd_sc_hd__o21ai_1_39/A1 sky130_fd_sc_hd__nor2b_1_66/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1033 sky130_fd_sc_hd__nand2_1_543/B sky130_fd_sc_hd__nor2_1_309/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1033/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_77 sky130_fd_sc_hd__dfxtp_1_501/Q sky130_fd_sc_hd__nor2b_1_77/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1044 sky130_fd_sc_hd__o32ai_1_10/A2 sky130_fd_sc_hd__fa_2_1293/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1044/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1055 sky130_fd_sc_hd__o22ai_1_405/A1 sky130_fd_sc_hd__fa_2_26/SUM
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_88 sky130_fd_sc_hd__fa_2_964/A sky130_fd_sc_hd__o31ai_1_4/A3
+ sky130_fd_sc_hd__nor2b_1_88/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1066 sky130_fd_sc_hd__nand2_1_524/B sky130_fd_sc_hd__fa_2_4/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1066/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_99 sky130_fd_sc_hd__a32o_1_1/B2 sky130_fd_sc_hd__nor2b_1_99/Y
+ sky130_fd_sc_hd__buf_2_262/X VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__xnor2_1_7 VSS VDD sky130_fd_sc_hd__xnor2_1_7/B sky130_fd_sc_hd__xnor2_1_7/Y
+ sky130_fd_sc_hd__xnor2_1_7/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_1077 sky130_fd_sc_hd__o22ai_1_418/A1 sky130_fd_sc_hd__fa_2_1285/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1077/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1088 sky130_fd_sc_hd__nor2_1_271/B sky130_fd_sc_hd__fa_2_1286/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1088/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1099 sky130_fd_sc_hd__nand2_1_497/B sky130_fd_sc_hd__nor2b_2_5/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1099/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_260 VDD VSS sky130_fd_sc_hd__dfxtp_1_260/Q sky130_fd_sc_hd__dfxtp_1_262/CLK
+ sky130_fd_sc_hd__and2_0_223/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_271 VDD VSS sky130_fd_sc_hd__dfxtp_1_271/Q sky130_fd_sc_hd__dfxtp_1_463/CLK
+ sky130_fd_sc_hd__and2_0_213/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_282 VDD VSS sky130_fd_sc_hd__dfxtp_1_282/Q sky130_fd_sc_hd__dfxtp_1_282/CLK
+ sky130_fd_sc_hd__nor3_1_26/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_293 VDD VSS sky130_fd_sc_hd__a22o_1_54/A1 sky130_fd_sc_hd__clkinv_4_31/Y
+ sky130_fd_sc_hd__nand2_1_123/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o22ai_1_2 sky130_fd_sc_hd__fa_2_87/A sky130_fd_sc_hd__fa_2_49/B
+ sky130_fd_sc_hd__o22ai_1_2/Y sky130_fd_sc_hd__ha_2_95/A sky130_fd_sc_hd__fa_2_66/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_110 sky130_fd_sc_hd__fa_2_113/B sky130_fd_sc_hd__fa_2_110/SUM
+ sky130_fd_sc_hd__fa_2_110/A sky130_fd_sc_hd__fa_2_110/B sky130_fd_sc_hd__fa_2_110/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_121 sky130_fd_sc_hd__maj3_1_4/B sky130_fd_sc_hd__maj3_1_5/A
+ sky130_fd_sc_hd__fa_2_121/A sky130_fd_sc_hd__fa_2_121/B sky130_fd_sc_hd__fa_2_122/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_132 sky130_fd_sc_hd__fa_2_130/B sky130_fd_sc_hd__fa_2_127/B
+ sky130_fd_sc_hd__fa_2_81/B sky130_fd_sc_hd__fa_2_91/A sky130_fd_sc_hd__fa_2_80/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_143 sky130_fd_sc_hd__fa_2_142/CIN sky130_fd_sc_hd__fa_2_143/SUM
+ sky130_fd_sc_hd__fa_2_143/A sky130_fd_sc_hd__fa_2_143/B sky130_fd_sc_hd__fa_2_143/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_154 sky130_fd_sc_hd__fa_2_153/B sky130_fd_sc_hd__fa_2_154/SUM
+ sky130_fd_sc_hd__ha_2_97/A sky130_fd_sc_hd__ha_2_104/B sky130_fd_sc_hd__fa_2_277/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_165 sky130_fd_sc_hd__fa_2_162/CIN sky130_fd_sc_hd__fa_2_167/CIN
+ sky130_fd_sc_hd__fa_2_274/A sky130_fd_sc_hd__fa_2_250/A sky130_fd_sc_hd__fa_2_165/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_176 sky130_fd_sc_hd__maj3_1_51/B sky130_fd_sc_hd__maj3_1_52/A
+ sky130_fd_sc_hd__fa_2_242/A sky130_fd_sc_hd__fa_2_176/B sky130_fd_sc_hd__fa_2_177/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_187 sky130_fd_sc_hd__fa_2_189/B sky130_fd_sc_hd__fa_2_187/SUM
+ sky130_fd_sc_hd__fa_2_281/A sky130_fd_sc_hd__fa_2_187/B sky130_fd_sc_hd__fa_2_187/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_198 sky130_fd_sc_hd__fa_2_202/CIN sky130_fd_sc_hd__fa_2_196/B
+ sky130_fd_sc_hd__fa_2_198/A sky130_fd_sc_hd__fa_2_198/B sky130_fd_sc_hd__fa_2_207/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o22ai_1_20 sky130_fd_sc_hd__fa_2_144/B sky130_fd_sc_hd__fa_2_266/B
+ sky130_fd_sc_hd__fa_2_271/A sky130_fd_sc_hd__ha_2_93/A sky130_fd_sc_hd__ha_2_97/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_31 sky130_fd_sc_hd__fa_2_554/A sky130_fd_sc_hd__fa_2_427/B
+ sky130_fd_sc_hd__xnor2_1_3/B sky130_fd_sc_hd__ha_2_125/A sky130_fd_sc_hd__ha_2_117/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_42 sky130_fd_sc_hd__fa_2_673/B sky130_fd_sc_hd__ha_2_132/B
+ sky130_fd_sc_hd__o22ai_1_42/Y sky130_fd_sc_hd__fa_2_672/A sky130_fd_sc_hd__ha_2_130/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_160 VDD VSS sky130_fd_sc_hd__buf_2_160/X sky130_fd_sc_hd__a22o_2_9/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_53 sky130_fd_sc_hd__fa_2_834/A sky130_fd_sc_hd__fa_2_823/B
+ sky130_fd_sc_hd__fa_2_783/A sky130_fd_sc_hd__ha_2_144/B sky130_fd_sc_hd__fa_2_826/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_171 VDD VSS sky130_fd_sc_hd__buf_2_171/X sky130_fd_sc_hd__buf_2_171/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_64 sky130_fd_sc_hd__o22ai_1_88/B1 sky130_fd_sc_hd__nand2_2_3/Y
+ sky130_fd_sc_hd__o22ai_1_64/Y sky130_fd_sc_hd__xnor2_1_39/Y sky130_fd_sc_hd__o22ai_1_78/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_182 VDD VSS sky130_fd_sc_hd__buf_2_182/X sky130_fd_sc_hd__buf_2_182/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_75 sky130_fd_sc_hd__o22ai_1_89/A1 sky130_fd_sc_hd__o22ai_1_88/B1
+ sky130_fd_sc_hd__o22ai_1_75/Y sky130_fd_sc_hd__xnor2_1_33/Y sky130_fd_sc_hd__o22ai_1_75/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_193 VDD VSS sky130_fd_sc_hd__buf_2_193/X sky130_fd_sc_hd__buf_2_193/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_86 sky130_fd_sc_hd__o22ai_1_89/A1 sky130_fd_sc_hd__o22ai_1_88/B1
+ sky130_fd_sc_hd__o22ai_1_86/Y sky130_fd_sc_hd__xnor2_1_55/Y sky130_fd_sc_hd__o22ai_1_86/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_97 sky130_fd_sc_hd__a21oi_1_93/Y sky130_fd_sc_hd__a21oi_1_92/Y
+ sky130_fd_sc_hd__o22ai_1_97/Y sky130_fd_sc_hd__nor2_2_9/B sky130_fd_sc_hd__nor2_1_76/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_4_11 VDD VSS sky130_fd_sc_hd__buf_4_11/X sky130_fd_sc_hd__buf_4_11/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_22 VDD VSS sky130_fd_sc_hd__buf_4_22/X sky130_fd_sc_hd__buf_8_28/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_33 VDD VSS sky130_fd_sc_hd__buf_4_33/X sky130_fd_sc_hd__buf_4_33/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_44 VDD VSS sky130_fd_sc_hd__buf_4_44/X sky130_fd_sc_hd__buf_4_44/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_55 VDD VSS sky130_fd_sc_hd__buf_4_55/X sky130_fd_sc_hd__buf_4_55/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_66 VDD VSS sky130_fd_sc_hd__buf_4_66/X sky130_fd_sc_hd__buf_4_66/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_77 VDD VSS sky130_fd_sc_hd__buf_4_77/X sky130_fd_sc_hd__buf_4_77/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_88 VDD VSS sky130_fd_sc_hd__buf_4_88/X sky130_fd_sc_hd__buf_4_88/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_99 VDD VSS sky130_fd_sc_hd__buf_4_99/X sky130_fd_sc_hd__buf_4_99/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_12_104 sky130_fd_sc_hd__buf_12_12/X sky130_fd_sc_hd__buf_12_104/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_115 sky130_fd_sc_hd__buf_12_94/X sky130_fd_sc_hd__buf_12_115/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_126 sky130_fd_sc_hd__buf_12_126/A sky130_fd_sc_hd__buf_12_126/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_137 sky130_fd_sc_hd__buf_12_137/A sky130_fd_sc_hd__buf_12_234/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_60 VSS VDD sky130_fd_sc_hd__clkbuf_1_60/X sky130_fd_sc_hd__clkbuf_1_60/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_148 sky130_fd_sc_hd__buf_12_148/A sky130_fd_sc_hd__buf_12_148/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_71 VSS VDD sky130_fd_sc_hd__clkbuf_1_71/X sky130_fd_sc_hd__nand3_1_23/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_159 sky130_fd_sc_hd__buf_8_72/X sky130_fd_sc_hd__buf_12_209/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_82 VSS VDD sky130_fd_sc_hd__nand4_1_5/A sky130_fd_sc_hd__a22oi_2_6/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_93 VSS VDD sky130_fd_sc_hd__buf_8_45/A sky130_fd_sc_hd__inv_2_3/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_4_7 sky130_fd_sc_hd__clkbuf_4_7/X sky130_fd_sc_hd__buf_2_10/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_1_304 sky130_fd_sc_hd__fa_2_273/A sky130_fd_sc_hd__ha_2_99/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_304/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_315 sky130_fd_sc_hd__fa_2_401/A sky130_fd_sc_hd__fa_2_393/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_315/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_326 sky130_fd_sc_hd__fa_2_531/B sky130_fd_sc_hd__ha_2_124/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_326/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_337 sky130_fd_sc_hd__fa_2_559/B sky130_fd_sc_hd__ha_2_169/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_337/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_348 sky130_fd_sc_hd__ha_2_126/A sky130_fd_sc_hd__fa_2_677/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_348/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_359 sky130_fd_sc_hd__fa_2_834/B sky130_fd_sc_hd__fa_2_835/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_359/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_201 sky130_fd_sc_hd__clkinv_1_622/Y sky130_fd_sc_hd__o22ai_1_172/Y
+ sky130_fd_sc_hd__a21oi_1_201/Y sky130_fd_sc_hd__nand2_1_331/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_212 sky130_fd_sc_hd__a21o_2_5/A2 sky130_fd_sc_hd__o22ai_1_192/Y
+ sky130_fd_sc_hd__a21oi_1_212/Y sky130_fd_sc_hd__fa_2_1048/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_223 sky130_fd_sc_hd__a211o_1_9/A1 sky130_fd_sc_hd__o22ai_1_198/Y
+ sky130_fd_sc_hd__a21oi_1_223/Y sky130_fd_sc_hd__nand2_1_332/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_234 sky130_fd_sc_hd__a21o_2_5/A2 sky130_fd_sc_hd__o21ai_1_269/Y
+ sky130_fd_sc_hd__a21oi_1_234/Y sky130_fd_sc_hd__fa_2_1084/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_245 sky130_fd_sc_hd__nor2_1_146/A sky130_fd_sc_hd__o21a_1_21/A1
+ sky130_fd_sc_hd__dfxtp_1_899/D sky130_fd_sc_hd__nor2_1_146/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_2_30 sky130_fd_sc_hd__buf_2_165/X sky130_fd_sc_hd__a22oi_2_30/A2
+ sky130_fd_sc_hd__nor2_4_7/Y sky130_fd_sc_hd__a22oi_2_30/B2 sky130_fd_sc_hd__nand4_1_63/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__a21oi_1_256 sky130_fd_sc_hd__nor2_1_157/A sky130_fd_sc_hd__nor2_1_157/Y
+ sky130_fd_sc_hd__dfxtp_1_879/D sky130_fd_sc_hd__nor2_1_157/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_267 sky130_fd_sc_hd__clkinv_1_819/Y sky130_fd_sc_hd__nor2_1_173/Y
+ sky130_fd_sc_hd__a21oi_1_267/Y sky130_fd_sc_hd__nor2b_1_104/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_278 sky130_fd_sc_hd__fa_2_1128/A sky130_fd_sc_hd__o22ai_1_248/Y
+ sky130_fd_sc_hd__a21oi_1_278/Y sky130_fd_sc_hd__nor3_1_38/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_289 sky130_fd_sc_hd__nand2_1_387/B sky130_fd_sc_hd__o22ai_1_255/Y
+ sky130_fd_sc_hd__a21oi_1_289/Y sky130_fd_sc_hd__o21ai_1_329/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_4_7 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_4_7/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_7/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_8_208 sky130_fd_sc_hd__buf_8_208/A sky130_fd_sc_hd__buf_8_208/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_219 sky130_fd_sc_hd__buf_8_219/A sky130_fd_sc_hd__buf_6_79/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nand2_1_250 sky130_fd_sc_hd__nand2_1_250/Y sky130_fd_sc_hd__nor2_1_49/B
+ sky130_fd_sc_hd__nor2_1_49/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_261 sky130_fd_sc_hd__o211ai_1_4/C1 sky130_fd_sc_hd__a211o_1_8/A2
+ sky130_fd_sc_hd__nand2_1_261/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_860 sky130_fd_sc_hd__nor2_4_15/B sky130_fd_sc_hd__nor2_4_14/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_860/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_272 sky130_fd_sc_hd__nand2_1_272/Y sky130_fd_sc_hd__a211o_1_3/A1
+ sky130_fd_sc_hd__a211o_1_5/A2 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_871 sky130_fd_sc_hd__nor2_1_188/A sky130_fd_sc_hd__nor2_1_189/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_871/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_283 sky130_fd_sc_hd__nor2_1_127/A sky130_fd_sc_hd__nand2_1_339/A
+ sky130_fd_sc_hd__nand2_2_6/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_882 sky130_fd_sc_hd__o22ai_1_285/A1 sky130_fd_sc_hd__nor2_1_210/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_882/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_294 sky130_fd_sc_hd__nand2_1_294/Y sky130_fd_sc_hd__nor2_1_112/B
+ sky130_fd_sc_hd__fa_2_1120/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_893 sky130_fd_sc_hd__nor2_1_205/B sky130_fd_sc_hd__xor2_1_185/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_893/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__mux2_2_0 VSS VDD sky130_fd_sc_hd__mux2_2_0/A1 sky130_fd_sc_hd__xor2_1_58/X
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_0/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__a21boi_0_0 sky130_fd_sc_hd__a22oi_1_336/Y sky130_fd_sc_hd__o21a_1_8/B1
+ sky130_fd_sc_hd__nor2_4_9/B sky130_fd_sc_hd__nor2_2_8/Y VSS VDD VDD VSS sky130_fd_sc_hd__a21boi_0
Xsky130_fd_sc_hd__fa_2_8 sky130_fd_sc_hd__fa_2_1/CIN sky130_fd_sc_hd__fa_2_8/SUM sky130_fd_sc_hd__fa_2_8/A
+ sky130_fd_sc_hd__fa_2_8/B sky130_fd_sc_hd__fa_2_8/CIN VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a211o_1_14 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_130/A sky130_fd_sc_hd__nand2_1_333/B
+ sky130_fd_sc_hd__o22ai_1_170/Y sky130_fd_sc_hd__o21ai_1_231/Y sky130_fd_sc_hd__nor2_1_127/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__a211o_1_25 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_272/A sky130_fd_sc_hd__nor2b_1_119/Y
+ sky130_fd_sc_hd__o22ai_1_354/Y sky130_fd_sc_hd__o21ai_1_402/Y sky130_fd_sc_hd__o22ai_1_353/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__clkinv_1_101 sky130_fd_sc_hd__inv_2_65/A sky130_fd_sc_hd__buf_8_88/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_101/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_112 sky130_fd_sc_hd__inv_16_3/A sky130_fd_sc_hd__clkinv_1_112/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_112/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_123 sky130_fd_sc_hd__nor3_1_16/C sky130_fd_sc_hd__nor3_2_6/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_123/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_134 sky130_fd_sc_hd__clkinv_2_12/A sky130_fd_sc_hd__clkinv_1_134/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_134/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_145 sky130_fd_sc_hd__clkinv_1_146/A sky130_fd_sc_hd__inv_2_96/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_145/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_156 sky130_fd_sc_hd__inv_2_87/A sky130_fd_sc_hd__clkinv_1_156/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_156/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_167 sky130_fd_sc_hd__inv_2_98/A sky130_fd_sc_hd__clkinv_1_167/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_167/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_178 sky130_fd_sc_hd__bufinv_8_7/A sky130_fd_sc_hd__buf_8_161/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_178/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_14 sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__ha_2_67/A
+ sky130_fd_sc_hd__a22o_1_14/X sky130_fd_sc_hd__dfxtp_1_4/Q sky130_fd_sc_hd__a22o_2_3/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_1_189 sky130_fd_sc_hd__nor3_1_21/C sky130_fd_sc_hd__nor3_2_9/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_189/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_25 sky130_fd_sc_hd__nor2_4_4/Y sky130_fd_sc_hd__ha_2_76/A
+ sky130_fd_sc_hd__a22o_1_25/X sky130_fd_sc_hd__a22o_1_25/B2 sky130_fd_sc_hd__a22o_2_6/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_36 sky130_fd_sc_hd__nor2_1_29/Y sky130_fd_sc_hd__nor3_1_31/Y
+ sky130_fd_sc_hd__a22o_1_36/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__a22o_1_36/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_47 sky130_fd_sc_hd__a22o_1_47/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_47/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__fa_2_953/SUM
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__o21ai_1_1 VSS VDD sky130_fd_sc_hd__o21ai_1_1/A2 sky130_fd_sc_hd__or2_0_0/A
+ sky130_fd_sc_hd__inv_8_1/Y sky130_fd_sc_hd__o21ai_1_1/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a22o_1_58 sky130_fd_sc_hd__a22o_1_58/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_58/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__nor4_1_9/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_69 sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__fa_2_995/A
+ sky130_fd_sc_hd__a22o_1_69/X sky130_fd_sc_hd__fa_2_997/A sky130_fd_sc_hd__nor2_2_8/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__bufbuf_16_0 sky130_fd_sc_hd__inv_2_9/Y sky130_fd_sc_hd__buf_6_13/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__nand4_1_8 sky130_fd_sc_hd__nand4_1_8/C sky130_fd_sc_hd__nand4_1_8/B
+ sky130_fd_sc_hd__nand4_1_8/Y sky130_fd_sc_hd__nand4_1_8/D sky130_fd_sc_hd__nand4_1_8/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nor2_1_250 sky130_fd_sc_hd__nor2_1_250/B sky130_fd_sc_hd__nor2_1_250/Y
+ sky130_fd_sc_hd__nor2_1_267/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_2_4 sky130_fd_sc_hd__clkinv_2_4/Y sky130_fd_sc_hd__ha_2_34/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_4/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__nor2_1_261 sky130_fd_sc_hd__o21a_1_55/A1 sky130_fd_sc_hd__nor2_1_261/Y
+ sky130_fd_sc_hd__nor2_1_261/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_272 sky130_fd_sc_hd__nor2_1_272/B sky130_fd_sc_hd__o21a_1_59/A1
+ sky130_fd_sc_hd__o21a_1_60/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_283 sky130_fd_sc_hd__nor2_1_283/B sky130_fd_sc_hd__o21a_1_67/A1
+ sky130_fd_sc_hd__nor2_1_283/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_294 sky130_fd_sc_hd__nor2_1_294/B sky130_fd_sc_hd__nor2_1_294/Y
+ sky130_fd_sc_hd__fa_2_7/SUM VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_490 sky130_fd_sc_hd__buf_12_490/A sky130_fd_sc_hd__buf_12_490/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_360 sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__nor2_4_13/Y
+ sky130_fd_sc_hd__fa_2_1089/A sky130_fd_sc_hd__fa_2_1090/A sky130_fd_sc_hd__a22oi_1_360/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_371 sky130_fd_sc_hd__clkinv_1_779/Y sky130_fd_sc_hd__nor3_1_38/B
+ sky130_fd_sc_hd__fa_2_1146/A sky130_fd_sc_hd__fa_2_1147/A sky130_fd_sc_hd__a22oi_1_371/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_382 sky130_fd_sc_hd__nor3_1_39/B sky130_fd_sc_hd__fa_2_1190/A
+ sky130_fd_sc_hd__xor2_1_209/A sky130_fd_sc_hd__clkinv_1_861/Y sky130_fd_sc_hd__a22oi_1_382/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_393 sky130_fd_sc_hd__nor2_1_265/Y sky130_fd_sc_hd__nor2_1_267/Y
+ sky130_fd_sc_hd__fa_2_1251/A sky130_fd_sc_hd__fa_2_1247/A sky130_fd_sc_hd__a22oi_1_393/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nand2_1_15 sky130_fd_sc_hd__nand3_1_15/A sky130_fd_sc_hd__nand2_1_9/A
+ sky130_fd_sc_hd__nand4_1_64/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_26 sky130_fd_sc_hd__or2_0_3/B sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__or2_1_1/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_37 sky130_fd_sc_hd__nand2_1_37/Y sky130_fd_sc_hd__xnor2_1_11/Y
+ sky130_fd_sc_hd__a21oi_2_0/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_690 sky130_fd_sc_hd__nor2_1_117/A sky130_fd_sc_hd__nor2_1_118/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_690/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_48 sky130_fd_sc_hd__nand2_1_48/Y sky130_fd_sc_hd__nor2_1_12/B
+ sky130_fd_sc_hd__xor2_1_19/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_59 sky130_fd_sc_hd__nand2_1_59/Y sky130_fd_sc_hd__nand2_1_4/B
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2_8_1 sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__nor2_8_1/A
+ sky130_fd_sc_hd__nor2_8_1/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_8
Xsky130_fd_sc_hd__xnor2_1_90 VSS VDD sky130_fd_sc_hd__o21a_1_9/B1 sky130_fd_sc_hd__xnor2_1_90/Y
+ sky130_fd_sc_hd__fa_2_1067/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__dfxtp_1_804 VDD VSS sky130_fd_sc_hd__fa_2_1056/A sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__mux2_2_65/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_815 VDD VSS sky130_fd_sc_hd__fa_2_1067/A sky130_fd_sc_hd__clkinv_4_25/Y
+ sky130_fd_sc_hd__mux2_2_43/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_826 VDD VSS sky130_fd_sc_hd__fa_2_1100/A sky130_fd_sc_hd__clkinv_8_59/Y
+ sky130_fd_sc_hd__and2_0_306/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_837 VDD VSS sky130_fd_sc_hd__nor2_1_139/A sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__o21bai_1_1/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_848 VDD VSS sky130_fd_sc_hd__mux2_2_57/A1 sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__o21ai_1_165/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_859 VDD VSS sky130_fd_sc_hd__mux2_2_66/A1 sky130_fd_sc_hd__clkinv_4_25/Y
+ sky130_fd_sc_hd__nor2_2_10/B VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_402 VSS VDD sky130_fd_sc_hd__clkbuf_1_402/X sky130_fd_sc_hd__clkbuf_1_402/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_413 VSS VDD sky130_fd_sc_hd__clkbuf_1_413/X sky130_fd_sc_hd__clkbuf_1_413/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_424 VSS VDD sky130_fd_sc_hd__clkbuf_1_424/X sky130_fd_sc_hd__clkbuf_1_535/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_435 VSS VDD sky130_fd_sc_hd__clkbuf_1_435/X sky130_fd_sc_hd__clkbuf_1_435/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_446 VSS VDD sky130_fd_sc_hd__a22oi_2_23/A2 sky130_fd_sc_hd__clkbuf_1_446/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_457 VSS VDD sky130_fd_sc_hd__clkbuf_1_457/X sky130_fd_sc_hd__clkbuf_1_457/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_468 VSS VDD sky130_fd_sc_hd__clkbuf_1_468/X sky130_fd_sc_hd__clkbuf_1_468/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_479 VSS VDD sky130_fd_sc_hd__nand4_1_53/D sky130_fd_sc_hd__a22oi_1_224/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_709 sky130_fd_sc_hd__fa_2_708/CIN sky130_fd_sc_hd__fa_2_709/SUM
+ sky130_fd_sc_hd__fa_2_709/A sky130_fd_sc_hd__fa_2_709/B sky130_fd_sc_hd__fa_2_709/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor2b_1_106 sky130_fd_sc_hd__or2_0_9/X sky130_fd_sc_hd__nor2b_1_106/Y
+ sky130_fd_sc_hd__buf_2_262/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_117 sky130_fd_sc_hd__and2_0_328/X sky130_fd_sc_hd__nor2b_1_117/Y
+ sky130_fd_sc_hd__buf_2_262/X VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_128 sky130_fd_sc_hd__nor3_1_41/Y sky130_fd_sc_hd__nor2b_1_128/Y
+ sky130_fd_sc_hd__buf_2_262/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_139 sky130_fd_sc_hd__o21ai_1_508/Y sky130_fd_sc_hd__nor2b_1_139/Y
+ sky130_fd_sc_hd__nor2b_1_142/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__buf_6_7 VDD VSS sky130_fd_sc_hd__buf_6_7/X sky130_fd_sc_hd__buf_6_7/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__clkinv_2_20 sky130_fd_sc_hd__buf_8_204/A sky130_fd_sc_hd__clkinv_2_20/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_20/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_31 sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__nor2_1_29/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_31/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_42 sky130_fd_sc_hd__dfxtp_1_93/D sky130_fd_sc_hd__clkinv_2_42/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_42/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__or2_1_2 sky130_fd_sc_hd__or2_1_2/A sky130_fd_sc_hd__or2_1_2/X sky130_fd_sc_hd__or2_1_2/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__or2_1
Xsky130_fd_sc_hd__o22ai_1_207 sky130_fd_sc_hd__nor2_2_13/B sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__o22ai_1_207/Y sky130_fd_sc_hd__a21oi_1_234/Y sky130_fd_sc_hd__a21boi_0_3/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__sdlclkp_4_5 sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__clkinv_8_69/A
+ sky130_fd_sc_hd__dfxtp_1_73/CLK sky130_fd_sc_hd__nor3_1_3/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__o22ai_1_218 sky130_fd_sc_hd__nand2_1_358/Y sky130_fd_sc_hd__nand2_1_357/Y
+ sky130_fd_sc_hd__o22ai_1_218/Y sky130_fd_sc_hd__nand2_1_371/B sky130_fd_sc_hd__o21ai_1_281/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_229 sky130_fd_sc_hd__nand2_1_360/Y sky130_fd_sc_hd__nand2_1_359/Y
+ sky130_fd_sc_hd__o22ai_1_229/Y sky130_fd_sc_hd__nand2_1_370/B sky130_fd_sc_hd__o21ai_1_280/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_1_8 sky130_fd_sc_hd__or4_1_1/C sky130_fd_sc_hd__nor2_1_8/Y
+ sky130_fd_sc_hd__nor2_1_8/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_190 sky130_fd_sc_hd__clkbuf_1_264/X sky130_fd_sc_hd__nor2_2_3/Y
+ sky130_fd_sc_hd__a22oi_1_190/B2 sky130_fd_sc_hd__clkbuf_4_127/X sky130_fd_sc_hd__nand4_1_42/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__o21ai_1_401 VSS VDD sky130_fd_sc_hd__a222oi_1_26/Y sky130_fd_sc_hd__nor2_1_265/A
+ sky130_fd_sc_hd__a21oi_1_384/Y sky130_fd_sc_hd__xor2_1_260/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_412 VSS VDD sky130_fd_sc_hd__o21ai_1_412/A2 sky130_fd_sc_hd__o22ai_1_379/A2
+ sky130_fd_sc_hd__a22oi_1_392/Y sky130_fd_sc_hd__o21ai_1_412/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_423 VSS VDD sky130_fd_sc_hd__a21oi_1_410/Y sky130_fd_sc_hd__nor2_1_257/A
+ sky130_fd_sc_hd__o21ai_1_425/B1 sky130_fd_sc_hd__o21ai_1_423/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_434 VSS VDD sky130_fd_sc_hd__o22ai_1_375/A2 sky130_fd_sc_hd__o21a_1_55/A2
+ sky130_fd_sc_hd__a21oi_1_415/Y sky130_fd_sc_hd__o21ai_1_434/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_445 VSS VDD sky130_fd_sc_hd__o22ai_1_406/A1 sky130_fd_sc_hd__nor2_1_289/Y
+ sky130_fd_sc_hd__or3_1_5/X sky130_fd_sc_hd__o21ai_1_445/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_456 VSS VDD sky130_fd_sc_hd__o22ai_1_418/A1 sky130_fd_sc_hd__o21a_1_68/A1
+ sky130_fd_sc_hd__a21oi_1_446/Y sky130_fd_sc_hd__o21ai_1_456/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_467 VSS VDD sky130_fd_sc_hd__o22ai_1_423/B1 sky130_fd_sc_hd__o21a_1_68/A1
+ sky130_fd_sc_hd__a21oi_1_457/Y sky130_fd_sc_hd__o21ai_1_467/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_478 VSS VDD sky130_fd_sc_hd__o22ai_1_429/B1 sky130_fd_sc_hd__o21a_1_68/A1
+ sky130_fd_sc_hd__a21oi_1_463/Y sky130_fd_sc_hd__o21ai_1_478/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_489 VSS VDD sky130_fd_sc_hd__nor2_1_299/A sky130_fd_sc_hd__o21a_1_68/X
+ sky130_fd_sc_hd__a211oi_1_38/Y sky130_fd_sc_hd__xor2_1_295/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_4_10 sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_2_7/A
+ sky130_fd_sc_hd__nor2_4_10/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__dfxtp_1_1007 VDD VSS sky130_fd_sc_hd__mux2_2_101/A0 sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__o22ai_1_232/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_16 VSS VDD sky130_fd_sc_hd__nor2b_1_50/Y sky130_fd_sc_hd__nand2_1_33/A
+ sky130_fd_sc_hd__nand2_1_33/Y sky130_fd_sc_hd__o21ai_1_4/A2 VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1018 VDD VSS sky130_fd_sc_hd__mux2_2_76/A1 sky130_fd_sc_hd__clkinv_8_46/Y
+ sky130_fd_sc_hd__a221oi_1_2/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_27 VSS VDD sky130_fd_sc_hd__a21oi_2_0/Y sky130_fd_sc_hd__nor2_1_13/B
+ sky130_fd_sc_hd__nand2_1_46/Y sky130_fd_sc_hd__o21ai_1_27/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_250 sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1225/B
+ sky130_fd_sc_hd__xor2_1_250/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_1029 VDD VSS sky130_fd_sc_hd__fa_2_840/A sky130_fd_sc_hd__dfxtp_1_1038/CLK
+ sky130_fd_sc_hd__o21a_1_38/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_38 VSS VDD sky130_fd_sc_hd__o21ai_1_38/A2 sky130_fd_sc_hd__o21ai_1_38/A1
+ sky130_fd_sc_hd__xor2_1_30/B sky130_fd_sc_hd__o21ai_1_38/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_601 VDD VSS sky130_fd_sc_hd__and2_0_211/A sky130_fd_sc_hd__dfxtp_1_601/CLK
+ sky130_fd_sc_hd__fa_2_1021/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_261 sky130_fd_sc_hd__xor2_1_267/B sky130_fd_sc_hd__fa_2_1253/B
+ sky130_fd_sc_hd__xor2_1_261/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o21ai_1_49 VSS VDD sky130_fd_sc_hd__o21ai_1_53/A2 sky130_fd_sc_hd__xnor2_1_52/Y
+ sky130_fd_sc_hd__a21oi_1_37/Y sky130_fd_sc_hd__o21ai_1_49/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_612 VDD VSS sky130_fd_sc_hd__fa_2_801/B sky130_fd_sc_hd__dfxtp_1_627/CLK
+ sky130_fd_sc_hd__a21oi_1_80/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_272 sky130_fd_sc_hd__fa_2_1242/A sky130_fd_sc_hd__xor2_1_272/X
+ sky130_fd_sc_hd__xor2_1_272/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_623 VDD VSS sky130_fd_sc_hd__ha_2_145/B sky130_fd_sc_hd__dfxtp_1_626/CLK
+ sky130_fd_sc_hd__a21oi_1_74/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_283 sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1288/B
+ sky130_fd_sc_hd__xor2_1_283/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_634 VDD VSS sky130_fd_sc_hd__fa_2_998/A sky130_fd_sc_hd__clkinv_8_44/Y
+ sky130_fd_sc_hd__and2_0_293/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_294 sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1277/B
+ sky130_fd_sc_hd__xor2_1_294/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_645 VDD VSS sky130_fd_sc_hd__fa_2_1009/A sky130_fd_sc_hd__clkinv_8_44/Y
+ sky130_fd_sc_hd__mux2_2_14/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_656 VDD VSS sky130_fd_sc_hd__fa_2_973/A sky130_fd_sc_hd__clkinv_8_41/Y
+ sky130_fd_sc_hd__and2_0_284/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_667 VDD VSS sky130_fd_sc_hd__fa_2_984/A sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__mux2_2_19/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_678 VDD VSS sky130_fd_sc_hd__fa_2_1017/A sky130_fd_sc_hd__clkinv_8_59/Y
+ sky130_fd_sc_hd__and2_0_270/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_689 VDD VSS sky130_fd_sc_hd__fa_2_1028/A sky130_fd_sc_hd__clkinv_4_26/Y
+ sky130_fd_sc_hd__and2_0_292/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_210 VSS VDD sky130_fd_sc_hd__buf_8_89/A sky130_fd_sc_hd__buf_8_67/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_221 VSS VDD sky130_fd_sc_hd__buf_8_107/A sky130_fd_sc_hd__buf_8_74/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_232 VSS VDD sky130_fd_sc_hd__clkbuf_1_232/X sky130_fd_sc_hd__clkbuf_1_232/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_243 VSS VDD sky130_fd_sc_hd__clkbuf_1_243/X sky130_fd_sc_hd__a22oi_1_122/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_254 VSS VDD sky130_fd_sc_hd__clkbuf_1_254/X sky130_fd_sc_hd__clkbuf_1_254/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_265 VSS VDD sky130_fd_sc_hd__clkbuf_1_265/X sky130_fd_sc_hd__nor3_2_6/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_276 VSS VDD sky130_fd_sc_hd__clkbuf_1_276/X sky130_fd_sc_hd__clkbuf_1_276/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_287 VSS VDD sky130_fd_sc_hd__clkbuf_1_287/X sky130_fd_sc_hd__clkbuf_1_287/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_298 VSS VDD sky130_fd_sc_hd__nand4_1_47/D sky130_fd_sc_hd__a22oi_1_207/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_506 sky130_fd_sc_hd__fa_2_507/B sky130_fd_sc_hd__fa_2_499/A
+ sky130_fd_sc_hd__ha_2_118/B sky130_fd_sc_hd__ha_2_122/B sky130_fd_sc_hd__fa_2_555/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_517 sky130_fd_sc_hd__fa_2_518/B sky130_fd_sc_hd__fa_2_509/A
+ sky130_fd_sc_hd__fa_2_546/A sky130_fd_sc_hd__ha_2_123/A sky130_fd_sc_hd__fa_2_502/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_528 sky130_fd_sc_hd__fa_2_530/CIN sky130_fd_sc_hd__fa_2_524/A
+ sky130_fd_sc_hd__fa_2_528/A sky130_fd_sc_hd__fa_2_528/B sky130_fd_sc_hd__fa_2_528/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_539 sky130_fd_sc_hd__fa_2_544/B sky130_fd_sc_hd__fa_2_539/SUM
+ sky130_fd_sc_hd__fa_2_539/A sky130_fd_sc_hd__fa_2_539/B sky130_fd_sc_hd__fa_2_539/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_4_4 VDD VSS sky130_fd_sc_hd__buf_4_4/X sky130_fd_sc_hd__buf_4_4/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__and2_0_230 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_230/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_847/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_241 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_241/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__or2_0_4/X sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_252 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_252/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__and2_0_252/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_263 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_263/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__fa_2_964/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_274 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_274/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__and2_0_274/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_285 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_285/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__and2_0_285/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_296 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_296/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_296/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__sdlclkp_2_2 sky130_fd_sc_hd__conb_1_8/LO sky130_fd_sc_hd__clkinv_4_5/Y
+ sky130_fd_sc_hd__clkinv_4_6/A sky130_fd_sc_hd__nand2b_1_0/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__nand3b_1_0 sky130_fd_sc_hd__nor2_4_1/Y sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__nand3b_1_0/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand3b_1
Xsky130_fd_sc_hd__o21ai_1_220 VSS VDD sky130_fd_sc_hd__a21oi_1_202/Y sky130_fd_sc_hd__nor2_1_127/A
+ sky130_fd_sc_hd__nand2_1_321/Y sky130_fd_sc_hd__o21ai_1_220/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_231 VSS VDD sky130_fd_sc_hd__o22ai_1_193/A1 sky130_fd_sc_hd__o21a_1_16/A2
+ sky130_fd_sc_hd__a21oi_1_205/Y sky130_fd_sc_hd__o21ai_1_231/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_242 VSS VDD sky130_fd_sc_hd__o21a_1_16/X sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__nand2_1_330/Y sky130_fd_sc_hd__xor2_1_91/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_60 sky130_fd_sc_hd__clkbuf_4_60/X sky130_fd_sc_hd__buf_2_35/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_253 VSS VDD sky130_fd_sc_hd__nand2_2_6/Y sky130_fd_sc_hd__o21ai_1_253/A1
+ sky130_fd_sc_hd__a21oi_1_219/Y sky130_fd_sc_hd__xor2_1_101/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_71 sky130_fd_sc_hd__clkbuf_4_71/X sky130_fd_sc_hd__buf_2_42/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_264 VSS VDD sky130_fd_sc_hd__a21oi_1_231/Y sky130_fd_sc_hd__nor2_1_127/A
+ sky130_fd_sc_hd__a21oi_1_229/Y sky130_fd_sc_hd__xor2_1_108/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_82 sky130_fd_sc_hd__clkbuf_4_82/X sky130_fd_sc_hd__clkbuf_4_82/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_275 VSS VDD sky130_fd_sc_hd__o22ai_1_197/A2 sky130_fd_sc_hd__o22ai_1_206/A1
+ sky130_fd_sc_hd__a22oi_1_370/Y sky130_fd_sc_hd__o21ai_1_275/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_93 sky130_fd_sc_hd__buf_2_38/A sky130_fd_sc_hd__inv_2_47/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_286 VSS VDD sky130_fd_sc_hd__nor2_1_148/B sky130_fd_sc_hd__o22ai_1_265/A2
+ sky130_fd_sc_hd__a22oi_1_372/Y sky130_fd_sc_hd__o21ai_1_286/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_297 VSS VDD sky130_fd_sc_hd__o21ai_1_306/A1 sky130_fd_sc_hd__nor2_1_180/A
+ sky130_fd_sc_hd__a21oi_1_271/Y sky130_fd_sc_hd__xor2_1_177/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2b_2_4 sky130_fd_sc_hd__o32ai_1_8/A1 sky130_fd_sc_hd__nor2b_2_4/A
+ sky130_fd_sc_hd__nor2b_2_4/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_2
Xsky130_fd_sc_hd__fa_2_1007 sky130_fd_sc_hd__fa_2_1008/CIN sky130_fd_sc_hd__mux2_2_18/A0
+ sky130_fd_sc_hd__fa_2_1007/A sky130_fd_sc_hd__xor2_1_69/X sky130_fd_sc_hd__fa_2_1007/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1018 sky130_fd_sc_hd__fa_2_1019/CIN sky130_fd_sc_hd__and2_0_271/A
+ sky130_fd_sc_hd__fa_2_1018/A sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_1018/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1029 sky130_fd_sc_hd__fa_2_1030/CIN sky130_fd_sc_hd__or2_0_5/B
+ sky130_fd_sc_hd__fa_2_1029/A sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_1029/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_16 sky130_fd_sc_hd__inv_2_16/A sky130_fd_sc_hd__inv_2_16/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_420 VDD VSS sky130_fd_sc_hd__fa_2_1040/B sky130_fd_sc_hd__dfxtp_1_425/CLK
+ sky130_fd_sc_hd__and2_0_127/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_27 sky130_fd_sc_hd__inv_2_27/A sky130_fd_sc_hd__inv_2_27/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_431 VDD VSS sky130_fd_sc_hd__dfxtp_1_431/Q sky130_fd_sc_hd__dfxtp_1_433/CLK
+ sky130_fd_sc_hd__nand2_1_102/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_442 VDD VSS sky130_fd_sc_hd__dfxtp_1_988/D sky130_fd_sc_hd__dfxtp_1_448/CLK
+ sky130_fd_sc_hd__nand2_1_80/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_38 sky130_fd_sc_hd__inv_2_38/A sky130_fd_sc_hd__inv_2_38/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_49 sky130_fd_sc_hd__ha_2_31/A sky130_fd_sc_hd__inv_2_50/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_453 VDD VSS sky130_fd_sc_hd__dfxtp_1_999/D sky130_fd_sc_hd__dfxtp_1_454/CLK
+ sky130_fd_sc_hd__nand2_1_58/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_464 VDD VSS sky130_fd_sc_hd__buf_2_6/A sky130_fd_sc_hd__dfxtp_1_472/CLK
+ sky130_fd_sc_hd__and2_0_151/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_475 VDD VSS sky130_fd_sc_hd__nor3_1_27/A sky130_fd_sc_hd__dfxtp_1_476/CLK
+ sky130_fd_sc_hd__and2_0_242/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_486 VDD VSS sky130_fd_sc_hd__dfxtp_1_486/Q sky130_fd_sc_hd__dfxtp_1_488/CLK
+ sky130_fd_sc_hd__nor2b_1_72/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_2_6 sky130_fd_sc_hd__nand2_2_6/Y sky130_fd_sc_hd__nand2_2_6/A
+ sky130_fd_sc_hd__nand2_2_6/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__dfxtp_1_497 VDD VSS sky130_fd_sc_hd__nor2b_1_86/A sky130_fd_sc_hd__dfxtp_1_502/CLK
+ sky130_fd_sc_hd__nor2b_1_78/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2b_1_12 sky130_fd_sc_hd__xnor2_1_33/B sky130_fd_sc_hd__ha_2_185/A
+ sky130_fd_sc_hd__ha_2_185/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__fa_2_303 sky130_fd_sc_hd__fa_2_300/CIN sky130_fd_sc_hd__nor2_1_212/A
+ sky130_fd_sc_hd__fa_2_303/A sky130_fd_sc_hd__fa_2_303/B sky130_fd_sc_hd__fa_2_303/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_314 sky130_fd_sc_hd__fa_2_310/CIN sky130_fd_sc_hd__or3_1_3/A
+ sky130_fd_sc_hd__fa_2_314/A sky130_fd_sc_hd__fa_2_314/B sky130_fd_sc_hd__fa_2_314/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_325 sky130_fd_sc_hd__fa_2_326/CIN sky130_fd_sc_hd__maj3_1_80/A
+ sky130_fd_sc_hd__ha_2_114/A sky130_fd_sc_hd__ha_2_112/B sky130_fd_sc_hd__ha_2_113/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_336 sky130_fd_sc_hd__fa_2_338/CIN sky130_fd_sc_hd__fa_2_334/A
+ sky130_fd_sc_hd__ha_2_116/B sky130_fd_sc_hd__ha_2_114/B sky130_fd_sc_hd__fa_2_425/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_347 sky130_fd_sc_hd__maj3_1_70/B sky130_fd_sc_hd__maj3_1_71/A
+ sky130_fd_sc_hd__fa_2_347/A sky130_fd_sc_hd__fa_2_347/B sky130_fd_sc_hd__fa_2_348/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_358 sky130_fd_sc_hd__fa_2_355/B sky130_fd_sc_hd__fa_2_358/SUM
+ sky130_fd_sc_hd__fa_2_404/A sky130_fd_sc_hd__ha_2_116/A sky130_fd_sc_hd__fa_2_395/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_369 sky130_fd_sc_hd__fa_2_370/CIN sky130_fd_sc_hd__fa_2_363/A
+ sky130_fd_sc_hd__fa_2_416/B sky130_fd_sc_hd__fa_2_409/A sky130_fd_sc_hd__fa_2_425/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_1_7 VDD VSS sky130_fd_sc_hd__and2_1_7/X sky130_fd_sc_hd__ha_2_59/A
+ sky130_fd_sc_hd__nor2_4_2/Y VDD VSS sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__diode_2_208 sig_frequency[7] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkinv_8_30 sky130_fd_sc_hd__clkinv_8_32/A sky130_fd_sc_hd__clkinv_8_30/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_30/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__diode_2_219 sig_amplitude[3] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkinv_8_41 sky130_fd_sc_hd__clkinv_8_41/Y sky130_fd_sc_hd__clkinv_8_43/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_41/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_52 sky130_fd_sc_hd__clkinv_8_53/A sky130_fd_sc_hd__clkinv_8_95/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_52/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_63 sky130_fd_sc_hd__clkinv_8_63/Y sky130_fd_sc_hd__clkinv_8_63/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_63/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_74 sky130_fd_sc_hd__clkinv_8_74/Y sky130_fd_sc_hd__clkinv_8_74/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_74/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_85 sky130_fd_sc_hd__clkinv_8_86/A sky130_fd_sc_hd__clkinv_8_85/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_96 sky130_fd_sc_hd__clkinv_4_2/A sky130_fd_sc_hd__clkinv_8_96/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_50 sky130_fd_sc_hd__buf_8_31/X sky130_fd_sc_hd__buf_12_50/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_61 sky130_fd_sc_hd__buf_12_61/A sky130_fd_sc_hd__buf_12_61/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_72 sky130_fd_sc_hd__buf_4_21/X sky130_fd_sc_hd__buf_12_72/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_83 sky130_fd_sc_hd__buf_4_13/X sky130_fd_sc_hd__buf_12_83/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_94 sky130_fd_sc_hd__buf_12_94/A sky130_fd_sc_hd__buf_12_94/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_2_1 VDD VSS sky130_fd_sc_hd__buf_2_1/X sky130_fd_sc_hd__buf_4_0/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1360 VDD VSS sky130_fd_sc_hd__fa_2_1282/A sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__mux2_2_246/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1371 VDD VSS sky130_fd_sc_hd__xor2_1_299/A sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__mux2_2_221/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1382 VDD VSS sky130_fd_sc_hd__fa_2_1321/A sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__mux2_2_247/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1393 VDD VSS sky130_fd_sc_hd__nor2_4_19/A sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__nor2b_1_129/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_12_308 sky130_fd_sc_hd__buf_8_163/X sky130_fd_sc_hd__buf_12_308/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_319 sky130_fd_sc_hd__buf_4_87/X sky130_fd_sc_hd__buf_12_319/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__fa_2_870 sky130_fd_sc_hd__fa_2_869/CIN sky130_fd_sc_hd__fa_2_870/SUM
+ sky130_fd_sc_hd__fa_2_870/A sky130_fd_sc_hd__fa_2_870/B sky130_fd_sc_hd__fa_2_870/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_881 sky130_fd_sc_hd__fa_2_880/CIN sky130_fd_sc_hd__nand2_1_41/B
+ sky130_fd_sc_hd__ha_2_152/A sky130_fd_sc_hd__fa_2_881/B sky130_fd_sc_hd__fa_2_881/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_892 sky130_fd_sc_hd__fa_2_891/CIN sky130_fd_sc_hd__fa_2_892/SUM
+ sky130_fd_sc_hd__fa_2_892/A sky130_fd_sc_hd__fa_2_892/B sky130_fd_sc_hd__fa_2_892/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_1 sky130_fd_sc_hd__inv_2_1/A sky130_fd_sc_hd__inv_2_1/Y VDD
+ VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__nor3_2_3 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__nor3_2_3/Y
+ sky130_fd_sc_hd__nor3_2_3/A sky130_fd_sc_hd__nor3_2_3/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_2
Xsky130_fd_sc_hd__clkinv_1_508 sky130_fd_sc_hd__a21oi_1_61/A1 sky130_fd_sc_hd__nor2_1_51/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_508/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_519 sky130_fd_sc_hd__nor2_1_58/B sky130_fd_sc_hd__fa_2_1036/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_519/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_11 sky130_fd_sc_hd__nor2_1_11/B sky130_fd_sc_hd__nor2_1_11/Y
+ sky130_fd_sc_hd__xor2_1_20/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_22 sky130_fd_sc_hd__nor2_1_22/B sky130_fd_sc_hd__nor2_1_22/Y
+ sky130_fd_sc_hd__nor2_1_22/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_33 sky130_fd_sc_hd__nor2_1_33/B sky130_fd_sc_hd__nor2_1_33/Y
+ sky130_fd_sc_hd__nor4_1_8/D VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_44 sky130_fd_sc_hd__nor2_1_44/B sky130_fd_sc_hd__nor2_1_44/Y
+ sky130_fd_sc_hd__nor2_1_53/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_55 sky130_fd_sc_hd__nor2_1_55/B sky130_fd_sc_hd__nor2_1_55/Y
+ sky130_fd_sc_hd__nor2_1_55/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_66 sky130_fd_sc_hd__nor2_1_66/B sky130_fd_sc_hd__o21a_1_4/A1
+ sky130_fd_sc_hd__o21a_1_5/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_170 VSS VDD sky130_fd_sc_hd__mux2_2_170/A1 sky130_fd_sc_hd__mux2_2_170/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_170/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_77 sky130_fd_sc_hd__nor2_1_79/Y sky130_fd_sc_hd__nor2_1_77/Y
+ sky130_fd_sc_hd__nor2_1_77/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_181 VSS VDD sky130_fd_sc_hd__mux2_2_181/A1 sky130_fd_sc_hd__mux2_2_181/A0
+ sky130_fd_sc_hd__nor2_8_1/A sky130_fd_sc_hd__mux2_2_181/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_88 sky130_fd_sc_hd__o21a_1_8/A2 sky130_fd_sc_hd__nor2_1_88/Y
+ sky130_fd_sc_hd__nor2_1_88/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_192 VSS VDD sky130_fd_sc_hd__mux2_2_192/A1 sky130_fd_sc_hd__mux2_2_192/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_192/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_99 sky130_fd_sc_hd__nor2_1_99/B sky130_fd_sc_hd__nor2_1_99/Y
+ sky130_fd_sc_hd__nor2_1_99/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_sram_2kbyte_1rw1r_32x512_8_7 sky130_fd_sc_hd__buf_4_32/X sky130_fd_sc_hd__buf_8_63/X
+ sky130_fd_sc_hd__buf_2_35/A sky130_fd_sc_hd__buf_4_34/X sky130_fd_sc_hd__inv_12_0/Y
+ sky130_fd_sc_hd__clkbuf_4_63/X sky130_fd_sc_hd__buf_2_36/A sky130_fd_sc_hd__buf_4_36/X
+ sky130_fd_sc_hd__clkbuf_1_198/X sky130_fd_sc_hd__clkbuf_1_201/X sky130_fd_sc_hd__buf_2_38/A
+ sky130_fd_sc_hd__buf_2_39/A sky130_fd_sc_hd__clkbuf_4_95/X sky130_fd_sc_hd__buf_2_40/A
+ sky130_fd_sc_hd__buf_2_41/A sky130_fd_sc_hd__buf_2_42/A sky130_fd_sc_hd__buf_4_32/X
+ sky130_fd_sc_hd__buf_8_63/X sky130_fd_sc_hd__buf_2_35/A sky130_fd_sc_hd__buf_4_34/X
+ sky130_fd_sc_hd__inv_12_0/Y sky130_fd_sc_hd__clkbuf_4_63/X sky130_fd_sc_hd__buf_2_36/A
+ sky130_fd_sc_hd__buf_4_36/X sky130_fd_sc_hd__buf_2_116/X sky130_fd_sc_hd__buf_2_117/X
+ sky130_fd_sc_hd__buf_2_38/A sky130_fd_sc_hd__buf_2_39/A sky130_fd_sc_hd__clkbuf_4_95/X
+ sky130_fd_sc_hd__buf_2_40/A sky130_fd_sc_hd__buf_2_41/A sky130_fd_sc_hd__buf_2_42/A
+ sky130_fd_sc_hd__buf_12_193/X sky130_fd_sc_hd__buf_12_215/X sky130_fd_sc_hd__buf_12_173/X
+ sky130_fd_sc_hd__buf_12_125/X sky130_fd_sc_hd__buf_12_264/X sky130_fd_sc_hd__buf_12_178/X
+ sky130_fd_sc_hd__buf_12_203/X sky130_fd_sc_hd__buf_12_254/X sky130_fd_sc_hd__buf_12_258/X
+ sky130_fd_sc_hd__buf_12_253/X sky130_fd_sc_hd__buf_12_138/X sky130_fd_sc_hd__buf_12_143/X
+ sky130_fd_sc_hd__buf_12_237/X sky130_fd_sc_hd__buf_12_241/X sky130_fd_sc_hd__buf_12_154/X
+ sky130_fd_sc_hd__buf_12_214/X sky130_fd_sc_hd__buf_12_195/X sky130_fd_sc_hd__buf_12_255/X
+ sky130_fd_sc_hd__buf_2_120/X sky130_fd_sc_hd__nand3_1_31/Y sky130_fd_sc_hd__buf_2_120/X
+ sky130_fd_sc_hd__clkinv_8_11/Y sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__buf_12_248/X
+ sky130_fd_sc_hd__buf_12_240/X sky130_fd_sc_hd__buf_12_246/X sky130_fd_sc_hd__buf_12_192/X
+ sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[0] sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[1]
+ sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[2] sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[3]
+ sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[4] sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[5]
+ sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[6] sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[7]
+ sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[8] sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[9]
+ sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[10] sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[11]
+ sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[12] sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[13]
+ sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[14] sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[15]
+ sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[16] sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[17]
+ sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[18] sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[19]
+ sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[20] sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[21]
+ sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[22] sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[23]
+ sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[24] sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[25]
+ sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[26] sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[27]
+ sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[28] sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[29]
+ sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[30] sky130_sram_2kbyte_1rw1r_32x512_8_7/dout0[31]
+ sky130_fd_sc_hd__clkbuf_1_139/A sky130_fd_sc_hd__clkbuf_1_140/A sky130_fd_sc_hd__clkbuf_1_141/A
+ sky130_fd_sc_hd__clkbuf_1_142/A sky130_fd_sc_hd__clkbuf_1_143/A sky130_fd_sc_hd__clkbuf_1_144/A
+ sky130_fd_sc_hd__clkbuf_1_145/A sky130_fd_sc_hd__buf_2_122/A sky130_fd_sc_hd__clkbuf_1_147/A
+ sky130_fd_sc_hd__clkbuf_1_148/A sky130_fd_sc_hd__clkbuf_1_149/A sky130_fd_sc_hd__clkbuf_1_251/A
+ sky130_fd_sc_hd__clkbuf_1_151/A sky130_fd_sc_hd__clkbuf_1_152/A sky130_fd_sc_hd__clkbuf_1_153/A
+ sky130_fd_sc_hd__clkbuf_1_154/A sky130_fd_sc_hd__a22oi_1_143/A2 sky130_fd_sc_hd__a22oi_1_139/A2
+ sky130_fd_sc_hd__a22oi_1_135/A2 sky130_fd_sc_hd__a22oi_1_131/A2 sky130_fd_sc_hd__a22oi_1_128/A2
+ sky130_fd_sc_hd__a22oi_1_124/A2 sky130_fd_sc_hd__a22oi_1_120/A2 sky130_fd_sc_hd__a22oi_1_116/A2
+ sky130_fd_sc_hd__a22oi_1_112/A2 sky130_fd_sc_hd__a22oi_1_108/A2 sky130_fd_sc_hd__a22oi_1_104/A2
+ sky130_fd_sc_hd__a22oi_1_100/A2 sky130_fd_sc_hd__a22oi_1_96/A2 sky130_fd_sc_hd__a22oi_1_92/A2
+ sky130_fd_sc_hd__a22oi_1_88/A2 sky130_fd_sc_hd__a22oi_1_84/A2 VDD VSS sky130_sram_2kbyte_1rw1r_32x512_8
Xsky130_fd_sc_hd__a21oi_1_405 sky130_fd_sc_hd__fa_2_1256/A sky130_fd_sc_hd__o22ai_1_368/Y
+ sky130_fd_sc_hd__a21oi_1_405/Y sky130_fd_sc_hd__clkinv_1_946/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_416 sky130_fd_sc_hd__fa_2_1248/A sky130_fd_sc_hd__o22ai_1_375/Y
+ sky130_fd_sc_hd__a21oi_1_416/Y sky130_fd_sc_hd__nor3_1_40/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_427 sky130_fd_sc_hd__nor2_1_275/A sky130_fd_sc_hd__o21a_1_61/A1
+ sky130_fd_sc_hd__a21oi_1_427/Y sky130_fd_sc_hd__nor2_1_275/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_438 sky130_fd_sc_hd__or3_1_5/C sky130_fd_sc_hd__o21ai_1_438/Y
+ sky130_fd_sc_hd__a21oi_1_438/Y sky130_fd_sc_hd__nor2_1_288/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_449 sky130_fd_sc_hd__nor2b_2_5/Y sky130_fd_sc_hd__o21ai_1_458/Y
+ sky130_fd_sc_hd__a21oi_1_449/Y sky130_fd_sc_hd__o21ai_1_467/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_8_107 sky130_fd_sc_hd__clkinv_8_114/A sky130_fd_sc_hd__clkinv_8_107/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_107/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_118 sky130_fd_sc_hd__clkinv_8_118/Y sky130_fd_sc_hd__clkinv_4_60/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_118/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_129 sky130_fd_sc_hd__clkinv_8_129/Y sky130_fd_sc_hd__clkinv_4_69/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_129/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__o21a_1_9 sky130_fd_sc_hd__o21a_1_9/X sky130_fd_sc_hd__o21a_1_9/A1
+ sky130_fd_sc_hd__o21a_1_9/B1 sky130_fd_sc_hd__o21a_1_9/A2 VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__maj3_1_130 sky130_fd_sc_hd__maj3_1_131/X sky130_fd_sc_hd__maj3_1_130/X
+ sky130_fd_sc_hd__maj3_1_130/B sky130_fd_sc_hd__maj3_1_130/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_141 sky130_fd_sc_hd__maj3_1_142/X sky130_fd_sc_hd__maj3_1_141/X
+ sky130_fd_sc_hd__maj3_1_141/B sky130_fd_sc_hd__maj3_1_141/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_410 sky130_fd_sc_hd__nand2_1_410/Y sky130_fd_sc_hd__nor2_1_203/B
+ sky130_fd_sc_hd__o31ai_1_7/A2 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_152 sky130_fd_sc_hd__maj3_1_153/X sky130_fd_sc_hd__maj3_1_152/X
+ sky130_fd_sc_hd__maj3_1_152/B sky130_fd_sc_hd__maj3_1_152/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_421 sky130_fd_sc_hd__nor2_1_209/B sky130_fd_sc_hd__nand2_1_421/B
+ sky130_fd_sc_hd__nor2_1_210/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_432 sky130_fd_sc_hd__nand2_1_432/Y sky130_fd_sc_hd__fa_2_1190/A
+ sky130_fd_sc_hd__nor3_1_39/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_443 sky130_fd_sc_hd__nor2_1_225/A sky130_fd_sc_hd__nor2b_2_3/A
+ sky130_fd_sc_hd__o32ai_1_5/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_390 sky130_fd_sc_hd__nand2_1_514/Y sky130_fd_sc_hd__nand2_1_513/Y
+ sky130_fd_sc_hd__o22ai_1_390/Y sky130_fd_sc_hd__o22ai_1_403/A1 sky130_fd_sc_hd__a21o_2_28/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_454 sky130_fd_sc_hd__o21a_1_50/B1 sky130_fd_sc_hd__fa_2_1256/A
+ sky130_fd_sc_hd__o21a_1_50/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_465 sky130_fd_sc_hd__nand2_1_465/Y sky130_fd_sc_hd__nand2_1_468/Y
+ sky130_fd_sc_hd__nand2_1_466/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_476 sky130_fd_sc_hd__nor2_1_255/B sky130_fd_sc_hd__nand2_1_476/B
+ sky130_fd_sc_hd__nor2_1_256/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_487 sky130_fd_sc_hd__nand2_1_487/Y sky130_fd_sc_hd__nand2_1_491/B
+ sky130_fd_sc_hd__o21ai_1_436/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_498 sky130_fd_sc_hd__o21a_1_56/B1 sky130_fd_sc_hd__fa_2_1291/A
+ sky130_fd_sc_hd__o21a_1_56/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_12 sky130_fd_sc_hd__ha_2_28/SUM sky130_fd_sc_hd__nor2b_1_12/Y
+ sky130_fd_sc_hd__or2_0_1/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_23 sky130_fd_sc_hd__ha_2_47/SUM sky130_fd_sc_hd__nor2b_1_23/Y
+ sky130_fd_sc_hd__or2_1_0/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_34 sky130_fd_sc_hd__ha_2_62/SUM sky130_fd_sc_hd__nor2b_1_34/Y
+ sky130_fd_sc_hd__or2_0_2/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1001 sky130_fd_sc_hd__o22ai_1_366/B1 sky130_fd_sc_hd__fa_2_1236/A
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_45 sky130_fd_sc_hd__ha_2_83/SUM sky130_fd_sc_hd__nor2b_1_45/Y
+ sky130_fd_sc_hd__or2_0_3/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1012 sky130_fd_sc_hd__nor2_1_242/B sky130_fd_sc_hd__fa_2_1245/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1012/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_56 sky130_fd_sc_hd__dfxtp_1_486/Q sky130_fd_sc_hd__nor2b_1_56/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1023 sky130_fd_sc_hd__o22ai_1_379/B1 sky130_fd_sc_hd__fa_2_1254/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1023/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_67 sky130_fd_sc_hd__o21ai_1_38/A1 sky130_fd_sc_hd__nor2b_1_67/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1034 sky130_fd_sc_hd__or2_0_12/B sky130_fd_sc_hd__nor2_1_310/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1034/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_78 sky130_fd_sc_hd__dfxtp_1_498/Q sky130_fd_sc_hd__nor2b_1_78/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1045 sky130_fd_sc_hd__nor2_1_281/A sky130_fd_sc_hd__nor2_1_282/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1045/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_89 sky130_fd_sc_hd__fa_2_957/A sky130_fd_sc_hd__or3_1_1/A
+ sky130_fd_sc_hd__nor2b_1_89/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1056 sky130_fd_sc_hd__o22ai_1_406/A1 sky130_fd_sc_hd__or3_1_5/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1056/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1067 sky130_fd_sc_hd__nand2_1_525/B sky130_fd_sc_hd__fa_2_6/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1067/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_8 VSS VDD sky130_fd_sc_hd__xnor2_1_8/B sky130_fd_sc_hd__xnor2_1_8/Y
+ sky130_fd_sc_hd__xnor2_1_9/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_1078 sky130_fd_sc_hd__nor2_1_276/B sky130_fd_sc_hd__fa_2_1278/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1078/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1089 sky130_fd_sc_hd__a21oi_1_461/B1 sky130_fd_sc_hd__nand2_1_542/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1089/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_250 VDD VSS sky130_fd_sc_hd__dfxtp_1_250/Q sky130_fd_sc_hd__dfxtp_1_262/CLK
+ sky130_fd_sc_hd__and2_0_202/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_261 VDD VSS sky130_fd_sc_hd__dfxtp_1_261/Q sky130_fd_sc_hd__dfxtp_1_262/CLK
+ sky130_fd_sc_hd__and2_0_183/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_272 VDD VSS sky130_fd_sc_hd__dfxtp_1_272/Q sky130_fd_sc_hd__dfxtp_1_472/CLK
+ sky130_fd_sc_hd__and2_0_212/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_283 VDD VSS sky130_fd_sc_hd__a22o_1_64/A1 sky130_fd_sc_hd__dfxtp_1_477/CLK
+ sky130_fd_sc_hd__nand2_1_143/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_294 VDD VSS sky130_fd_sc_hd__a22o_1_53/A1 sky130_fd_sc_hd__clkinv_4_31/Y
+ sky130_fd_sc_hd__nand2_1_121/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o22ai_1_3 sky130_fd_sc_hd__ha_2_95/B sky130_fd_sc_hd__fa_2_76/B
+ sky130_fd_sc_hd__o22ai_1_3/Y sky130_fd_sc_hd__ha_2_91/B sky130_fd_sc_hd__fa_2_139/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_100 sky130_fd_sc_hd__fa_2_97/B sky130_fd_sc_hd__fa_2_93/B sky130_fd_sc_hd__fa_2_87/A
+ sky130_fd_sc_hd__ha_2_96/B sky130_fd_sc_hd__fa_2_87/B VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_111 sky130_fd_sc_hd__fa_2_110/A sky130_fd_sc_hd__fa_2_104/B
+ sky130_fd_sc_hd__fa_2_82/A sky130_fd_sc_hd__fa_2_45/A sky130_fd_sc_hd__fa_2_76/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_122 sky130_fd_sc_hd__fa_2_125/B sky130_fd_sc_hd__fa_2_122/SUM
+ sky130_fd_sc_hd__fa_2_122/A sky130_fd_sc_hd__fa_2_122/B sky130_fd_sc_hd__fa_2_122/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_133 sky130_fd_sc_hd__fa_2_26/A sky130_fd_sc_hd__fa_2_27/B sky130_fd_sc_hd__fa_2_133/A
+ sky130_fd_sc_hd__fa_2_133/B sky130_fd_sc_hd__fa_2_137/SUM VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_144 sky130_fd_sc_hd__xnor2_1_1/A sky130_fd_sc_hd__fa_2_144/SUM
+ sky130_fd_sc_hd__fa_2_2/A sky130_fd_sc_hd__fa_2_144/B sky130_fd_sc_hd__fa_2_144/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_155 sky130_fd_sc_hd__fa_2_151/B sky130_fd_sc_hd__fa_2_155/SUM
+ sky130_fd_sc_hd__fa_2_2/A sky130_fd_sc_hd__fa_2_242/A sky130_fd_sc_hd__fa_2_274/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_166 sky130_fd_sc_hd__fa_2_162/A sky130_fd_sc_hd__fa_2_167/A
+ sky130_fd_sc_hd__fa_2_209/B sky130_fd_sc_hd__fa_2_5/A sky130_fd_sc_hd__fa_2_144/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_177 sky130_fd_sc_hd__fa_2_178/A sky130_fd_sc_hd__fa_2_177/SUM
+ sky130_fd_sc_hd__ha_2_104/B sky130_fd_sc_hd__fa_2_31/A sky130_fd_sc_hd__fa_2_266/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_188 sky130_fd_sc_hd__fa_2_190/B sky130_fd_sc_hd__fa_2_186/A
+ sky130_fd_sc_hd__fa_2_5/B sky130_fd_sc_hd__fa_2_15/B sky130_fd_sc_hd__fa_2_277/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_199 sky130_fd_sc_hd__fa_2_198/A sky130_fd_sc_hd__fa_2_193/B
+ sky130_fd_sc_hd__ha_2_107/A sky130_fd_sc_hd__fa_2_247/A sky130_fd_sc_hd__fa_2_250/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor3_2_10 sky130_fd_sc_hd__nor2_2_4/A sky130_fd_sc_hd__nor3_2_10/Y
+ sky130_fd_sc_hd__nor3_2_10/A sky130_fd_sc_hd__nor3_2_10/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_2
Xsky130_fd_sc_hd__o22ai_1_10 sky130_fd_sc_hd__fa_2_2/B sky130_fd_sc_hd__fa_2_91/B
+ sky130_fd_sc_hd__fa_2_129/A sky130_fd_sc_hd__ha_2_93/A sky130_fd_sc_hd__ha_2_97/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_21 sky130_fd_sc_hd__fa_2_412/A sky130_fd_sc_hd__fa_2_286/B
+ sky130_fd_sc_hd__xnor2_1_2/B sky130_fd_sc_hd__ha_2_116/A sky130_fd_sc_hd__ha_2_108/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_32 sky130_fd_sc_hd__fa_2_535/A sky130_fd_sc_hd__fa_2_537/A
+ sky130_fd_sc_hd__o22ai_1_32/Y sky130_fd_sc_hd__ha_2_123/A sky130_fd_sc_hd__fa_2_543/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_150 VDD VSS sky130_fd_sc_hd__buf_4_100/A sky130_fd_sc_hd__buf_6_52/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_43 sky130_fd_sc_hd__fa_2_677/A sky130_fd_sc_hd__ha_2_131/B
+ sky130_fd_sc_hd__o22ai_1_43/Y sky130_fd_sc_hd__fa_2_678/B sky130_fd_sc_hd__ha_2_126/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_161 VDD VSS sky130_fd_sc_hd__buf_8_201/A sky130_fd_sc_hd__buf_2_161/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_54 sky130_fd_sc_hd__fa_2_835/B sky130_fd_sc_hd__ha_2_140/A
+ sky130_fd_sc_hd__o22ai_1_54/Y sky130_fd_sc_hd__fa_2_807/B sky130_fd_sc_hd__fa_2_834/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_172 VDD VSS sky130_fd_sc_hd__buf_2_172/X sky130_fd_sc_hd__buf_2_172/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_65 sky130_fd_sc_hd__o22ai_1_88/B1 sky130_fd_sc_hd__nand2_2_3/Y
+ sky130_fd_sc_hd__o22ai_1_65/Y sky130_fd_sc_hd__xnor2_1_41/Y sky130_fd_sc_hd__o22ai_1_79/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_183 VDD VSS sky130_fd_sc_hd__buf_2_183/X sky130_fd_sc_hd__buf_2_183/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_76 sky130_fd_sc_hd__o22ai_1_89/A1 sky130_fd_sc_hd__o22ai_1_88/B1
+ sky130_fd_sc_hd__o22ai_1_76/Y sky130_fd_sc_hd__xnor2_1_35/Y sky130_fd_sc_hd__o22ai_1_76/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_194 VDD VSS sky130_fd_sc_hd__buf_2_194/X sky130_fd_sc_hd__buf_2_194/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_87 sky130_fd_sc_hd__o22ai_1_89/A1 sky130_fd_sc_hd__o22ai_1_88/B1
+ sky130_fd_sc_hd__o22ai_1_87/Y sky130_fd_sc_hd__xnor2_1_57/Y sky130_fd_sc_hd__o22ai_1_87/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_98 sky130_fd_sc_hd__nor2_1_76/A sky130_fd_sc_hd__nor2_2_9/B
+ sky130_fd_sc_hd__o22ai_1_98/Y sky130_fd_sc_hd__a21oi_1_95/Y sky130_fd_sc_hd__a222oi_1_0/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__dfxtp_1_1190 VDD VSS sky130_fd_sc_hd__fa_2_943/A sky130_fd_sc_hd__clkinv_4_24/Y
+ sky130_fd_sc_hd__o21a_1_43/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_4_12 VDD VSS sky130_fd_sc_hd__buf_4_12/X sky130_fd_sc_hd__buf_4_12/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_23 VDD VSS sky130_fd_sc_hd__buf_4_23/X sky130_fd_sc_hd__buf_8_52/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_34 VDD VSS sky130_fd_sc_hd__buf_4_34/X sky130_fd_sc_hd__buf_4_34/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_45 VDD VSS sky130_fd_sc_hd__buf_4_45/X sky130_fd_sc_hd__buf_8_75/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_56 VDD VSS sky130_fd_sc_hd__buf_4_56/X sky130_fd_sc_hd__buf_4_56/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_67 VDD VSS sky130_fd_sc_hd__buf_4_67/X sky130_fd_sc_hd__buf_4_67/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_78 VDD VSS sky130_fd_sc_hd__buf_4_78/X sky130_fd_sc_hd__buf_4_79/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_89 VDD VSS sky130_fd_sc_hd__buf_4_89/X sky130_fd_sc_hd__buf_4_89/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_12_105 sky130_fd_sc_hd__buf_12_9/X sky130_fd_sc_hd__buf_12_105/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_116 sky130_fd_sc_hd__buf_12_116/A sky130_fd_sc_hd__buf_12_117/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_127 sky130_fd_sc_hd__buf_12_127/A sky130_fd_sc_hd__buf_12_172/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_50 VSS VDD sky130_fd_sc_hd__clkbuf_1_50/X sky130_fd_sc_hd__clkbuf_1_50/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_138 sky130_fd_sc_hd__inv_2_71/Y sky130_fd_sc_hd__buf_12_138/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_61 VSS VDD sky130_fd_sc_hd__clkbuf_1_61/X sky130_fd_sc_hd__clkbuf_1_61/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_149 sky130_fd_sc_hd__inv_2_73/Y sky130_fd_sc_hd__buf_12_236/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_72 VSS VDD sky130_fd_sc_hd__nand4_1_15/A sky130_fd_sc_hd__a22oi_1_83/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_83 VSS VDD sky130_fd_sc_hd__nand4_1_4/A sky130_fd_sc_hd__a22oi_2_5/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_94 VSS VDD sky130_fd_sc_hd__buf_12_11/A sky130_fd_sc_hd__ha_2_14/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_4_8 sky130_fd_sc_hd__clkbuf_4_8/X sky130_fd_sc_hd__nor3_2_2/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_1_305 sky130_fd_sc_hd__fa_2_266/B sky130_fd_sc_hd__ha_2_93/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_305/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_316 sky130_fd_sc_hd__fa_2_395/A sky130_fd_sc_hd__ha_2_114/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_316/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_327 sky130_fd_sc_hd__fa_2_566/B sky130_fd_sc_hd__fa_2_546/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_327/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_338 sky130_fd_sc_hd__fa_2_558/B sky130_fd_sc_hd__ha_2_119/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_338/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_349 sky130_fd_sc_hd__ha_2_132/A sky130_fd_sc_hd__fa_2_686/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_349/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_202 sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__o21ai_1_228/Y
+ sky130_fd_sc_hd__a21oi_1_202/Y sky130_fd_sc_hd__fa_2_1063/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_213 sky130_fd_sc_hd__fa_2_1054/A sky130_fd_sc_hd__o22ai_1_193/Y
+ sky130_fd_sc_hd__a21oi_1_213/Y sky130_fd_sc_hd__nor2_4_12/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_224 sky130_fd_sc_hd__nand2_1_333/A sky130_fd_sc_hd__o22ai_1_199/Y
+ sky130_fd_sc_hd__a21oi_1_224/Y sky130_fd_sc_hd__a211o_1_9/A1 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_235 sky130_fd_sc_hd__a21o_2_5/A2 sky130_fd_sc_hd__o21ai_1_271/Y
+ sky130_fd_sc_hd__a21oi_1_235/Y sky130_fd_sc_hd__fa_2_1080/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_2_20 sky130_fd_sc_hd__nor3_2_7/Y sky130_fd_sc_hd__a22oi_2_20/A2
+ sky130_fd_sc_hd__nor3_2_8/Y sky130_fd_sc_hd__a22oi_2_20/B2 sky130_fd_sc_hd__nand4_1_54/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__a21oi_1_246 sky130_fd_sc_hd__o21a_1_22/B1 sky130_fd_sc_hd__nor2_1_147/Y
+ sky130_fd_sc_hd__dfxtp_1_898/D sky130_fd_sc_hd__nor2_1_147/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_257 sky130_fd_sc_hd__nor3_1_38/B sky130_fd_sc_hd__nor2b_1_105/Y
+ sky130_fd_sc_hd__a21oi_1_257/Y sky130_fd_sc_hd__nor2b_1_104/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_268 sky130_fd_sc_hd__fa_2_1136/A sky130_fd_sc_hd__o22ai_1_243/Y
+ sky130_fd_sc_hd__a21oi_1_268/Y sky130_fd_sc_hd__clkinv_1_779/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_279 sky130_fd_sc_hd__nor3_1_38/A sky130_fd_sc_hd__o22ai_1_251/Y
+ sky130_fd_sc_hd__a21oi_1_279/Y sky130_fd_sc_hd__fa_2_1127/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_4_8 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkinv_4_8/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_8/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__buf_8_209 sky130_fd_sc_hd__buf_8_209/A sky130_fd_sc_hd__buf_8_209/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nand2_1_240 sky130_fd_sc_hd__o21ai_1_84/B1 sky130_fd_sc_hd__nor2_1_59/B
+ sky130_fd_sc_hd__nor2_1_59/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_251 sky130_fd_sc_hd__o21a_1_1/B1 sky130_fd_sc_hd__fa_2_990/A
+ sky130_fd_sc_hd__o21a_1_1/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_850 sky130_fd_sc_hd__nor2_1_151/B sky130_fd_sc_hd__fa_2_1153/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_850/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_262 sky130_fd_sc_hd__o211ai_1_5/C1 sky130_fd_sc_hd__a211o_1_6/A1
+ sky130_fd_sc_hd__nand2_1_262/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_861 sky130_fd_sc_hd__clkinv_1_861/Y sky130_fd_sc_hd__o21a_1_42/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_861/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_273 sky130_fd_sc_hd__nand2_1_273/Y sky130_fd_sc_hd__nor2_4_9/B
+ sky130_fd_sc_hd__nor2_1_74/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_872 sky130_fd_sc_hd__nor2_1_190/A sky130_fd_sc_hd__nor2_1_191/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_872/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_284 sky130_fd_sc_hd__nand2_1_284/Y sky130_fd_sc_hd__nor2_2_11/B
+ sky130_fd_sc_hd__nor2_2_11/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_883 sky130_fd_sc_hd__o22ai_1_287/A1 sky130_fd_sc_hd__nor2_1_211/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_883/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_295 sky130_fd_sc_hd__nand2_1_295/Y sky130_fd_sc_hd__nor2_1_111/B
+ sky130_fd_sc_hd__fa_2_1118/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_894 sky130_fd_sc_hd__o31ai_1_8/A3 sky130_fd_sc_hd__xnor2_1_2/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_894/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__mux2_2_1 VSS VDD sky130_fd_sc_hd__mux2_2_1/A1 sky130_fd_sc_hd__mux2_2_1/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_1/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__a21boi_0_1 sky130_fd_sc_hd__a21oi_1_126/Y sky130_fd_sc_hd__a21boi_0_1/Y
+ sky130_fd_sc_hd__fa_2_996/A sky130_fd_sc_hd__a21o_2_3/A2 VSS VDD VDD VSS sky130_fd_sc_hd__a21boi_0
Xsky130_fd_sc_hd__fa_2_1190 sky130_fd_sc_hd__xor2_1_186/B sky130_fd_sc_hd__mux2_2_127/A0
+ sky130_fd_sc_hd__fa_2_1190/A sky130_fd_sc_hd__fa_2_1190/B sky130_fd_sc_hd__fa_2_1190/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_9 sky130_fd_sc_hd__fa_2_0/A sky130_fd_sc_hd__fa_2_1/B sky130_fd_sc_hd__fa_2_9/A
+ sky130_fd_sc_hd__fa_2_9/B sky130_fd_sc_hd__fa_2_9/CIN VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a211o_1_15 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_161/A sky130_fd_sc_hd__nor2b_1_105/Y
+ sky130_fd_sc_hd__o22ai_1_237/Y sky130_fd_sc_hd__o21ai_1_316/Y sky130_fd_sc_hd__o22ai_1_236/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__a211o_1_26 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_268/A sky130_fd_sc_hd__o21ai_1_402/Y
+ sky130_fd_sc_hd__nor2_1_250/Y sky130_fd_sc_hd__nor2b_2_4/Y sky130_fd_sc_hd__o22ai_1_355/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__clkinv_1_102 sky130_fd_sc_hd__inv_2_66/A sky130_fd_sc_hd__buf_8_94/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_102/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_113 sky130_fd_sc_hd__bufinv_8_1/A sky130_fd_sc_hd__buf_8_101/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_113/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_124 sky130_fd_sc_hd__nor3_1_17/C sky130_fd_sc_hd__nor3_2_6/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_124/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_135 sky130_fd_sc_hd__clkinv_2_13/A sky130_fd_sc_hd__clkinv_1_135/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_135/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_146 sky130_fd_sc_hd__clkinv_1_167/A sky130_fd_sc_hd__clkinv_1_146/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_146/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_157 sky130_fd_sc_hd__inv_2_88/A sky130_fd_sc_hd__and2_2_1/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_157/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_168 sky130_fd_sc_hd__inv_2_99/A sky130_fd_sc_hd__clkinv_2_15/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_168/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_179 sky130_fd_sc_hd__buf_8_146/A sky130_fd_sc_hd__bufinv_8_7/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_179/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_15 sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__xor2_1_6/B
+ sky130_fd_sc_hd__nand3_4_1/B sky130_fd_sc_hd__dfxtp_1_12/Q sky130_fd_sc_hd__a22o_2_3/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_26 sky130_fd_sc_hd__nor2_4_4/Y sky130_fd_sc_hd__ha_2_78/A
+ sky130_fd_sc_hd__buf_2_238/A sky130_fd_sc_hd__a22o_1_26/B2 sky130_fd_sc_hd__a22o_2_6/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_37 sky130_fd_sc_hd__a22o_1_37/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_37/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__xnor2_1_32/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__o21ai_1_2 VSS VDD sky130_fd_sc_hd__nor3_2_1/A sky130_fd_sc_hd__nor2_1_2/Y
+ sky130_fd_sc_hd__nor3_1_3/A sky130_fd_sc_hd__o21ai_1_2/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a22o_1_48 sky130_fd_sc_hd__a22o_1_48/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_48/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__fa_2_954/SUM
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_59 sky130_fd_sc_hd__a22o_1_59/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_59/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__nor4_1_11/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__bufbuf_16_1 sky130_fd_sc_hd__buf_8_2/A sky130_fd_sc_hd__buf_6_14/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__nand4_1_9 sky130_fd_sc_hd__nand4_1_9/C sky130_fd_sc_hd__nand4_1_9/B
+ sky130_fd_sc_hd__nand4_1_9/Y sky130_fd_sc_hd__nand4_1_9/D sky130_fd_sc_hd__nand4_1_9/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nor2_1_240 sky130_fd_sc_hd__nor2_1_240/B sky130_fd_sc_hd__nor2_1_240/Y
+ sky130_fd_sc_hd__o21a_1_54/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_251 sky130_fd_sc_hd__nor2_1_251/B sky130_fd_sc_hd__nor2_1_251/Y
+ sky130_fd_sc_hd__nor2_1_251/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_2_5 sky130_fd_sc_hd__clkinv_2_5/Y sky130_fd_sc_hd__ha_2_39/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_5/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__nor2_1_262 sky130_fd_sc_hd__nor2_1_268/A sky130_fd_sc_hd__nor2_1_262/Y
+ sky130_fd_sc_hd__nor2_1_263/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_273 sky130_fd_sc_hd__nor2_1_273/B sky130_fd_sc_hd__o21a_1_60/A1
+ sky130_fd_sc_hd__nor2_1_273/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_284 sky130_fd_sc_hd__nor2_1_284/B sky130_fd_sc_hd__nor2_1_284/Y
+ sky130_fd_sc_hd__nor2_1_284/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_295 sky130_fd_sc_hd__nor2_1_295/B sky130_fd_sc_hd__nor2_1_295/Y
+ sky130_fd_sc_hd__fa_2_0/SUM VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_480 sky130_fd_sc_hd__buf_12_480/A sky130_fd_sc_hd__buf_12_480/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_491 sky130_fd_sc_hd__buf_12_491/A sky130_fd_sc_hd__buf_12_491/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_350 sky130_fd_sc_hd__fa_2_1064/A sky130_fd_sc_hd__o21a_1_9/A2
+ sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__nor2_2_12/Y sky130_fd_sc_hd__a22oi_1_350/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_361 sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__nor2_2_12/Y
+ sky130_fd_sc_hd__fa_2_1089/A sky130_fd_sc_hd__fa_2_1091/A sky130_fd_sc_hd__a22oi_1_361/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_372 sky130_fd_sc_hd__clkinv_1_779/Y sky130_fd_sc_hd__nor3_1_38/B
+ sky130_fd_sc_hd__fa_2_1128/A sky130_fd_sc_hd__fa_2_1129/A sky130_fd_sc_hd__a22oi_1_372/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_383 sky130_fd_sc_hd__fa_2_1181/A sky130_fd_sc_hd__nor2_1_224/Y
+ sky130_fd_sc_hd__nor2_1_222/Y sky130_fd_sc_hd__fa_2_1177/A sky130_fd_sc_hd__a22oi_1_383/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_394 sky130_fd_sc_hd__nor2_1_265/Y sky130_fd_sc_hd__nor2_1_267/Y
+ sky130_fd_sc_hd__fa_2_1250/A sky130_fd_sc_hd__fa_2_1246/A sky130_fd_sc_hd__a22oi_1_394/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nand2_1_16 sky130_fd_sc_hd__nor3_1_2/C sky130_fd_sc_hd__nor3_1_4/B
+ sky130_fd_sc_hd__nand2_1_19/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_27 sky130_fd_sc_hd__nor2_4_8/B sky130_fd_sc_hd__nor3_2_9/B
+ sky130_fd_sc_hd__nor3_2_8/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_680 sky130_fd_sc_hd__nor2_1_108/B sky130_fd_sc_hd__fa_2_1112/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_680/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_38 sky130_fd_sc_hd__nand2_1_38/Y sky130_fd_sc_hd__nand2_1_38/B
+ sky130_fd_sc_hd__a21oi_2_0/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_49 sky130_fd_sc_hd__nand2_1_49/Y sky130_fd_sc_hd__xor2_1_18/B
+ sky130_fd_sc_hd__maj3_1_2/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_691 sky130_fd_sc_hd__a32o_1_1/A3 sky130_fd_sc_hd__nor2_1_139/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_691/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_8_2 sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__nor2_8_2/A
+ sky130_fd_sc_hd__nor2_8_2/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_8
Xsky130_fd_sc_hd__sdlclkp_2_10 sky130_fd_sc_hd__conb_1_20/LO sky130_fd_sc_hd__clkinv_8_62/Y
+ sky130_fd_sc_hd__dfxtp_1_526/CLK sky130_fd_sc_hd__o21ai_1_32/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__xnor2_1_80 VSS VDD sky130_fd_sc_hd__xnor2_1_81/B sky130_fd_sc_hd__xnor2_1_80/Y
+ sky130_fd_sc_hd__xnor2_1_80/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_91 VSS VDD sky130_fd_sc_hd__xnor2_1_91/B sky130_fd_sc_hd__xnor2_1_91/Y
+ sky130_fd_sc_hd__fa_2_1139/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__dfxtp_1_805 VDD VSS sky130_fd_sc_hd__fa_2_1057/A sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__mux2_2_63/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_816 VDD VSS sky130_fd_sc_hd__fa_2_1068/A sky130_fd_sc_hd__clkinv_4_25/Y
+ sky130_fd_sc_hd__mux2_2_41/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_827 VDD VSS sky130_fd_sc_hd__fa_2_1101/A sky130_fd_sc_hd__clkinv_8_59/Y
+ sky130_fd_sc_hd__and2_0_310/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_838 VDD VSS sky130_fd_sc_hd__nand2_1_339/B sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__nor2b_1_103/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_849 VDD VSS sky130_fd_sc_hd__mux2_2_55/A1 sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__o21ai_1_166/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_403 VSS VDD sky130_fd_sc_hd__clkbuf_1_403/X sky130_fd_sc_hd__clkbuf_1_403/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_414 VSS VDD sky130_fd_sc_hd__clkbuf_1_414/X sky130_fd_sc_hd__clkbuf_1_414/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_425 VSS VDD sky130_fd_sc_hd__clkbuf_1_425/X sky130_fd_sc_hd__clkbuf_1_425/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_436 VSS VDD sky130_fd_sc_hd__clkbuf_1_436/X sky130_fd_sc_hd__clkbuf_1_436/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_447 VSS VDD sky130_fd_sc_hd__a22oi_2_21/A2 sky130_fd_sc_hd__clkbuf_1_447/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_458 VSS VDD sky130_fd_sc_hd__clkbuf_1_458/X sky130_fd_sc_hd__clkbuf_1_458/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_469 VSS VDD sky130_fd_sc_hd__clkbuf_1_469/X sky130_fd_sc_hd__clkbuf_1_469/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__nor2b_1_107 sky130_fd_sc_hd__nor3_1_38/Y sky130_fd_sc_hd__nor2b_1_107/Y
+ sky130_fd_sc_hd__buf_2_262/X VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_118 sky130_fd_sc_hd__o22ai_1_266/Y sky130_fd_sc_hd__nor2b_1_118/Y
+ sky130_fd_sc_hd__buf_2_262/X VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_129 sky130_fd_sc_hd__nor2_1_285/Y sky130_fd_sc_hd__nor2b_1_129/Y
+ sky130_fd_sc_hd__buf_2_262/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__buf_6_8 VDD VSS sky130_fd_sc_hd__buf_6_8/X sky130_fd_sc_hd__buf_6_8/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__clkinv_2_10 sky130_fd_sc_hd__clkinv_2_10/Y sky130_fd_sc_hd__clkinv_2_10/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_10/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_21 sky130_fd_sc_hd__buf_8_202/A sky130_fd_sc_hd__clkinv_2_21/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_21/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_32 sky130_fd_sc_hd__clkinv_4_22/A sky130_fd_sc_hd__clkinv_2_32/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_32/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_43 sky130_fd_sc_hd__buf_6_52/A sky130_fd_sc_hd__clkinv_2_43/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_43/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__o22ai_1_208 sky130_fd_sc_hd__nor2_2_13/B sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__o22ai_1_208/Y sky130_fd_sc_hd__a21oi_1_238/Y sky130_fd_sc_hd__a21boi_0_4/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__sdlclkp_4_6 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__clkinv_8_112/A
+ sky130_fd_sc_hd__dfxtp_1_26/CLK sky130_fd_sc_hd__nor3_1_2/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__o22ai_1_219 sky130_fd_sc_hd__nand2_1_358/Y sky130_fd_sc_hd__nand2_1_357/Y
+ sky130_fd_sc_hd__o22ai_1_219/Y sky130_fd_sc_hd__o22ai_1_232/A1 sky130_fd_sc_hd__a21o_2_10/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_1_9 sky130_fd_sc_hd__nor2_1_9/B sky130_fd_sc_hd__nor2_1_9/Y
+ sky130_fd_sc_hd__nor2_1_9/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_180 sky130_fd_sc_hd__clkbuf_1_351/X sky130_fd_sc_hd__clkbuf_1_353/X
+ sky130_fd_sc_hd__clkbuf_4_117/X sky130_fd_sc_hd__a22oi_1_180/A2 sky130_fd_sc_hd__nand4_1_40/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_191 sky130_fd_sc_hd__clkbuf_1_265/X sky130_fd_sc_hd__clkbuf_1_266/X
+ sky130_fd_sc_hd__clkbuf_1_271/X sky130_fd_sc_hd__a22oi_1_191/A2 sky130_fd_sc_hd__a22oi_1_191/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22o_4_0 sky130_fd_sc_hd__a22o_4_0/B1 sky130_fd_sc_hd__a22o_4_0/B2
+ sky130_fd_sc_hd__a22o_4_0/X sky130_fd_sc_hd__ha_2_88/A sky130_fd_sc_hd__or2_1_1/B
+ VSS VDD VSS VDD sky130_fd_sc_hd__a22o_4
Xsky130_fd_sc_hd__o21ai_1_402 VSS VDD sky130_fd_sc_hd__o22ai_1_361/A1 sky130_fd_sc_hd__o21a_1_55/A1
+ sky130_fd_sc_hd__a21oi_1_386/Y sky130_fd_sc_hd__o21ai_1_402/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_413 VSS VDD sky130_fd_sc_hd__o22ai_1_366/B1 sky130_fd_sc_hd__o21a_1_55/A1
+ sky130_fd_sc_hd__a21oi_1_397/Y sky130_fd_sc_hd__o21ai_1_413/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_424 VSS VDD sky130_fd_sc_hd__o22ai_1_372/B1 sky130_fd_sc_hd__o21a_1_55/A1
+ sky130_fd_sc_hd__a21oi_1_403/Y sky130_fd_sc_hd__o21ai_1_424/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_435 VSS VDD sky130_fd_sc_hd__nor2_1_257/A sky130_fd_sc_hd__o21a_1_55/X
+ sky130_fd_sc_hd__a211oi_1_31/Y sky130_fd_sc_hd__xor2_1_250/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_446 VSS VDD sky130_fd_sc_hd__nor2_1_290/Y sky130_fd_sc_hd__or3_1_5/C
+ sky130_fd_sc_hd__nor2_1_287/A sky130_fd_sc_hd__o21ai_1_446/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_457 VSS VDD sky130_fd_sc_hd__nor2_1_309/A sky130_fd_sc_hd__a21oi_1_458/Y
+ sky130_fd_sc_hd__a21oi_1_449/Y sky130_fd_sc_hd__xor2_1_311/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_468 VSS VDD sky130_fd_sc_hd__nor2_1_299/A sky130_fd_sc_hd__o21ai_1_468/A1
+ sky130_fd_sc_hd__a211oi_1_34/Y sky130_fd_sc_hd__xor2_1_316/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_479 VSS VDD sky130_fd_sc_hd__o22ai_1_433/A1 sky130_fd_sc_hd__nor2_1_280/B
+ sky130_fd_sc_hd__o21ai_1_479/B1 sky130_fd_sc_hd__o21ai_1_479/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_4_11 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__or2_0_7/A
+ sky130_fd_sc_hd__xor2_1_88/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__dfxtp_1_1008 VDD VSS sky130_fd_sc_hd__mux2_2_98/A0 sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__o22ai_1_231/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_17 VSS VDD sky130_fd_sc_hd__nor4_1_4/C sky130_fd_sc_hd__xor2_1_9/A
+ sky130_fd_sc_hd__nor4_1_4/B sky130_fd_sc_hd__o31ai_1_1/B1 VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_240 sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1235/B
+ sky130_fd_sc_hd__xor2_1_240/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_1019 VDD VSS sky130_fd_sc_hd__ha_2_146/A sky130_fd_sc_hd__dfxtp_1_1026/CLK
+ sky130_fd_sc_hd__o32ai_1_4/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_28 VSS VDD sky130_fd_sc_hd__a21oi_2_0/Y sky130_fd_sc_hd__o21ai_1_28/A1
+ sky130_fd_sc_hd__nand2_1_47/Y sky130_fd_sc_hd__o21ai_1_28/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_251 sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__xor2_1_251/X
+ sky130_fd_sc_hd__xor2_1_251/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o21ai_1_39 VSS VDD sky130_fd_sc_hd__o21ai_1_39/A2 sky130_fd_sc_hd__o21ai_1_39/A1
+ sky130_fd_sc_hd__o21ai_1_39/B1 sky130_fd_sc_hd__o21ai_1_39/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_602 VDD VSS sky130_fd_sc_hd__and2_0_212/A sky130_fd_sc_hd__dfxtp_1_606/CLK
+ sky130_fd_sc_hd__fa_2_1022/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_262 sky130_fd_sc_hd__xor2_1_267/B sky130_fd_sc_hd__fa_2_1252/B
+ sky130_fd_sc_hd__xor2_1_262/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_613 VDD VSS sky130_fd_sc_hd__fa_2_807/B sky130_fd_sc_hd__dfxtp_1_627/CLK
+ sky130_fd_sc_hd__o21a_1_7/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_273 sky130_fd_sc_hd__xor2_1_273/B sky130_fd_sc_hd__xor2_1_273/X
+ sky130_fd_sc_hd__xor2_1_274/X VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_624 VDD VSS sky130_fd_sc_hd__fa_2_834/A sky130_fd_sc_hd__dfxtp_1_627/CLK
+ sky130_fd_sc_hd__o21a_1_2/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_284 sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1287/B
+ sky130_fd_sc_hd__xor2_1_284/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_635 VDD VSS sky130_fd_sc_hd__fa_2_999/A sky130_fd_sc_hd__clkinv_8_44/Y
+ sky130_fd_sc_hd__mux2_2_36/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_295 sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1276/B
+ sky130_fd_sc_hd__xor2_1_295/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_646 VDD VSS sky130_fd_sc_hd__fa_2_1010/A sky130_fd_sc_hd__clkinv_8_44/Y
+ sky130_fd_sc_hd__mux2_2_12/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_657 VDD VSS sky130_fd_sc_hd__fa_2_974/A sky130_fd_sc_hd__clkinv_8_41/Y
+ sky130_fd_sc_hd__and2_0_288/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_668 VDD VSS sky130_fd_sc_hd__fa_2_985/A sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__mux2_2_17/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_679 VDD VSS sky130_fd_sc_hd__fa_2_1018/A sky130_fd_sc_hd__clkinv_8_59/Y
+ sky130_fd_sc_hd__and2_0_271/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_200 VSS VDD sky130_fd_sc_hd__clkbuf_1_200/X sky130_fd_sc_hd__clkbuf_1_200/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_211 VSS VDD sky130_fd_sc_hd__buf_8_96/A sky130_fd_sc_hd__buf_12_127/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_222 VSS VDD sky130_fd_sc_hd__buf_8_72/A sky130_fd_sc_hd__ha_2_44/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_233 VSS VDD sky130_fd_sc_hd__clkbuf_4_61/A sky130_fd_sc_hd__inv_12_0/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_244 VSS VDD sky130_fd_sc_hd__clkbuf_1_244/X sky130_fd_sc_hd__a22oi_1_102/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_255 VSS VDD sky130_fd_sc_hd__clkbuf_1_255/X sky130_fd_sc_hd__clkbuf_1_256/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_266 VSS VDD sky130_fd_sc_hd__clkbuf_1_266/X sky130_fd_sc_hd__nor3_2_5/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_277 VSS VDD sky130_fd_sc_hd__clkbuf_1_277/X sky130_fd_sc_hd__clkbuf_1_277/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_288 VSS VDD sky130_fd_sc_hd__clkbuf_1_288/X sky130_fd_sc_hd__clkbuf_1_288/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_299 VSS VDD sky130_fd_sc_hd__nand4_1_46/D sky130_fd_sc_hd__a22oi_1_203/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_507 sky130_fd_sc_hd__fa_2_509/CIN sky130_fd_sc_hd__fa_2_504/A
+ sky130_fd_sc_hd__fa_2_507/A sky130_fd_sc_hd__fa_2_507/B sky130_fd_sc_hd__fa_2_515/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_518 sky130_fd_sc_hd__fa_2_520/CIN sky130_fd_sc_hd__fa_2_513/A
+ sky130_fd_sc_hd__fa_2_518/A sky130_fd_sc_hd__fa_2_518/B sky130_fd_sc_hd__fa_2_518/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_529 sky130_fd_sc_hd__maj3_1_88/B sky130_fd_sc_hd__maj3_1_89/A
+ sky130_fd_sc_hd__fa_2_529/A sky130_fd_sc_hd__fa_2_529/B sky130_fd_sc_hd__fa_2_530/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_4_5 VDD VSS sky130_fd_sc_hd__buf_4_5/X sky130_fd_sc_hd__buf_4_5/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__and2_0_220 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_220/X sky130_fd_sc_hd__and2_0_235/B
+ sky130_fd_sc_hd__and2_0_220/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_231 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_231/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_848/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_242 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_242/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__o21ai_1_3/Y sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_253 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_253/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__xnor2_1_30/Y sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_264 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_264/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__fa_2_966/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_275 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_275/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__and2_0_275/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_286 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_286/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__fa_2_996/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_297 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_297/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_297/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__sdlclkp_2_3 sky130_fd_sc_hd__conb_1_9/LO sky130_fd_sc_hd__clkinv_8_9/Y
+ sky130_fd_sc_hd__dfxtp_1_143/CLK sky130_fd_sc_hd__or2_0_1/X VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__o21ai_1_210 VSS VDD sky130_fd_sc_hd__o21ai_1_210/A2 sky130_fd_sc_hd__o22ai_1_206/A1
+ sky130_fd_sc_hd__a22oi_1_348/Y sky130_fd_sc_hd__o21ai_1_210/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_221 VSS VDD sky130_fd_sc_hd__nor2_1_134/Y sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__a21oi_1_195/Y sky130_fd_sc_hd__xor2_1_125/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_232 VSS VDD sky130_fd_sc_hd__o21a_1_16/A2 sky130_fd_sc_hd__nor2_1_114/B
+ sky130_fd_sc_hd__a22oi_1_354/Y sky130_fd_sc_hd__o21ai_1_232/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_50 sky130_fd_sc_hd__nand4_1_7/D sky130_fd_sc_hd__a22oi_1_52/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_243 VSS VDD sky130_fd_sc_hd__a21oi_1_226/Y sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__nand2_1_330/Y sky130_fd_sc_hd__xor2_1_92/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_61 sky130_fd_sc_hd__clkbuf_4_61/X sky130_fd_sc_hd__clkbuf_4_61/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_254 VSS VDD sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__nor2_1_140/B
+ sky130_fd_sc_hd__nand2_1_335/Y sky130_fd_sc_hd__o21ai_1_254/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_72 sky130_fd_sc_hd__clkbuf_4_72/X sky130_fd_sc_hd__nor3_1_13/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_265 VSS VDD sky130_fd_sc_hd__o21ai_1_265/A2 sky130_fd_sc_hd__o22ai_1_206/A1
+ sky130_fd_sc_hd__a22oi_1_362/Y sky130_fd_sc_hd__o21ai_1_265/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_83 sky130_fd_sc_hd__clkbuf_4_83/X sky130_fd_sc_hd__clkbuf_4_83/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_276 VSS VDD sky130_fd_sc_hd__nor2_1_161/Y sky130_fd_sc_hd__or3_1_2/C
+ sky130_fd_sc_hd__xnor2_1_93/Y sky130_fd_sc_hd__o21ai_1_276/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_94 sky130_fd_sc_hd__buf_2_39/A sky130_fd_sc_hd__inv_2_48/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_287 VSS VDD sky130_fd_sc_hd__xor2_1_140/X sky130_fd_sc_hd__xnor2_1_3/Y
+ sky130_fd_sc_hd__xnor2_1_93/Y sky130_fd_sc_hd__o21ai_1_287/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_298 VSS VDD sky130_fd_sc_hd__nor3_1_38/A sky130_fd_sc_hd__nor2_1_173/A
+ sky130_fd_sc_hd__nand2_1_380/Y sky130_fd_sc_hd__o21ai_1_298/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2b_2_5 sky130_fd_sc_hd__o32ai_1_11/A1 sky130_fd_sc_hd__nor2b_2_5/A
+ sky130_fd_sc_hd__nor2b_2_5/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_2
Xsky130_fd_sc_hd__fa_2_1008 sky130_fd_sc_hd__fa_2_1009/CIN sky130_fd_sc_hd__mux2_2_16/A0
+ sky130_fd_sc_hd__fa_2_1008/A sky130_fd_sc_hd__xor2_1_68/X sky130_fd_sc_hd__fa_2_1008/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1019 sky130_fd_sc_hd__fa_2_1020/CIN sky130_fd_sc_hd__and2_0_272/A
+ sky130_fd_sc_hd__fa_2_1019/A sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_1019/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_410 VDD VSS sky130_fd_sc_hd__ha_2_185/B sky130_fd_sc_hd__dfxtp_1_411/CLK
+ sky130_fd_sc_hd__and2_0_195/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_17 sky130_fd_sc_hd__inv_2_17/A sky130_fd_sc_hd__buf_8_6/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_421 VDD VSS sky130_fd_sc_hd__nor2_1_50/A sky130_fd_sc_hd__dfxtp_1_424/CLK
+ sky130_fd_sc_hd__and2_0_122/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_28 sky130_fd_sc_hd__inv_2_28/A sky130_fd_sc_hd__inv_2_28/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_432 VDD VSS sky130_fd_sc_hd__dfxtp_1_432/Q sky130_fd_sc_hd__dfxtp_1_433/CLK
+ sky130_fd_sc_hd__nand2_1_100/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_39 sky130_fd_sc_hd__inv_2_39/A sky130_fd_sc_hd__inv_2_39/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_443 VDD VSS sky130_fd_sc_hd__dfxtp_1_989/D sky130_fd_sc_hd__dfxtp_1_448/CLK
+ sky130_fd_sc_hd__nand2_1_78/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_454 VDD VSS sky130_fd_sc_hd__dfxtp_1_454/Q sky130_fd_sc_hd__dfxtp_1_454/CLK
+ sky130_fd_sc_hd__nand2_1_56/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_465 VDD VSS sky130_fd_sc_hd__clkbuf_1_9/A sky130_fd_sc_hd__dfxtp_1_472/CLK
+ sky130_fd_sc_hd__and2_0_146/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_476 VDD VSS sky130_fd_sc_hd__nor3_1_27/B sky130_fd_sc_hd__dfxtp_1_476/CLK
+ sky130_fd_sc_hd__and2_0_240/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_487 VDD VSS sky130_fd_sc_hd__nor2_1_37/B sky130_fd_sc_hd__dfxtp_1_488/CLK
+ sky130_fd_sc_hd__nor2b_1_71/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_498 VDD VSS sky130_fd_sc_hd__dfxtp_1_498/Q sky130_fd_sc_hd__dfxtp_1_502/CLK
+ sky130_fd_sc_hd__nor2b_1_83/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2b_1_13 sky130_fd_sc_hd__nand2b_1_13/Y sky130_fd_sc_hd__nor2_2_9/B
+ sky130_fd_sc_hd__nor2_4_9/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__fa_2_304 sky130_fd_sc_hd__fa_2_300/B sky130_fd_sc_hd__fa_2_303/B
+ sky130_fd_sc_hd__fa_2_304/A sky130_fd_sc_hd__fa_2_304/B sky130_fd_sc_hd__fa_2_304/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_315 sky130_fd_sc_hd__fa_2_312/CIN sky130_fd_sc_hd__fa_2_317/A
+ sky130_fd_sc_hd__fa_2_404/B sky130_fd_sc_hd__fa_2_413/A sky130_fd_sc_hd__fa_2_389/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_326 sky130_fd_sc_hd__maj3_1_78/B sky130_fd_sc_hd__maj3_1_79/A
+ sky130_fd_sc_hd__fa_2_360/B sky130_fd_sc_hd__fa_2_416/B sky130_fd_sc_hd__fa_2_326/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_337 sky130_fd_sc_hd__maj3_1_73/B sky130_fd_sc_hd__maj3_1_74/A
+ sky130_fd_sc_hd__fa_2_337/A sky130_fd_sc_hd__fa_2_337/B sky130_fd_sc_hd__fa_2_338/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_348 sky130_fd_sc_hd__fa_2_352/B sky130_fd_sc_hd__fa_2_348/SUM
+ sky130_fd_sc_hd__fa_2_348/A sky130_fd_sc_hd__fa_2_348/B sky130_fd_sc_hd__fa_2_348/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_359 sky130_fd_sc_hd__fa_2_357/B sky130_fd_sc_hd__fa_2_353/B
+ sky130_fd_sc_hd__fa_2_409/A sky130_fd_sc_hd__fa_2_401/A sky130_fd_sc_hd__ha_2_112/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_8_20 sky130_fd_sc_hd__clkinv_8_21/A sky130_fd_sc_hd__clkinv_8_20/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_20/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__diode_2_209 sig_frequency[7] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkinv_8_31 sky130_fd_sc_hd__clkinv_8_31/Y sky130_fd_sc_hd__clkinv_8_32/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_31/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_42 sky130_fd_sc_hd__clkinv_8_42/Y sky130_fd_sc_hd__clkinv_8_43/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_42/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_53 sky130_fd_sc_hd__clkinv_8_56/A sky130_fd_sc_hd__clkinv_8_53/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_64 sky130_fd_sc_hd__clkinv_8_64/Y sky130_fd_sc_hd__clkinv_8_65/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_64/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_75 sky130_fd_sc_hd__clkinv_8_75/Y sky130_fd_sc_hd__clkinv_8_75/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_75/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_86 sky130_fd_sc_hd__clkinv_8_87/A sky130_fd_sc_hd__clkinv_8_86/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_40 sky130_fd_sc_hd__buf_8_39/X sky130_fd_sc_hd__buf_12_40/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_8_97 sky130_fd_sc_hd__clkinv_8_98/A sky130_fd_sc_hd__clkinv_8_97/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_97/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_51 sky130_fd_sc_hd__buf_8_33/X sky130_fd_sc_hd__buf_12_89/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_62 sky130_fd_sc_hd__buf_4_14/X sky130_fd_sc_hd__buf_12_62/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_73 sky130_fd_sc_hd__buf_4_25/X sky130_fd_sc_hd__buf_8_59/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_84 sky130_fd_sc_hd__buf_8_58/X sky130_fd_sc_hd__buf_12_84/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_95 sky130_fd_sc_hd__buf_12_95/A sky130_fd_sc_hd__buf_12_95/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_2_2 VDD VSS sky130_fd_sc_hd__buf_6_2/A sky130_fd_sc_hd__buf_2_2/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1350 VDD VSS sky130_fd_sc_hd__fa_2_1309/A sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__mux2_2_224/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1361 VDD VSS sky130_fd_sc_hd__fa_2_1283/A sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__mux2_2_243/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1372 VDD VSS sky130_fd_sc_hd__fa_2_1311/B sky130_fd_sc_hd__clkinv_8_102/Y
+ sky130_fd_sc_hd__mux2_2_267/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1383 VDD VSS sky130_fd_sc_hd__fa_2_1322/A sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__mux2_2_244/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1394 VDD VSS sky130_fd_sc_hd__mux2_2_261/A0 sky130_fd_sc_hd__clkinv_8_75/Y
+ sky130_fd_sc_hd__nor2_1_287/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_12_309 sky130_fd_sc_hd__buf_8_165/X sky130_fd_sc_hd__buf_8_172/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__fa_2_860 sky130_fd_sc_hd__fa_2_859/CIN sky130_fd_sc_hd__fa_2_860/SUM
+ sky130_fd_sc_hd__fa_2_860/A sky130_fd_sc_hd__fa_2_860/B sky130_fd_sc_hd__fa_2_860/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_871 sky130_fd_sc_hd__fa_2_870/CIN sky130_fd_sc_hd__fa_2_871/SUM
+ sky130_fd_sc_hd__fa_2_871/A sky130_fd_sc_hd__fa_2_871/B sky130_fd_sc_hd__fa_2_871/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_882 sky130_fd_sc_hd__fa_2_881/CIN sky130_fd_sc_hd__nand2_1_42/B
+ sky130_fd_sc_hd__ha_2_153/A sky130_fd_sc_hd__fa_2_882/B sky130_fd_sc_hd__fa_2_882/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_893 sky130_fd_sc_hd__fa_2_892/CIN sky130_fd_sc_hd__fa_2_893/SUM
+ sky130_fd_sc_hd__fa_2_893/A sky130_fd_sc_hd__fa_2_893/B sky130_fd_sc_hd__fa_2_893/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_2 sky130_fd_sc_hd__inv_2_2/A sky130_fd_sc_hd__inv_2_2/Y VDD
+ VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__nor3_2_4 sky130_fd_sc_hd__nor3_2_4/C sky130_fd_sc_hd__nor3_2_4/Y
+ sky130_fd_sc_hd__nor3_2_4/A sky130_fd_sc_hd__nor3_2_4/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_2
Xsky130_fd_sc_hd__clkinv_1_509 sky130_fd_sc_hd__o21ai_1_76/A1 sky130_fd_sc_hd__o21ai_1_83/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_509/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_12 sky130_fd_sc_hd__nor2_1_12/B sky130_fd_sc_hd__nor2_1_12/Y
+ sky130_fd_sc_hd__xor2_1_19/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_23 sky130_fd_sc_hd__nor2_1_23/B sky130_fd_sc_hd__nor2_1_23/Y
+ sky130_fd_sc_hd__nor2_1_23/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_34 sky130_fd_sc_hd__nor2_1_34/B sky130_fd_sc_hd__nor2_1_34/Y
+ sky130_fd_sc_hd__nor4_1_8/C VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_45 sky130_fd_sc_hd__nor2_1_45/B sky130_fd_sc_hd__nor2_1_45/Y
+ sky130_fd_sc_hd__nor2_1_52/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_56 sky130_fd_sc_hd__nor2_1_56/B sky130_fd_sc_hd__nor2_1_56/Y
+ sky130_fd_sc_hd__nor2_1_56/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_160 VSS VDD sky130_fd_sc_hd__mux2_2_160/A1 sky130_fd_sc_hd__mux2_2_160/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_160/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_67 sky130_fd_sc_hd__nor2_1_67/B sky130_fd_sc_hd__o21a_1_5/A1
+ sky130_fd_sc_hd__nor2_1_67/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_171 VSS VDD sky130_fd_sc_hd__mux2_2_171/A1 sky130_fd_sc_hd__mux2_2_171/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_171/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_78 sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_1_78/Y
+ sky130_fd_sc_hd__nor2_1_78/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_182 VSS VDD sky130_fd_sc_hd__mux2_2_182/A1 sky130_fd_sc_hd__mux2_2_182/A0
+ sky130_fd_sc_hd__nor2_8_1/A sky130_fd_sc_hd__mux2_2_182/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_89 sky130_fd_sc_hd__or2_0_6/B sky130_fd_sc_hd__nor2_1_89/Y
+ sky130_fd_sc_hd__nor2_1_89/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_193 VSS VDD sky130_fd_sc_hd__mux2_2_193/A1 sky130_fd_sc_hd__mux2_2_193/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_193/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_sram_2kbyte_1rw1r_32x512_8_8 sky130_fd_sc_hd__clkbuf_4_102/X sky130_fd_sc_hd__clkbuf_4_103/X
+ sky130_fd_sc_hd__clkbuf_4_104/X sky130_fd_sc_hd__clkbuf_4_105/X sky130_fd_sc_hd__inv_8_0/Y
+ sky130_fd_sc_hd__buf_6_88/X sky130_fd_sc_hd__buf_2_285/A sky130_fd_sc_hd__buf_6_89/X
+ sky130_fd_sc_hd__clkbuf_4_227/A sky130_fd_sc_hd__buf_6_84/X sky130_fd_sc_hd__buf_4_122/X
+ sky130_fd_sc_hd__buf_4_121/X sky130_fd_sc_hd__buf_6_85/X sky130_fd_sc_hd__nand2_1_566/B
+ sky130_fd_sc_hd__nand2_1_567/B sky130_fd_sc_hd__clkbuf_4_109/X sky130_fd_sc_hd__clkbuf_4_102/X
+ sky130_fd_sc_hd__clkbuf_4_103/X sky130_fd_sc_hd__clkbuf_4_104/X sky130_fd_sc_hd__clkbuf_4_105/X
+ sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__buf_6_88/X sky130_fd_sc_hd__buf_2_285/X
+ sky130_fd_sc_hd__buf_6_89/X sky130_fd_sc_hd__clkbuf_4_227/X sky130_fd_sc_hd__buf_6_84/X
+ sky130_fd_sc_hd__buf_4_122/X sky130_fd_sc_hd__buf_4_121/X sky130_fd_sc_hd__buf_6_85/X
+ sky130_fd_sc_hd__nand2_1_566/B sky130_fd_sc_hd__nand2_1_567/B sky130_fd_sc_hd__clkbuf_4_109/X
+ sky130_fd_sc_hd__buf_12_366/X sky130_fd_sc_hd__buf_8_174/X sky130_fd_sc_hd__buf_12_344/X
+ sky130_fd_sc_hd__buf_12_356/X sky130_fd_sc_hd__buf_12_323/X sky130_fd_sc_hd__buf_12_292/X
+ sky130_fd_sc_hd__buf_12_353/X sky130_fd_sc_hd__buf_12_313/X sky130_fd_sc_hd__buf_12_302/X
+ sky130_fd_sc_hd__buf_12_365/X sky130_fd_sc_hd__buf_12_267/X sky130_fd_sc_hd__buf_12_321/X
+ sky130_fd_sc_hd__buf_12_278/X sky130_fd_sc_hd__buf_12_299/X sky130_fd_sc_hd__buf_12_290/X
+ sky130_fd_sc_hd__buf_12_310/X sky130_fd_sc_hd__buf_12_364/X sky130_fd_sc_hd__buf_12_367/X
+ sky130_fd_sc_hd__clkbuf_1_322/X sky130_fd_sc_hd__buf_2_125/X sky130_fd_sc_hd__clkbuf_1_322/X
+ sky130_fd_sc_hd__clkinv_2_19/Y sky130_fd_sc_hd__clkinv_8_129/Y sky130_fd_sc_hd__buf_8_177/X
+ sky130_fd_sc_hd__buf_8_178/X sky130_fd_sc_hd__buf_12_371/X sky130_fd_sc_hd__buf_12_361/X
+ sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[0] sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[1]
+ sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[2] sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[3]
+ sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[4] sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[5]
+ sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[6] sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[7]
+ sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[8] sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[9]
+ sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[10] sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[11]
+ sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[12] sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[13]
+ sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[14] sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[15]
+ sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[16] sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[17]
+ sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[18] sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[19]
+ sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[20] sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[21]
+ sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[22] sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[23]
+ sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[24] sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[25]
+ sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[26] sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[27]
+ sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[28] sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[29]
+ sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[30] sky130_sram_2kbyte_1rw1r_32x512_8_8/dout0[31]
+ sky130_fd_sc_hd__a22oi_1_209/B2 sky130_fd_sc_hd__a22oi_1_205/B2 sky130_fd_sc_hd__a22oi_1_201/B2
+ sky130_fd_sc_hd__a22oi_1_197/B2 sky130_fd_sc_hd__a22oi_1_193/B2 sky130_fd_sc_hd__a22oi_1_189/B2
+ sky130_fd_sc_hd__a22oi_1_185/B2 sky130_fd_sc_hd__a22oi_1_181/B2 sky130_fd_sc_hd__a22oi_1_177/B2
+ sky130_fd_sc_hd__a22oi_1_173/B2 sky130_fd_sc_hd__a22oi_1_169/B2 sky130_fd_sc_hd__a22oi_1_165/B2
+ sky130_fd_sc_hd__a22oi_1_161/B2 sky130_fd_sc_hd__a22oi_1_157/B2 sky130_fd_sc_hd__a22oi_1_153/B2
+ sky130_fd_sc_hd__a22oi_1_149/B2 sky130_fd_sc_hd__clkbuf_4_122/A sky130_fd_sc_hd__clkbuf_4_123/A
+ sky130_fd_sc_hd__clkbuf_4_124/A sky130_fd_sc_hd__clkbuf_4_125/A sky130_fd_sc_hd__clkbuf_4_126/A
+ sky130_fd_sc_hd__clkbuf_4_127/A sky130_fd_sc_hd__clkbuf_4_128/A sky130_fd_sc_hd__clkbuf_4_129/A
+ sky130_fd_sc_hd__clkbuf_4_130/A sky130_fd_sc_hd__clkbuf_4_131/A sky130_fd_sc_hd__clkbuf_4_132/A
+ sky130_fd_sc_hd__clkbuf_4_133/A sky130_fd_sc_hd__clkbuf_4_134/A sky130_fd_sc_hd__clkbuf_4_135/A
+ sky130_fd_sc_hd__clkbuf_4_136/A sky130_fd_sc_hd__clkbuf_4_137/A VDD VSS sky130_sram_2kbyte_1rw1r_32x512_8
Xsky130_fd_sc_hd__a21oi_1_406 sky130_fd_sc_hd__o21ai_1_430/Y sky130_fd_sc_hd__o21ai_1_425/Y
+ sky130_fd_sc_hd__a21oi_1_406/Y sky130_fd_sc_hd__nor2b_1_119/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_417 sky130_fd_sc_hd__clkinv_1_946/Y sky130_fd_sc_hd__o22ai_1_377/Y
+ sky130_fd_sc_hd__a21oi_1_417/Y sky130_fd_sc_hd__fa_2_1257/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_428 sky130_fd_sc_hd__nor2_1_276/A sky130_fd_sc_hd__nor2_1_276/Y
+ sky130_fd_sc_hd__a21oi_1_428/Y sky130_fd_sc_hd__nor2_1_276/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_439 sky130_fd_sc_hd__or3_1_5/C sky130_fd_sc_hd__o21ai_1_446/Y
+ sky130_fd_sc_hd__a21oi_1_439/Y sky130_fd_sc_hd__nor2_1_290/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_8_108 sky130_fd_sc_hd__clkinv_4_55/A sky130_fd_sc_hd__clkinv_8_114/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_108/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_119 sky130_fd_sc_hd__clkinv_8_120/A sky130_fd_sc_hd__clkinv_8_89/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_119/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__maj3_1_120 sky130_fd_sc_hd__maj3_1_121/X sky130_fd_sc_hd__maj3_1_120/X
+ sky130_fd_sc_hd__maj3_1_120/B sky130_fd_sc_hd__maj3_1_120/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_400 sky130_fd_sc_hd__nor2_1_191/A sky130_fd_sc_hd__fa_2_1175/A
+ sky130_fd_sc_hd__fa_2_1174/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_131 sky130_fd_sc_hd__maj3_1_132/X sky130_fd_sc_hd__maj3_1_131/X
+ sky130_fd_sc_hd__maj3_1_131/B sky130_fd_sc_hd__maj3_1_131/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_411 sky130_fd_sc_hd__nand2_1_411/Y sky130_fd_sc_hd__xor2_1_185/B
+ sky130_fd_sc_hd__o31ai_1_8/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_142 sky130_fd_sc_hd__maj3_1_143/X sky130_fd_sc_hd__maj3_1_142/X
+ sky130_fd_sc_hd__maj3_1_142/B sky130_fd_sc_hd__maj3_1_142/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_422 sky130_fd_sc_hd__nor2_1_210/B sky130_fd_sc_hd__nand2_1_422/B
+ sky130_fd_sc_hd__nor2_1_211/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_153 sky130_fd_sc_hd__maj3_1_154/X sky130_fd_sc_hd__maj3_1_153/X
+ sky130_fd_sc_hd__maj3_1_153/B sky130_fd_sc_hd__maj3_1_153/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_433 sky130_fd_sc_hd__nand2_1_433/Y sky130_fd_sc_hd__nor2b_1_112/Y
+ sky130_fd_sc_hd__o21ai_1_355/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_380 sky130_fd_sc_hd__a21oi_1_437/Y sky130_fd_sc_hd__nand2_1_497/B
+ sky130_fd_sc_hd__o22ai_1_380/Y sky130_fd_sc_hd__nor3_1_41/C sky130_fd_sc_hd__o32ai_1_11/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_444 sky130_fd_sc_hd__o32ai_1_8/A3 sky130_fd_sc_hd__nor2_4_18/B
+ sky130_fd_sc_hd__nor2_4_18/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_391 sky130_fd_sc_hd__nand2_1_514/Y sky130_fd_sc_hd__nand2_1_513/Y
+ sky130_fd_sc_hd__o22ai_1_391/Y sky130_fd_sc_hd__nand2_1_528/B sky130_fd_sc_hd__o21ai_1_444/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_455 sky130_fd_sc_hd__o21a_1_51/B1 sky130_fd_sc_hd__fa_2_1254/A
+ sky130_fd_sc_hd__o21a_1_51/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_466 sky130_fd_sc_hd__nand2_1_466/Y sky130_fd_sc_hd__inv_2_139/Y
+ sky130_fd_sc_hd__nand2_1_466/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_477 sky130_fd_sc_hd__nand2_1_477/Y sky130_fd_sc_hd__xor2_1_254/A
+ sky130_fd_sc_hd__nor2_1_267/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_488 sky130_fd_sc_hd__nand2_1_488/Y sky130_fd_sc_hd__nand2_1_491/B
+ sky130_fd_sc_hd__o21ai_1_431/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_499 sky130_fd_sc_hd__o21a_1_57/B1 sky130_fd_sc_hd__fa_2_1289/A
+ sky130_fd_sc_hd__o21a_1_57/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_13 sky130_fd_sc_hd__ha_2_24/SUM sky130_fd_sc_hd__nor2b_1_13/Y
+ sky130_fd_sc_hd__or2_0_1/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_24 sky130_fd_sc_hd__nor2_4_1/Y sky130_fd_sc_hd__and2_0_61/A
+ sky130_fd_sc_hd__ha_2_59/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_35 sky130_fd_sc_hd__ha_2_69/SUM sky130_fd_sc_hd__nor2b_1_35/Y
+ sky130_fd_sc_hd__or2_0_2/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1002 sky130_fd_sc_hd__nor2_1_230/B sky130_fd_sc_hd__fa_2_1233/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1002/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_46 sky130_fd_sc_hd__ha_2_82/SUM sky130_fd_sc_hd__nor2b_1_46/Y
+ sky130_fd_sc_hd__or2_0_3/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1013 sky130_fd_sc_hd__o22ai_1_376/A1 sky130_fd_sc_hd__nor2_1_267/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1013/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_57 sky130_fd_sc_hd__nor2b_1_85/A sky130_fd_sc_hd__nor2b_1_57/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1024 sky130_fd_sc_hd__nor2_1_238/B sky130_fd_sc_hd__fa_2_1251/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1024/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_68 sky130_fd_sc_hd__nand2_1_223/A sky130_fd_sc_hd__nor2b_1_68/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1035 sky130_fd_sc_hd__o22ai_1_436/A2 sky130_fd_sc_hd__nor3_1_41/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1035/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1046 sky130_fd_sc_hd__nor2_1_283/A sky130_fd_sc_hd__nor2_1_284/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1046/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_79 sky130_fd_sc_hd__o21ai_1_35/A1 sky130_fd_sc_hd__nor2b_1_79/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1057 sky130_fd_sc_hd__nor2_1_287/A sky130_fd_sc_hd__nor2_1_286/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1057/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1068 sky130_fd_sc_hd__nand2_1_526/B sky130_fd_sc_hd__fa_2_1/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1068/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xnor2_1_9 VSS VDD sky130_fd_sc_hd__xnor2_1_9/B sky130_fd_sc_hd__xnor2_1_9/Y
+ sky130_fd_sc_hd__xnor2_1_9/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_1079 sky130_fd_sc_hd__nor2_1_303/A sky130_fd_sc_hd__fa_2_1290/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1079/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_240 VDD VSS sky130_fd_sc_hd__fa_2_869/A sky130_fd_sc_hd__dfxtp_1_277/CLK
+ sky130_fd_sc_hd__and2_0_182/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_251 VDD VSS sky130_fd_sc_hd__inv_2_45/A sky130_fd_sc_hd__dfxtp_1_262/CLK
+ sky130_fd_sc_hd__and2_0_203/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_262 VDD VSS sky130_fd_sc_hd__dfxtp_1_262/Q sky130_fd_sc_hd__dfxtp_1_262/CLK
+ sky130_fd_sc_hd__and2_0_225/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_273 VDD VSS sky130_fd_sc_hd__dfxtp_1_273/Q sky130_fd_sc_hd__dfxtp_1_463/CLK
+ sky130_fd_sc_hd__and2_0_211/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_284 VDD VSS sky130_fd_sc_hd__a22o_1_63/A1 sky130_fd_sc_hd__dfxtp_1_477/CLK
+ sky130_fd_sc_hd__nand2_1_141/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_295 VDD VSS sky130_fd_sc_hd__a22o_1_52/A1 sky130_fd_sc_hd__clkinv_4_31/Y
+ sky130_fd_sc_hd__nand2_1_119/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o22ai_1_4 sky130_fd_sc_hd__ha_2_99/A sky130_fd_sc_hd__fa_2_87/B
+ sky130_fd_sc_hd__fa_2_55/B sky130_fd_sc_hd__ha_2_99/B sky130_fd_sc_hd__fa_2_92/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_101 sky130_fd_sc_hd__fa_2_102/CIN sky130_fd_sc_hd__fa_2_95/A
+ sky130_fd_sc_hd__ha_2_95/B sky130_fd_sc_hd__fa_2_45/A sky130_fd_sc_hd__fa_2_92/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_112 sky130_fd_sc_hd__fa_2_114/B sky130_fd_sc_hd__fa_2_109/A
+ sky130_fd_sc_hd__fa_2_139/B sky130_fd_sc_hd__fa_2_112/B sky130_fd_sc_hd__ha_2_97/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_123 sky130_fd_sc_hd__fa_2_122/A sky130_fd_sc_hd__fa_2_118/A
+ sky130_fd_sc_hd__fa_2_81/B sky130_fd_sc_hd__fa_2_76/A sky130_fd_sc_hd__fa_2_92/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_134 sky130_fd_sc_hd__fa_2_133/B sky130_fd_sc_hd__fa_2_134/SUM
+ sky130_fd_sc_hd__fa_2_134/A sky130_fd_sc_hd__fa_2_134/B sky130_fd_sc_hd__fa_2_138/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_145 sky130_fd_sc_hd__fa_2_144/CIN sky130_fd_sc_hd__nor2_1_251/A
+ sky130_fd_sc_hd__fa_2_238/B sky130_fd_sc_hd__fa_2_145/B sky130_fd_sc_hd__fa_2_145/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_156 sky130_fd_sc_hd__fa_2_149/B sky130_fd_sc_hd__fa_2_148/B
+ sky130_fd_sc_hd__fa_2_2/A sky130_fd_sc_hd__fa_2_242/B sky130_fd_sc_hd__fa_2_250/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_167 sky130_fd_sc_hd__fa_2_161/A sky130_fd_sc_hd__fa_2_164/B
+ sky130_fd_sc_hd__fa_2_167/A sky130_fd_sc_hd__fa_2_167/B sky130_fd_sc_hd__fa_2_167/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_178 sky130_fd_sc_hd__maj3_1_50/B sky130_fd_sc_hd__maj3_1_51/A
+ sky130_fd_sc_hd__fa_2_178/A sky130_fd_sc_hd__fa_2_178/B sky130_fd_sc_hd__o22ai_1_13/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_189 sky130_fd_sc_hd__maj3_1_46/B sky130_fd_sc_hd__maj3_1_47/A
+ sky130_fd_sc_hd__fa_2_189/A sky130_fd_sc_hd__fa_2_189/B sky130_fd_sc_hd__fa_2_190/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o22ai_1_11 sky130_fd_sc_hd__fa_2_261/A sky130_fd_sc_hd__fa_2_144/B
+ sky130_fd_sc_hd__xnor2_1_1/B sky130_fd_sc_hd__ha_2_97/A sky130_fd_sc_hd__fa_2_5/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_22 sky130_fd_sc_hd__fa_2_393/A sky130_fd_sc_hd__fa_2_395/A
+ sky130_fd_sc_hd__maj3_1_79/B sky130_fd_sc_hd__ha_2_114/A sky130_fd_sc_hd__fa_2_401/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_140 VDD VSS sky130_fd_sc_hd__buf_2_140/X sky130_fd_sc_hd__buf_2_140/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_33 sky130_fd_sc_hd__ha_2_123/B sky130_fd_sc_hd__fa_2_551/A
+ sky130_fd_sc_hd__o22ai_1_33/Y sky130_fd_sc_hd__ha_2_119/B sky130_fd_sc_hd__fa_2_555/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_151 VDD VSS sky130_fd_sc_hd__buf_6_54/A sky130_fd_sc_hd__buf_6_53/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_44 sky130_fd_sc_hd__fa_2_659/A sky130_fd_sc_hd__ha_2_128/A
+ sky130_fd_sc_hd__fa_2_638/A sky130_fd_sc_hd__ha_2_133/B sky130_fd_sc_hd__fa_2_683/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_162 VDD VSS sky130_fd_sc_hd__buf_2_162/X sky130_fd_sc_hd__buf_2_162/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_55 sky130_fd_sc_hd__ha_2_143/A sky130_fd_sc_hd__ha_2_142/B
+ sky130_fd_sc_hd__fa_2_810/B sky130_fd_sc_hd__fa_2_806/A sky130_fd_sc_hd__ha_2_141/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_173 VDD VSS sky130_fd_sc_hd__buf_2_173/X sky130_fd_sc_hd__buf_2_173/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_66 sky130_fd_sc_hd__o22ai_1_88/B1 sky130_fd_sc_hd__nand2_2_3/Y
+ sky130_fd_sc_hd__o22ai_1_66/Y sky130_fd_sc_hd__xnor2_1_43/Y sky130_fd_sc_hd__o22ai_1_80/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_184 VDD VSS sky130_fd_sc_hd__buf_2_184/X sky130_fd_sc_hd__buf_2_184/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_77 sky130_fd_sc_hd__o22ai_1_89/A1 sky130_fd_sc_hd__o22ai_1_88/B1
+ sky130_fd_sc_hd__o22ai_1_77/Y sky130_fd_sc_hd__xnor2_1_37/Y sky130_fd_sc_hd__o22ai_1_77/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_195 VDD VSS sky130_fd_sc_hd__buf_2_195/X sky130_fd_sc_hd__buf_2_195/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_88 sky130_fd_sc_hd__o22ai_1_89/A1 sky130_fd_sc_hd__o22ai_1_88/B1
+ sky130_fd_sc_hd__o22ai_1_88/Y sky130_fd_sc_hd__xnor2_1_59/Y sky130_fd_sc_hd__o22ai_1_88/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_99 sky130_fd_sc_hd__o22ai_1_99/A2 sky130_fd_sc_hd__a21oi_1_97/Y
+ sky130_fd_sc_hd__o22ai_1_99/Y sky130_fd_sc_hd__nor2_1_76/A sky130_fd_sc_hd__nor2_2_9/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__dfxtp_1_1180 VDD VSS sky130_fd_sc_hd__fa_2_933/A sky130_fd_sc_hd__dfxtp_1_1180/CLK
+ sky130_fd_sc_hd__a21oi_1_366/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1191 VDD VSS sky130_fd_sc_hd__xor2_1_26/B sky130_fd_sc_hd__clkinv_4_24/Y
+ sky130_fd_sc_hd__xnor2_1_97/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_4_13 VDD VSS sky130_fd_sc_hd__buf_4_13/X sky130_fd_sc_hd__buf_4_13/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_24 VDD VSS sky130_fd_sc_hd__buf_4_24/X sky130_fd_sc_hd__buf_8_21/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_35 VDD VSS sky130_fd_sc_hd__buf_4_35/X sky130_fd_sc_hd__buf_4_35/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_46 VDD VSS sky130_fd_sc_hd__buf_4_46/X sky130_fd_sc_hd__buf_8_78/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_57 VDD VSS sky130_fd_sc_hd__buf_4_57/X sky130_fd_sc_hd__buf_4_57/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_68 VDD VSS sky130_fd_sc_hd__buf_4_68/X sky130_fd_sc_hd__inv_2_83/Y
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_79 VDD VSS sky130_fd_sc_hd__buf_4_79/X sky130_fd_sc_hd__buf_4_79/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_12_106 sky130_fd_sc_hd__buf_12_86/X sky130_fd_sc_hd__buf_12_106/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_117 sky130_fd_sc_hd__buf_12_117/A sky130_fd_sc_hd__buf_12_117/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_40 VSS VDD sky130_fd_sc_hd__clkbuf_1_40/X sky130_fd_sc_hd__clkbuf_1_40/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_128 sky130_fd_sc_hd__buf_12_128/A sky130_fd_sc_hd__buf_12_148/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_51 VSS VDD sky130_fd_sc_hd__clkbuf_1_51/X sky130_fd_sc_hd__clkbuf_1_51/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_139 sky130_fd_sc_hd__inv_2_70/Y sky130_fd_sc_hd__buf_12_139/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_62 VSS VDD sky130_fd_sc_hd__clkbuf_1_62/X sky130_fd_sc_hd__clkbuf_1_62/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_73 VSS VDD sky130_fd_sc_hd__nand4_1_14/A sky130_fd_sc_hd__a22oi_1_79/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_84 VSS VDD sky130_fd_sc_hd__nand4_1_3/A sky130_fd_sc_hd__a22oi_1_42/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_690 sky130_fd_sc_hd__fa_2_692/CIN sky130_fd_sc_hd__fa_2_684/A
+ sky130_fd_sc_hd__fa_2_701/B sky130_fd_sc_hd__ha_2_134/A sky130_fd_sc_hd__fa_2_686/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_95 VSS VDD sky130_fd_sc_hd__buf_8_44/A sky130_fd_sc_hd__ha_2_18/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_4_9 sky130_fd_sc_hd__clkbuf_4_9/X sky130_fd_sc_hd__nor3_1_5/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_1_306 sky130_fd_sc_hd__fa_2_265/B sky130_fd_sc_hd__ha_2_91/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_306/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_317 sky130_fd_sc_hd__fa_2_422/B sky130_fd_sc_hd__ha_2_112/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_317/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_328 sky130_fd_sc_hd__fa_2_567/B sky130_fd_sc_hd__ha_2_125/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_328/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_339 sky130_fd_sc_hd__fa_2_683/B sky130_fd_sc_hd__fa_2_659/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_339/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_203 sky130_fd_sc_hd__clkinv_1_711/Y sky130_fd_sc_hd__o22ai_1_173/Y
+ sky130_fd_sc_hd__a21oi_1_203/Y sky130_fd_sc_hd__nand2_1_331/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_214 sky130_fd_sc_hd__clkinv_1_729/Y sky130_fd_sc_hd__clkinv_1_726/Y
+ sky130_fd_sc_hd__a21oi_1_214/Y sky130_fd_sc_hd__nand2_1_333/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_225 sky130_fd_sc_hd__a21o_2_5/X sky130_fd_sc_hd__o22ai_1_200/Y
+ sky130_fd_sc_hd__a21oi_1_225/Y sky130_fd_sc_hd__nand2_1_331/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_2_10 sky130_fd_sc_hd__nor2_4_5/Y sky130_fd_sc_hd__a22oi_2_10/A2
+ sky130_fd_sc_hd__a22oi_2_9/B1 sky130_fd_sc_hd__clkbuf_4_32/X sky130_fd_sc_hd__a22oi_2_10/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__a21oi_1_236 sky130_fd_sc_hd__clkinv_1_747/Y sky130_fd_sc_hd__o22ai_1_208/Y
+ sky130_fd_sc_hd__a21oi_1_236/Y sky130_fd_sc_hd__nand2_1_331/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_2_21 sky130_fd_sc_hd__buf_2_165/X sky130_fd_sc_hd__a22oi_2_21/A2
+ sky130_fd_sc_hd__nor2_4_7/Y sky130_fd_sc_hd__a22oi_2_21/B2 sky130_fd_sc_hd__nand4_1_55/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__a21oi_1_247 sky130_fd_sc_hd__nor2_1_148/A sky130_fd_sc_hd__o21a_1_22/A1
+ sky130_fd_sc_hd__dfxtp_1_896/D sky130_fd_sc_hd__nor2_1_148/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_258 sky130_fd_sc_hd__or3_1_2/C sky130_fd_sc_hd__o21ai_1_276/Y
+ sky130_fd_sc_hd__dfxtp_1_972/D sky130_fd_sc_hd__nor2_1_161/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_269 sky130_fd_sc_hd__nor2b_1_104/Y sky130_fd_sc_hd__o21ai_1_296/Y
+ sky130_fd_sc_hd__a21oi_1_269/Y sky130_fd_sc_hd__o21ai_1_305/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_4_9 sky130_fd_sc_hd__clkinv_4_9/A sky130_fd_sc_hd__clkinv_4_9/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_9/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__nand2_1_230 sky130_fd_sc_hd__xnor2_1_36/B sky130_fd_sc_hd__o21ai_1_80/B1
+ sky130_fd_sc_hd__o21ai_1_87/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_241 sky130_fd_sc_hd__o21ai_1_85/B1 sky130_fd_sc_hd__nor2_1_58/B
+ sky130_fd_sc_hd__nor2_1_58/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_840 sky130_fd_sc_hd__nor2_1_178/A sky130_fd_sc_hd__xor2_1_163/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_840/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_252 sky130_fd_sc_hd__o21a_1_2/B1 sky130_fd_sc_hd__fa_2_988/A
+ sky130_fd_sc_hd__o21a_1_2/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_851 sky130_fd_sc_hd__o21ai_1_328/A1 sky130_fd_sc_hd__fa_2_1154/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_851/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_263 sky130_fd_sc_hd__o211ai_1_5/B1 sky130_fd_sc_hd__nand2_1_282/B
+ sky130_fd_sc_hd__xor2_1_60/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_862 sky130_fd_sc_hd__o22ai_1_318/A2 sky130_fd_sc_hd__nor2_2_16/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_862/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_274 sky130_fd_sc_hd__nand2_1_274/Y sky130_fd_sc_hd__a211o_1_6/A1
+ sky130_fd_sc_hd__o21ai_1_136/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_873 sky130_fd_sc_hd__o32ai_1_4/A3 sky130_fd_sc_hd__fa_2_1192/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_873/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_285 sky130_fd_sc_hd__nand2_1_285/Y sky130_fd_sc_hd__nor2_1_141/B
+ sky130_fd_sc_hd__nor2_2_10/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_884 sky130_fd_sc_hd__o22ai_1_289/A1 sky130_fd_sc_hd__nor2_1_212/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_884/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_296 sky130_fd_sc_hd__nand2_1_296/Y sky130_fd_sc_hd__nor2_1_110/B
+ sky130_fd_sc_hd__fa_2_1116/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_895 sky130_fd_sc_hd__nand2_1_419/B sky130_fd_sc_hd__fa_2_286/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_895/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand4_1_80 sky130_fd_sc_hd__buf_2_252/A sky130_fd_sc_hd__or2_0_12/A
+ sky130_fd_sc_hd__nand4_1_80/Y sky130_fd_sc_hd__or2_0_10/A sky130_fd_sc_hd__or2_0_4/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__mux2_2_2 VSS VDD sky130_fd_sc_hd__mux2_2_2/A1 sky130_fd_sc_hd__xor2_1_32/X
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_2/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__a21boi_0_2 sky130_fd_sc_hd__a22oi_1_360/Y sky130_fd_sc_hd__o21a_1_16/B1
+ sky130_fd_sc_hd__xor2_1_88/A sky130_fd_sc_hd__nor2_2_12/Y VSS VDD VDD VSS sky130_fd_sc_hd__a21boi_0
Xsky130_fd_sc_hd__fa_2_1180 sky130_fd_sc_hd__fa_2_1181/CIN sky130_fd_sc_hd__mux2_2_150/A1
+ sky130_fd_sc_hd__fa_2_1180/A sky130_fd_sc_hd__fa_2_1180/B sky130_fd_sc_hd__fa_2_1180/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1191 sky130_fd_sc_hd__fa_2_1192/CIN sky130_fd_sc_hd__and2_0_325/A
+ sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__fa_2_1191/B sky130_fd_sc_hd__xor2_1_227/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a211o_1_16 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_157/A sky130_fd_sc_hd__o21ai_1_316/Y
+ sky130_fd_sc_hd__nor2_1_164/Y sky130_fd_sc_hd__nor2b_1_104/Y sky130_fd_sc_hd__o22ai_1_238/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__a211o_1_27 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_296/A sky130_fd_sc_hd__nor2b_1_126/Y
+ sky130_fd_sc_hd__o22ai_1_408/Y sky130_fd_sc_hd__o21ai_1_478/Y sky130_fd_sc_hd__o22ai_1_407/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__clkinv_1_103 sky130_fd_sc_hd__inv_2_67/A sky130_fd_sc_hd__ha_2_33/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_103/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_114 sky130_fd_sc_hd__clkinv_1_114/Y sky130_fd_sc_hd__bufinv_8_1/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_114/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_125 sky130_fd_sc_hd__nand3_2_4/C sky130_fd_sc_hd__nand3_2_3/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_125/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_136 sky130_fd_sc_hd__clkinv_2_14/A sky130_fd_sc_hd__clkinv_1_136/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_136/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_147 sky130_fd_sc_hd__clkinv_1_148/A sky130_fd_sc_hd__and2_1_4/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_147/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_158 sky130_fd_sc_hd__inv_2_89/A sky130_fd_sc_hd__and2_1_4/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_158/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_169 sky130_fd_sc_hd__clkinv_1_170/A sky130_fd_sc_hd__clkinv_1_169/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_169/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_16 sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__ha_2_60/A
+ sky130_fd_sc_hd__nand3_4_0/B sky130_fd_sc_hd__dfxtp_1_11/Q sky130_fd_sc_hd__a22o_2_3/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_27 sky130_fd_sc_hd__or2_1_1/B sky130_fd_sc_hd__xor2_1_8/B
+ sky130_fd_sc_hd__a22o_1_27/X sky130_fd_sc_hd__a22o_1_27/B2 sky130_fd_sc_hd__a22o_4_0/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_38 sky130_fd_sc_hd__a22o_1_38/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_38/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__fa_2_944/SUM
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_49 sky130_fd_sc_hd__a22o_1_49/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_49/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__fa_2_955/SUM
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__o21ai_1_3 VSS VDD sky130_fd_sc_hd__o21ai_1_4/Y sky130_fd_sc_hd__inv_4_1/A
+ sky130_fd_sc_hd__o21ai_1_3/B1 sky130_fd_sc_hd__o21ai_1_3/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__bufbuf_16_2 sky130_fd_sc_hd__buf_8_54/A sky130_fd_sc_hd__buf_6_15/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__nor2_1_230 sky130_fd_sc_hd__nor2_1_230/B sky130_fd_sc_hd__o21a_1_46/A1
+ sky130_fd_sc_hd__o21a_1_47/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_241 sky130_fd_sc_hd__nor2_1_241/B sky130_fd_sc_hd__o21a_1_54/A1
+ sky130_fd_sc_hd__nor2_1_241/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_252 sky130_fd_sc_hd__nor2_1_252/B sky130_fd_sc_hd__nor2_1_252/Y
+ sky130_fd_sc_hd__nor2_1_252/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_2_6 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkinv_2_6/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_6/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__nor2_1_263 sky130_fd_sc_hd__nor3_1_40/A sky130_fd_sc_hd__nor2_1_263/Y
+ sky130_fd_sc_hd__nor2_1_263/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_274 sky130_fd_sc_hd__nor2_1_274/B sky130_fd_sc_hd__nor2_1_274/Y
+ sky130_fd_sc_hd__o21a_1_61/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_285 sky130_fd_sc_hd__nor2_1_285/B sky130_fd_sc_hd__nor2_1_285/Y
+ sky130_fd_sc_hd__nor2_4_19/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_296 sky130_fd_sc_hd__nor2_1_296/B sky130_fd_sc_hd__nor2_1_296/Y
+ sky130_fd_sc_hd__fa_2_8/SUM VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_470 sky130_fd_sc_hd__buf_6_80/X sky130_fd_sc_hd__buf_12_470/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_481 sky130_fd_sc_hd__buf_12_481/A sky130_fd_sc_hd__buf_12_481/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_340 sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_2_7/Y
+ sky130_fd_sc_hd__fa_2_1000/A sky130_fd_sc_hd__fa_2_1001/A sky130_fd_sc_hd__a22oi_1_340/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_492 sky130_fd_sc_hd__buf_12_492/A sky130_fd_sc_hd__buf_12_517/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_351 sky130_fd_sc_hd__nor2_2_12/Y sky130_fd_sc_hd__fa_2_1067/A
+ sky130_fd_sc_hd__xor2_1_87/A sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__a22oi_1_351/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_362 sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__nor2_4_13/Y
+ sky130_fd_sc_hd__fa_2_1072/A sky130_fd_sc_hd__fa_2_1073/A sky130_fd_sc_hd__a22oi_1_362/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_373 sky130_fd_sc_hd__nor2_1_180/Y sky130_fd_sc_hd__nor2_1_182/Y
+ sky130_fd_sc_hd__fa_2_1131/A sky130_fd_sc_hd__fa_2_1127/A sky130_fd_sc_hd__a22oi_1_373/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_384 sky130_fd_sc_hd__clkinv_1_861/Y sky130_fd_sc_hd__nor3_1_39/B
+ sky130_fd_sc_hd__fa_2_1189/A sky130_fd_sc_hd__fa_2_1190/A sky130_fd_sc_hd__a22oi_1_384/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_395 sky130_fd_sc_hd__a22oi_1_400/B1 sky130_fd_sc_hd__nor3_1_41/B
+ sky130_fd_sc_hd__fa_2_1299/A sky130_fd_sc_hd__fa_2_1300/A sky130_fd_sc_hd__a22oi_1_395/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nand2_1_17 sky130_fd_sc_hd__nand3_1_17/C sky130_fd_sc_hd__nor3_1_4/B
+ sky130_fd_sc_hd__o21ai_1_0/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_670 sky130_fd_sc_hd__o21ai_1_194/A1 sky130_fd_sc_hd__nand2_1_296/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_670/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_28 sky130_fd_sc_hd__nor2_2_5/B sky130_fd_sc_hd__nor3_2_10/B
+ sky130_fd_sc_hd__nor3_2_10/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_681 sky130_fd_sc_hd__nor2_1_102/B sky130_fd_sc_hd__fa_2_1113/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_681/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_39 sky130_fd_sc_hd__nand2_1_39/Y sky130_fd_sc_hd__nand2_1_39/B
+ sky130_fd_sc_hd__a21oi_2_0/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_692 sky130_fd_sc_hd__o21ai_1_209/A2 sky130_fd_sc_hd__fa_2_1074/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_692/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__sdlclkp_2_11 sky130_fd_sc_hd__conb_1_24/LO sky130_fd_sc_hd__clkinv_8_96/A
+ sky130_fd_sc_hd__dfxtp_1_744/CLK sky130_fd_sc_hd__or2_0_8/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__xnor2_1_70 VSS VDD sky130_fd_sc_hd__xnor2_1_70/B sky130_fd_sc_hd__xnor2_1_70/Y
+ sky130_fd_sc_hd__nor2_1_94/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_81 VSS VDD sky130_fd_sc_hd__xnor2_1_81/B sky130_fd_sc_hd__xnor2_1_81/Y
+ sky130_fd_sc_hd__xnor2_1_81/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_92 VSS VDD sky130_fd_sc_hd__xnor2_1_92/B sky130_fd_sc_hd__xnor2_1_92/Y
+ sky130_fd_sc_hd__fa_2_1157/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__dfxtp_1_806 VDD VSS sky130_fd_sc_hd__fa_2_1058/A sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__mux2_2_61/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_817 VDD VSS sky130_fd_sc_hd__xor2_1_87/A sky130_fd_sc_hd__clkinv_4_25/Y
+ sky130_fd_sc_hd__mux2_2_40/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_828 VDD VSS sky130_fd_sc_hd__fa_2_1102/A sky130_fd_sc_hd__clkinv_8_54/Y
+ sky130_fd_sc_hd__and2_0_315/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_839 VDD VSS sky130_fd_sc_hd__nor2_4_12/B sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__nor2b_1_99/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_404 VSS VDD sky130_fd_sc_hd__clkbuf_1_404/X sky130_fd_sc_hd__clkbuf_1_404/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_415 VSS VDD sky130_fd_sc_hd__clkbuf_1_415/X sky130_fd_sc_hd__clkbuf_1_415/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_426 VSS VDD sky130_fd_sc_hd__clkbuf_1_426/X sky130_fd_sc_hd__clkbuf_1_426/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_437 VSS VDD sky130_fd_sc_hd__clkbuf_1_437/X sky130_fd_sc_hd__clkbuf_1_437/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_448 VSS VDD sky130_fd_sc_hd__clkbuf_1_448/X sky130_fd_sc_hd__clkbuf_1_448/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_459 VSS VDD sky130_fd_sc_hd__clkbuf_1_459/X sky130_fd_sc_hd__clkbuf_1_459/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__nor2b_1_108 sky130_fd_sc_hd__nor2_1_158/Y sky130_fd_sc_hd__nor2b_1_108/Y
+ sky130_fd_sc_hd__buf_2_262/X VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_119 sky130_fd_sc_hd__nor2b_2_4/A sky130_fd_sc_hd__nor2b_1_119/Y
+ sky130_fd_sc_hd__o32ai_1_8/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__buf_6_9 VDD VSS sky130_fd_sc_hd__buf_6_9/X sky130_fd_sc_hd__buf_6_9/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__clkinv_2_11 sky130_fd_sc_hd__clkinv_2_11/Y sky130_fd_sc_hd__clkinv_2_11/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_11/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_22 sky130_fd_sc_hd__clkinv_2_22/Y sky130_fd_sc_hd__nand3_1_39/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_22/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_33 sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__nor2_8_0/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_33/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkbuf_4_220 sky130_fd_sc_hd__a22o_1_8/A1 sig_amplitude[6] VSS VDD
+ VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_2_44 sky130_fd_sc_hd__clkinv_8_79/A clk VSS VDD VDD VSS VSS
+ sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__o22ai_1_209 sky130_fd_sc_hd__a21oi_1_257/Y sky130_fd_sc_hd__nand2_1_341/B
+ sky130_fd_sc_hd__o22ai_1_209/Y sky130_fd_sc_hd__nor3_1_38/C sky130_fd_sc_hd__o32ai_1_2/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__sdlclkp_4_7 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__clkinv_8_112/A
+ sky130_fd_sc_hd__dfxtp_1_29/CLK sky130_fd_sc_hd__nor3_1_2/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__a22oi_1_170 sky130_fd_sc_hd__clkbuf_1_264/X sky130_fd_sc_hd__nor2_2_3/Y
+ sky130_fd_sc_hd__a22oi_1_170/B2 sky130_fd_sc_hd__clkbuf_4_132/X sky130_fd_sc_hd__nand4_1_37/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_181 sky130_fd_sc_hd__clkbuf_4_111/X sky130_fd_sc_hd__clkbuf_4_112/X
+ sky130_fd_sc_hd__a22oi_1_181/B2 sky130_fd_sc_hd__clkbuf_1_289/X sky130_fd_sc_hd__a22oi_1_181/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_192 sky130_fd_sc_hd__clkbuf_1_351/X sky130_fd_sc_hd__clkbuf_1_353/X
+ sky130_fd_sc_hd__clkinv_2_10/Y sky130_fd_sc_hd__a22oi_1_192/A2 sky130_fd_sc_hd__nand4_1_43/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__o21ai_1_403 VSS VDD sky130_fd_sc_hd__nor2_1_267/A sky130_fd_sc_hd__a21oi_1_398/Y
+ sky130_fd_sc_hd__a21oi_1_389/Y sky130_fd_sc_hd__xor2_1_266/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_414 VSS VDD sky130_fd_sc_hd__nor2_1_257/A sky130_fd_sc_hd__o21ai_1_414/A1
+ sky130_fd_sc_hd__a211oi_1_27/Y sky130_fd_sc_hd__xor2_1_271/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_425 VSS VDD sky130_fd_sc_hd__o22ai_1_376/A1 sky130_fd_sc_hd__nor2_1_238/B
+ sky130_fd_sc_hd__o21ai_1_425/B1 sky130_fd_sc_hd__o21ai_1_425/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_436 VSS VDD sky130_fd_sc_hd__o22ai_1_375/A2 sky130_fd_sc_hd__o21ai_1_436/A1
+ sky130_fd_sc_hd__a21oi_1_417/Y sky130_fd_sc_hd__o21ai_1_436/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_447 VSS VDD sky130_fd_sc_hd__nor2_1_283/B sky130_fd_sc_hd__o22ai_1_436/A2
+ sky130_fd_sc_hd__a22oi_1_395/Y sky130_fd_sc_hd__o21ai_1_447/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_458 VSS VDD sky130_fd_sc_hd__nor2_1_301/B sky130_fd_sc_hd__nor2_1_299/A
+ sky130_fd_sc_hd__a21oi_1_450/Y sky130_fd_sc_hd__o21ai_1_458/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_469 VSS VDD sky130_fd_sc_hd__o22ai_1_432/A2 sky130_fd_sc_hd__nor2_1_274/B
+ sky130_fd_sc_hd__a21oi_1_459/Y sky130_fd_sc_hd__o21ai_1_469/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_4_12 sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__nor2_4_13/A
+ sky130_fd_sc_hd__nor2_4_12/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__xor2_1_230 sky130_fd_sc_hd__xor2_1_275/B sky130_fd_sc_hd__xor2_1_230/X
+ sky130_fd_sc_hd__xor2_1_275/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_1009 VDD VSS sky130_fd_sc_hd__mux2_2_95/A0 sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__o22ai_1_230/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_241 sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1234/B
+ sky130_fd_sc_hd__xor2_1_241/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o21ai_1_18 VSS VDD sky130_fd_sc_hd__a21oi_2_0/Y sky130_fd_sc_hd__maj3_1_0/C
+ sky130_fd_sc_hd__nand2_1_37/Y sky130_fd_sc_hd__o21ai_1_18/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_252 sky130_fd_sc_hd__xor2_1_252/B sky130_fd_sc_hd__xor2_1_252/X
+ sky130_fd_sc_hd__xor2_1_253/X VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o21ai_1_29 VSS VDD sky130_fd_sc_hd__xor2_1_18/B sky130_fd_sc_hd__maj3_1_2/X
+ sky130_fd_sc_hd__o21ai_1_29/B1 sky130_fd_sc_hd__o21ai_1_29/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_603 VDD VSS sky130_fd_sc_hd__and2_0_213/A sky130_fd_sc_hd__dfxtp_1_606/CLK
+ sky130_fd_sc_hd__fa_2_1023/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_263 sky130_fd_sc_hd__xor2_1_267/B sky130_fd_sc_hd__fa_2_1251/B
+ sky130_fd_sc_hd__xor2_1_263/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_614 VDD VSS sky130_fd_sc_hd__fa_2_812/B sky130_fd_sc_hd__dfxtp_1_627/CLK
+ sky130_fd_sc_hd__a21oi_1_79/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_274 sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__xor2_1_274/X
+ sky130_fd_sc_hd__nor2_8_1/B VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_625 VDD VSS sky130_fd_sc_hd__ha_2_145/A sky130_fd_sc_hd__dfxtp_1_626/CLK
+ sky130_fd_sc_hd__a21oi_1_73/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_285 sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1286/B
+ sky130_fd_sc_hd__xor2_1_285/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_636 VDD VSS sky130_fd_sc_hd__fa_2_1000/A sky130_fd_sc_hd__clkinv_8_44/Y
+ sky130_fd_sc_hd__mux2_2_34/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_296 sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__xor2_1_296/X
+ sky130_fd_sc_hd__xor2_1_296/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_647 VDD VSS sky130_fd_sc_hd__fa_2_1011/A sky130_fd_sc_hd__clkinv_8_44/Y
+ sky130_fd_sc_hd__mux2_2_10/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_658 VDD VSS sky130_fd_sc_hd__fa_2_975/A sky130_fd_sc_hd__clkinv_8_41/Y
+ sky130_fd_sc_hd__and2_0_289/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_669 VDD VSS sky130_fd_sc_hd__fa_2_986/A sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__mux2_2_15/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_201 VSS VDD sky130_fd_sc_hd__clkbuf_1_201/X sky130_fd_sc_hd__inv_2_46/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_212 VSS VDD sky130_fd_sc_hd__buf_12_129/A sky130_fd_sc_hd__buf_8_79/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_223 VSS VDD sky130_fd_sc_hd__buf_12_145/A sky130_fd_sc_hd__clkbuf_1_235/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_234 VSS VDD sky130_fd_sc_hd__buf_4_41/A sky130_fd_sc_hd__buf_12_152/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_245 VSS VDD sky130_fd_sc_hd__clkbuf_1_246/A sky130_fd_sc_hd__buf_4_55/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_256 VSS VDD sky130_fd_sc_hd__clkbuf_1_256/X sky130_fd_sc_hd__clkbuf_1_257/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_267 VSS VDD sky130_fd_sc_hd__clkbuf_1_267/X sky130_fd_sc_hd__clkbuf_1_267/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_278 VSS VDD sky130_fd_sc_hd__clkbuf_1_278/X sky130_fd_sc_hd__clkbuf_1_278/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_289 VSS VDD sky130_fd_sc_hd__clkbuf_1_289/X sky130_fd_sc_hd__clkbuf_1_289/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_508 sky130_fd_sc_hd__maj3_1_92/B sky130_fd_sc_hd__maj3_1_93/A
+ sky130_fd_sc_hd__fa_2_508/A sky130_fd_sc_hd__fa_2_508/B sky130_fd_sc_hd__fa_2_509/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_519 sky130_fd_sc_hd__maj3_1_90/B sky130_fd_sc_hd__maj3_1_91/A
+ sky130_fd_sc_hd__fa_2_519/A sky130_fd_sc_hd__fa_2_519/B sky130_fd_sc_hd__fa_2_520/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_90 VDD VSS sky130_fd_sc_hd__buf_2_90/X sky130_fd_sc_hd__buf_2_90/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_4_6 VDD VSS sky130_fd_sc_hd__buf_4_6/X sky130_fd_sc_hd__buf_4_6/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__and2_0_210 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_210/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_210/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_221 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_221/X sky130_fd_sc_hd__and2_0_235/B
+ sky130_fd_sc_hd__and2_0_221/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_232 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_232/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_849/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_243 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_243/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__and2_0_243/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_254 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_254/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__o31ai_1_3/Y sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_265 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_265/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__fa_2_965/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_276 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_276/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__fa_2_970/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_287 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_287/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__fa_2_997/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_298 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_298/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_298/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__sdlclkp_2_4 sky130_fd_sc_hd__conb_1_10/LO sky130_fd_sc_hd__clkinv_4_63/Y
+ sky130_fd_sc_hd__dfxtp_1_158/CLK sky130_fd_sc_hd__nand2b_1_1/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__o21ai_1_200 VSS VDD sky130_fd_sc_hd__xnor2_1_84/A sky130_fd_sc_hd__nor2_1_111/Y
+ sky130_fd_sc_hd__nand2_1_295/Y sky130_fd_sc_hd__xnor2_1_86/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_211 VSS VDD sky130_fd_sc_hd__a21oi_1_200/Y sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__nand2_1_317/Y sky130_fd_sc_hd__xor2_1_115/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_222 VSS VDD sky130_fd_sc_hd__o22ai_1_173/A2 sky130_fd_sc_hd__nor2_1_127/A
+ sky130_fd_sc_hd__nand2_1_321/Y sky130_fd_sc_hd__o21ai_1_222/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_40 sky130_fd_sc_hd__clkbuf_4_40/X sky130_fd_sc_hd__clkbuf_4_40/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_233 VSS VDD sky130_fd_sc_hd__o22ai_1_204/B1 sky130_fd_sc_hd__nand4_1_86/A
+ sky130_fd_sc_hd__a21oi_1_207/Y sky130_fd_sc_hd__o21ai_1_233/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_51 sky130_fd_sc_hd__nand4_1_6/D sky130_fd_sc_hd__a22oi_1_49/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_244 VSS VDD sky130_fd_sc_hd__nor2_1_127/A sky130_fd_sc_hd__a21oi_1_226/Y
+ sky130_fd_sc_hd__a21oi_1_214/Y sky130_fd_sc_hd__xor2_1_96/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_62 sky130_fd_sc_hd__clkbuf_4_64/A sky130_fd_sc_hd__dfxtp_1_252/Q
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_255 VSS VDD sky130_fd_sc_hd__nor2_1_136/A sky130_fd_sc_hd__o22ai_1_206/B1
+ sky130_fd_sc_hd__a22oi_1_358/Y sky130_fd_sc_hd__o21ai_1_255/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_73 sky130_fd_sc_hd__clkbuf_4_73/X sky130_fd_sc_hd__nor2_1_4/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_266 VSS VDD sky130_fd_sc_hd__o21ai_1_271/A2 sky130_fd_sc_hd__o22ai_1_206/B1
+ sky130_fd_sc_hd__a22oi_1_363/Y sky130_fd_sc_hd__a21o_2_5/B1 VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_84 sky130_fd_sc_hd__clkbuf_4_84/X sky130_fd_sc_hd__clkbuf_4_84/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_277 VSS VDD sky130_fd_sc_hd__nand2_1_367/B sky130_fd_sc_hd__a21o_2_6/B1
+ sky130_fd_sc_hd__o31ai_1_6/A2 sky130_fd_sc_hd__o21ai_1_277/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_95 sky130_fd_sc_hd__clkbuf_4_95/X sky130_fd_sc_hd__clkinv_1_76/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_288 VSS VDD sky130_fd_sc_hd__o22ai_1_244/A1 sky130_fd_sc_hd__nor2_1_182/A
+ sky130_fd_sc_hd__nand2_1_373/Y sky130_fd_sc_hd__xor2_1_165/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_299 VSS VDD sky130_fd_sc_hd__a222oi_1_7/Y sky130_fd_sc_hd__nor2_1_182/A
+ sky130_fd_sc_hd__a22oi_1_373/Y sky130_fd_sc_hd__o21ai_1_299/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__buf_8_190 sky130_fd_sc_hd__inv_2_105/Y sky130_fd_sc_hd__buf_8_190/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__fa_2_1009 sky130_fd_sc_hd__fa_2_1010/CIN sky130_fd_sc_hd__mux2_2_14/A0
+ sky130_fd_sc_hd__fa_2_1009/A sky130_fd_sc_hd__xor2_1_67/X sky130_fd_sc_hd__fa_2_1009/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_400 VDD VSS sky130_fd_sc_hd__nor2_1_58/A sky130_fd_sc_hd__dfxtp_1_424/CLK
+ sky130_fd_sc_hd__and2_0_148/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_411 VDD VSS sky130_fd_sc_hd__nor2_1_55/A sky130_fd_sc_hd__dfxtp_1_411/CLK
+ sky130_fd_sc_hd__and2_0_194/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_18 sky130_fd_sc_hd__inv_2_18/A sky130_fd_sc_hd__inv_2_18/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_422 VDD VSS sky130_fd_sc_hd__fa_2_1042/B sky130_fd_sc_hd__dfxtp_1_424/CLK
+ sky130_fd_sc_hd__and2_0_117/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_29 sky130_fd_sc_hd__inv_2_29/A sky130_fd_sc_hd__inv_2_29/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_433 VDD VSS sky130_fd_sc_hd__dfxtp_1_433/Q sky130_fd_sc_hd__dfxtp_1_433/CLK
+ sky130_fd_sc_hd__nand2_1_98/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_444 VDD VSS sky130_fd_sc_hd__dfxtp_1_990/D sky130_fd_sc_hd__dfxtp_1_448/CLK
+ sky130_fd_sc_hd__nand2_1_76/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_455 VDD VSS sky130_fd_sc_hd__xnor2_1_96/A sky130_fd_sc_hd__dfxtp_1_457/CLK
+ sky130_fd_sc_hd__nand2_1_54/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_466 VDD VSS sky130_fd_sc_hd__clkbuf_1_8/A sky130_fd_sc_hd__dfxtp_1_473/CLK
+ sky130_fd_sc_hd__and2_0_141/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_477 VDD VSS sky130_fd_sc_hd__a22o_1_65/A1 sky130_fd_sc_hd__dfxtp_1_477/CLK
+ sky130_fd_sc_hd__nand2_1_145/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_488 VDD VSS sky130_fd_sc_hd__nand3_1_48/C sky130_fd_sc_hd__dfxtp_1_488/CLK
+ sky130_fd_sc_hd__nor2b_1_70/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_499 VDD VSS sky130_fd_sc_hd__nor2b_1_87/A sky130_fd_sc_hd__dfxtp_1_502/CLK
+ sky130_fd_sc_hd__nor2b_1_64/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2b_1_14 sky130_fd_sc_hd__xnor2_1_63/B sky130_fd_sc_hd__ha_2_201/B
+ sky130_fd_sc_hd__ha_2_201/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__fa_2_305 sky130_fd_sc_hd__fa_2_302/B sky130_fd_sc_hd__fa_2_304/B
+ sky130_fd_sc_hd__ha_2_116/B sky130_fd_sc_hd__ha_2_113/B sky130_fd_sc_hd__fa_2_413/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_316 sky130_fd_sc_hd__fa_2_313/B sky130_fd_sc_hd__fa_2_317/CIN
+ sky130_fd_sc_hd__fa_2_316/A sky130_fd_sc_hd__fa_2_316/B sky130_fd_sc_hd__fa_2_316/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_327 sky130_fd_sc_hd__maj3_1_77/B sky130_fd_sc_hd__maj3_1_78/A
+ sky130_fd_sc_hd__fa_2_393/A sky130_fd_sc_hd__fa_2_327/B sky130_fd_sc_hd__fa_2_328/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_338 sky130_fd_sc_hd__fa_2_340/B sky130_fd_sc_hd__fa_2_338/SUM
+ sky130_fd_sc_hd__fa_2_404/B sky130_fd_sc_hd__fa_2_338/B sky130_fd_sc_hd__fa_2_338/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_349 sky130_fd_sc_hd__fa_2_353/CIN sky130_fd_sc_hd__fa_2_347/B
+ sky130_fd_sc_hd__fa_2_349/A sky130_fd_sc_hd__fa_2_349/B sky130_fd_sc_hd__fa_2_358/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_8_10 sky130_fd_sc_hd__clkinv_8_2/A sky130_fd_sc_hd__clkinv_4_7/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_10/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_21 sky130_fd_sc_hd__clkinv_8_22/A sky130_fd_sc_hd__clkinv_8_21/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_21/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_32 sky130_fd_sc_hd__clkinv_8_32/Y sky130_fd_sc_hd__clkinv_8_32/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_43 sky130_fd_sc_hd__clkinv_8_43/Y sky130_fd_sc_hd__clkinv_8_43/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_43/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_54 sky130_fd_sc_hd__clkinv_8_54/Y sky130_fd_sc_hd__clkinv_8_56/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_54/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_65 sky130_fd_sc_hd__clkinv_8_65/Y sky130_fd_sc_hd__clkinv_8_65/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_65/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_76 sky130_fd_sc_hd__clkinv_8_78/A sky130_fd_sc_hd__clkinv_8_76/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_76/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_30 sky130_fd_sc_hd__buf_8_43/X sky130_fd_sc_hd__buf_6_18/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_8_87 sky130_fd_sc_hd__clkinv_8_88/A sky130_fd_sc_hd__clkinv_8_87/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_87/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_41 sky130_fd_sc_hd__buf_8_50/X sky130_fd_sc_hd__buf_12_41/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_8_98 sky130_fd_sc_hd__clkinv_8_99/A sky130_fd_sc_hd__clkinv_8_98/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_98/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_52 sky130_fd_sc_hd__buf_8_35/X sky130_fd_sc_hd__buf_12_52/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_63 sky130_fd_sc_hd__buf_6_15/X sky130_fd_sc_hd__buf_12_99/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_74 sky130_fd_sc_hd__buf_4_17/X sky130_fd_sc_hd__buf_12_74/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_85 sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__buf_12_85/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_96 sky130_fd_sc_hd__buf_12_96/A sky130_fd_sc_hd__buf_12_96/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_2_3 VDD VSS sky130_fd_sc_hd__buf_4_5/A sky130_fd_sc_hd__buf_4_4/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1340 VDD VSS sky130_fd_sc_hd__fa_2_1299/A sky130_fd_sc_hd__clkinv_8_70/Y
+ sky130_fd_sc_hd__mux2_2_248/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1351 VDD VSS sky130_fd_sc_hd__fa_2_1310/A sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__mux2_2_222/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1362 VDD VSS sky130_fd_sc_hd__fa_2_1284/A sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__mux2_2_240/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1373 VDD VSS sky130_fd_sc_hd__fa_2_1312/A sky130_fd_sc_hd__clkinv_8_102/Y
+ sky130_fd_sc_hd__mux2_2_266/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1384 VDD VSS sky130_fd_sc_hd__fa_2_1323/A sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__mux2_2_241/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1395 VDD VSS sky130_fd_sc_hd__mux2_2_258/A0 sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__a21oi_1_438/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_850 sky130_fd_sc_hd__xnor2_1_9/B sky130_fd_sc_hd__fa_2_850/SUM
+ sky130_fd_sc_hd__fa_2_850/A sky130_fd_sc_hd__fa_2_850/B sky130_fd_sc_hd__fa_2_850/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_861 sky130_fd_sc_hd__fa_2_860/CIN sky130_fd_sc_hd__fa_2_861/SUM
+ sky130_fd_sc_hd__fa_2_861/A sky130_fd_sc_hd__fa_2_861/B sky130_fd_sc_hd__fa_2_861/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_872 sky130_fd_sc_hd__fa_2_871/CIN sky130_fd_sc_hd__fa_2_872/SUM
+ sky130_fd_sc_hd__fa_2_872/A sky130_fd_sc_hd__fa_2_872/B sky130_fd_sc_hd__fa_2_872/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_883 sky130_fd_sc_hd__fa_2_882/CIN sky130_fd_sc_hd__nand2_1_43/B
+ sky130_fd_sc_hd__ha_2_154/A sky130_fd_sc_hd__fa_2_883/B sky130_fd_sc_hd__fa_2_883/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_894 sky130_fd_sc_hd__fa_2_893/CIN sky130_fd_sc_hd__fa_2_894/SUM
+ sky130_fd_sc_hd__fa_2_894/A sky130_fd_sc_hd__fa_2_894/B sky130_fd_sc_hd__fa_2_894/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_3 sky130_fd_sc_hd__inv_2_3/A sky130_fd_sc_hd__inv_2_3/Y VDD
+ VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__nor3_2_5 sky130_fd_sc_hd__nor3_2_6/B sky130_fd_sc_hd__nor3_2_5/Y
+ sky130_fd_sc_hd__nor3_2_5/A sky130_fd_sc_hd__nor3_2_6/A VDD VSS VSS VDD sky130_fd_sc_hd__nor3_2
Xsky130_fd_sc_hd__nor2_1_13 sky130_fd_sc_hd__nor2_1_13/B sky130_fd_sc_hd__nor2_1_13/Y
+ sky130_fd_sc_hd__xor2_1_21/X VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_24 sky130_fd_sc_hd__nor2_1_24/B sky130_fd_sc_hd__nor2_1_24/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_35 sky130_fd_sc_hd__or4_1_2/X sky130_fd_sc_hd__nor2_1_35/Y
+ sky130_fd_sc_hd__nor4_1_6/C VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_46 sky130_fd_sc_hd__nor2_1_46/B sky130_fd_sc_hd__nor2_1_46/Y
+ sky130_fd_sc_hd__nor2_1_51/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_150 VSS VDD sky130_fd_sc_hd__mux2_2_150/A1 sky130_fd_sc_hd__mux2_2_150/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_150/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_57 sky130_fd_sc_hd__nor2_1_57/B sky130_fd_sc_hd__nor2_1_57/Y
+ sky130_fd_sc_hd__nor2_1_57/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_161 VSS VDD sky130_fd_sc_hd__mux2_2_161/A1 sky130_fd_sc_hd__mux2_2_161/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_161/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_68 sky130_fd_sc_hd__nor2_1_68/B sky130_fd_sc_hd__nor2_1_68/Y
+ sky130_fd_sc_hd__o21a_1_6/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_172 VSS VDD sky130_fd_sc_hd__mux2_2_172/A1 sky130_fd_sc_hd__xor2_1_252/X
+ sky130_fd_sc_hd__nor2_8_1/A sky130_fd_sc_hd__mux2_2_172/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_79 sky130_fd_sc_hd__nor2_1_79/B sky130_fd_sc_hd__nor2_1_79/Y
+ sky130_fd_sc_hd__nor2_1_79/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_183 VSS VDD sky130_fd_sc_hd__mux2_2_183/A1 sky130_fd_sc_hd__mux2_2_183/A0
+ sky130_fd_sc_hd__nor2_8_1/A sky130_fd_sc_hd__mux2_2_183/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_194 VSS VDD sky130_fd_sc_hd__mux2_2_194/A1 sky130_fd_sc_hd__mux2_2_194/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_194/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_sram_2kbyte_1rw1r_32x512_8_9 sky130_fd_sc_hd__buf_4_56/X sky130_fd_sc_hd__buf_4_57/X
+ sky130_fd_sc_hd__buf_4_58/X sky130_fd_sc_hd__clkbuf_4_106/X sky130_fd_sc_hd__clkbuf_4_155/X
+ sky130_fd_sc_hd__buf_4_59/X sky130_fd_sc_hd__buf_4_60/X sky130_fd_sc_hd__buf_4_61/X
+ sky130_fd_sc_hd__buf_4_62/X sky130_fd_sc_hd__clkbuf_4_107/X sky130_fd_sc_hd__buf_4_63/X
+ sky130_fd_sc_hd__buf_4_64/X sky130_fd_sc_hd__buf_4_65/X sky130_fd_sc_hd__buf_4_66/X
+ sky130_fd_sc_hd__clkbuf_4_108/X sky130_fd_sc_hd__buf_4_67/X sky130_fd_sc_hd__buf_4_56/X
+ sky130_fd_sc_hd__buf_4_57/X sky130_fd_sc_hd__buf_4_58/X sky130_fd_sc_hd__clkbuf_4_106/X
+ sky130_fd_sc_hd__clkbuf_4_155/X sky130_fd_sc_hd__buf_4_59/X sky130_fd_sc_hd__buf_4_60/X
+ sky130_fd_sc_hd__buf_4_61/X sky130_fd_sc_hd__buf_4_62/X sky130_fd_sc_hd__clkbuf_4_107/X
+ sky130_fd_sc_hd__buf_4_63/X sky130_fd_sc_hd__buf_4_64/X sky130_fd_sc_hd__buf_4_65/X
+ sky130_fd_sc_hd__buf_4_66/X sky130_fd_sc_hd__clkbuf_4_108/X sky130_fd_sc_hd__buf_4_67/X
+ sky130_fd_sc_hd__buf_12_312/X sky130_fd_sc_hd__buf_12_285/X sky130_fd_sc_hd__buf_12_355/X
+ sky130_fd_sc_hd__buf_12_343/X sky130_fd_sc_hd__buf_12_334/X sky130_fd_sc_hd__buf_12_288/X
+ sky130_fd_sc_hd__buf_12_346/X sky130_fd_sc_hd__buf_12_333/X sky130_fd_sc_hd__buf_12_369/X
+ sky130_fd_sc_hd__buf_12_345/X sky130_fd_sc_hd__buf_12_336/X sky130_fd_sc_hd__buf_12_286/X
+ sky130_fd_sc_hd__buf_12_359/X sky130_fd_sc_hd__buf_12_273/X sky130_fd_sc_hd__buf_12_289/X
+ sky130_fd_sc_hd__buf_12_340/X sky130_fd_sc_hd__buf_12_341/X sky130_fd_sc_hd__buf_12_329/X
+ sky130_fd_sc_hd__buf_2_133/X sky130_fd_sc_hd__clkbuf_4_110/X sky130_fd_sc_hd__buf_2_133/X
+ sky130_fd_sc_hd__clkinv_4_12/Y sky130_fd_sc_hd__clkinv_4_14/Y sky130_fd_sc_hd__buf_12_328/X
+ sky130_fd_sc_hd__buf_12_301/X sky130_fd_sc_hd__buf_12_327/X sky130_fd_sc_hd__buf_12_342/X
+ sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[0] sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[1]
+ sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[2] sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[3]
+ sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[4] sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[5]
+ sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[6] sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[7]
+ sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[8] sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[9]
+ sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[10] sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[11]
+ sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[12] sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[13]
+ sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[14] sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[15]
+ sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[16] sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[17]
+ sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[18] sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[19]
+ sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[20] sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[21]
+ sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[22] sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[23]
+ sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[24] sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[25]
+ sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[26] sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[27]
+ sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[28] sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[29]
+ sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[30] sky130_sram_2kbyte_1rw1r_32x512_8_9/dout0[31]
+ sky130_fd_sc_hd__clkbuf_4_113/A sky130_fd_sc_hd__clkbuf_4_114/A sky130_fd_sc_hd__clkinv_1_130/A
+ sky130_fd_sc_hd__clkinv_1_131/A sky130_fd_sc_hd__clkinv_1_132/A sky130_fd_sc_hd__clkbuf_4_115/A
+ sky130_fd_sc_hd__clkbuf_4_116/A sky130_fd_sc_hd__clkbuf_4_117/A sky130_fd_sc_hd__clkinv_1_133/A
+ sky130_fd_sc_hd__clkbuf_4_118/A sky130_fd_sc_hd__clkinv_1_134/A sky130_fd_sc_hd__clkinv_1_135/A
+ sky130_fd_sc_hd__clkinv_1_136/A sky130_fd_sc_hd__clkbuf_4_119/A sky130_fd_sc_hd__clkbuf_4_120/A
+ sky130_fd_sc_hd__clkbuf_4_121/A sky130_fd_sc_hd__clkbuf_1_282/A sky130_fd_sc_hd__clkbuf_1_283/A
+ sky130_fd_sc_hd__clkbuf_1_284/A sky130_fd_sc_hd__clkbuf_1_285/A sky130_fd_sc_hd__clkbuf_1_286/A
+ sky130_fd_sc_hd__clkbuf_1_287/A sky130_fd_sc_hd__clkbuf_1_288/A sky130_fd_sc_hd__clkbuf_1_289/A
+ sky130_fd_sc_hd__clkbuf_1_290/A sky130_fd_sc_hd__clkbuf_1_291/A sky130_fd_sc_hd__clkbuf_1_292/A
+ sky130_fd_sc_hd__clkbuf_1_293/A sky130_fd_sc_hd__clkbuf_1_294/A sky130_fd_sc_hd__clkbuf_1_295/A
+ sky130_fd_sc_hd__clkbuf_1_296/A sky130_fd_sc_hd__clkbuf_1_297/A VDD VSS sky130_sram_2kbyte_1rw1r_32x512_8
Xsky130_fd_sc_hd__a21oi_1_407 sky130_fd_sc_hd__nor2b_2_4/Y sky130_fd_sc_hd__o21ai_1_427/Y
+ sky130_fd_sc_hd__a21oi_1_407/Y sky130_fd_sc_hd__o21ai_1_434/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_418 sky130_fd_sc_hd__nor3_1_40/A sky130_fd_sc_hd__o22ai_1_378/Y
+ sky130_fd_sc_hd__a21oi_1_418/Y sky130_fd_sc_hd__fa_2_1247/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_429 sky130_fd_sc_hd__o21a_1_63/B1 sky130_fd_sc_hd__o21a_1_62/A1
+ sky130_fd_sc_hd__a21oi_1_429/Y sky130_fd_sc_hd__nor2_1_277/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkinv_8_109 sky130_fd_sc_hd__clkinv_8_47/A sky130_fd_sc_hd__clkinv_8_68/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__maj3_1_110 sky130_fd_sc_hd__maj3_1_111/X sky130_fd_sc_hd__maj3_1_110/X
+ sky130_fd_sc_hd__maj3_1_110/B sky130_fd_sc_hd__maj3_1_110/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_121 sky130_fd_sc_hd__maj3_1_122/X sky130_fd_sc_hd__maj3_1_121/X
+ sky130_fd_sc_hd__maj3_1_121/B sky130_fd_sc_hd__maj3_1_121/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_132 sky130_fd_sc_hd__maj3_1_133/X sky130_fd_sc_hd__maj3_1_132/X
+ sky130_fd_sc_hd__maj3_1_132/B sky130_fd_sc_hd__maj3_1_132/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_401 sky130_fd_sc_hd__xnor2_1_95/B sky130_fd_sc_hd__fa_2_1207/A
+ sky130_fd_sc_hd__o21a_1_36/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_143 sky130_fd_sc_hd__maj3_1_144/X sky130_fd_sc_hd__maj3_1_143/X
+ sky130_fd_sc_hd__maj3_1_143/B sky130_fd_sc_hd__maj3_1_143/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_412 sky130_fd_sc_hd__nand2_1_412/Y sky130_fd_sc_hd__nor2_1_205/B
+ sky130_fd_sc_hd__o31ai_1_8/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_90 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_90/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_90/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_154 sky130_fd_sc_hd__maj3_1_155/X sky130_fd_sc_hd__maj3_1_154/X
+ sky130_fd_sc_hd__maj3_1_154/B sky130_fd_sc_hd__maj3_1_154/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_423 sky130_fd_sc_hd__nor2_1_211/B sky130_fd_sc_hd__nand2_1_423/B
+ sky130_fd_sc_hd__nor2_1_212/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_370 sky130_fd_sc_hd__o32ai_1_8/A3 sky130_fd_sc_hd__o22ai_1_373/B1
+ sky130_fd_sc_hd__o22ai_1_370/Y sky130_fd_sc_hd__nor2_1_263/A sky130_fd_sc_hd__o21a_1_55/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_434 sky130_fd_sc_hd__nand2_1_434/Y sky130_fd_sc_hd__xor2_1_208/A
+ sky130_fd_sc_hd__nor2_1_224/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_381 sky130_fd_sc_hd__nand2_1_514/Y sky130_fd_sc_hd__o21ai_1_439/Y
+ sky130_fd_sc_hd__o22ai_1_381/Y sky130_fd_sc_hd__nand2_1_523/B sky130_fd_sc_hd__nand2_1_513/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_445 sky130_fd_sc_hd__nor2_1_267/A sky130_fd_sc_hd__nand2_1_445/B
+ sky130_fd_sc_hd__o32ai_1_8/B2 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_392 sky130_fd_sc_hd__nand2_1_514/Y sky130_fd_sc_hd__nand2_1_513/Y
+ sky130_fd_sc_hd__o22ai_1_392/Y sky130_fd_sc_hd__o22ai_1_405/A1 sky130_fd_sc_hd__a21o_2_29/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_456 sky130_fd_sc_hd__o21a_1_52/B1 sky130_fd_sc_hd__fa_2_1252/A
+ sky130_fd_sc_hd__o21a_1_52/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_467 sky130_fd_sc_hd__nand2_1_467/Y sky130_fd_sc_hd__nand2_1_468/Y
+ sky130_fd_sc_hd__nand2_1_469/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_478 sky130_fd_sc_hd__nand2_1_478/Y sky130_fd_sc_hd__nand2_1_491/B
+ sky130_fd_sc_hd__o21ai_1_409/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_489 sky130_fd_sc_hd__nand2_1_489/Y sky130_fd_sc_hd__nand2_1_491/B
+ sky130_fd_sc_hd__o21ai_1_434/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_14 sky130_fd_sc_hd__ha_2_40/SUM sky130_fd_sc_hd__nor2b_1_14/Y
+ sky130_fd_sc_hd__or2_1_0/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_25 sky130_fd_sc_hd__xor2_1_6/X sky130_fd_sc_hd__nor2b_1_25/Y
+ sky130_fd_sc_hd__or2_0_2/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_36 sky130_fd_sc_hd__ha_2_67/SUM sky130_fd_sc_hd__nor2b_1_36/Y
+ sky130_fd_sc_hd__or2_0_2/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1003 sky130_fd_sc_hd__nor2_1_229/B sky130_fd_sc_hd__fa_2_1235/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1003/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_47 sky130_fd_sc_hd__ha_2_86/SUM sky130_fd_sc_hd__nor2b_1_47/Y
+ sky130_fd_sc_hd__or2_0_3/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1014 sky130_fd_sc_hd__nand2_1_445/B sky130_fd_sc_hd__nor2b_2_4/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1014/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_58 sky130_fd_sc_hd__nand2b_1_7/B sky130_fd_sc_hd__nor2b_1_58/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1025 sky130_fd_sc_hd__o21a_1_55/A2 sky130_fd_sc_hd__fa_2_1253/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1025/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_69 sky130_fd_sc_hd__nor2b_1_86/A sky130_fd_sc_hd__nor2b_1_69/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1036 sky130_fd_sc_hd__nor3_1_41/B sky130_fd_sc_hd__o32ai_1_11/A3
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1047 sky130_fd_sc_hd__o31ai_1_11/B1 sky130_fd_sc_hd__a221oi_1_5/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1047/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1058 sky130_fd_sc_hd__nor2_1_290/A sky130_fd_sc_hd__or3_1_5/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1058/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1069 sky130_fd_sc_hd__nand2_1_527/B sky130_fd_sc_hd__fa_2_16/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1069/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_230 VDD VSS sky130_fd_sc_hd__nor3_2_10/A sky130_fd_sc_hd__clkinv_8_102/Y
+ sky130_fd_sc_hd__a22o_1_27/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_241 VDD VSS sky130_fd_sc_hd__fa_2_868/A sky130_fd_sc_hd__dfxtp_1_277/CLK
+ sky130_fd_sc_hd__and2_0_168/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_252 VDD VSS sky130_fd_sc_hd__dfxtp_1_252/Q sky130_fd_sc_hd__dfxtp_1_262/CLK
+ sky130_fd_sc_hd__and2_0_216/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_263 VDD VSS sky130_fd_sc_hd__xnor2_1_10/A sky130_fd_sc_hd__dfxtp_1_266/CLK
+ sky130_fd_sc_hd__and2_0_227/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_274 VDD VSS sky130_fd_sc_hd__dfxtp_1_274/Q sky130_fd_sc_hd__dfxtp_1_463/CLK
+ sky130_fd_sc_hd__and2_0_210/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_285 VDD VSS sky130_fd_sc_hd__a22o_1_62/A1 sky130_fd_sc_hd__dfxtp_1_477/CLK
+ sky130_fd_sc_hd__nand2_1_139/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_296 VDD VSS sky130_fd_sc_hd__and2_0_256/A sky130_fd_sc_hd__clkinv_4_31/Y
+ sky130_fd_sc_hd__nand2_1_117/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o22ai_1_5 sky130_fd_sc_hd__ha_2_94/B sky130_fd_sc_hd__fa_2_92/B
+ sky130_fd_sc_hd__fa_2_70/B sky130_fd_sc_hd__ha_2_99/A sky130_fd_sc_hd__fa_2_45/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_102 sky130_fd_sc_hd__fa_2_104/CIN sky130_fd_sc_hd__fa_2_98/A
+ sky130_fd_sc_hd__fa_2_49/B sky130_fd_sc_hd__fa_2_102/B sky130_fd_sc_hd__fa_2_102/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_113 sky130_fd_sc_hd__maj3_1_6/B sky130_fd_sc_hd__maj3_1_7/A
+ sky130_fd_sc_hd__fa_2_113/A sky130_fd_sc_hd__fa_2_113/B sky130_fd_sc_hd__fa_2_114/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_124 sky130_fd_sc_hd__fa_2_125/A sky130_fd_sc_hd__fa_2_121/A
+ sky130_fd_sc_hd__fa_2_96/A sky130_fd_sc_hd__fa_2_91/B sky130_fd_sc_hd__fa_2_124/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_135 sky130_fd_sc_hd__fa_2_134/B sky130_fd_sc_hd__fa_2_135/SUM
+ sky130_fd_sc_hd__fa_2_86/A sky130_fd_sc_hd__fa_2_92/B sky130_fd_sc_hd__fa_2_49/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_146 sky130_fd_sc_hd__fa_2_145/CIN sky130_fd_sc_hd__fa_2_146/SUM
+ sky130_fd_sc_hd__fa_2_146/A sky130_fd_sc_hd__fa_2_146/B sky130_fd_sc_hd__fa_2_146/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_157 sky130_fd_sc_hd__fa_2_146/A sky130_fd_sc_hd__fa_2_149/A
+ sky130_fd_sc_hd__ha_2_97/A sky130_fd_sc_hd__fa_2_15/B sky130_fd_sc_hd__fa_2_238/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_168 sky130_fd_sc_hd__fa_2_164/CIN sky130_fd_sc_hd__nor2_1_256/A
+ sky130_fd_sc_hd__fa_2_168/A sky130_fd_sc_hd__fa_2_168/B sky130_fd_sc_hd__fa_2_168/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_179 sky130_fd_sc_hd__fa_2_180/A sky130_fd_sc_hd__fa_2_178/B
+ sky130_fd_sc_hd__fa_2_32/A sky130_fd_sc_hd__fa_2_273/A sky130_fd_sc_hd__fa_2_265/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o22ai_1_12 sky130_fd_sc_hd__fa_2_242/A sky130_fd_sc_hd__fa_2_283/A
+ sky130_fd_sc_hd__maj3_1_53/B sky130_fd_sc_hd__fa_2_32/A sky130_fd_sc_hd__fa_2_250/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_130 VDD VSS sky130_fd_sc_hd__buf_8_131/A sky130_fd_sc_hd__and2_1_6/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_23 sky130_fd_sc_hd__ha_2_114/B sky130_fd_sc_hd__fa_2_409/A
+ sky130_fd_sc_hd__o22ai_1_23/Y sky130_fd_sc_hd__ha_2_110/B sky130_fd_sc_hd__fa_2_413/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_141 VDD VSS sky130_fd_sc_hd__buf_6_51/A sky130_fd_sc_hd__buf_2_275/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_34 sky130_fd_sc_hd__ha_2_121/B sky130_fd_sc_hd__fa_2_567/A
+ sky130_fd_sc_hd__fa_2_490/B sky130_fd_sc_hd__ha_2_118/B sky130_fd_sc_hd__fa_2_564/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_152 VDD VSS sky130_fd_sc_hd__buf_4_101/A sky130_fd_sc_hd__buf_6_55/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_45 sky130_fd_sc_hd__fa_2_700/A sky130_fd_sc_hd__fa_2_689/B
+ sky130_fd_sc_hd__fa_2_649/A sky130_fd_sc_hd__ha_2_134/B sky130_fd_sc_hd__fa_2_692/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_163 VDD VSS sky130_fd_sc_hd__buf_2_163/X sky130_fd_sc_hd__nand3_2_8/Y
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_56 sky130_fd_sc_hd__fa_2_833/A sky130_fd_sc_hd__fa_2_834/B
+ sky130_fd_sc_hd__fa_2_703/B sky130_fd_sc_hd__fa_2_835/B sky130_fd_sc_hd__fa_2_832/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_174 VDD VSS sky130_fd_sc_hd__buf_2_174/X sky130_fd_sc_hd__buf_2_174/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_67 sky130_fd_sc_hd__o22ai_1_88/B1 sky130_fd_sc_hd__nand2_2_3/Y
+ sky130_fd_sc_hd__o22ai_1_67/Y sky130_fd_sc_hd__xnor2_1_45/Y sky130_fd_sc_hd__o22ai_1_81/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_185 VDD VSS sky130_fd_sc_hd__buf_2_185/X sky130_fd_sc_hd__buf_2_185/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_78 sky130_fd_sc_hd__o22ai_1_89/A1 sky130_fd_sc_hd__o22ai_1_88/B1
+ sky130_fd_sc_hd__o22ai_1_78/Y sky130_fd_sc_hd__xnor2_1_39/Y sky130_fd_sc_hd__o22ai_1_78/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_196 VDD VSS sky130_fd_sc_hd__buf_2_196/X sky130_fd_sc_hd__buf_2_196/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_89 sky130_fd_sc_hd__o21ai_1_81/Y sky130_fd_sc_hd__nand2_2_3/Y
+ sky130_fd_sc_hd__o22ai_1_89/Y sky130_fd_sc_hd__o22ai_1_89/A1 sky130_fd_sc_hd__o21ai_1_74/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__dfxtp_1_1170 VDD VSS sky130_fd_sc_hd__fa_2_854/B sky130_fd_sc_hd__dfxtp_1_1184/CLK
+ sky130_fd_sc_hd__o21a_1_51/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1181 VDD VSS sky130_fd_sc_hd__fa_2_934/A sky130_fd_sc_hd__dfxtp_1_1184/CLK
+ sky130_fd_sc_hd__a21oi_1_365/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1192 VDD VSS sky130_fd_sc_hd__or2_0_11/A sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__nor2b_1_120/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_4_14 VDD VSS sky130_fd_sc_hd__buf_4_14/X sky130_fd_sc_hd__buf_8_10/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_25 VDD VSS sky130_fd_sc_hd__buf_4_25/X sky130_fd_sc_hd__buf_8_1/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_36 VDD VSS sky130_fd_sc_hd__buf_4_36/X sky130_fd_sc_hd__buf_4_36/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_47 VDD VSS sky130_fd_sc_hd__buf_4_47/X sky130_fd_sc_hd__buf_4_47/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_58 VDD VSS sky130_fd_sc_hd__buf_4_58/X sky130_fd_sc_hd__buf_4_58/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_69 VDD VSS sky130_fd_sc_hd__buf_4_69/X sky130_fd_sc_hd__buf_4_69/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__clkbuf_1_30 VSS VDD sky130_fd_sc_hd__clkbuf_1_30/X sky130_fd_sc_hd__clkbuf_1_30/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_107 sky130_fd_sc_hd__buf_12_77/X sky130_fd_sc_hd__buf_12_107/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_118 sky130_fd_sc_hd__buf_12_95/X sky130_fd_sc_hd__buf_12_118/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_41 VSS VDD sky130_fd_sc_hd__clkbuf_1_41/X sky130_fd_sc_hd__clkbuf_1_41/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_129 sky130_fd_sc_hd__buf_12_129/A sky130_fd_sc_hd__buf_12_129/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_52 VSS VDD sky130_fd_sc_hd__clkbuf_1_52/X sky130_fd_sc_hd__clkbuf_1_52/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_63 VSS VDD sky130_fd_sc_hd__clkbuf_1_63/X sky130_fd_sc_hd__clkbuf_1_63/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_74 VSS VDD sky130_fd_sc_hd__nand4_1_13/A sky130_fd_sc_hd__a22oi_1_75/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_680 sky130_fd_sc_hd__fa_2_577/A sky130_fd_sc_hd__fa_2_578/B
+ sky130_fd_sc_hd__fa_2_680/A sky130_fd_sc_hd__fa_2_680/B sky130_fd_sc_hd__fa_2_685/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_85 VSS VDD sky130_fd_sc_hd__nand4_1_2/A sky130_fd_sc_hd__a22oi_1_38/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_691 sky130_fd_sc_hd__fa_2_574/A sky130_fd_sc_hd__fa_2_575/B
+ sky130_fd_sc_hd__fa_2_691/A sky130_fd_sc_hd__fa_2_691/B sky130_fd_sc_hd__fa_2_695/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_96 VSS VDD sky130_fd_sc_hd__buf_8_13/A sky130_fd_sc_hd__ha_2_11/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkinv_1_307 sky130_fd_sc_hd__fa_2_404/B sky130_fd_sc_hd__ha_2_113/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_307/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_318 sky130_fd_sc_hd__fa_2_417/A sky130_fd_sc_hd__fa_2_360/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_318/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_329 sky130_fd_sc_hd__fa_2_566/A sky130_fd_sc_hd__ha_2_124/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_329/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_204 sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__o21ai_1_230/Y
+ sky130_fd_sc_hd__a21oi_1_204/Y sky130_fd_sc_hd__o21a_1_9/A2 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_215 sky130_fd_sc_hd__a211o_1_9/A1 sky130_fd_sc_hd__o21ai_1_246/Y
+ sky130_fd_sc_hd__a21oi_1_215/Y sky130_fd_sc_hd__o21ai_1_254/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__or2_0_10 sky130_fd_sc_hd__or2_0_10/A sky130_fd_sc_hd__or2_0_10/X
+ sky130_fd_sc_hd__or2_0_10/B VSS VDD VSS VDD sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__a21oi_1_226 sky130_fd_sc_hd__fa_2_1088/A sky130_fd_sc_hd__o21ai_1_261/Y
+ sky130_fd_sc_hd__a21oi_1_226/Y sky130_fd_sc_hd__nor2_4_12/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_2_11 sky130_fd_sc_hd__nor2_4_5/Y sky130_fd_sc_hd__a22oi_2_11/A2
+ sky130_fd_sc_hd__a22oi_2_9/B1 sky130_fd_sc_hd__clkbuf_4_31/X sky130_fd_sc_hd__a22oi_2_11/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__a21oi_1_237 sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__a22o_1_75/X
+ sky130_fd_sc_hd__a21oi_1_237/Y sky130_fd_sc_hd__fa_2_1069/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_2_22 sky130_fd_sc_hd__a22oi_2_25/A1 sky130_fd_sc_hd__a22oi_2_22/A2
+ sky130_fd_sc_hd__a22oi_2_25/B1 sky130_fd_sc_hd__a22oi_2_22/B2 sky130_fd_sc_hd__nand4_1_56/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__a21oi_1_248 sky130_fd_sc_hd__nor2_1_149/A sky130_fd_sc_hd__nor2_1_149/Y
+ sky130_fd_sc_hd__dfxtp_1_895/D sky130_fd_sc_hd__nor2_1_149/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_259 sky130_fd_sc_hd__or3_1_2/C sky130_fd_sc_hd__o21ai_1_284/Y
+ sky130_fd_sc_hd__a21oi_1_259/Y sky130_fd_sc_hd__nor2_1_163/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nand2_1_220 sky130_fd_sc_hd__o21ai_1_36/B1 sky130_fd_sc_hd__o22ai_1_58/A2
+ sky130_fd_sc_hd__fa_2_947/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_231 sky130_fd_sc_hd__xnor2_1_40/B sky130_fd_sc_hd__o21ai_1_79/B1
+ sky130_fd_sc_hd__o21ai_1_86/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_830 sky130_fd_sc_hd__o22ai_1_251/A1 sky130_fd_sc_hd__fa_2_1130/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_830/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_242 sky130_fd_sc_hd__o21ai_1_86/B1 sky130_fd_sc_hd__nor2_1_57/B
+ sky130_fd_sc_hd__nor2_1_57/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_841 sky130_fd_sc_hd__o22ai_1_258/B1 sky130_fd_sc_hd__fa_2_1150/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_841/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_253 sky130_fd_sc_hd__o21a_1_3/B1 sky130_fd_sc_hd__fa_2_986/A
+ sky130_fd_sc_hd__o21a_1_3/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_852 sky130_fd_sc_hd__nor2_1_154/B sky130_fd_sc_hd__fa_2_1147/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_852/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_264 sky130_fd_sc_hd__nand2_1_264/Y sky130_fd_sc_hd__xor2_1_60/A
+ sky130_fd_sc_hd__nand2_1_264/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_863 sky130_fd_sc_hd__nand2_1_439/B sky130_fd_sc_hd__nor2_1_224/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_863/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_275 sky130_fd_sc_hd__nand2_1_275/Y sky130_fd_sc_hd__a211o_1_8/A2
+ sky130_fd_sc_hd__nand2_1_275/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_874 sky130_fd_sc_hd__o32ai_1_4/A2 sky130_fd_sc_hd__fa_2_1191/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_874/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_286 sky130_fd_sc_hd__a22o_1_73/B2 sky130_fd_sc_hd__xnor2_1_63/B
+ sky130_fd_sc_hd__xnor2_1_62/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_885 sky130_fd_sc_hd__o22ai_1_291/A1 sky130_fd_sc_hd__nor2_1_213/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_885/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_297 sky130_fd_sc_hd__nand2_1_297/Y sky130_fd_sc_hd__nor2_1_109/B
+ sky130_fd_sc_hd__fa_2_1114/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_896 sky130_fd_sc_hd__nand2_1_420/B sky130_fd_sc_hd__fa_2_288/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_896/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand4_1_70 sky130_fd_sc_hd__nand4_1_70/C sky130_fd_sc_hd__nand4_1_70/B
+ sky130_fd_sc_hd__nand2_1_9/B sky130_fd_sc_hd__nand4_1_70/D sky130_fd_sc_hd__nand4_1_70/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_81 sky130_fd_sc_hd__or2_0_11/A sky130_fd_sc_hd__or2_0_8/A
+ sky130_fd_sc_hd__nand4_1_81/Y sky130_fd_sc_hd__or2_0_6/A sky130_fd_sc_hd__or2_0_9/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__mux2_2_3 VSS VDD sky130_fd_sc_hd__mux2_2_3/A1 sky130_fd_sc_hd__mux2_2_3/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_3/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__a21boi_0_3 sky130_fd_sc_hd__a21oi_1_233/Y sky130_fd_sc_hd__a21boi_0_3/Y
+ sky130_fd_sc_hd__fa_2_1072/A sky130_fd_sc_hd__a21o_2_5/A2 VSS VDD VDD VSS sky130_fd_sc_hd__a21boi_0
Xsky130_fd_sc_hd__fa_2_1170 sky130_fd_sc_hd__fa_2_1171/CIN sky130_fd_sc_hd__mux2_2_97/A1
+ sky130_fd_sc_hd__fa_2_1170/A sky130_fd_sc_hd__fa_2_1172/B sky130_fd_sc_hd__fa_2_1170/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1181 sky130_fd_sc_hd__fa_2_1182/CIN sky130_fd_sc_hd__mux2_2_147/A1
+ sky130_fd_sc_hd__fa_2_1181/A sky130_fd_sc_hd__fa_2_1181/B sky130_fd_sc_hd__fa_2_1181/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1192 sky130_fd_sc_hd__fa_2_1193/CIN sky130_fd_sc_hd__and2_0_326/A
+ sky130_fd_sc_hd__fa_2_1192/A sky130_fd_sc_hd__fa_2_1192/B sky130_fd_sc_hd__fa_2_1192/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a211o_1_17 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_182/A sky130_fd_sc_hd__nor2b_1_105/Y
+ sky130_fd_sc_hd__o22ai_1_240/Y sky130_fd_sc_hd__o21ai_1_294/Y sky130_fd_sc_hd__o22ai_1_239/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__a211o_1_28 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_292/A sky130_fd_sc_hd__o21ai_1_478/Y
+ sky130_fd_sc_hd__nor2_1_291/Y sky130_fd_sc_hd__nor2b_2_5/Y sky130_fd_sc_hd__o22ai_1_409/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__clkinv_1_104 sky130_fd_sc_hd__buf_8_70/A sky130_fd_sc_hd__inv_2_68/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_104/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_115 sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__buf_8_79/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_115/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_126 sky130_fd_sc_hd__nand3_2_4/B sky130_fd_sc_hd__and2_0_37/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_126/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_137 sky130_fd_sc_hd__clkinv_1_138/A sky130_fd_sc_hd__inv_2_74/Y
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_148 sky130_fd_sc_hd__buf_8_142/A sky130_fd_sc_hd__clkinv_1_148/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_148/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_159 sky130_fd_sc_hd__inv_2_90/A sky130_fd_sc_hd__buf_2_134/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_159/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_17 sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__ha_2_69/B
+ sky130_fd_sc_hd__a22o_1_17/X sky130_fd_sc_hd__dfxtp_1_1/Q sky130_fd_sc_hd__a22o_2_3/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_28 sky130_fd_sc_hd__or2_1_1/B sky130_fd_sc_hd__ha_2_80/A
+ sky130_fd_sc_hd__a22o_1_28/X sky130_fd_sc_hd__a22o_1_28/B2 sky130_fd_sc_hd__a22o_4_0/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_39 sky130_fd_sc_hd__a22o_1_39/A1 sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a22o_1_39/X sky130_fd_sc_hd__a21o_2_2/A2 sky130_fd_sc_hd__fa_2_945/SUM
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__o21ai_1_4 VSS VDD sky130_fd_sc_hd__o21ai_1_4/A2 sky130_fd_sc_hd__or4_1_0/A
+ sky130_fd_sc_hd__a21oi_1_2/Y sky130_fd_sc_hd__o21ai_1_4/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__bufbuf_16_3 sky130_fd_sc_hd__bufbuf_16_3/A sky130_fd_sc_hd__buf_12_259/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__nor2_1_220 sky130_fd_sc_hd__nor3_1_39/A sky130_fd_sc_hd__nor2_1_220/Y
+ sky130_fd_sc_hd__nor2_1_220/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_231 sky130_fd_sc_hd__nor2_1_231/B sky130_fd_sc_hd__o21a_1_47/A1
+ sky130_fd_sc_hd__nor2_1_231/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_242 sky130_fd_sc_hd__nor2_1_242/B sky130_fd_sc_hd__nor2_1_242/Y
+ sky130_fd_sc_hd__nor2_1_242/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_253 sky130_fd_sc_hd__nor2_1_253/B sky130_fd_sc_hd__nor2_1_253/Y
+ sky130_fd_sc_hd__nor2_1_253/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_2_7 sky130_fd_sc_hd__clkinv_2_7/Y sky130_fd_sc_hd__clkinv_2_7/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_7/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__nor2_1_264 sky130_fd_sc_hd__nor2_1_264/B sky130_fd_sc_hd__nor2_1_264/Y
+ sky130_fd_sc_hd__nor2_1_267/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_275 sky130_fd_sc_hd__nor2_1_275/B sky130_fd_sc_hd__o21a_1_61/A1
+ sky130_fd_sc_hd__nor2_1_275/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_286 sky130_fd_sc_hd__nor2_1_290/A sky130_fd_sc_hd__nor2_1_286/Y
+ sky130_fd_sc_hd__nor2_1_286/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_297 sky130_fd_sc_hd__nor2_1_297/B sky130_fd_sc_hd__nor2_1_297/Y
+ sky130_fd_sc_hd__fa_2_19/SUM VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_460 sky130_fd_sc_hd__buf_6_67/X sky130_fd_sc_hd__buf_12_460/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_471 sky130_fd_sc_hd__buf_6_82/X sky130_fd_sc_hd__buf_12_477/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_330 sky130_fd_sc_hd__fa_2_986/A sky130_fd_sc_hd__fa_2_988/A
+ sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__a22oi_1_330/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_482 sky130_fd_sc_hd__buf_12_482/A sky130_fd_sc_hd__buf_12_482/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_341 sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_2_7/Y
+ sky130_fd_sc_hd__fa_2_1006/A sky130_fd_sc_hd__fa_2_1007/A sky130_fd_sc_hd__a22oi_1_341/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_493 sky130_fd_sc_hd__buf_12_493/A sky130_fd_sc_hd__buf_12_493/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_352 sky130_fd_sc_hd__fa_2_1065/A sky130_fd_sc_hd__fa_2_1063/A
+ sky130_fd_sc_hd__nor2_2_12/Y sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__nand3_1_50/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_363 sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__nor2_2_12/Y
+ sky130_fd_sc_hd__fa_2_1080/A sky130_fd_sc_hd__fa_2_1083/A sky130_fd_sc_hd__a22oi_1_363/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_374 sky130_fd_sc_hd__nor3_1_38/B sky130_fd_sc_hd__fa_2_1139/A
+ sky130_fd_sc_hd__xor2_1_164/A sky130_fd_sc_hd__clkinv_1_779/Y sky130_fd_sc_hd__a22oi_1_374/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_385 sky130_fd_sc_hd__nor2_1_222/Y sky130_fd_sc_hd__nor2_1_224/Y
+ sky130_fd_sc_hd__fa_2_1200/A sky130_fd_sc_hd__fa_2_1196/A sky130_fd_sc_hd__a22oi_1_385/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_396 sky130_fd_sc_hd__a22oi_1_400/B1 sky130_fd_sc_hd__nor3_1_41/B
+ sky130_fd_sc_hd__fa_2_1281/A sky130_fd_sc_hd__fa_2_1282/A sky130_fd_sc_hd__a22oi_1_396/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nand2_1_18 sky130_fd_sc_hd__nor3_2_1/B sky130_fd_sc_hd__nor3_1_1/B
+ sky130_fd_sc_hd__nor3_1_3/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_660 sky130_fd_sc_hd__nor2_1_92/B sky130_fd_sc_hd__nand2_1_301/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_660/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_671 sky130_fd_sc_hd__clkinv_1_671/Y sky130_fd_sc_hd__nor2_1_97/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_671/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_29 sky130_fd_sc_hd__buf_2_244/A sky130_fd_sc_hd__nor2_1_6/Y
+ sky130_fd_sc_hd__or2_1_2/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_682 sky130_fd_sc_hd__nor2_1_109/B sky130_fd_sc_hd__fa_2_1114/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_682/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_693 sky130_fd_sc_hd__o21ai_1_210/A2 sky130_fd_sc_hd__fa_2_1078/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_693/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand3_1_0 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__nand3_1_0/A
+ sky130_fd_sc_hd__nand3_1_0/C sky130_fd_sc_hd__nand3_1_0/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__sdlclkp_2_12 sky130_fd_sc_hd__conb_1_29/LO sky130_fd_sc_hd__clkinv_4_33/Y
+ sky130_fd_sc_hd__dfxtp_1_1458/CLK sky130_fd_sc_hd__nand2b_1_18/Y VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__xnor2_1_60 VSS VDD sky130_fd_sc_hd__xnor2_1_60/B sky130_fd_sc_hd__xnor2_1_60/Y
+ sky130_fd_sc_hd__xnor2_1_60/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_71 VSS VDD sky130_fd_sc_hd__xnor2_1_71/B sky130_fd_sc_hd__xnor2_1_71/Y
+ sky130_fd_sc_hd__nor2_1_94/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_82 VSS VDD sky130_fd_sc_hd__xnor2_1_82/B sky130_fd_sc_hd__xnor2_1_82/Y
+ sky130_fd_sc_hd__nor2_1_97/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_93 VSS VDD sky130_fd_sc_hd__xor2_1_185/A sky130_fd_sc_hd__xnor2_1_93/Y
+ sky130_fd_sc_hd__xnor2_1_96/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__dfxtp_1_807 VDD VSS sky130_fd_sc_hd__fa_2_1059/A sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__mux2_2_59/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_818 VDD VSS sky130_fd_sc_hd__fa_2_1092/B sky130_fd_sc_hd__clkinv_8_59/Y
+ sky130_fd_sc_hd__and2_0_294/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_829 VDD VSS sky130_fd_sc_hd__fa_2_1103/A sky130_fd_sc_hd__clkinv_8_54/Y
+ sky130_fd_sc_hd__and2_0_316/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_405 VSS VDD sky130_fd_sc_hd__clkbuf_1_405/X sky130_fd_sc_hd__clkbuf_1_405/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_416 VSS VDD sky130_fd_sc_hd__clkbuf_1_416/X sky130_fd_sc_hd__clkbuf_1_416/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_427 VSS VDD sky130_fd_sc_hd__clkbuf_1_427/X sky130_fd_sc_hd__clkbuf_1_427/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_438 VSS VDD sky130_fd_sc_hd__clkbuf_1_438/X sky130_fd_sc_hd__clkbuf_1_438/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_449 VSS VDD sky130_fd_sc_hd__clkbuf_1_449/X sky130_fd_sc_hd__clkbuf_1_449/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__nor2b_1_109 sky130_fd_sc_hd__o32ai_1_2/Y sky130_fd_sc_hd__nor2b_1_109/Y
+ sky130_fd_sc_hd__buf_2_262/X VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__diode_2_190 sky130_fd_sc_hd__buf_2_153/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkinv_2_12 sky130_fd_sc_hd__clkinv_2_12/Y sky130_fd_sc_hd__clkinv_2_12/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_12/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkbuf_4_210 sky130_fd_sc_hd__clkbuf_4_210/X sky130_fd_sc_hd__clkbuf_4_210/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_2_23 sky130_fd_sc_hd__clkinv_2_23/Y sky130_fd_sc_hd__clkinv_2_23/A
+ VSS VDD VDD VSS VSS sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_34 sky130_fd_sc_hd__clkinv_2_35/A sky130_fd_sc_hd__clkinv_4_60/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_34/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkbuf_4_221 sky130_fd_sc_hd__a22o_1_7/A1 sig_amplitude[5] VSS VDD
+ VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_2_45 sky130_fd_sc_hd__clkinv_4_54/A sky130_fd_sc_hd__clkinv_4_53/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_45/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__sdlclkp_4_8 sky130_fd_sc_hd__conb_1_4/LO sky130_fd_sc_hd__clkinv_8_112/A
+ sky130_fd_sc_hd__dfxtp_1_9/CLK sky130_fd_sc_hd__buf_6_86/X VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__buf_12_290 sky130_fd_sc_hd__buf_12_290/A sky130_fd_sc_hd__buf_12_290/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_160 sky130_fd_sc_hd__clkbuf_1_351/X sky130_fd_sc_hd__clkbuf_1_353/X
+ sky130_fd_sc_hd__clkinv_2_14/Y sky130_fd_sc_hd__a22oi_1_160/A2 sky130_fd_sc_hd__nand4_1_35/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_171 sky130_fd_sc_hd__clkbuf_1_265/X sky130_fd_sc_hd__clkbuf_1_266/X
+ sky130_fd_sc_hd__clkbuf_1_276/X sky130_fd_sc_hd__a22oi_1_171/A2 sky130_fd_sc_hd__a22oi_1_171/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_182 sky130_fd_sc_hd__clkbuf_1_264/X sky130_fd_sc_hd__nor2_2_3/Y
+ sky130_fd_sc_hd__a22oi_1_182/B2 sky130_fd_sc_hd__clkbuf_4_129/X sky130_fd_sc_hd__nand4_1_40/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_193 sky130_fd_sc_hd__clkbuf_4_111/X sky130_fd_sc_hd__clkbuf_4_112/X
+ sky130_fd_sc_hd__a22oi_1_193/B2 sky130_fd_sc_hd__clkbuf_1_286/X sky130_fd_sc_hd__a22oi_1_193/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_490 sky130_fd_sc_hd__o21ai_1_76/B1 sky130_fd_sc_hd__nor2_1_60/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_490/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_404 VSS VDD sky130_fd_sc_hd__nor2_1_259/B sky130_fd_sc_hd__nor2_1_257/A
+ sky130_fd_sc_hd__a21oi_1_390/Y sky130_fd_sc_hd__o21ai_1_404/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_415 VSS VDD sky130_fd_sc_hd__o22ai_1_375/A2 sky130_fd_sc_hd__nor2_1_232/B
+ sky130_fd_sc_hd__a21oi_1_399/Y sky130_fd_sc_hd__o21ai_1_415/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_426 VSS VDD sky130_fd_sc_hd__a21oi_1_416/Y sky130_fd_sc_hd__nor2_1_267/A
+ sky130_fd_sc_hd__a21oi_1_407/Y sky130_fd_sc_hd__xor2_1_245/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_437 VSS VDD sky130_fd_sc_hd__o22ai_1_375/A2 sky130_fd_sc_hd__nor2_1_240/B
+ sky130_fd_sc_hd__a21oi_1_418/Y sky130_fd_sc_hd__o21ai_1_437/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_448 VSS VDD sky130_fd_sc_hd__nor2_1_275/B sky130_fd_sc_hd__o22ai_1_436/A2
+ sky130_fd_sc_hd__a22oi_1_396/Y sky130_fd_sc_hd__o21ai_1_448/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_459 VSS VDD sky130_fd_sc_hd__o21ai_1_468/A1 sky130_fd_sc_hd__nor2_1_307/A
+ sky130_fd_sc_hd__a21oi_1_451/Y sky130_fd_sc_hd__xor2_1_312/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_4_13 sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__nor2_4_13/A
+ sky130_fd_sc_hd__nor2_4_13/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__xor2_1_220 sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__fa_2_1198/B
+ sky130_fd_sc_hd__xor2_1_220/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_231 sky130_fd_sc_hd__xor2_1_231/B sky130_fd_sc_hd__xor2_1_231/X
+ sky130_fd_sc_hd__xor2_1_232/X VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__o21ai_1_19 VSS VDD sky130_fd_sc_hd__a21oi_2_0/Y sky130_fd_sc_hd__maj3_1_1/B
+ sky130_fd_sc_hd__nand2_1_38/Y sky130_fd_sc_hd__o21ai_1_19/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_242 sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1233/B
+ sky130_fd_sc_hd__xor2_1_242/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_253 sky130_fd_sc_hd__xor2_1_254/X sky130_fd_sc_hd__xor2_1_253/X
+ sky130_fd_sc_hd__xor2_1_253/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_604 VDD VSS sky130_fd_sc_hd__and2_0_214/A sky130_fd_sc_hd__dfxtp_1_606/CLK
+ sky130_fd_sc_hd__fa_2_1024/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_264 sky130_fd_sc_hd__xor2_1_267/B sky130_fd_sc_hd__fa_2_1250/B
+ sky130_fd_sc_hd__xor2_1_264/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_615 VDD VSS sky130_fd_sc_hd__fa_2_806/A sky130_fd_sc_hd__dfxtp_1_626/CLK
+ sky130_fd_sc_hd__o21a_1_6/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_275 sky130_fd_sc_hd__xor2_1_275/B sky130_fd_sc_hd__xor2_1_275/X
+ sky130_fd_sc_hd__xor2_1_275/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_626 VDD VSS sky130_fd_sc_hd__fa_2_835/B sky130_fd_sc_hd__dfxtp_1_626/CLK
+ sky130_fd_sc_hd__o21a_1_1/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_286 sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1285/B
+ sky130_fd_sc_hd__xor2_1_286/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_637 VDD VSS sky130_fd_sc_hd__fa_2_1001/A sky130_fd_sc_hd__clkinv_8_44/Y
+ sky130_fd_sc_hd__mux2_2_32/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_297 sky130_fd_sc_hd__xor2_1_297/B sky130_fd_sc_hd__xor2_1_297/X
+ sky130_fd_sc_hd__xor2_1_298/X VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_648 VDD VSS sky130_fd_sc_hd__fa_2_1012/A sky130_fd_sc_hd__clkinv_8_44/Y
+ sky130_fd_sc_hd__mux2_2_8/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_659 VDD VSS sky130_fd_sc_hd__fa_2_976/A sky130_fd_sc_hd__clkinv_8_41/Y
+ sky130_fd_sc_hd__mux2_2_37/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_202 VSS VDD sky130_fd_sc_hd__nand4_1_21/B sky130_fd_sc_hd__a22oi_1_106/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_213 VSS VDD sky130_fd_sc_hd__buf_12_130/A sky130_fd_sc_hd__buf_8_80/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_224 VSS VDD sky130_fd_sc_hd__buf_12_144/A sky130_fd_sc_hd__clkbuf_1_236/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_235 VSS VDD sky130_fd_sc_hd__clkbuf_1_235/X sky130_fd_sc_hd__buf_8_84/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_246 VSS VDD sky130_fd_sc_hd__buf_8_97/A sky130_fd_sc_hd__clkbuf_1_246/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_257 VSS VDD sky130_fd_sc_hd__clkbuf_1_257/X sky130_fd_sc_hd__clkbuf_1_259/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_268 VSS VDD sky130_fd_sc_hd__clkbuf_1_268/X sky130_fd_sc_hd__clkbuf_1_268/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_279 VSS VDD sky130_fd_sc_hd__clkbuf_1_279/X sky130_fd_sc_hd__clkbuf_1_279/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_509 sky130_fd_sc_hd__fa_2_513/B sky130_fd_sc_hd__fa_2_509/SUM
+ sky130_fd_sc_hd__fa_2_509/A sky130_fd_sc_hd__fa_2_509/B sky130_fd_sc_hd__fa_2_509/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_80 VDD VSS sky130_fd_sc_hd__buf_2_80/X sky130_fd_sc_hd__buf_2_80/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_91 VDD VSS sky130_fd_sc_hd__buf_2_91/X sky130_fd_sc_hd__buf_2_91/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_4_7 VDD VSS sky130_fd_sc_hd__buf_4_7/X sky130_fd_sc_hd__buf_4_7/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__and2_0_200 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_200/X sky130_fd_sc_hd__and2_0_235/B
+ sky130_fd_sc_hd__and2_0_200/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_211 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_211/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_211/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_222 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_222/X sky130_fd_sc_hd__and2_0_235/B
+ sky130_fd_sc_hd__and2_0_222/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_233 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_233/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__ha_2_146/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_244 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_244/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__xnor2_1_31/Y sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_255 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_255/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__xor2_1_30/X sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_266 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_266/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__fa_2_969/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_277 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_277/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__fa_2_993/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_288 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_288/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__fa_2_974/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_299 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_299/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_299/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__sdlclkp_2_5 sky130_fd_sc_hd__conb_1_13/LO sky130_fd_sc_hd__clkinv_8_112/A
+ sky130_fd_sc_hd__dfxtp_1_197/CLK sky130_fd_sc_hd__or2_0_2/X VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__o21ai_1_201 VSS VDD sky130_fd_sc_hd__xnor2_1_80/A sky130_fd_sc_hd__nor2_1_110/Y
+ sky130_fd_sc_hd__nand2_1_296/Y sky130_fd_sc_hd__xnor2_1_82/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_212 VSS VDD sky130_fd_sc_hd__a222oi_1_2/Y sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__nand2_1_317/Y sky130_fd_sc_hd__xor2_1_116/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_30 sky130_fd_sc_hd__clkbuf_4_30/X sky130_fd_sc_hd__clkbuf_4_30/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_223 VSS VDD sky130_fd_sc_hd__nor2_1_129/Y sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__a21oi_1_196/Y sky130_fd_sc_hd__xor2_1_126/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_41 sky130_fd_sc_hd__a22oi_2_4/B2 sky130_fd_sc_hd__clkbuf_4_41/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_234 VSS VDD sky130_fd_sc_hd__nor2_1_119/B sky130_fd_sc_hd__o21a_1_16/A2
+ sky130_fd_sc_hd__a21oi_1_208/Y sky130_fd_sc_hd__o21ai_1_234/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_52 sky130_fd_sc_hd__nand4_1_5/D sky130_fd_sc_hd__a22oi_1_46/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_245 VSS VDD sky130_fd_sc_hd__nor2_1_123/B sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__a21oi_1_215/Y sky130_fd_sc_hd__xor2_1_97/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_63 sky130_fd_sc_hd__clkbuf_4_63/X sky130_fd_sc_hd__clkbuf_4_64/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_256 VSS VDD sky130_fd_sc_hd__nor2_1_138/A sky130_fd_sc_hd__o22ai_1_206/A1
+ sky130_fd_sc_hd__a22oi_1_359/Y sky130_fd_sc_hd__o21ai_1_256/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_74 sky130_fd_sc_hd__clkbuf_4_74/X sky130_fd_sc_hd__clkbuf_4_74/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_267 VSS VDD sky130_fd_sc_hd__o22ai_1_197/B2 sky130_fd_sc_hd__o22ai_1_206/A1
+ sky130_fd_sc_hd__a22oi_1_364/Y sky130_fd_sc_hd__o21ai_1_267/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_85 sky130_fd_sc_hd__clkbuf_4_85/X sky130_fd_sc_hd__clkbuf_4_85/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_278 VSS VDD sky130_fd_sc_hd__nand2_1_368/B sky130_fd_sc_hd__a21o_2_7/B1
+ sky130_fd_sc_hd__a21o_2_6/A2 sky130_fd_sc_hd__o21ai_1_278/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_96 sky130_fd_sc_hd__buf_6_22/A sky130_fd_sc_hd__buf_6_21/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_289 VSS VDD sky130_fd_sc_hd__a222oi_1_6/Y sky130_fd_sc_hd__nor2_1_182/A
+ sky130_fd_sc_hd__nand2_1_373/Y sky130_fd_sc_hd__xor2_1_166/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__buf_8_180 sky130_fd_sc_hd__inv_2_124/Y sky130_fd_sc_hd__buf_8_180/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_191 sky130_fd_sc_hd__a22o_2_7/X sky130_fd_sc_hd__buf_8_222/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_401 VDD VSS sky130_fd_sc_hd__fa_2_1037/A sky130_fd_sc_hd__dfxtp_1_424/CLK
+ sky130_fd_sc_hd__and2_0_144/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_412 VDD VSS sky130_fd_sc_hd__fa_2_1032/B sky130_fd_sc_hd__dfxtp_1_419/CLK
+ sky130_fd_sc_hd__and2_0_193/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__inv_2_19 sky130_fd_sc_hd__inv_2_19/A sky130_fd_sc_hd__buf_8_4/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfxtp_1_423 VDD VSS sky130_fd_sc_hd__nor2_1_49/A sky130_fd_sc_hd__dfxtp_1_424/CLK
+ sky130_fd_sc_hd__and2_0_112/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_434 VDD VSS sky130_fd_sc_hd__dfxtp_1_434/Q sky130_fd_sc_hd__dfxtp_1_452/CLK
+ sky130_fd_sc_hd__nand2_1_96/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_445 VDD VSS sky130_fd_sc_hd__dfxtp_1_991/D sky130_fd_sc_hd__dfxtp_1_448/CLK
+ sky130_fd_sc_hd__nand2_1_74/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_456 VDD VSS sky130_fd_sc_hd__xor2_1_185/A sky130_fd_sc_hd__dfxtp_1_457/CLK
+ sky130_fd_sc_hd__nand2_1_52/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_467 VDD VSS sky130_fd_sc_hd__clkbuf_1_7/A sky130_fd_sc_hd__dfxtp_1_473/CLK
+ sky130_fd_sc_hd__and2_0_136/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_478 VDD VSS sky130_fd_sc_hd__xor2_1_30/B sky130_fd_sc_hd__dfxtp_1_483/CLK
+ sky130_fd_sc_hd__nor2b_1_67/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_489 VDD VSS sky130_fd_sc_hd__dfxtp_1_489/Q sky130_fd_sc_hd__dfxtp_1_496/CLK
+ sky130_fd_sc_hd__nor2b_1_76/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2b_1_15 sky130_fd_sc_hd__xnor2_1_62/B sky130_fd_sc_hd__ha_2_201/A
+ sky130_fd_sc_hd__ha_2_201/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__fa_2_306 sky130_fd_sc_hd__fa_2_303/CIN sky130_fd_sc_hd__fa_2_306/SUM
+ sky130_fd_sc_hd__fa_2_306/A sky130_fd_sc_hd__fa_2_306/B sky130_fd_sc_hd__fa_2_306/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_317 sky130_fd_sc_hd__fa_2_310/A sky130_fd_sc_hd__fa_2_314/B
+ sky130_fd_sc_hd__fa_2_317/A sky130_fd_sc_hd__fa_2_317/B sky130_fd_sc_hd__fa_2_317/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_328 sky130_fd_sc_hd__fa_2_329/A sky130_fd_sc_hd__fa_2_328/SUM
+ sky130_fd_sc_hd__ha_2_114/B sky130_fd_sc_hd__ha_2_113/B sky130_fd_sc_hd__fa_2_417/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_339 sky130_fd_sc_hd__fa_2_341/B sky130_fd_sc_hd__fa_2_337/A
+ sky130_fd_sc_hd__fa_2_404/A sky130_fd_sc_hd__ha_2_116/B sky130_fd_sc_hd__fa_2_422/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_8_11 sky130_fd_sc_hd__clkinv_8_11/Y sky130_fd_sc_hd__clkinv_4_2/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_22 sky130_fd_sc_hd__clkinv_8_23/A sky130_fd_sc_hd__clkinv_8_22/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_22/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_33 sky130_fd_sc_hd__clkinv_8_33/Y sky130_fd_sc_hd__clkinv_8_33/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_33/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_44 sky130_fd_sc_hd__clkinv_8_44/Y sky130_fd_sc_hd__clkinv_8_44/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_44/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_55 sky130_fd_sc_hd__clkinv_8_55/Y sky130_fd_sc_hd__clkinv_8_56/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_55/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_66 sky130_fd_sc_hd__clkinv_8_66/Y sky130_fd_sc_hd__clkinv_8_67/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_66/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_20 sky130_fd_sc_hd__buf_12_20/A sky130_fd_sc_hd__buf_12_20/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_8_77 sky130_fd_sc_hd__clkinv_8_77/Y sky130_fd_sc_hd__clkinv_8_78/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_77/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_31 sky130_fd_sc_hd__buf_8_11/X sky130_fd_sc_hd__buf_12_31/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_8_88 sky130_fd_sc_hd__clkinv_8_89/A sky130_fd_sc_hd__clkinv_8_88/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_88/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_42 sky130_fd_sc_hd__buf_8_55/X sky130_fd_sc_hd__buf_12_42/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_8_99 sky130_fd_sc_hd__clkinv_8_99/Y sky130_fd_sc_hd__clkinv_8_99/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_99/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_53 sky130_fd_sc_hd__buf_8_42/X sky130_fd_sc_hd__buf_12_53/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_64 sky130_fd_sc_hd__buf_4_29/X sky130_fd_sc_hd__buf_12_64/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_75 sky130_fd_sc_hd__buf_4_28/X sky130_fd_sc_hd__buf_12_75/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_86 sky130_fd_sc_hd__buf_6_17/X sky130_fd_sc_hd__buf_12_86/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_97 sky130_fd_sc_hd__buf_12_97/A sky130_fd_sc_hd__buf_12_97/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_2_4 VDD VSS sky130_fd_sc_hd__buf_4_7/A sky130_fd_sc_hd__buf_4_6/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1330 VDD VSS sky130_fd_sc_hd__fa_2_914/A sky130_fd_sc_hd__dfxtp_1_1332/CLK
+ sky130_fd_sc_hd__a21oi_1_421/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1341 VDD VSS sky130_fd_sc_hd__fa_2_1300/A sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__mux2_2_245/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1352 VDD VSS sky130_fd_sc_hd__xor2_1_298/A sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__mux2_2_220/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1363 VDD VSS sky130_fd_sc_hd__fa_2_1285/A sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__mux2_2_238/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1374 VDD VSS sky130_fd_sc_hd__fa_2_1313/A sky130_fd_sc_hd__clkinv_8_102/Y
+ sky130_fd_sc_hd__mux2_2_265/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1385 VDD VSS sky130_fd_sc_hd__fa_2_1324/A sky130_fd_sc_hd__clkinv_8_75/Y
+ sky130_fd_sc_hd__nand2_1_517/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1396 VDD VSS sky130_fd_sc_hd__mux2_2_255/A0 sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__o22ai_1_393/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_990 VDD VSS sky130_fd_sc_hd__mux2_2_121/A0 sky130_fd_sc_hd__clkinv_8_64/Y
+ sky130_fd_sc_hd__dfxtp_1_990/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_840 sky130_fd_sc_hd__fa_2_839/CIN sky130_fd_sc_hd__fa_2_840/SUM
+ sky130_fd_sc_hd__fa_2_840/A sky130_fd_sc_hd__fa_2_840/B sky130_fd_sc_hd__fa_2_840/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_851 sky130_fd_sc_hd__fa_2_850/CIN sky130_fd_sc_hd__fa_2_851/SUM
+ sky130_fd_sc_hd__fa_2_851/A sky130_fd_sc_hd__fa_2_851/B sky130_fd_sc_hd__fa_2_851/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_862 sky130_fd_sc_hd__fa_2_861/CIN sky130_fd_sc_hd__fa_2_862/SUM
+ sky130_fd_sc_hd__fa_2_862/A sky130_fd_sc_hd__fa_2_862/B sky130_fd_sc_hd__fa_2_862/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_873 sky130_fd_sc_hd__fa_2_872/CIN sky130_fd_sc_hd__fa_2_873/SUM
+ sky130_fd_sc_hd__fa_2_873/A sky130_fd_sc_hd__fa_2_873/B sky130_fd_sc_hd__fa_2_873/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_884 sky130_fd_sc_hd__fa_2_883/CIN sky130_fd_sc_hd__nand2_1_44/B
+ sky130_fd_sc_hd__ha_2_155/A sky130_fd_sc_hd__fa_2_884/B sky130_fd_sc_hd__fa_2_884/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_895 sky130_fd_sc_hd__fa_2_894/CIN sky130_fd_sc_hd__fa_2_895/SUM
+ sky130_fd_sc_hd__fa_2_895/A sky130_fd_sc_hd__fa_2_895/B sky130_fd_sc_hd__fa_2_895/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_4 sky130_fd_sc_hd__inv_2_4/A sky130_fd_sc_hd__inv_2_4/Y VDD
+ VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__nor3_2_6 sky130_fd_sc_hd__nor3_2_6/C sky130_fd_sc_hd__nor3_2_6/Y
+ sky130_fd_sc_hd__nor3_2_6/A sky130_fd_sc_hd__nor3_2_6/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_2
Xsky130_fd_sc_hd__nor2_1_14 sky130_fd_sc_hd__or2_0_0/B sky130_fd_sc_hd__nor2_1_14/Y
+ sky130_fd_sc_hd__inv_4_1/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_25 sky130_fd_sc_hd__nor2_1_25/B sky130_fd_sc_hd__nor2_1_25/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_36 sky130_fd_sc_hd__nor2_1_36/B sky130_fd_sc_hd__nor3_1_34/C
+ sky130_fd_sc_hd__nor2_1_36/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_140 VSS VDD sky130_fd_sc_hd__xor2_1_228/X sky130_fd_sc_hd__nand2_1_416/B
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_140/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_47 sky130_fd_sc_hd__nor2_1_47/B sky130_fd_sc_hd__nor2_1_47/Y
+ sky130_fd_sc_hd__nor2_1_50/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_151 VSS VDD sky130_fd_sc_hd__mux2_2_151/A1 sky130_fd_sc_hd__mux2_2_151/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_151/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_58 sky130_fd_sc_hd__nor2_1_58/B sky130_fd_sc_hd__nor2_1_58/Y
+ sky130_fd_sc_hd__nor2_1_58/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_162 VSS VDD sky130_fd_sc_hd__mux2_2_162/A1 sky130_fd_sc_hd__mux2_2_162/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_162/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_69 sky130_fd_sc_hd__nor2_1_69/B sky130_fd_sc_hd__o21a_1_6/A1
+ sky130_fd_sc_hd__o21a_1_7/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_173 VSS VDD sky130_fd_sc_hd__mux2_2_173/A1 sky130_fd_sc_hd__xor2_1_231/X
+ sky130_fd_sc_hd__nor2_8_1/A sky130_fd_sc_hd__mux2_2_173/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_184 VSS VDD sky130_fd_sc_hd__mux2_2_184/A1 sky130_fd_sc_hd__mux2_2_184/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_184/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_195 VSS VDD sky130_fd_sc_hd__mux2_2_195/A1 sky130_fd_sc_hd__mux2_2_195/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_195/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__a21oi_1_408 sky130_fd_sc_hd__nor2_1_267/Y sky130_fd_sc_hd__nor2_1_262/Y
+ sky130_fd_sc_hd__a21oi_1_408/Y sky130_fd_sc_hd__fa_2_1250/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_419 sky130_fd_sc_hd__fa_2_1252/A sky130_fd_sc_hd__o22ai_1_379/Y
+ sky130_fd_sc_hd__o21a_1_55/B1 sky130_fd_sc_hd__nor2_2_17/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__maj3_1_100 sky130_fd_sc_hd__maj3_1_101/X sky130_fd_sc_hd__maj3_1_99/C
+ sky130_fd_sc_hd__maj3_1_100/B sky130_fd_sc_hd__maj3_1_100/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_111 sky130_fd_sc_hd__maj3_1_112/X sky130_fd_sc_hd__maj3_1_111/X
+ sky130_fd_sc_hd__maj3_1_111/B sky130_fd_sc_hd__maj3_1_111/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_122 sky130_fd_sc_hd__maj3_1_123/X sky130_fd_sc_hd__maj3_1_122/X
+ sky130_fd_sc_hd__maj3_1_122/B sky130_fd_sc_hd__maj3_1_122/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_402 sky130_fd_sc_hd__o21a_1_37/B1 sky130_fd_sc_hd__fa_2_1205/A
+ sky130_fd_sc_hd__o21a_1_37/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_133 sky130_fd_sc_hd__maj3_1_134/X sky130_fd_sc_hd__maj3_1_133/X
+ sky130_fd_sc_hd__maj3_1_133/B sky130_fd_sc_hd__maj3_1_133/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__and2_0_80 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_80/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__and2_0_80/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_413 sky130_fd_sc_hd__nand2_1_413/Y sky130_fd_sc_hd__nand2_1_416/Y
+ sky130_fd_sc_hd__nand2_1_414/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_144 sky130_fd_sc_hd__maj3_1_145/X sky130_fd_sc_hd__maj3_1_144/X
+ sky130_fd_sc_hd__maj3_1_144/B sky130_fd_sc_hd__maj3_1_144/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_360 sky130_fd_sc_hd__o22ai_1_379/A2 sky130_fd_sc_hd__o22ai_1_361/A1
+ sky130_fd_sc_hd__o22ai_1_360/Y sky130_fd_sc_hd__nor2_1_231/B sky130_fd_sc_hd__o32ai_1_8/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_91 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_91/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_91/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_424 sky130_fd_sc_hd__nor2_1_212/B sky130_fd_sc_hd__nand2_1_424/B
+ sky130_fd_sc_hd__nor2_1_213/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_155 sky130_fd_sc_hd__maj3_1_156/X sky130_fd_sc_hd__maj3_1_155/X
+ sky130_fd_sc_hd__maj3_1_155/B sky130_fd_sc_hd__maj3_1_155/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_371 sky130_fd_sc_hd__o22ai_1_379/A2 sky130_fd_sc_hd__o22ai_1_379/B1
+ sky130_fd_sc_hd__o22ai_1_371/Y sky130_fd_sc_hd__o21a_1_55/A2 sky130_fd_sc_hd__o22ai_1_375/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_435 sky130_fd_sc_hd__nand2_1_435/Y sky130_fd_sc_hd__nand2_1_439/B
+ sky130_fd_sc_hd__o21ai_1_382/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_382 sky130_fd_sc_hd__nand2_1_514/Y sky130_fd_sc_hd__nand2_1_513/Y
+ sky130_fd_sc_hd__o22ai_1_382/Y sky130_fd_sc_hd__o22ai_1_395/A1 sky130_fd_sc_hd__a21o_2_24/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_446 sky130_fd_sc_hd__xnor2_1_97/B sky130_fd_sc_hd__fa_2_1240/A
+ sky130_fd_sc_hd__o21a_1_43/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_393 sky130_fd_sc_hd__nand2_1_514/Y sky130_fd_sc_hd__nand2_1_513/Y
+ sky130_fd_sc_hd__o22ai_1_393/Y sky130_fd_sc_hd__o22ai_1_406/A1 sky130_fd_sc_hd__o21ai_1_445/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_457 sky130_fd_sc_hd__o21a_1_53/B1 sky130_fd_sc_hd__fa_2_1250/A
+ sky130_fd_sc_hd__o21a_1_53/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_468 sky130_fd_sc_hd__nand2_1_468/Y sky130_fd_sc_hd__nand2_1_468/B
+ sky130_fd_sc_hd__nor2_8_1/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_479 sky130_fd_sc_hd__nand2_1_479/Y sky130_fd_sc_hd__nand2_1_491/B
+ sky130_fd_sc_hd__o21ai_1_413/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_15 sky130_fd_sc_hd__xor2_1_4/X sky130_fd_sc_hd__nor2b_1_15/Y
+ sky130_fd_sc_hd__or2_1_0/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_26 sky130_fd_sc_hd__nor2b_1_26/B_N sky130_fd_sc_hd__nor2b_1_26/Y
+ sky130_fd_sc_hd__or2_0_2/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_37 sky130_fd_sc_hd__nor2_4_0/Y sky130_fd_sc_hd__and2_0_84/A
+ sky130_fd_sc_hd__ha_2_79/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1004 sky130_fd_sc_hd__a21oi_1_401/B1 sky130_fd_sc_hd__nand2_1_490/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1004/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_48 sky130_fd_sc_hd__ha_2_85/SUM sky130_fd_sc_hd__nor2b_1_48/Y
+ sky130_fd_sc_hd__or2_0_3/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1015 sky130_fd_sc_hd__o32ai_1_8/B2 sky130_fd_sc_hd__o32ai_1_8/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1015/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_59 sky130_fd_sc_hd__dfxtp_1_493/Q sky130_fd_sc_hd__nor2b_1_59/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1026 sky130_fd_sc_hd__nor2_1_243/B sky130_fd_sc_hd__o21bai_1_4/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1026/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1037 sky130_fd_sc_hd__nor2_1_299/A sky130_fd_sc_hd__nor2b_1_126/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1037/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1048 sky130_fd_sc_hd__o31ai_1_12/B1 sky130_fd_sc_hd__a21oi_1_442/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1048/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_90 sky130_fd_sc_hd__ha_2_33/A sky130_fd_sc_hd__buf_8_90/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__clkinv_1_1059 sky130_fd_sc_hd__o32ai_1_10/B2 sky130_fd_sc_hd__fa_2_1295/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1059/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_220 VDD VSS sky130_fd_sc_hd__ha_2_83/A sky130_fd_sc_hd__dfxtp_1_223/CLK
+ sky130_fd_sc_hd__nor2b_1_45/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_231 VDD VSS sky130_fd_sc_hd__xor2_1_14/A sky130_fd_sc_hd__dfxtp_1_472/CLK
+ sky130_fd_sc_hd__and2_0_163/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_242 VDD VSS sky130_fd_sc_hd__fa_2_867/A sky130_fd_sc_hd__dfxtp_1_277/CLK
+ sky130_fd_sc_hd__and2_0_172/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_253 VDD VSS sky130_fd_sc_hd__dfxtp_1_253/Q sky130_fd_sc_hd__dfxtp_1_258/CLK
+ sky130_fd_sc_hd__and2_0_217/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_264 VDD VSS sky130_fd_sc_hd__dfxtp_1_264/Q sky130_fd_sc_hd__dfxtp_1_313/CLK
+ sky130_fd_sc_hd__and2_0_224/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_275 VDD VSS sky130_fd_sc_hd__dfxtp_1_275/Q sky130_fd_sc_hd__dfxtp_1_462/CLK
+ sky130_fd_sc_hd__and2_0_209/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_286 VDD VSS sky130_fd_sc_hd__a22o_1_61/A1 sky130_fd_sc_hd__dfxtp_1_477/CLK
+ sky130_fd_sc_hd__nand2_1_137/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_297 VDD VSS sky130_fd_sc_hd__xor2_1_27/A sky130_fd_sc_hd__dfxtp_1_477/CLK
+ sky130_fd_sc_hd__nand2_1_115/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o22ai_1_6 sky130_fd_sc_hd__ha_2_91/B sky130_fd_sc_hd__fa_2_80/B
+ sky130_fd_sc_hd__fa_2_90/A sky130_fd_sc_hd__fa_2_5/A sky130_fd_sc_hd__fa_2_76/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_103 sky130_fd_sc_hd__maj3_1_8/B sky130_fd_sc_hd__maj3_1_9/A
+ sky130_fd_sc_hd__fa_2_103/A sky130_fd_sc_hd__fa_2_103/B sky130_fd_sc_hd__fa_2_104/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_114 sky130_fd_sc_hd__fa_2_117/B sky130_fd_sc_hd__fa_2_114/SUM
+ sky130_fd_sc_hd__fa_2_114/A sky130_fd_sc_hd__fa_2_114/B sky130_fd_sc_hd__o22ai_1_7/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_125 sky130_fd_sc_hd__fa_2_28/A sky130_fd_sc_hd__maj3_1_4/A
+ sky130_fd_sc_hd__fa_2_125/A sky130_fd_sc_hd__fa_2_125/B sky130_fd_sc_hd__fa_2_127/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_136 sky130_fd_sc_hd__fa_2_22/A sky130_fd_sc_hd__fa_2_26/B sky130_fd_sc_hd__fa_2_136/A
+ sky130_fd_sc_hd__fa_2_136/B sky130_fd_sc_hd__fa_2_141/SUM VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_147 sky130_fd_sc_hd__fa_2_145/B sky130_fd_sc_hd__fa_2_146/B
+ sky130_fd_sc_hd__fa_2_5/A sky130_fd_sc_hd__fa_2_5/B sky130_fd_sc_hd__fa_2_144/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_158 sky130_fd_sc_hd__fa_2_150/CIN sky130_fd_sc_hd__fa_2_158/SUM
+ sky130_fd_sc_hd__fa_2_158/A sky130_fd_sc_hd__fa_2_158/B sky130_fd_sc_hd__fa_2_158/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_169 sky130_fd_sc_hd__fa_2_168/CIN sky130_fd_sc_hd__or3_1_4/A
+ sky130_fd_sc_hd__fa_2_169/A sky130_fd_sc_hd__fa_2_169/B sky130_fd_sc_hd__fa_2_169/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_120 VDD VSS sky130_fd_sc_hd__buf_2_120/X sky130_fd_sc_hd__buf_2_120/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_13 sky130_fd_sc_hd__ha_2_104/B sky130_fd_sc_hd__fa_2_258/A
+ sky130_fd_sc_hd__o22ai_1_13/Y sky130_fd_sc_hd__ha_2_91/B sky130_fd_sc_hd__fa_2_281/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_131 VDD VSS sky130_fd_sc_hd__inv_2_85/A sky130_fd_sc_hd__and2_1_7/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_24 sky130_fd_sc_hd__ha_2_112/B sky130_fd_sc_hd__fa_2_425/A
+ sky130_fd_sc_hd__fa_2_348/B sky130_fd_sc_hd__ha_2_109/B sky130_fd_sc_hd__fa_2_422/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_142 VDD VSS sky130_fd_sc_hd__buf_2_142/X sky130_fd_sc_hd__buf_6_51/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_35 sky130_fd_sc_hd__ha_2_122/B sky130_fd_sc_hd__fa_2_564/B
+ sky130_fd_sc_hd__fa_2_505/B sky130_fd_sc_hd__ha_2_121/B sky130_fd_sc_hd__fa_2_546/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_153 VDD VSS sky130_fd_sc_hd__buf_4_102/A sky130_fd_sc_hd__buf_2_153/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_46 sky130_fd_sc_hd__fa_2_701/B sky130_fd_sc_hd__ha_2_130/A
+ sky130_fd_sc_hd__o22ai_1_46/Y sky130_fd_sc_hd__fa_2_673/B sky130_fd_sc_hd__fa_2_700/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_164 VDD VSS sky130_fd_sc_hd__buf_2_164/X sky130_fd_sc_hd__nor3_1_21/Y
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_57 sky130_fd_sc_hd__ha_2_157/B sky130_fd_sc_hd__ha_2_157/A
+ sky130_fd_sc_hd__o22ai_1_57/Y sky130_fd_sc_hd__nor4_1_4/C sky130_fd_sc_hd__o22ai_1_57/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_175 VDD VSS sky130_fd_sc_hd__buf_2_175/X sky130_fd_sc_hd__buf_2_175/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_68 sky130_fd_sc_hd__o22ai_1_88/B1 sky130_fd_sc_hd__nand2_2_3/Y
+ sky130_fd_sc_hd__o22ai_1_68/Y sky130_fd_sc_hd__xnor2_1_47/Y sky130_fd_sc_hd__o22ai_1_82/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_186 VDD VSS sky130_fd_sc_hd__buf_2_186/X sky130_fd_sc_hd__buf_2_186/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_79 sky130_fd_sc_hd__o22ai_1_89/A1 sky130_fd_sc_hd__o22ai_1_88/B1
+ sky130_fd_sc_hd__o22ai_1_79/Y sky130_fd_sc_hd__xnor2_1_41/Y sky130_fd_sc_hd__o22ai_1_79/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_197 VDD VSS sky130_fd_sc_hd__buf_2_197/X sky130_fd_sc_hd__buf_2_197/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1160 VDD VSS sky130_fd_sc_hd__ha_2_147/B sky130_fd_sc_hd__dfxtp_1_1179/CLK
+ sky130_fd_sc_hd__o32ai_1_7/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1171 VDD VSS sky130_fd_sc_hd__fa_2_853/B sky130_fd_sc_hd__dfxtp_1_1184/CLK
+ sky130_fd_sc_hd__a21oi_1_370/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1182 VDD VSS sky130_fd_sc_hd__fa_2_935/A sky130_fd_sc_hd__clkinv_4_24/Y
+ sky130_fd_sc_hd__o21a_1_47/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1193 VDD VSS sky130_fd_sc_hd__fa_2_1242/B sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__and2_0_330/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_4_15 VDD VSS sky130_fd_sc_hd__buf_4_15/X sky130_fd_sc_hd__buf_8_38/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_26 VDD VSS sky130_fd_sc_hd__buf_4_26/X sky130_fd_sc_hd__buf_8_22/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_37 VDD VSS sky130_fd_sc_hd__buf_4_37/X sky130_fd_sc_hd__buf_4_37/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_48 VDD VSS sky130_fd_sc_hd__buf_4_48/X sky130_fd_sc_hd__buf_8_99/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_59 VDD VSS sky130_fd_sc_hd__buf_4_59/X sky130_fd_sc_hd__buf_6_88/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__clkbuf_1_20 VSS VDD sky130_fd_sc_hd__clkbuf_1_20/X sky130_fd_sc_hd__clkbuf_1_20/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_108 sky130_fd_sc_hd__buf_12_76/X sky130_fd_sc_hd__buf_12_114/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_31 VSS VDD sky130_fd_sc_hd__clkbuf_1_31/X sky130_fd_sc_hd__clkbuf_1_31/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_119 sky130_fd_sc_hd__buf_12_119/A sky130_fd_sc_hd__buf_12_119/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_42 VSS VDD sky130_fd_sc_hd__clkbuf_1_42/X sky130_fd_sc_hd__clkbuf_1_42/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_53 VSS VDD sky130_fd_sc_hd__clkbuf_1_53/X sky130_fd_sc_hd__clkbuf_1_53/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_64 VSS VDD sky130_fd_sc_hd__clkbuf_1_64/X sky130_fd_sc_hd__clkbuf_1_64/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_670 sky130_fd_sc_hd__fa_2_579/A sky130_fd_sc_hd__fa_2_580/B
+ sky130_fd_sc_hd__fa_2_670/A sky130_fd_sc_hd__fa_2_670/B sky130_fd_sc_hd__fa_2_676/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_75 VSS VDD sky130_fd_sc_hd__nand4_1_12/A sky130_fd_sc_hd__a22oi_1_71/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_681 sky130_fd_sc_hd__fa_2_680/B sky130_fd_sc_hd__fa_2_681/SUM
+ sky130_fd_sc_hd__fa_2_681/A sky130_fd_sc_hd__fa_2_681/B sky130_fd_sc_hd__fa_2_681/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_86 VSS VDD sky130_fd_sc_hd__nand4_1_1/A sky130_fd_sc_hd__a22oi_1_34/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_692 sky130_fd_sc_hd__fa_2_691/B sky130_fd_sc_hd__fa_2_692/SUM
+ sky130_fd_sc_hd__fa_2_692/A sky130_fd_sc_hd__fa_2_700/B sky130_fd_sc_hd__fa_2_692/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_97 VSS VDD sky130_fd_sc_hd__buf_8_20/A sky130_fd_sc_hd__ha_2_13/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkinv_1_308 sky130_fd_sc_hd__fa_2_412/A sky130_fd_sc_hd__ha_2_108/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_308/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_319 sky130_fd_sc_hd__fa_2_417/B sky130_fd_sc_hd__ha_2_112/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_319/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_205 sky130_fd_sc_hd__fa_2_1054/A sky130_fd_sc_hd__o22ai_1_174/Y
+ sky130_fd_sc_hd__a21oi_1_205/Y sky130_fd_sc_hd__nor2_4_13/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_216 sky130_fd_sc_hd__clkinv_1_727/Y sky130_fd_sc_hd__o21ai_1_248/Y
+ sky130_fd_sc_hd__a21oi_1_216/Y sky130_fd_sc_hd__a211o_1_9/A1 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__or2_0_11 sky130_fd_sc_hd__or2_0_11/A sky130_fd_sc_hd__or2_0_11/X
+ sky130_fd_sc_hd__or2_0_11/B VSS VDD VSS VDD sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__a21oi_1_227 sky130_fd_sc_hd__a21o_2_4/X sky130_fd_sc_hd__o22ai_1_201/Y
+ sky130_fd_sc_hd__a21oi_1_227/Y sky130_fd_sc_hd__nand2_1_333/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_2_12 sky130_fd_sc_hd__a22oi_2_12/A1 sky130_fd_sc_hd__a22oi_2_12/A2
+ sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__buf_2_70/X sky130_fd_sc_hd__a22oi_2_12/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__a21oi_1_238 sky130_fd_sc_hd__fa_2_1081/A sky130_fd_sc_hd__o21ai_1_273/Y
+ sky130_fd_sc_hd__a21oi_1_238/Y sky130_fd_sc_hd__nor2_4_12/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_2_23 sky130_fd_sc_hd__buf_2_165/X sky130_fd_sc_hd__a22oi_2_23/A2
+ sky130_fd_sc_hd__nor2_4_7/Y sky130_fd_sc_hd__a22oi_2_23/B2 sky130_fd_sc_hd__nand4_1_56/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__a21oi_1_249 sky130_fd_sc_hd__o21a_1_24/B1 sky130_fd_sc_hd__o21a_1_23/A1
+ sky130_fd_sc_hd__dfxtp_1_891/D sky130_fd_sc_hd__nor2_1_150/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nand2_1_210 sky130_fd_sc_hd__nand2_1_210/Y sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__or4_1_2/C VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_221 sky130_fd_sc_hd__o22ai_1_59/B2 sky130_fd_sc_hd__o21ai_1_39/B1
+ sky130_fd_sc_hd__o21ai_1_39/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_820 sky130_fd_sc_hd__o22ai_1_244/A1 sky130_fd_sc_hd__o21ai_1_298/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_820/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_232 sky130_fd_sc_hd__xnor2_1_44/B sky130_fd_sc_hd__o21ai_1_78/B1
+ sky130_fd_sc_hd__o21ai_1_85/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_831 sky130_fd_sc_hd__nor2_1_147/B sky130_fd_sc_hd__fa_2_1128/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_831/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_243 sky130_fd_sc_hd__o21ai_1_87/B1 sky130_fd_sc_hd__nor2_1_56/B
+ sky130_fd_sc_hd__nor2_1_56/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_190 sky130_fd_sc_hd__o21a_1_16/A2 sky130_fd_sc_hd__nor2_1_115/B
+ sky130_fd_sc_hd__nor2_1_134/B sky130_fd_sc_hd__o22ai_1_190/A1 sky130_fd_sc_hd__o22ai_1_206/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_842 sky130_fd_sc_hd__o22ai_1_259/B1 sky130_fd_sc_hd__fa_2_1157/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_842/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_254 sky130_fd_sc_hd__o21a_1_4/B1 sky130_fd_sc_hd__fa_2_984/A
+ sky130_fd_sc_hd__o21a_1_4/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_853 sky130_fd_sc_hd__o22ai_1_264/A1 sky130_fd_sc_hd__fa_2_1148/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_853/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_265 sky130_fd_sc_hd__o211ai_1_6/C1 sky130_fd_sc_hd__fa_2_988/A
+ sky130_fd_sc_hd__nor2_4_10/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_864 sky130_fd_sc_hd__or2_0_10/B sky130_fd_sc_hd__nor2_1_225/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_864/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_276 sky130_fd_sc_hd__nand2_1_276/Y sky130_fd_sc_hd__a211o_1_8/A2
+ sky130_fd_sc_hd__nand2_1_276/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_875 sky130_fd_sc_hd__nor2_1_196/A sky130_fd_sc_hd__nor2_1_197/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_875/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_287 sky130_fd_sc_hd__xnor2_1_65/B sky130_fd_sc_hd__nand2_1_287/B
+ sky130_fd_sc_hd__nand2_1_300/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_886 sky130_fd_sc_hd__o22ai_1_292/A1 sky130_fd_sc_hd__or3_1_3/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_886/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand4_1_60 sky130_fd_sc_hd__nand4_1_60/C sky130_fd_sc_hd__nand4_1_60/B
+ sky130_fd_sc_hd__nand4_1_60/Y sky130_fd_sc_hd__nand4_1_60/D sky130_fd_sc_hd__nand4_1_60/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand2_1_298 sky130_fd_sc_hd__nand2_1_298/Y sky130_fd_sc_hd__nor2_1_108/B
+ sky130_fd_sc_hd__fa_2_1112/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_897 sky130_fd_sc_hd__nand2_1_421/B sky130_fd_sc_hd__fa_2_292/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_897/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand4_1_71 sky130_fd_sc_hd__nand4_1_71/C sky130_fd_sc_hd__nand4_1_71/B
+ sky130_fd_sc_hd__nand2_1_8/B sky130_fd_sc_hd__nand4_1_71/D sky130_fd_sc_hd__nand4_1_71/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_82 sky130_fd_sc_hd__xnor2_1_13/Y sky130_fd_sc_hd__xnor2_1_14/Y
+ sky130_fd_sc_hd__nor3_1_28/A sky130_fd_sc_hd__xnor2_1_12/Y sky130_fd_sc_hd__nor4_1_3/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__conb_1_20 sky130_fd_sc_hd__conb_1_20/LO sky130_fd_sc_hd__conb_1_20/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__mux2_2_4 VSS VDD sky130_fd_sc_hd__mux2_2_4/A1 sky130_fd_sc_hd__mux2_2_4/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_4/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__a21boi_0_4 sky130_fd_sc_hd__a21oi_1_237/Y sky130_fd_sc_hd__a21boi_0_4/Y
+ sky130_fd_sc_hd__fa_2_1071/A sky130_fd_sc_hd__a21o_2_5/A2 VSS VDD VDD VSS sky130_fd_sc_hd__a21boi_0
Xsky130_fd_sc_hd__fa_2_1160 sky130_fd_sc_hd__fa_2_1161/CIN sky130_fd_sc_hd__mux2_2_121/A1
+ sky130_fd_sc_hd__fa_2_1160/A sky130_fd_sc_hd__fa_2_1172/B sky130_fd_sc_hd__fa_2_1160/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1171 sky130_fd_sc_hd__fa_2_1172/CIN sky130_fd_sc_hd__nand2_1_362/A
+ sky130_fd_sc_hd__fa_2_1171/A sky130_fd_sc_hd__fa_2_1172/B sky130_fd_sc_hd__fa_2_1171/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1182 sky130_fd_sc_hd__fa_2_1183/CIN sky130_fd_sc_hd__mux2_2_144/A1
+ sky130_fd_sc_hd__fa_2_1182/A sky130_fd_sc_hd__fa_2_1182/B sky130_fd_sc_hd__fa_2_1182/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1193 sky130_fd_sc_hd__fa_2_1194/CIN sky130_fd_sc_hd__mux2_2_164/A1
+ sky130_fd_sc_hd__fa_2_1193/A sky130_fd_sc_hd__fa_2_1193/B sky130_fd_sc_hd__fa_2_1193/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a211o_1_18 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_178/A sky130_fd_sc_hd__o21ai_1_294/Y
+ sky130_fd_sc_hd__nor2_1_165/Y sky130_fd_sc_hd__nor2b_1_104/Y sky130_fd_sc_hd__o22ai_1_241/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__a211o_1_29 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_317/A sky130_fd_sc_hd__nor2b_1_126/Y
+ sky130_fd_sc_hd__o22ai_1_411/Y sky130_fd_sc_hd__o21ai_1_456/Y sky130_fd_sc_hd__o22ai_1_410/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o2bb2ai_1_0 sky130_fd_sc_hd__maj3_1_1/C sky130_fd_sc_hd__o22ai_1_0/B2
+ sky130_fd_sc_hd__xnor2_1_19/Y sky130_fd_sc_hd__nor2_1_10/Y sky130_fd_sc_hd__o22ai_1_0/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__clkinv_1_105 sky130_fd_sc_hd__clkinv_1_106/A sky130_fd_sc_hd__ha_2_39/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_105/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_116 sky130_fd_sc_hd__bufinv_8_2/A sky130_fd_sc_hd__buf_8_87/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_116/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_127 sky130_fd_sc_hd__nand3_1_35/C sky130_fd_sc_hd__nand3_4_1/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_127/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_138 sky130_fd_sc_hd__clkinv_1_139/A sky130_fd_sc_hd__clkinv_1_138/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_138/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_149 sky130_fd_sc_hd__clkinv_1_150/A sky130_fd_sc_hd__and2_2_1/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_149/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_18 sky130_fd_sc_hd__nor2_4_4/Y sky130_fd_sc_hd__ha_2_72/A
+ sky130_fd_sc_hd__a22o_1_18/X sky130_fd_sc_hd__a22o_1_18/B2 sky130_fd_sc_hd__a22o_2_6/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_29 sky130_fd_sc_hd__or2_1_1/B sky130_fd_sc_hd__ha_2_82/A
+ sky130_fd_sc_hd__buf_2_158/A sky130_fd_sc_hd__a22o_1_29/B2 sky130_fd_sc_hd__a22o_4_0/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__o21ai_1_5 VSS VDD sky130_fd_sc_hd__xor2_1_11/X sky130_fd_sc_hd__nor2_1_21/A
+ sky130_fd_sc_hd__a21oi_1_3/Y sky130_fd_sc_hd__o21ai_1_5/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__bufbuf_16_4 sky130_fd_sc_hd__buf_8_72/A sky130_fd_sc_hd__buf_12_164/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__nor2_1_210 sky130_fd_sc_hd__nor2_1_210/B sky130_fd_sc_hd__nor2_1_210/Y
+ sky130_fd_sc_hd__nor2_1_210/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_221 sky130_fd_sc_hd__nor2_1_221/B sky130_fd_sc_hd__nor2_1_221/Y
+ sky130_fd_sc_hd__nor2_1_224/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_232 sky130_fd_sc_hd__nor2_1_232/B sky130_fd_sc_hd__nor2_1_232/Y
+ sky130_fd_sc_hd__o21a_1_48/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_243 sky130_fd_sc_hd__nor2_1_243/B sky130_fd_sc_hd__nor2_1_243/Y
+ sky130_fd_sc_hd__nor2_4_18/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_254 sky130_fd_sc_hd__nor2_1_254/B sky130_fd_sc_hd__nor2_1_254/Y
+ sky130_fd_sc_hd__nor2_1_254/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_2_8 sky130_fd_sc_hd__clkinv_2_8/Y sky130_fd_sc_hd__clkinv_2_8/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_8/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__nor2_1_265 sky130_fd_sc_hd__o21a_1_55/A1 sky130_fd_sc_hd__nor2_1_265/Y
+ sky130_fd_sc_hd__nor2_1_265/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_276 sky130_fd_sc_hd__nor2_1_276/B sky130_fd_sc_hd__nor2_1_276/Y
+ sky130_fd_sc_hd__nor2_1_276/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_287 sky130_fd_sc_hd__nor2_1_290/A sky130_fd_sc_hd__nor2_1_287/Y
+ sky130_fd_sc_hd__nor2_1_287/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_298 sky130_fd_sc_hd__or3_1_5/X sky130_fd_sc_hd__nor2_1_298/Y
+ sky130_fd_sc_hd__fa_2_26/SUM VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_450 sky130_fd_sc_hd__buf_6_70/X sky130_fd_sc_hd__buf_12_502/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_461 sky130_fd_sc_hd__buf_12_461/A sky130_fd_sc_hd__buf_12_461/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_320 sky130_fd_sc_hd__nor3_1_25/Y sky130_fd_sc_hd__nor2_2_5/Y
+ sky130_fd_sc_hd__buf_2_203/X sky130_fd_sc_hd__clkbuf_1_458/X sky130_fd_sc_hd__nand4_1_79/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_472 sky130_fd_sc_hd__buf_6_79/X sky130_fd_sc_hd__buf_12_483/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_331 sky130_fd_sc_hd__clkinv_1_545/Y sky130_fd_sc_hd__a211o_1_7/A2
+ sky130_fd_sc_hd__nand2_1_264/A sky130_fd_sc_hd__a211o_1_6/A1 sky130_fd_sc_hd__o211ai_1_8/C1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_483 sky130_fd_sc_hd__buf_12_483/A sky130_fd_sc_hd__buf_12_516/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_342 sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_2_7/Y
+ sky130_fd_sc_hd__fa_2_998/A sky130_fd_sc_hd__fa_2_999/A sky130_fd_sc_hd__a22oi_1_342/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_494 sky130_fd_sc_hd__buf_12_494/A sky130_fd_sc_hd__buf_12_494/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_353 sky130_fd_sc_hd__clkinv_1_705/Y sky130_fd_sc_hd__nand2_1_333/B
+ sky130_fd_sc_hd__nand2_1_321/A sky130_fd_sc_hd__o21ai_1_233/Y sky130_fd_sc_hd__a22oi_1_353/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_364 sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__nor2_4_13/Y
+ sky130_fd_sc_hd__fa_2_1076/A sky130_fd_sc_hd__fa_2_1077/A sky130_fd_sc_hd__a22oi_1_364/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_375 sky130_fd_sc_hd__fa_2_1130/A sky130_fd_sc_hd__nor2_1_182/Y
+ sky130_fd_sc_hd__nor2_1_180/Y sky130_fd_sc_hd__fa_2_1126/A sky130_fd_sc_hd__a22oi_1_375/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_386 sky130_fd_sc_hd__nor2_1_222/Y sky130_fd_sc_hd__nor2_1_224/Y
+ sky130_fd_sc_hd__fa_2_1199/A sky130_fd_sc_hd__fa_2_1195/A sky130_fd_sc_hd__a22oi_1_386/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_397 sky130_fd_sc_hd__nor2_1_307/Y sky130_fd_sc_hd__nor2_1_309/Y
+ sky130_fd_sc_hd__fa_2_1284/A sky130_fd_sc_hd__fa_2_1280/A sky130_fd_sc_hd__a22oi_1_397/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_650 sky130_fd_sc_hd__nor2_1_97/B sky130_fd_sc_hd__nand2_1_306/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_650/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_19 sky130_fd_sc_hd__nor3_1_4/A sky130_fd_sc_hd__nor3_2_1/A
+ sky130_fd_sc_hd__nand2_1_19/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_661 sky130_fd_sc_hd__clkinv_1_661/Y sky130_fd_sc_hd__nor2_1_92/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_661/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_672 sky130_fd_sc_hd__o21ai_1_193/A1 sky130_fd_sc_hd__nand2_1_295/Y
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_683 sky130_fd_sc_hd__nor2_1_101/B sky130_fd_sc_hd__fa_2_1115/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_683/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_694 sky130_fd_sc_hd__clkinv_1_694/Y sky130_fd_sc_hd__nand2_1_320/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_694/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand3_1_1 sky130_fd_sc_hd__nand3_1_1/Y sky130_fd_sc_hd__nand3_1_1/A
+ sky130_fd_sc_hd__nand3_1_1/C sky130_fd_sc_hd__nand3_1_1/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__sdlclkp_2_13 sky130_fd_sc_hd__conb_1_29/LO sky130_fd_sc_hd__clkinv_8_17/A
+ sky130_fd_sc_hd__dfxtp_1_1461/CLK sky130_fd_sc_hd__nand2b_1_18/Y VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__xnor2_1_50 VSS VDD sky130_fd_sc_hd__xnor2_1_50/B sky130_fd_sc_hd__xnor2_1_50/Y
+ sky130_fd_sc_hd__nor2_1_46/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_61 VSS VDD sky130_fd_sc_hd__o21a_1_1/B1 sky130_fd_sc_hd__xnor2_1_61/Y
+ sky130_fd_sc_hd__fa_2_991/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_72 VSS VDD sky130_fd_sc_hd__xnor2_1_73/B sky130_fd_sc_hd__xnor2_1_72/Y
+ sky130_fd_sc_hd__xnor2_1_72/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_83 VSS VDD sky130_fd_sc_hd__xnor2_1_83/B sky130_fd_sc_hd__xnor2_1_83/Y
+ sky130_fd_sc_hd__nor2_1_97/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_94 VSS VDD sky130_fd_sc_hd__xnor2_1_94/B sky130_fd_sc_hd__xnor2_1_94/Y
+ sky130_fd_sc_hd__fa_2_1190/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__dfxtp_1_808 VDD VSS sky130_fd_sc_hd__fa_2_1060/A sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__mux2_2_57/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_819 VDD VSS sky130_fd_sc_hd__fa_2_1093/A sky130_fd_sc_hd__clkinv_8_59/Y
+ sky130_fd_sc_hd__and2_0_295/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_406 VSS VDD sky130_fd_sc_hd__clkbuf_1_406/X sky130_fd_sc_hd__clkbuf_1_406/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_417 VSS VDD sky130_fd_sc_hd__clkbuf_1_417/X sky130_fd_sc_hd__clkbuf_1_417/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_428 VSS VDD sky130_fd_sc_hd__clkbuf_1_428/X sky130_fd_sc_hd__clkbuf_1_428/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_439 VSS VDD sky130_fd_sc_hd__a22oi_2_30/A2 sky130_fd_sc_hd__clkbuf_1_439/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o32ai_1_0 sky130_fd_sc_hd__o32ai_1_0/A2 sky130_fd_sc_hd__o32ai_1_0/Y
+ sky130_fd_sc_hd__fa_2_1124/A sky130_fd_sc_hd__o32ai_1_0/A3 sky130_fd_sc_hd__o32ai_1_0/B2
+ sky130_fd_sc_hd__fa_2_1123/A VDD VSS VSS VDD sky130_fd_sc_hd__o32ai_1
Xsky130_fd_sc_hd__diode_2_180 sky130_fd_sc_hd__a22o_4_0/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_191 sky130_fd_sc_hd__buf_2_144/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkinv_2_13 sky130_fd_sc_hd__clkinv_2_13/Y sky130_fd_sc_hd__clkinv_2_13/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_13/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkbuf_4_200 sky130_fd_sc_hd__nand4_1_68/D sky130_fd_sc_hd__a22oi_1_273/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_2_24 sky130_fd_sc_hd__nand4_1_75/D sky130_fd_sc_hd__clkinv_2_24/A
+ VSS VDD VDD VSS VSS sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkbuf_4_211 sky130_fd_sc_hd__clkbuf_4_211/X sky130_fd_sc_hd__a21oi_1_16/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_2_35 sky130_fd_sc_hd__clkinv_2_35/Y sky130_fd_sc_hd__clkinv_2_35/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_35/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkbuf_4_222 sky130_fd_sc_hd__a22oi_1_7/A2 sig_amplitude[4] VSS
+ VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_2_46 sky130_fd_sc_hd__clkinv_4_56/A sky130_fd_sc_hd__clkinv_2_47/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_46/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__sdlclkp_4_9 sky130_fd_sc_hd__conb_1_4/LO sky130_fd_sc_hd__clkinv_8_112/A
+ sky130_fd_sc_hd__dfxtp_1_8/CLK sky130_fd_sc_hd__buf_6_86/X VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__buf_12_280 sky130_fd_sc_hd__inv_2_101/Y sky130_fd_sc_hd__buf_12_363/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_291 sky130_fd_sc_hd__buf_6_40/X sky130_fd_sc_hd__buf_12_291/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_150 sky130_fd_sc_hd__clkbuf_1_264/X sky130_fd_sc_hd__nor2_2_3/Y
+ sky130_fd_sc_hd__a22oi_1_150/B2 sky130_fd_sc_hd__clkbuf_4_137/X sky130_fd_sc_hd__nand4_1_32/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_161 sky130_fd_sc_hd__clkbuf_4_111/X sky130_fd_sc_hd__clkbuf_4_112/X
+ sky130_fd_sc_hd__a22oi_1_161/B2 sky130_fd_sc_hd__clkbuf_1_294/X sky130_fd_sc_hd__a22oi_1_161/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_172 sky130_fd_sc_hd__clkbuf_1_351/X sky130_fd_sc_hd__clkbuf_1_353/X
+ sky130_fd_sc_hd__clkbuf_4_118/X sky130_fd_sc_hd__a22oi_1_172/A2 sky130_fd_sc_hd__nand4_1_38/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_183 sky130_fd_sc_hd__clkbuf_1_265/X sky130_fd_sc_hd__clkbuf_1_266/X
+ sky130_fd_sc_hd__clkbuf_1_273/X sky130_fd_sc_hd__a22oi_1_183/A2 sky130_fd_sc_hd__a22oi_1_183/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_194 sky130_fd_sc_hd__clkbuf_1_264/X sky130_fd_sc_hd__nor2_2_3/Y
+ sky130_fd_sc_hd__a22oi_1_194/B2 sky130_fd_sc_hd__clkbuf_4_126/X sky130_fd_sc_hd__nand4_1_43/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_480 sky130_fd_sc_hd__o22ai_1_85/B2 sky130_fd_sc_hd__ha_2_174/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_480/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_491 sky130_fd_sc_hd__nor2_1_46/B sky130_fd_sc_hd__nand2_1_248/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_491/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_405 VSS VDD sky130_fd_sc_hd__o21ai_1_414/A1 sky130_fd_sc_hd__nor2_1_265/A
+ sky130_fd_sc_hd__a21oi_1_391/Y sky130_fd_sc_hd__xor2_1_267/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_416 VSS VDD sky130_fd_sc_hd__nor2_1_229/B sky130_fd_sc_hd__o21a_1_55/A1
+ sky130_fd_sc_hd__a21oi_1_400/Y sky130_fd_sc_hd__o21ai_1_416/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_427 VSS VDD sky130_fd_sc_hd__a211oi_1_30/Y sky130_fd_sc_hd__nor2_1_257/A
+ sky130_fd_sc_hd__a21oi_1_408/Y sky130_fd_sc_hd__o21ai_1_427/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_438 VSS VDD sky130_fd_sc_hd__nor2_1_288/Y sky130_fd_sc_hd__or3_1_5/C
+ sky130_fd_sc_hd__nor2_1_286/A sky130_fd_sc_hd__o21ai_1_438/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_449 VSS VDD sky130_fd_sc_hd__xor2_1_275/X sky130_fd_sc_hd__xnor2_1_0/Y
+ sky130_fd_sc_hd__nor2_1_286/A sky130_fd_sc_hd__o21ai_1_449/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_4_14 sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__nor2_4_15/A
+ sky130_fd_sc_hd__nor2_4_14/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__xor2_1_210 sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__fa_2_1208/B
+ sky130_fd_sc_hd__xor2_1_210/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_221 sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__fa_2_1197/B
+ sky130_fd_sc_hd__xor2_1_221/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_232 sky130_fd_sc_hd__xor2_1_233/X sky130_fd_sc_hd__xor2_1_232/X
+ sky130_fd_sc_hd__xor2_1_254/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_243 sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1232/B
+ sky130_fd_sc_hd__xor2_1_243/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_254 sky130_fd_sc_hd__xor2_1_267/B sky130_fd_sc_hd__xor2_1_254/X
+ sky130_fd_sc_hd__xor2_1_254/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_605 VDD VSS sky130_fd_sc_hd__and2_0_215/A sky130_fd_sc_hd__dfxtp_1_606/CLK
+ sky130_fd_sc_hd__fa_2_1025/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_265 sky130_fd_sc_hd__xor2_1_267/B sky130_fd_sc_hd__fa_2_1249/B
+ sky130_fd_sc_hd__xor2_1_265/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_616 VDD VSS sky130_fd_sc_hd__fa_2_811/A sky130_fd_sc_hd__dfxtp_1_627/CLK
+ sky130_fd_sc_hd__a21oi_1_78/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_276 sky130_fd_sc_hd__xor2_1_276/B sky130_fd_sc_hd__xor2_1_276/X
+ sky130_fd_sc_hd__xor2_1_277/X VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_627 VDD VSS sky130_fd_sc_hd__fa_2_833/A sky130_fd_sc_hd__dfxtp_1_627/CLK
+ sky130_fd_sc_hd__xnor2_1_61/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_287 sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1284/B
+ sky130_fd_sc_hd__xor2_1_287/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_638 VDD VSS sky130_fd_sc_hd__fa_2_1002/A sky130_fd_sc_hd__clkinv_8_44/Y
+ sky130_fd_sc_hd__mux2_2_29/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_298 sky130_fd_sc_hd__xor2_1_299/X sky130_fd_sc_hd__xor2_1_298/X
+ sky130_fd_sc_hd__xor2_1_298/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_649 VDD VSS sky130_fd_sc_hd__fa_2_1013/A sky130_fd_sc_hd__clkinv_8_44/Y
+ sky130_fd_sc_hd__mux2_2_6/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_203 VSS VDD sky130_fd_sc_hd__buf_8_87/A sky130_fd_sc_hd__buf_12_133/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_214 VSS VDD sky130_fd_sc_hd__buf_12_137/A sky130_fd_sc_hd__inv_2_50/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_225 VSS VDD sky130_fd_sc_hd__buf_8_110/A sky130_fd_sc_hd__buf_2_121/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_236 VSS VDD sky130_fd_sc_hd__clkbuf_1_236/X sky130_fd_sc_hd__buf_8_92/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_247 VSS VDD sky130_fd_sc_hd__clkbuf_1_247/X sky130_fd_sc_hd__clkbuf_1_247/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_258 VSS VDD sky130_fd_sc_hd__clkbuf_4_74/A sky130_fd_sc_hd__clkbuf_1_258/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_269 VSS VDD sky130_fd_sc_hd__clkbuf_1_269/X sky130_fd_sc_hd__clkbuf_1_269/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_2_70 VDD VSS sky130_fd_sc_hd__buf_2_70/X sky130_fd_sc_hd__buf_2_70/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_81 VDD VSS sky130_fd_sc_hd__buf_2_81/X sky130_fd_sc_hd__buf_2_81/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_92 VDD VSS sky130_fd_sc_hd__buf_2_92/X sky130_fd_sc_hd__buf_2_92/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_4_8 VDD VSS sky130_fd_sc_hd__buf_4_8/X sky130_fd_sc_hd__buf_4_8/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__and2_0_201 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_201/X sky130_fd_sc_hd__and2_0_235/B
+ sky130_fd_sc_hd__and2_0_201/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_212 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_212/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_212/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_223 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_223/X sky130_fd_sc_hd__and2_0_235/B
+ sky130_fd_sc_hd__and2_0_223/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_234 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_234/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_234/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_245 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_245/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__and2_0_245/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_256 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_256/X sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__and2_0_256/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_267 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_267/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__fa_2_968/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_278 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_278/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__fa_2_971/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_289 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_289/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__fa_2_975/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__sdlclkp_2_6 sky130_fd_sc_hd__conb_1_15/LO sky130_fd_sc_hd__clkinv_8_100/Y
+ sky130_fd_sc_hd__dfxtp_1_223/CLK sky130_fd_sc_hd__or2_0_3/X VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__a22o_2_0 sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__ha_2_64/A
+ sky130_fd_sc_hd__a22o_2_0/X sky130_fd_sc_hd__dfxtp_1_7/Q sky130_fd_sc_hd__a22o_2_3/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_2
Xsky130_fd_sc_hd__o21ai_1_202 VSS VDD sky130_fd_sc_hd__xnor2_1_76/A sky130_fd_sc_hd__nor2_1_109/Y
+ sky130_fd_sc_hd__nand2_1_297/Y sky130_fd_sc_hd__xnor2_1_78/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_20 sky130_fd_sc_hd__clkbuf_4_20/X sky130_fd_sc_hd__clkbuf_4_20/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_213 VSS VDD sky130_fd_sc_hd__a21oi_1_204/Y sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__nand2_1_317/Y sky130_fd_sc_hd__xor2_1_117/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_31 sky130_fd_sc_hd__clkbuf_4_31/X sky130_fd_sc_hd__clkbuf_4_31/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_224 VSS VDD sky130_fd_sc_hd__a21oi_1_197/Y sky130_fd_sc_hd__nor2_1_126/A
+ sky130_fd_sc_hd__nand2_1_321/Y sky130_fd_sc_hd__o21ai_1_224/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_42 sky130_fd_sc_hd__nand4_1_15/D sky130_fd_sc_hd__a22oi_1_80/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_235 VSS VDD sky130_fd_sc_hd__o22ai_1_204/B1 sky130_fd_sc_hd__nand4_1_86/B
+ sky130_fd_sc_hd__a21oi_1_209/Y sky130_fd_sc_hd__o21ai_1_235/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_53 sky130_fd_sc_hd__nand4_1_4/D sky130_fd_sc_hd__a22oi_1_43/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_246 VSS VDD sky130_fd_sc_hd__a21oi_1_220/Y sky130_fd_sc_hd__nor2_1_127/A
+ sky130_fd_sc_hd__nand2b_1_16/Y sky130_fd_sc_hd__o21ai_1_246/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_64 sky130_fd_sc_hd__clkbuf_4_64/X sky130_fd_sc_hd__clkbuf_4_64/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_257 VSS VDD sky130_fd_sc_hd__o21ai_1_271/A2 sky130_fd_sc_hd__o21a_1_16/A2
+ sky130_fd_sc_hd__a21oi_1_222/Y sky130_fd_sc_hd__a211o_1_9/A2 VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_75 sky130_fd_sc_hd__clkbuf_4_75/X sky130_fd_sc_hd__clkbuf_4_75/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_268 VSS VDD sky130_fd_sc_hd__nor2_1_126/A sky130_fd_sc_hd__a21oi_1_235/Y
+ sky130_fd_sc_hd__a21oi_1_232/Y sky130_fd_sc_hd__xor2_1_110/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_86 sky130_fd_sc_hd__clkbuf_4_86/X sky130_fd_sc_hd__clkbuf_4_86/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_279 VSS VDD sky130_fd_sc_hd__nand2_1_369/B sky130_fd_sc_hd__a21o_2_8/B1
+ sky130_fd_sc_hd__a21o_2_7/A2 sky130_fd_sc_hd__o21ai_1_279/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_97 sky130_fd_sc_hd__inv_2_73/A sky130_fd_sc_hd__clkbuf_4_97/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_8_170 sky130_fd_sc_hd__buf_8_170/A sky130_fd_sc_hd__buf_8_170/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_181 sky130_fd_sc_hd__buf_8_186/A sky130_fd_sc_hd__buf_8_220/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_192 sky130_fd_sc_hd__buf_8_192/A sky130_fd_sc_hd__buf_8_223/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_402 VDD VSS sky130_fd_sc_hd__nor2_1_59/A sky130_fd_sc_hd__dfxtp_1_424/CLK
+ sky130_fd_sc_hd__and2_0_138/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_413 VDD VSS sky130_fd_sc_hd__nor2_1_54/A sky130_fd_sc_hd__dfxtp_1_419/CLK
+ sky130_fd_sc_hd__and2_0_192/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_424 VDD VSS sky130_fd_sc_hd__fa_2_1044/B sky130_fd_sc_hd__dfxtp_1_424/CLK
+ sky130_fd_sc_hd__and2_0_104/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_435 VDD VSS sky130_fd_sc_hd__dfxtp_1_435/Q sky130_fd_sc_hd__dfxtp_1_452/CLK
+ sky130_fd_sc_hd__nand2_1_94/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_446 VDD VSS sky130_fd_sc_hd__dfxtp_1_992/D sky130_fd_sc_hd__dfxtp_1_448/CLK
+ sky130_fd_sc_hd__nand2_1_72/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_457 VDD VSS sky130_fd_sc_hd__xor2_1_185/B sky130_fd_sc_hd__dfxtp_1_457/CLK
+ sky130_fd_sc_hd__nand2_1_50/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_468 VDD VSS sky130_fd_sc_hd__buf_6_3/A sky130_fd_sc_hd__dfxtp_1_473/CLK
+ sky130_fd_sc_hd__and2_0_131/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_479 VDD VSS sky130_fd_sc_hd__o21ai_1_38/A1 sky130_fd_sc_hd__dfxtp_1_483/CLK
+ sky130_fd_sc_hd__nor2b_1_81/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2b_1_16 sky130_fd_sc_hd__nand2b_1_16/Y sky130_fd_sc_hd__nor2_2_13/B
+ sky130_fd_sc_hd__xor2_1_88/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__fa_2_307 sky130_fd_sc_hd__fa_2_304/CIN sky130_fd_sc_hd__fa_2_309/CIN
+ sky130_fd_sc_hd__fa_2_424/A sky130_fd_sc_hd__fa_2_401/A sky130_fd_sc_hd__fa_2_307/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_318 sky130_fd_sc_hd__fa_2_314/CIN sky130_fd_sc_hd__or3_1_3/C
+ sky130_fd_sc_hd__fa_2_318/A sky130_fd_sc_hd__fa_2_318/B sky130_fd_sc_hd__fa_2_318/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_329 sky130_fd_sc_hd__maj3_1_76/B sky130_fd_sc_hd__maj3_1_77/A
+ sky130_fd_sc_hd__fa_2_329/A sky130_fd_sc_hd__fa_2_329/B sky130_fd_sc_hd__o22ai_1_23/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_8_12 sky130_fd_sc_hd__clkinv_8_12/Y sky130_fd_sc_hd__clkinv_4_8/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_12/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_23 sky130_fd_sc_hd__clkinv_8_24/A sky130_fd_sc_hd__clkinv_8_23/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_23/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_34 sky130_fd_sc_hd__clkinv_8_35/A sky130_fd_sc_hd__clkinv_8_34/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_45 sky130_fd_sc_hd__clkinv_8_45/Y sky130_fd_sc_hd__clkinv_8_59/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_56 sky130_fd_sc_hd__clkinv_8_56/Y sky130_fd_sc_hd__clkinv_8_56/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_10 sky130_fd_sc_hd__buf_12_10/A sky130_fd_sc_hd__buf_12_91/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_8_67 sky130_fd_sc_hd__clkinv_8_67/Y sky130_fd_sc_hd__clkinv_8_67/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_67/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_21 sky130_fd_sc_hd__inv_2_30/Y sky130_fd_sc_hd__buf_12_21/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_8_78 sky130_fd_sc_hd__clkinv_8_78/Y sky130_fd_sc_hd__clkinv_8_78/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_78/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_32 sky130_fd_sc_hd__buf_8_54/X sky130_fd_sc_hd__buf_12_96/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_8_89 sky130_fd_sc_hd__clkinv_8_90/A sky130_fd_sc_hd__clkinv_8_89/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_43 sky130_fd_sc_hd__buf_8_46/X sky130_fd_sc_hd__buf_12_43/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_54 sky130_fd_sc_hd__buf_8_29/X sky130_fd_sc_hd__buf_12_54/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_65 sky130_fd_sc_hd__buf_4_31/X sky130_fd_sc_hd__buf_12_65/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_76 sky130_fd_sc_hd__buf_4_19/X sky130_fd_sc_hd__buf_12_76/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_87 sky130_fd_sc_hd__buf_6_18/X sky130_fd_sc_hd__buf_12_87/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_98 sky130_fd_sc_hd__buf_12_98/A sky130_fd_sc_hd__buf_12_98/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_2_5 VDD VSS sky130_fd_sc_hd__buf_2_5/X sky130_fd_sc_hd__buf_6_7/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1320 VDD VSS sky130_fd_sc_hd__fa_2_904/A sky130_fd_sc_hd__dfxtp_1_1322/CLK
+ sky130_fd_sc_hd__o21a_1_61/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1331 VDD VSS sky130_fd_sc_hd__fa_2_915/A sky130_fd_sc_hd__dfxtp_1_1332/CLK
+ sky130_fd_sc_hd__o21a_1_56/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1342 VDD VSS sky130_fd_sc_hd__fa_2_1301/A sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__mux2_2_242/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1353 VDD VSS sky130_fd_sc_hd__fa_2_1275/B sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__and2_0_334/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1364 VDD VSS sky130_fd_sc_hd__fa_2_1286/A sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__mux2_2_235/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1375 VDD VSS sky130_fd_sc_hd__fa_2_1314/A sky130_fd_sc_hd__clkinv_8_102/Y
+ sky130_fd_sc_hd__mux2_2_264/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1386 VDD VSS sky130_fd_sc_hd__fa_2_1325/A sky130_fd_sc_hd__clkinv_8_75/Y
+ sky130_fd_sc_hd__nand2_1_519/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1397 VDD VSS sky130_fd_sc_hd__mux2_2_252/A0 sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__o22ai_1_392/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_980 VDD VSS sky130_fd_sc_hd__mux2_2_91/A0 sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__o22ai_1_215/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_991 VDD VSS sky130_fd_sc_hd__mux2_2_120/A0 sky130_fd_sc_hd__clkinv_8_64/Y
+ sky130_fd_sc_hd__dfxtp_1_991/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_830 sky130_fd_sc_hd__fa_2_706/A sky130_fd_sc_hd__fa_2_707/B
+ sky130_fd_sc_hd__fa_2_834/B sky130_fd_sc_hd__fa_2_830/B sky130_fd_sc_hd__fa_2_833/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_190 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_190/A sky130_fd_sc_hd__ha_2_189/A
+ sky130_fd_sc_hd__ha_2_190/SUM sky130_fd_sc_hd__ha_2_190/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_841 sky130_fd_sc_hd__fa_2_840/CIN sky130_fd_sc_hd__fa_2_841/SUM
+ sky130_fd_sc_hd__fa_2_841/A sky130_fd_sc_hd__fa_2_841/B sky130_fd_sc_hd__fa_2_841/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_852 sky130_fd_sc_hd__fa_2_851/CIN sky130_fd_sc_hd__fa_2_852/SUM
+ sky130_fd_sc_hd__fa_2_852/A sky130_fd_sc_hd__fa_2_852/B sky130_fd_sc_hd__fa_2_852/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_863 sky130_fd_sc_hd__fa_2_862/CIN sky130_fd_sc_hd__fa_2_863/SUM
+ sky130_fd_sc_hd__fa_2_863/A sky130_fd_sc_hd__fa_2_863/B sky130_fd_sc_hd__fa_2_863/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_874 sky130_fd_sc_hd__fa_2_873/CIN sky130_fd_sc_hd__fa_2_874/SUM
+ sky130_fd_sc_hd__fa_2_874/A sky130_fd_sc_hd__fa_2_874/B sky130_fd_sc_hd__fa_2_874/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_885 sky130_fd_sc_hd__fa_2_884/CIN sky130_fd_sc_hd__nand2_1_45/B
+ sky130_fd_sc_hd__ha_2_156/A sky130_fd_sc_hd__fa_2_885/B sky130_fd_sc_hd__fa_2_885/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_896 sky130_fd_sc_hd__fa_2_895/CIN sky130_fd_sc_hd__fa_2_896/SUM
+ sky130_fd_sc_hd__fa_2_896/A sky130_fd_sc_hd__fa_2_896/B sky130_fd_sc_hd__fa_2_896/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_5 sky130_fd_sc_hd__inv_2_5/A sky130_fd_sc_hd__inv_2_5/Y VDD
+ VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__nor3_2_7 sky130_fd_sc_hd__nor3_2_9/B sky130_fd_sc_hd__nor3_2_7/Y
+ sky130_fd_sc_hd__nor3_2_9/A sky130_fd_sc_hd__nor3_2_8/A VDD VSS VSS VDD sky130_fd_sc_hd__nor3_2
Xsky130_fd_sc_hd__nor2_1_15 sky130_fd_sc_hd__inv_4_1/A sky130_fd_sc_hd__nor2_1_15/Y
+ sky130_fd_sc_hd__ha_2_167/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_26 sky130_fd_sc_hd__nor2_1_26/B sky130_fd_sc_hd__nor2_1_26/Y
+ sky130_fd_sc_hd__nor3_1_31/C VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_130 VSS VDD sky130_fd_sc_hd__mux2_2_130/A1 sky130_fd_sc_hd__mux2_2_130/A0
+ sky130_fd_sc_hd__mux2_2_135/S sky130_fd_sc_hd__mux2_2_130/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_37 sky130_fd_sc_hd__nor2_1_37/B sky130_fd_sc_hd__nor3_1_36/C
+ sky130_fd_sc_hd__nor2_1_37/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_141 VSS VDD sky130_fd_sc_hd__mux2_2_141/A1 sky130_fd_sc_hd__mux2_2_141/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_141/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_48 sky130_fd_sc_hd__nor2_1_48/B sky130_fd_sc_hd__nor2_1_48/Y
+ sky130_fd_sc_hd__nor2_1_49/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_152 VSS VDD sky130_fd_sc_hd__mux2_2_152/A1 sky130_fd_sc_hd__mux2_2_152/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_152/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_59 sky130_fd_sc_hd__nor2_1_59/B sky130_fd_sc_hd__nor2_1_59/Y
+ sky130_fd_sc_hd__nor2_1_59/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_163 VSS VDD sky130_fd_sc_hd__mux2_2_163/A1 sky130_fd_sc_hd__mux2_2_163/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_163/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_174 VSS VDD sky130_fd_sc_hd__mux2_2_174/A1 sky130_fd_sc_hd__mux2_2_174/A0
+ sky130_fd_sc_hd__nor2_8_1/A sky130_fd_sc_hd__mux2_2_174/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_185 VSS VDD sky130_fd_sc_hd__mux2_2_185/A1 sky130_fd_sc_hd__mux2_2_185/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_185/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_196 VSS VDD sky130_fd_sc_hd__mux2_2_196/A1 sky130_fd_sc_hd__mux2_2_196/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_196/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__a21oi_1_409 sky130_fd_sc_hd__nand2_1_491/B sky130_fd_sc_hd__o22ai_1_369/Y
+ sky130_fd_sc_hd__a21oi_1_409/Y sky130_fd_sc_hd__o21ai_1_437/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__maj3_1_101 sky130_fd_sc_hd__maj3_1_102/X sky130_fd_sc_hd__maj3_1_101/X
+ sky130_fd_sc_hd__maj3_1_101/B sky130_fd_sc_hd__maj3_1_101/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_112 sky130_fd_sc_hd__maj3_1_113/X sky130_fd_sc_hd__maj3_1_112/X
+ sky130_fd_sc_hd__maj3_1_112/B sky130_fd_sc_hd__maj3_1_112/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_123 sky130_fd_sc_hd__maj3_1_124/X sky130_fd_sc_hd__maj3_1_123/X
+ sky130_fd_sc_hd__maj3_1_123/B sky130_fd_sc_hd__maj3_1_123/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__and2_0_70 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_75/A sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__ha_2_78/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_134 sky130_fd_sc_hd__fa_2_624/B sky130_fd_sc_hd__maj3_1_134/X
+ sky130_fd_sc_hd__ha_2_132/B sky130_fd_sc_hd__maj3_1_134/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_403 sky130_fd_sc_hd__o21a_1_38/B1 sky130_fd_sc_hd__fa_2_1203/A
+ sky130_fd_sc_hd__o21a_1_38/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_350 sky130_fd_sc_hd__nor2_1_268/A sky130_fd_sc_hd__nor2_1_265/A
+ sky130_fd_sc_hd__o22ai_1_350/Y sky130_fd_sc_hd__a21boi_1_6/Y sky130_fd_sc_hd__nor2_1_249/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_81 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_81/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__and2_0_81/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_145 sky130_fd_sc_hd__maj3_1_146/X sky130_fd_sc_hd__maj3_1_145/X
+ sky130_fd_sc_hd__maj3_1_145/B sky130_fd_sc_hd__maj3_1_145/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_414 sky130_fd_sc_hd__nand2_1_414/Y sky130_fd_sc_hd__mux2_2_171/S
+ sky130_fd_sc_hd__nand2_1_414/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_361 sky130_fd_sc_hd__o22ai_1_379/A2 sky130_fd_sc_hd__nor2_1_228/B
+ sky130_fd_sc_hd__o22ai_1_361/Y sky130_fd_sc_hd__o22ai_1_361/A1 sky130_fd_sc_hd__o32ai_1_8/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_92 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_92/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_92/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_156 sky130_fd_sc_hd__maj3_1_157/X sky130_fd_sc_hd__maj3_1_156/X
+ sky130_fd_sc_hd__maj3_1_156/B sky130_fd_sc_hd__maj3_1_156/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_425 sky130_fd_sc_hd__nand2_1_425/Y sky130_fd_sc_hd__xor2_1_209/A
+ sky130_fd_sc_hd__nor2_1_224/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_372 sky130_fd_sc_hd__o22ai_1_379/A2 sky130_fd_sc_hd__o22ai_1_372/B1
+ sky130_fd_sc_hd__o22ai_1_372/Y sky130_fd_sc_hd__nor2_1_239/B sky130_fd_sc_hd__o32ai_1_8/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_436 sky130_fd_sc_hd__nand2_1_436/Y sky130_fd_sc_hd__nand2_1_439/B
+ sky130_fd_sc_hd__o21ai_1_377/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_383 sky130_fd_sc_hd__nand2_1_514/Y sky130_fd_sc_hd__nand2_1_513/Y
+ sky130_fd_sc_hd__o22ai_1_383/Y sky130_fd_sc_hd__nand2_1_524/B sky130_fd_sc_hd__o21ai_1_440/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_447 sky130_fd_sc_hd__o21a_1_44/B1 sky130_fd_sc_hd__fa_2_1238/A
+ sky130_fd_sc_hd__o21a_1_44/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_394 sky130_fd_sc_hd__nand2_1_516/Y sky130_fd_sc_hd__o21ai_1_439/Y
+ sky130_fd_sc_hd__o22ai_1_394/Y sky130_fd_sc_hd__nand2_1_523/B sky130_fd_sc_hd__nand2_1_515/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_458 sky130_fd_sc_hd__o21a_1_54/B1 sky130_fd_sc_hd__fa_2_1247/A
+ sky130_fd_sc_hd__o21a_1_54/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_469 sky130_fd_sc_hd__nand2_1_469/Y sky130_fd_sc_hd__inv_2_139/Y
+ sky130_fd_sc_hd__nand2_1_469/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_16 sky130_fd_sc_hd__clkinv_1_61/Y sky130_fd_sc_hd__nor2b_1_16/Y
+ sky130_fd_sc_hd__or2_1_0/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_27 sky130_fd_sc_hd__ha_2_66/SUM sky130_fd_sc_hd__nor2b_1_27/Y
+ sky130_fd_sc_hd__or2_0_2/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1005 sky130_fd_sc_hd__o21ai_1_419/A2 sky130_fd_sc_hd__o21ai_1_430/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1005/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2b_1_38 sky130_fd_sc_hd__nor2b_1_38/B_N sky130_fd_sc_hd__nor2b_1_38/Y
+ sky130_fd_sc_hd__or2_0_3/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_49 sky130_fd_sc_hd__ha_2_84/SUM sky130_fd_sc_hd__nor2b_1_49/Y
+ sky130_fd_sc_hd__or2_0_3/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1016 sky130_fd_sc_hd__nor2_1_268/B sky130_fd_sc_hd__o21ai_1_436/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1016/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1027 sky130_fd_sc_hd__nor2_2_18/B sky130_fd_sc_hd__nor2_4_19/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1027/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1038 sky130_fd_sc_hd__nor2_1_307/A sky130_fd_sc_hd__nor2b_2_5/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1038/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_80 sky130_fd_sc_hd__ha_2_32/A sky130_fd_sc_hd__buf_8_80/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__clkinv_1_1049 sky130_fd_sc_hd__nor2_1_288/B sky130_fd_sc_hd__xor2_1_275/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1049/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_91 sky130_fd_sc_hd__buf_8_91/A sky130_fd_sc_hd__buf_8_91/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_210 VDD VSS sky130_fd_sc_hd__ha_2_71/A sky130_fd_sc_hd__dfxtp_1_212/CLK
+ sky130_fd_sc_hd__and2_0_83/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_221 VDD VSS sky130_fd_sc_hd__ha_2_82/A sky130_fd_sc_hd__dfxtp_1_223/CLK
+ sky130_fd_sc_hd__nor2b_1_46/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_232 VDD VSS sky130_fd_sc_hd__fa_2_877/A sky130_fd_sc_hd__dfxtp_1_472/CLK
+ sky130_fd_sc_hd__and2_0_179/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_243 VDD VSS sky130_fd_sc_hd__fa_2_866/A sky130_fd_sc_hd__dfxtp_1_277/CLK
+ sky130_fd_sc_hd__and2_0_173/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_254 VDD VSS sky130_fd_sc_hd__buf_2_118/A sky130_fd_sc_hd__dfxtp_1_258/CLK
+ sky130_fd_sc_hd__and2_0_235/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_265 VDD VSS sky130_fd_sc_hd__dfxtp_1_265/Q sky130_fd_sc_hd__dfxtp_1_266/CLK
+ sky130_fd_sc_hd__and2_0_234/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_276 VDD VSS sky130_fd_sc_hd__dfxtp_1_276/Q sky130_fd_sc_hd__dfxtp_1_463/CLK
+ sky130_fd_sc_hd__and2_0_208/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_287 VDD VSS sky130_fd_sc_hd__a22o_1_60/A1 sky130_fd_sc_hd__clkinv_4_31/Y
+ sky130_fd_sc_hd__nand2_1_135/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_298 VDD VSS sky130_fd_sc_hd__a22o_1_51/A1 sky130_fd_sc_hd__dfxtp_1_304/CLK
+ sky130_fd_sc_hd__and2_0_100/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o22ai_1_7 sky130_fd_sc_hd__fa_2_82/A sky130_fd_sc_hd__fa_2_2/B sky130_fd_sc_hd__o22ai_1_7/Y
+ sky130_fd_sc_hd__ha_2_97/A sky130_fd_sc_hd__fa_2_91/A VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_104 sky130_fd_sc_hd__fa_2_109/B sky130_fd_sc_hd__fa_2_104/SUM
+ sky130_fd_sc_hd__fa_2_104/A sky130_fd_sc_hd__fa_2_104/B sky130_fd_sc_hd__fa_2_104/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_115 sky130_fd_sc_hd__fa_2_116/CIN sky130_fd_sc_hd__fa_2_110/B
+ sky130_fd_sc_hd__fa_2_2/A sky130_fd_sc_hd__fa_2_91/B sky130_fd_sc_hd__fa_2_49/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_126 sky130_fd_sc_hd__fa_2_29/A sky130_fd_sc_hd__fa_2_28/B sky130_fd_sc_hd__fa_2_126/A
+ sky130_fd_sc_hd__fa_2_126/B sky130_fd_sc_hd__fa_2_130/SUM VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_137 sky130_fd_sc_hd__fa_2_136/B sky130_fd_sc_hd__fa_2_137/SUM
+ sky130_fd_sc_hd__fa_2_137/A sky130_fd_sc_hd__fa_2_137/B sky130_fd_sc_hd__fa_2_137/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_148 sky130_fd_sc_hd__fa_2_149/CIN sky130_fd_sc_hd__fa_2_148/SUM
+ sky130_fd_sc_hd__fa_2_148/A sky130_fd_sc_hd__fa_2_148/B sky130_fd_sc_hd__fa_2_148/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_159 sky130_fd_sc_hd__fa_2_152/B sky130_fd_sc_hd__fa_2_160/CIN
+ sky130_fd_sc_hd__fa_2_5/B sky130_fd_sc_hd__fa_2_32/A sky130_fd_sc_hd__fa_2_258/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_110 VDD VSS sky130_fd_sc_hd__buf_2_110/X sky130_fd_sc_hd__buf_2_110/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_121 VDD VSS sky130_fd_sc_hd__buf_2_121/X sky130_fd_sc_hd__buf_2_121/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_14 sky130_fd_sc_hd__ha_2_99/A sky130_fd_sc_hd__fa_2_273/A
+ sky130_fd_sc_hd__fa_2_197/B sky130_fd_sc_hd__ha_2_107/A sky130_fd_sc_hd__fa_2_277/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_1320 sky130_fd_sc_hd__fa_2_1321/CIN sky130_fd_sc_hd__mux2_2_250/A1
+ sky130_fd_sc_hd__fa_2_1320/A sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1320/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_132 VDD VSS sky130_fd_sc_hd__buf_2_132/X sky130_fd_sc_hd__buf_2_132/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_25 sky130_fd_sc_hd__ha_2_113/B sky130_fd_sc_hd__fa_2_422/B
+ sky130_fd_sc_hd__fa_2_363/B sky130_fd_sc_hd__ha_2_112/B sky130_fd_sc_hd__fa_2_404/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_143 VDD VSS sky130_fd_sc_hd__buf_2_143/X sky130_fd_sc_hd__buf_2_143/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_36 sky130_fd_sc_hd__ha_2_119/B sky130_fd_sc_hd__fa_2_554/A
+ sky130_fd_sc_hd__fa_2_525/A sky130_fd_sc_hd__ha_2_117/B sky130_fd_sc_hd__fa_2_551/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_154 VDD VSS sky130_fd_sc_hd__buf_4_103/A sky130_fd_sc_hd__buf_6_56/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_47 sky130_fd_sc_hd__ha_2_133/A sky130_fd_sc_hd__ha_2_132/B
+ sky130_fd_sc_hd__fa_2_676/B sky130_fd_sc_hd__fa_2_672/A sky130_fd_sc_hd__ha_2_131/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_165 VDD VSS sky130_fd_sc_hd__buf_2_165/X sky130_fd_sc_hd__buf_2_165/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_58 sky130_fd_sc_hd__o22ai_1_58/A2 sky130_fd_sc_hd__fa_2_948/A
+ sky130_fd_sc_hd__o22ai_1_58/Y sky130_fd_sc_hd__fa_2_947/A sky130_fd_sc_hd__o22ai_1_58/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_176 VDD VSS sky130_fd_sc_hd__buf_2_176/X sky130_fd_sc_hd__buf_2_176/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_69 sky130_fd_sc_hd__o22ai_1_88/B1 sky130_fd_sc_hd__nand2_2_3/Y
+ sky130_fd_sc_hd__o22ai_1_69/Y sky130_fd_sc_hd__xnor2_1_49/Y sky130_fd_sc_hd__o22ai_1_83/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_187 VDD VSS sky130_fd_sc_hd__buf_2_187/X sky130_fd_sc_hd__buf_2_187/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_198 VDD VSS sky130_fd_sc_hd__buf_2_198/X sky130_fd_sc_hd__buf_2_198/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1150 VDD VSS sky130_fd_sc_hd__mux2_2_143/A0 sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__o22ai_1_287/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1161 VDD VSS sky130_fd_sc_hd__fa_2_863/B sky130_fd_sc_hd__dfxtp_1_1179/CLK
+ sky130_fd_sc_hd__a21oi_1_376/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1172 VDD VSS sky130_fd_sc_hd__fa_2_852/B sky130_fd_sc_hd__dfxtp_1_1184/CLK
+ sky130_fd_sc_hd__o21a_1_50/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1183 VDD VSS sky130_fd_sc_hd__fa_2_936/A sky130_fd_sc_hd__clkinv_4_24/Y
+ sky130_fd_sc_hd__a21oi_1_364/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1194 VDD VSS sky130_fd_sc_hd__fa_2_1243/A sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__and2_0_332/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_4_16 VDD VSS sky130_fd_sc_hd__buf_4_16/X sky130_fd_sc_hd__buf_8_15/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_27 VDD VSS sky130_fd_sc_hd__buf_4_27/X sky130_fd_sc_hd__buf_8_24/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_38 VDD VSS sky130_fd_sc_hd__buf_4_38/X sky130_fd_sc_hd__buf_4_38/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_49 VDD VSS sky130_fd_sc_hd__buf_4_49/X sky130_fd_sc_hd__buf_8_67/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__clkbuf_1_10 VSS VDD sky130_fd_sc_hd__buf_4_8/A sky130_fd_sc_hd__clkbuf_4_2/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_21 VSS VDD sky130_fd_sc_hd__clkbuf_1_21/X sky130_fd_sc_hd__clkbuf_1_21/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_32 VSS VDD sky130_fd_sc_hd__clkbuf_1_32/X sky130_fd_sc_hd__clkbuf_1_32/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_109 sky130_fd_sc_hd__buf_12_64/X sky130_fd_sc_hd__buf_12_109/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkbuf_1_43 VSS VDD sky130_fd_sc_hd__clkbuf_1_43/X sky130_fd_sc_hd__clkbuf_1_43/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_54 VSS VDD sky130_fd_sc_hd__clkbuf_1_54/X sky130_fd_sc_hd__clkbuf_1_54/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_660 sky130_fd_sc_hd__fa_2_582/A sky130_fd_sc_hd__maj3_1_108/A
+ sky130_fd_sc_hd__fa_2_660/A sky130_fd_sc_hd__fa_2_660/B sky130_fd_sc_hd__fa_2_662/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_65 VSS VDD sky130_fd_sc_hd__clkbuf_1_65/X sky130_fd_sc_hd__clkbuf_1_65/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_671 sky130_fd_sc_hd__fa_2_670/B sky130_fd_sc_hd__fa_2_671/SUM
+ sky130_fd_sc_hd__fa_2_671/A sky130_fd_sc_hd__fa_2_671/B sky130_fd_sc_hd__fa_2_671/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_76 VSS VDD sky130_fd_sc_hd__nand4_1_11/A sky130_fd_sc_hd__a22oi_1_67/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_682 sky130_fd_sc_hd__fa_2_681/A sky130_fd_sc_hd__fa_2_676/A
+ sky130_fd_sc_hd__fa_2_700/B sky130_fd_sc_hd__fa_2_695/A sky130_fd_sc_hd__ha_2_129/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_87 VSS VDD sky130_fd_sc_hd__nand4_1_0/A sky130_fd_sc_hd__a22oi_2_4/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_693 sky130_fd_sc_hd__fa_2_691/A sky130_fd_sc_hd__fa_2_687/A
+ sky130_fd_sc_hd__fa_2_699/A sky130_fd_sc_hd__ha_2_133/B sky130_fd_sc_hd__fa_2_659/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_98 VSS VDD sky130_fd_sc_hd__buf_8_40/A sky130_fd_sc_hd__clkbuf_1_98/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkinv_1_309 sky130_fd_sc_hd__fa_2_286/B sky130_fd_sc_hd__ha_2_116/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_309/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_206 sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__o21ai_1_232/Y
+ sky130_fd_sc_hd__a21oi_1_206/Y sky130_fd_sc_hd__fa_2_1061/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_217 sky130_fd_sc_hd__clkinv_1_728/Y sky130_fd_sc_hd__o21ai_1_250/Y
+ sky130_fd_sc_hd__a21oi_1_217/Y sky130_fd_sc_hd__nand2_1_333/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__or2_0_12 sky130_fd_sc_hd__or2_0_12/A sky130_fd_sc_hd__or2_0_12/X
+ sky130_fd_sc_hd__or2_0_12/B VSS VDD VSS VDD sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__a21oi_1_228 sky130_fd_sc_hd__clkinv_1_747/Y sky130_fd_sc_hd__o22ai_1_203/Y
+ sky130_fd_sc_hd__a21oi_1_228/Y sky130_fd_sc_hd__nand2_1_333/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_2_13 sky130_fd_sc_hd__nor3_2_7/Y sky130_fd_sc_hd__a22oi_2_13/A2
+ sky130_fd_sc_hd__nor3_2_8/Y sky130_fd_sc_hd__a22oi_2_13/B2 sky130_fd_sc_hd__nand4_1_48/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__a21oi_1_239 sky130_fd_sc_hd__a21o_2_5/A2 sky130_fd_sc_hd__o21ai_1_274/Y
+ sky130_fd_sc_hd__a21oi_1_239/Y sky130_fd_sc_hd__fa_2_1075/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_2_24 sky130_fd_sc_hd__a22oi_2_25/A1 sky130_fd_sc_hd__a22oi_2_24/A2
+ sky130_fd_sc_hd__a22oi_2_25/B1 sky130_fd_sc_hd__a22oi_2_24/B2 sky130_fd_sc_hd__nand4_1_57/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__nand2_1_200 sky130_fd_sc_hd__fa_2_702/B sky130_fd_sc_hd__fa_2_832/A
+ sky130_fd_sc_hd__fa_2_834/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_211 sky130_fd_sc_hd__nor4_1_5/D sky130_fd_sc_hd__nor3_1_31/B
+ sky130_fd_sc_hd__nand3_1_45/C VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_810 sky130_fd_sc_hd__nor2_1_148/B sky130_fd_sc_hd__fa_2_1126/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_810/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_222 sky130_fd_sc_hd__nand3_1_48/B sky130_fd_sc_hd__o221ai_1_1/A2
+ sky130_fd_sc_hd__fa_2_959/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_821 sky130_fd_sc_hd__nor2_1_173/A sky130_fd_sc_hd__xor2_1_164/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_821/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_233 sky130_fd_sc_hd__xnor2_1_48/B sky130_fd_sc_hd__o21ai_1_77/B1
+ sky130_fd_sc_hd__o21ai_1_84/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_180 sky130_fd_sc_hd__o22ai_1_206/B1 sky130_fd_sc_hd__o22ai_1_193/A1
+ sky130_fd_sc_hd__o22ai_1_180/Y sky130_fd_sc_hd__o22ai_1_194/B1 sky130_fd_sc_hd__o22ai_1_206/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_832 sky130_fd_sc_hd__o21ai_1_306/A1 sky130_fd_sc_hd__o21ai_1_308/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_832/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_244 sky130_fd_sc_hd__nand2_1_244/Y sky130_fd_sc_hd__nor2_1_55/B
+ sky130_fd_sc_hd__nor2_1_55/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_191 sky130_fd_sc_hd__o22ai_1_204/B1 sky130_fd_sc_hd__nor2_1_116/B
+ sky130_fd_sc_hd__nor2_1_134/A sky130_fd_sc_hd__o22ai_1_191/A1 sky130_fd_sc_hd__o22ai_1_206/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_843 sky130_fd_sc_hd__nor2_1_150/B sky130_fd_sc_hd__fa_2_1155/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_843/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_255 sky130_fd_sc_hd__o21a_1_5/B1 sky130_fd_sc_hd__fa_2_982/A
+ sky130_fd_sc_hd__o21a_1_5/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_854 sky130_fd_sc_hd__nor2_1_155/B sky130_fd_sc_hd__fa_2_1146/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_854/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_266 sky130_fd_sc_hd__o211ai_1_6/B1 sky130_fd_sc_hd__nor2_2_7/Y
+ sky130_fd_sc_hd__fa_2_989/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_865 sky130_fd_sc_hd__o22ai_1_322/A2 sky130_fd_sc_hd__nor3_1_39/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_865/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_277 sky130_fd_sc_hd__nand2_1_277/Y sky130_fd_sc_hd__nand2_1_282/B
+ sky130_fd_sc_hd__nor2_4_9/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_876 sky130_fd_sc_hd__nor2_1_198/A sky130_fd_sc_hd__nor2_1_199/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_876/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand4_1_50 sky130_fd_sc_hd__nand4_1_50/C sky130_fd_sc_hd__nand4_1_50/B
+ sky130_fd_sc_hd__buf_2_271/A sky130_fd_sc_hd__nand4_1_50/D sky130_fd_sc_hd__nand4_1_50/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand2_1_288 sky130_fd_sc_hd__xnor2_1_69/B sky130_fd_sc_hd__nand2_1_288/B
+ sky130_fd_sc_hd__nand2_1_299/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_887 sky130_fd_sc_hd__o31ai_1_8/A1 sky130_fd_sc_hd__o31ai_1_7/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_887/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand4_1_61 sky130_fd_sc_hd__nand4_1_61/C sky130_fd_sc_hd__nand4_1_61/B
+ sky130_fd_sc_hd__nand4_1_61/Y sky130_fd_sc_hd__nand4_1_61/D sky130_fd_sc_hd__nand4_1_61/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand2_1_299 sky130_fd_sc_hd__nand2_1_299/Y sky130_fd_sc_hd__nor2_1_107/B
+ sky130_fd_sc_hd__fa_2_1110/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_898 sky130_fd_sc_hd__nand2_1_422/B sky130_fd_sc_hd__fa_2_285/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_898/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand4_1_72 sky130_fd_sc_hd__nand4_1_72/C sky130_fd_sc_hd__nand4_1_72/B
+ sky130_fd_sc_hd__nand2_1_7/B sky130_fd_sc_hd__nand4_1_72/D sky130_fd_sc_hd__nand4_1_72/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_83 sky130_fd_sc_hd__xnor2_1_16/Y sky130_fd_sc_hd__xnor2_1_17/Y
+ sky130_fd_sc_hd__nor4_1_3/D sky130_fd_sc_hd__xnor2_1_15/Y sky130_fd_sc_hd__nand4_1_83/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__conb_1_10 sky130_fd_sc_hd__conb_1_10/LO sky130_fd_sc_hd__conb_1_10/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_21 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__conb_1_21/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__mux2_2_5 VSS VDD sky130_fd_sc_hd__mux2_2_5/A1 sky130_fd_sc_hd__mux2_2_5/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_5/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1150 sky130_fd_sc_hd__fa_2_1151/CIN sky130_fd_sc_hd__mux2_2_93/A1
+ sky130_fd_sc_hd__fa_2_1150/A sky130_fd_sc_hd__fa_2_1150/B sky130_fd_sc_hd__fa_2_1150/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1161 sky130_fd_sc_hd__fa_2_1162/CIN sky130_fd_sc_hd__mux2_2_120/A1
+ sky130_fd_sc_hd__fa_2_1161/A sky130_fd_sc_hd__fa_2_1172/B sky130_fd_sc_hd__fa_2_1161/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1172 sky130_fd_sc_hd__xor2_1_183/B sky130_fd_sc_hd__nand2_1_365/A
+ sky130_fd_sc_hd__fa_2_1172/A sky130_fd_sc_hd__fa_2_1172/B sky130_fd_sc_hd__fa_2_1172/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1183 sky130_fd_sc_hd__fa_2_1184/CIN sky130_fd_sc_hd__mux2_2_142/A1
+ sky130_fd_sc_hd__fa_2_1183/A sky130_fd_sc_hd__fa_2_1183/B sky130_fd_sc_hd__fa_2_1183/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1194 sky130_fd_sc_hd__fa_2_1195/CIN sky130_fd_sc_hd__mux2_2_161/A1
+ sky130_fd_sc_hd__fa_2_1194/A sky130_fd_sc_hd__fa_2_1194/B sky130_fd_sc_hd__fa_2_1194/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a211o_1_19 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_206/A sky130_fd_sc_hd__nor2b_1_112/Y
+ sky130_fd_sc_hd__o22ai_1_294/Y sky130_fd_sc_hd__o21ai_1_370/Y sky130_fd_sc_hd__o22ai_1_293/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o2bb2ai_1_1 sky130_fd_sc_hd__o2bb2ai_1_1/Y sky130_fd_sc_hd__nor2_1_18/Y
+ sky130_fd_sc_hd__ha_2_153/SUM sky130_fd_sc_hd__o21ai_1_31/A1 sky130_fd_sc_hd__nor2_1_12/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_490 sky130_fd_sc_hd__fa_2_494/B sky130_fd_sc_hd__fa_2_490/SUM
+ sky130_fd_sc_hd__fa_2_490/A sky130_fd_sc_hd__fa_2_490/B sky130_fd_sc_hd__fa_2_490/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_1_106 sky130_fd_sc_hd__buf_12_133/A sky130_fd_sc_hd__clkinv_1_106/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_106/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_117 sky130_fd_sc_hd__bufinv_8_3/A sky130_fd_sc_hd__buf_8_83/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_117/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_128 sky130_fd_sc_hd__nand3_4_1/C sky130_fd_sc_hd__nand3_4_0/B
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_139 sky130_fd_sc_hd__buf_12_268/A sky130_fd_sc_hd__clkinv_1_139/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_139/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_19 sky130_fd_sc_hd__nor2_4_4/Y sky130_fd_sc_hd__ha_2_73/A
+ sky130_fd_sc_hd__a22o_1_19/X sky130_fd_sc_hd__a22o_1_19/B2 sky130_fd_sc_hd__a22o_2_6/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__o21ai_1_6 VSS VDD sky130_fd_sc_hd__nor2_1_9/Y sky130_fd_sc_hd__or4_1_1/A
+ sky130_fd_sc_hd__o21ai_1_6/B1 sky130_fd_sc_hd__o21ai_1_6/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__bufbuf_16_5 sky130_fd_sc_hd__buf_2_240/X sky130_fd_sc_hd__buf_12_416/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__nor2_1_200 sky130_fd_sc_hd__nor2_1_200/B sky130_fd_sc_hd__nor2_1_200/Y
+ sky130_fd_sc_hd__nor2_4_16/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_211 sky130_fd_sc_hd__nor2_1_211/B sky130_fd_sc_hd__nor2_1_211/Y
+ sky130_fd_sc_hd__nor2_1_211/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_222 sky130_fd_sc_hd__o21a_1_42/A1 sky130_fd_sc_hd__nor2_1_222/Y
+ sky130_fd_sc_hd__nor2_1_222/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_233 sky130_fd_sc_hd__nor2_1_233/B sky130_fd_sc_hd__o21a_1_48/A1
+ sky130_fd_sc_hd__nor2_1_233/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_244 sky130_fd_sc_hd__nor2_1_248/A sky130_fd_sc_hd__nor2_1_244/Y
+ sky130_fd_sc_hd__xnor2_1_99/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_255 sky130_fd_sc_hd__nor2_1_255/B sky130_fd_sc_hd__nor2_1_255/Y
+ sky130_fd_sc_hd__nor2_1_255/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_2_9 sky130_fd_sc_hd__clkinv_2_9/Y sky130_fd_sc_hd__clkinv_2_9/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_9/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__nor2_1_266 sky130_fd_sc_hd__o21a_1_55/A1 sky130_fd_sc_hd__nor2_1_266/Y
+ sky130_fd_sc_hd__nor2_1_266/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_277 sky130_fd_sc_hd__nor2_1_277/B sky130_fd_sc_hd__o21a_1_62/A1
+ sky130_fd_sc_hd__o21a_1_63/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_288 sky130_fd_sc_hd__nor2_1_288/B sky130_fd_sc_hd__nor2_1_288/Y
+ sky130_fd_sc_hd__nor2_1_290/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_299 sky130_fd_sc_hd__nor2_1_299/B sky130_fd_sc_hd__nor2_1_299/Y
+ sky130_fd_sc_hd__nor2_1_299/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_440 sky130_fd_sc_hd__buf_4_113/X sky130_fd_sc_hd__buf_12_440/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_451 sky130_fd_sc_hd__buf_12_451/A sky130_fd_sc_hd__buf_12_480/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_310 sky130_fd_sc_hd__clkbuf_1_378/X sky130_fd_sc_hd__clkbuf_1_379/X
+ sky130_fd_sc_hd__buf_2_220/X sky130_fd_sc_hd__buf_2_189/X sky130_fd_sc_hd__nand4_1_77/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_462 sky130_fd_sc_hd__buf_6_73/X sky130_fd_sc_hd__buf_12_503/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_321 sky130_fd_sc_hd__inv_4_1/Y sky130_fd_sc_hd__nor2_1_16/Y
+ sky130_fd_sc_hd__o21ai_1_4/Y sky130_fd_sc_hd__dfxtp_1_0/Q sky130_fd_sc_hd__o211ai_1_1/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_473 sky130_fd_sc_hd__buf_12_473/A sky130_fd_sc_hd__buf_12_473/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_332 sky130_fd_sc_hd__a21oi_1_94/A1 sky130_fd_sc_hd__a211o_1_6/A2
+ sky130_fd_sc_hd__nand2_1_264/A sky130_fd_sc_hd__a211o_1_3/A1 sky130_fd_sc_hd__o211ai_1_9/C1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_484 sky130_fd_sc_hd__buf_12_484/A sky130_fd_sc_hd__buf_12_484/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_343 sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_2_7/Y
+ sky130_fd_sc_hd__fa_2_1002/A sky130_fd_sc_hd__fa_2_1003/A sky130_fd_sc_hd__a22oi_1_343/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_495 sky130_fd_sc_hd__buf_12_495/A sky130_fd_sc_hd__buf_12_495/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_354 sky130_fd_sc_hd__fa_2_1062/A sky130_fd_sc_hd__fa_2_1064/A
+ sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__nor2_2_12/Y sky130_fd_sc_hd__a22oi_1_354/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_365 sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__nor2_4_13/Y
+ sky130_fd_sc_hd__fa_2_1082/A sky130_fd_sc_hd__fa_2_1083/A sky130_fd_sc_hd__a22oi_1_365/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_376 sky130_fd_sc_hd__clkinv_1_779/Y sky130_fd_sc_hd__nor3_1_38/B
+ sky130_fd_sc_hd__fa_2_1138/A sky130_fd_sc_hd__fa_2_1139/A sky130_fd_sc_hd__a22oi_1_376/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_387 sky130_fd_sc_hd__clkinv_1_946/Y sky130_fd_sc_hd__nor3_1_40/B
+ sky130_fd_sc_hd__fa_2_1248/A sky130_fd_sc_hd__fa_2_1249/A sky130_fd_sc_hd__a22oi_1_387/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_398 sky130_fd_sc_hd__nor3_1_41/B sky130_fd_sc_hd__fa_2_1292/A
+ sky130_fd_sc_hd__xor2_1_299/A sky130_fd_sc_hd__a22oi_1_400/B1 sky130_fd_sc_hd__a22oi_1_398/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_640 sky130_fd_sc_hd__o22ai_1_158/B2 sky130_fd_sc_hd__ha_2_191/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_640/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_651 sky130_fd_sc_hd__nand2_1_291/B sky130_fd_sc_hd__nor2_1_110/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_651/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_662 sky130_fd_sc_hd__o21ai_1_198/A1 sky130_fd_sc_hd__nand2_1_300/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_662/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_673 sky130_fd_sc_hd__clkinv_1_673/Y sky130_fd_sc_hd__nor2_1_99/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_673/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_684 sky130_fd_sc_hd__nor2_1_110/B sky130_fd_sc_hd__fa_2_1116/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_684/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_695 sky130_fd_sc_hd__clkinv_1_695/Y sky130_fd_sc_hd__a21oi_1_197/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_695/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand3_1_2 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__nand3_1_2/A
+ sky130_fd_sc_hd__nand3_1_2/C sky130_fd_sc_hd__nand3_1_2/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__xnor2_1_40 VSS VDD sky130_fd_sc_hd__xnor2_1_40/B sky130_fd_sc_hd__xnor2_1_40/Y
+ sky130_fd_sc_hd__xnor2_1_40/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_51 VSS VDD sky130_fd_sc_hd__xnor2_1_52/B sky130_fd_sc_hd__xnor2_1_51/Y
+ sky130_fd_sc_hd__xnor2_1_51/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_62 VSS VDD sky130_fd_sc_hd__xnor2_1_62/B sky130_fd_sc_hd__xnor2_1_62/Y
+ sky130_fd_sc_hd__nor2_1_92/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_73 VSS VDD sky130_fd_sc_hd__xnor2_1_73/B sky130_fd_sc_hd__xnor2_1_73/Y
+ sky130_fd_sc_hd__xnor2_1_73/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_84 VSS VDD sky130_fd_sc_hd__xnor2_1_85/B sky130_fd_sc_hd__xnor2_1_84/Y
+ sky130_fd_sc_hd__xnor2_1_84/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_95 VSS VDD sky130_fd_sc_hd__xnor2_1_95/B sky130_fd_sc_hd__xnor2_1_95/Y
+ sky130_fd_sc_hd__fa_2_1208/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__dfxtp_1_809 VDD VSS sky130_fd_sc_hd__fa_2_1061/A sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__mux2_2_55/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_407 VSS VDD sky130_fd_sc_hd__clkbuf_1_407/X sky130_fd_sc_hd__clkbuf_1_407/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_418 VSS VDD sky130_fd_sc_hd__clkbuf_1_418/X sky130_fd_sc_hd__buf_2_250/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_429 VSS VDD sky130_fd_sc_hd__clkbuf_1_429/X sky130_fd_sc_hd__clkbuf_1_429/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o32ai_1_1 sky130_fd_sc_hd__o32ai_1_1/A2 sky130_fd_sc_hd__o32ai_1_1/Y
+ sky130_fd_sc_hd__fa_2_1142/A sky130_fd_sc_hd__o32ai_1_1/A3 sky130_fd_sc_hd__o32ai_1_1/B2
+ sky130_fd_sc_hd__fa_2_1141/A VDD VSS VSS VDD sky130_fd_sc_hd__o32ai_1
Xsky130_fd_sc_hd__diode_2_170 sky130_fd_sc_hd__clkbuf_4_181/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_181 sky130_fd_sc_hd__buf_2_246/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_192 sky130_fd_sc_hd__inv_2_136/Y VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkinv_2_14 sky130_fd_sc_hd__clkinv_2_14/Y sky130_fd_sc_hd__clkinv_2_14/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_14/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkbuf_4_201 sky130_fd_sc_hd__nand4_1_65/D sky130_fd_sc_hd__a22oi_1_261/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_212 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__nor2_1_90/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_2_25 sky130_fd_sc_hd__nand4_1_74/D sky130_fd_sc_hd__clkinv_2_25/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_25/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_36 sky130_fd_sc_hd__clkinv_4_24/A sky130_fd_sc_hd__clkinv_2_36/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_36/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkbuf_4_223 sky130_fd_sc_hd__a22oi_1_9/A2 sig_amplitude[3] VSS
+ VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_2_47 sky130_fd_sc_hd__clkinv_2_48/A sky130_fd_sc_hd__clkinv_2_47/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_47/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__buf_12_270 sky130_fd_sc_hd__inv_2_88/Y sky130_fd_sc_hd__buf_12_270/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_281 sky130_fd_sc_hd__inv_2_103/Y sky130_fd_sc_hd__buf_12_355/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_140 sky130_fd_sc_hd__a22oi_1_97/B1 sky130_fd_sc_hd__a22oi_1_97/A1
+ sky130_fd_sc_hd__clkbuf_1_155/X sky130_fd_sc_hd__clkbuf_4_75/X sky130_fd_sc_hd__nand4_1_30/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_292 sky130_fd_sc_hd__buf_8_170/X sky130_fd_sc_hd__buf_12_292/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_151 sky130_fd_sc_hd__clkbuf_1_265/X sky130_fd_sc_hd__clkbuf_1_266/X
+ sky130_fd_sc_hd__clkbuf_1_280/X sky130_fd_sc_hd__a22oi_1_151/A2 sky130_fd_sc_hd__a22oi_1_151/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_162 sky130_fd_sc_hd__clkbuf_1_264/X sky130_fd_sc_hd__nor2_2_3/Y
+ sky130_fd_sc_hd__a22oi_1_162/B2 sky130_fd_sc_hd__clkbuf_4_134/X sky130_fd_sc_hd__nand4_1_35/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_173 sky130_fd_sc_hd__clkbuf_4_111/X sky130_fd_sc_hd__clkbuf_4_112/X
+ sky130_fd_sc_hd__a22oi_1_173/B2 sky130_fd_sc_hd__clkbuf_1_291/X sky130_fd_sc_hd__a22oi_1_173/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_184 sky130_fd_sc_hd__clkbuf_1_351/X sky130_fd_sc_hd__clkbuf_1_353/X
+ sky130_fd_sc_hd__clkbuf_4_116/X sky130_fd_sc_hd__a22oi_1_184/A2 sky130_fd_sc_hd__nand4_1_41/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_195 sky130_fd_sc_hd__clkbuf_1_265/X sky130_fd_sc_hd__clkbuf_1_266/X
+ sky130_fd_sc_hd__clkbuf_1_270/X sky130_fd_sc_hd__a22oi_1_195/A2 sky130_fd_sc_hd__a22oi_1_195/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_470 sky130_fd_sc_hd__o21ai_1_53/A2 sky130_fd_sc_hd__nor2_2_6/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_470/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_481 sky130_fd_sc_hd__o22ai_1_86/B2 sky130_fd_sc_hd__ha_2_173/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_481/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_492 sky130_fd_sc_hd__o21ai_1_77/B1 sky130_fd_sc_hd__nor2_1_59/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_492/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_406 VSS VDD sky130_fd_sc_hd__nor3_1_40/A sky130_fd_sc_hd__nor2_1_258/A
+ sky130_fd_sc_hd__nand2_1_484/Y sky130_fd_sc_hd__o21ai_1_406/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_417 VSS VDD sky130_fd_sc_hd__a21oi_1_410/Y sky130_fd_sc_hd__nor2_1_267/A
+ sky130_fd_sc_hd__nand2_1_486/Y sky130_fd_sc_hd__xor2_1_234/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_428 VSS VDD sky130_fd_sc_hd__o21a_1_55/X sky130_fd_sc_hd__nor2_1_265/A
+ sky130_fd_sc_hd__a21oi_1_409/Y sky130_fd_sc_hd__xor2_1_246/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_439 VSS VDD sky130_fd_sc_hd__nand2_1_523/B sky130_fd_sc_hd__nor2_1_293/Y
+ sky130_fd_sc_hd__o31ai_1_12/A2 sky130_fd_sc_hd__o21ai_1_439/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_4_15 sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__nor2_4_15/A
+ sky130_fd_sc_hd__nor2_4_15/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__xor2_1_200 sky130_fd_sc_hd__fa_2_1173/A sky130_fd_sc_hd__fa_2_1179/B
+ sky130_fd_sc_hd__xor2_1_200/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_211 sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__fa_2_1207/B
+ sky130_fd_sc_hd__xor2_1_211/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_222 sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__fa_2_1196/B
+ sky130_fd_sc_hd__xor2_1_222/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_233 sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__xor2_1_233/X
+ sky130_fd_sc_hd__xor2_1_253/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_244 sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1231/B
+ sky130_fd_sc_hd__xor2_1_244/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_255 sky130_fd_sc_hd__xor2_1_267/B sky130_fd_sc_hd__fa_2_1259/B
+ sky130_fd_sc_hd__xor2_1_255/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_606 VDD VSS sky130_fd_sc_hd__and2_0_226/A sky130_fd_sc_hd__dfxtp_1_606/CLK
+ sky130_fd_sc_hd__fa_2_1026/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_266 sky130_fd_sc_hd__xor2_1_267/B sky130_fd_sc_hd__fa_2_1248/B
+ sky130_fd_sc_hd__xor2_1_266/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_617 VDD VSS sky130_fd_sc_hd__ha_2_143/A sky130_fd_sc_hd__dfxtp_1_627/CLK
+ sky130_fd_sc_hd__a21oi_1_77/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_277 sky130_fd_sc_hd__xor2_1_278/X sky130_fd_sc_hd__xor2_1_277/X
+ sky130_fd_sc_hd__xor2_1_299/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_288 sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1283/B
+ sky130_fd_sc_hd__xor2_1_288/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_628 VDD VSS sky130_fd_sc_hd__or2_0_6/A sky130_fd_sc_hd__clkinv_4_25/Y
+ sky130_fd_sc_hd__nor2b_1_91/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_639 VDD VSS sky130_fd_sc_hd__fa_2_1003/A sky130_fd_sc_hd__clkinv_8_44/Y
+ sky130_fd_sc_hd__mux2_2_26/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_299 sky130_fd_sc_hd__nor2_4_20/Y sky130_fd_sc_hd__xor2_1_299/X
+ sky130_fd_sc_hd__xor2_1_299/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_204 VSS VDD sky130_fd_sc_hd__buf_8_103/A sky130_fd_sc_hd__buf_6_20/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_215 VSS VDD sky130_fd_sc_hd__buf_12_131/A sky130_fd_sc_hd__buf_2_47/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_226 VSS VDD sky130_fd_sc_hd__buf_8_111/A sky130_fd_sc_hd__buf_6_21/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_237 VSS VDD sky130_fd_sc_hd__clkinv_1_112/A sky130_fd_sc_hd__buf_8_65/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_248 VSS VDD sky130_fd_sc_hd__clkbuf_1_248/X sky130_fd_sc_hd__clkbuf_1_249/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_259 VSS VDD sky130_fd_sc_hd__clkbuf_1_259/X sky130_fd_sc_hd__clkbuf_1_260/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_2_60 VDD VSS sky130_fd_sc_hd__buf_2_60/X sky130_fd_sc_hd__buf_2_60/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_71 VDD VSS sky130_fd_sc_hd__buf_2_71/X sky130_fd_sc_hd__buf_2_71/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_82 VDD VSS sky130_fd_sc_hd__buf_2_82/X sky130_fd_sc_hd__buf_2_82/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_93 VDD VSS sky130_fd_sc_hd__buf_2_93/X sky130_fd_sc_hd__buf_2_93/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_4_9 VDD VSS sky130_fd_sc_hd__buf_4_9/X sky130_fd_sc_hd__buf_4_9/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__diode_2_0 sky130_fd_sc_hd__clkbuf_4_23/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__and2_0_202 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_202/X sky130_fd_sc_hd__and2_0_235/B
+ sky130_fd_sc_hd__and2_0_202/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_213 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_213/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_213/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_224 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_224/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_224/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_235 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_235/X sky130_fd_sc_hd__and2_0_235/B
+ sky130_fd_sc_hd__and2_0_235/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_246 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_246/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__and2_0_246/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_257 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_257/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__fa_2_958/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_268 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_268/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__fa_2_967/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_279 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_279/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__fa_2_994/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__sdlclkp_2_7 sky130_fd_sc_hd__conb_1_16/LO sky130_fd_sc_hd__clkinv_8_104/A
+ sky130_fd_sc_hd__dfxtp_1_282/CLK sky130_fd_sc_hd__a21oi_1_15/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__a22o_2_1 sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__ha_2_66/A
+ sky130_fd_sc_hd__a22o_2_1/X sky130_fd_sc_hd__dfxtp_1_5/Q sky130_fd_sc_hd__a22o_2_3/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_2
Xsky130_fd_sc_hd__o31ai_1_0 sky130_fd_sc_hd__o31ai_1_0/Y sky130_fd_sc_hd__xor2_1_9/X
+ sky130_fd_sc_hd__ha_2_167/B sky130_fd_sc_hd__o31ai_1_0/A3 sky130_fd_sc_hd__o31ai_1_0/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__o31ai_1
Xsky130_fd_sc_hd__clkbuf_4_10 sky130_fd_sc_hd__clkbuf_4_10/X sky130_fd_sc_hd__clkbuf_4_10/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_203 VSS VDD sky130_fd_sc_hd__xnor2_1_72/A sky130_fd_sc_hd__nor2_1_108/Y
+ sky130_fd_sc_hd__nand2_1_298/Y sky130_fd_sc_hd__xnor2_1_74/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_21 sky130_fd_sc_hd__clkbuf_4_21/X sky130_fd_sc_hd__clkbuf_4_21/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_214 VSS VDD sky130_fd_sc_hd__a21oi_1_197/Y sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__nand2_1_317/Y sky130_fd_sc_hd__xor2_1_118/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_32 sky130_fd_sc_hd__clkbuf_4_32/X sky130_fd_sc_hd__clkbuf_4_32/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_225 VSS VDD sky130_fd_sc_hd__o21ai_1_225/A2 sky130_fd_sc_hd__o22ai_1_206/B1
+ sky130_fd_sc_hd__a22oi_1_349/Y sky130_fd_sc_hd__o21ai_1_225/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_43 sky130_fd_sc_hd__nand4_1_14/D sky130_fd_sc_hd__a22oi_1_76/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_236 VSS VDD sky130_fd_sc_hd__nor2_1_117/B sky130_fd_sc_hd__o21a_1_16/A2
+ sky130_fd_sc_hd__a21oi_1_210/Y sky130_fd_sc_hd__o21ai_1_236/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_54 sky130_fd_sc_hd__nand4_1_3/D sky130_fd_sc_hd__a22oi_1_39/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_247 VSS VDD sky130_fd_sc_hd__nor2_1_127/A sky130_fd_sc_hd__a211oi_1_8/Y
+ sky130_fd_sc_hd__a21oi_1_216/Y sky130_fd_sc_hd__xor2_1_98/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_65 sky130_fd_sc_hd__buf_2_36/A sky130_fd_sc_hd__dfxtp_1_253/Q
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_258 VSS VDD sky130_fd_sc_hd__a21oi_1_235/Y sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__a21oi_1_223/Y sky130_fd_sc_hd__xor2_1_102/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_76 sky130_fd_sc_hd__clkbuf_4_76/X sky130_fd_sc_hd__clkbuf_4_76/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_269 VSS VDD sky130_fd_sc_hd__o22ai_1_206/B2 sky130_fd_sc_hd__o22ai_1_206/A1
+ sky130_fd_sc_hd__a22oi_1_365/Y sky130_fd_sc_hd__o21ai_1_269/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_87 sky130_fd_sc_hd__clkbuf_4_87/X sky130_fd_sc_hd__clkbuf_4_87/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_98 sky130_fd_sc_hd__buf_12_150/A sky130_fd_sc_hd__buf_6_20/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__nor2_4_0 sky130_fd_sc_hd__nor2_4_0/Y sky130_fd_sc_hd__nor2_4_4/A
+ sky130_fd_sc_hd__inv_2_0/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__buf_8_160 sky130_fd_sc_hd__buf_8_160/A sky130_fd_sc_hd__buf_8_160/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_171 sky130_fd_sc_hd__buf_8_171/A sky130_fd_sc_hd__buf_6_48/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_182 sky130_fd_sc_hd__buf_8_204/A sky130_fd_sc_hd__buf_8_221/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_193 sky130_fd_sc_hd__inv_2_122/Y sky130_fd_sc_hd__buf_8_193/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_403 VDD VSS sky130_fd_sc_hd__fa_2_1039/A sky130_fd_sc_hd__dfxtp_1_424/CLK
+ sky130_fd_sc_hd__and2_0_134/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_414 VDD VSS sky130_fd_sc_hd__fa_2_1034/B sky130_fd_sc_hd__dfxtp_1_419/CLK
+ sky130_fd_sc_hd__and2_0_159/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_425 VDD VSS sky130_fd_sc_hd__nor2_2_6/A sky130_fd_sc_hd__dfxtp_1_425/CLK
+ sky130_fd_sc_hd__and2_0_102/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_436 VDD VSS sky130_fd_sc_hd__dfxtp_1_436/Q sky130_fd_sc_hd__dfxtp_1_452/CLK
+ sky130_fd_sc_hd__nand2_1_92/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_447 VDD VSS sky130_fd_sc_hd__dfxtp_1_993/D sky130_fd_sc_hd__dfxtp_1_448/CLK
+ sky130_fd_sc_hd__nand2_1_70/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_458 VDD VSS sky130_fd_sc_hd__dfxtp_1_458/Q sky130_fd_sc_hd__dfxtp_1_473/CLK
+ sky130_fd_sc_hd__and2_0_175/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_469 VDD VSS sky130_fd_sc_hd__clkbuf_1_5/A sky130_fd_sc_hd__dfxtp_1_473/CLK
+ sky130_fd_sc_hd__and2_0_126/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2b_1_17 sky130_fd_sc_hd__nand2b_1_17/Y sky130_fd_sc_hd__nor2_1_314/Y
+ sky130_fd_sc_hd__nor4_1_13/C VDD VSS VSS VDD sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__fa_2_308 sky130_fd_sc_hd__fa_2_304/A sky130_fd_sc_hd__fa_2_309/A
+ sky130_fd_sc_hd__fa_2_360/B sky130_fd_sc_hd__ha_2_108/B sky130_fd_sc_hd__fa_2_286/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_319 sky130_fd_sc_hd__fa_2_316/CIN sky130_fd_sc_hd__fa_2_320/CIN
+ sky130_fd_sc_hd__fa_2_424/B sky130_fd_sc_hd__fa_2_417/A sky130_fd_sc_hd__fa_2_401/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_8_13 sky130_fd_sc_hd__clkinv_8_13/Y sky130_fd_sc_hd__clkinv_8_13/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_13/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_24 sky130_fd_sc_hd__clkinv_8_25/A sky130_fd_sc_hd__clkinv_8_24/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_35 sky130_fd_sc_hd__clkinv_8_36/A sky130_fd_sc_hd__clkinv_8_35/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_35/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_46 sky130_fd_sc_hd__clkinv_8_46/Y sky130_fd_sc_hd__clkinv_8_74/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_57 sky130_fd_sc_hd__clkinv_8_58/A sky130_fd_sc_hd__clkinv_8_95/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_11 sky130_fd_sc_hd__buf_12_11/A sky130_fd_sc_hd__buf_12_90/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_8_68 sky130_fd_sc_hd__clkinv_8_68/Y sky130_fd_sc_hd__clkinv_8_68/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_22 sky130_fd_sc_hd__buf_8_19/X sky130_fd_sc_hd__buf_12_22/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_8_79 sky130_fd_sc_hd__clkinv_8_80/A sky130_fd_sc_hd__clkinv_8_79/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_33 sky130_fd_sc_hd__buf_8_49/X sky130_fd_sc_hd__buf_12_33/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_44 sky130_fd_sc_hd__buf_8_48/X sky130_fd_sc_hd__buf_12_44/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_55 sky130_fd_sc_hd__buf_8_34/X sky130_fd_sc_hd__buf_12_55/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_66 sky130_fd_sc_hd__buf_4_23/X sky130_fd_sc_hd__buf_12_66/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_77 sky130_fd_sc_hd__buf_6_14/X sky130_fd_sc_hd__buf_12_77/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_88 sky130_fd_sc_hd__buf_12_88/A sky130_fd_sc_hd__buf_12_88/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_99 sky130_fd_sc_hd__buf_12_99/A sky130_fd_sc_hd__buf_12_99/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_2_6 VDD VSS sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__buf_2_6/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1310 VDD VSS sky130_fd_sc_hd__fa_2_841/B sky130_fd_sc_hd__dfxtp_1_1326/CLK
+ sky130_fd_sc_hd__a21oi_1_431/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1321 VDD VSS sky130_fd_sc_hd__fa_2_905/A sky130_fd_sc_hd__dfxtp_1_1326/CLK
+ sky130_fd_sc_hd__a21oi_1_426/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1332 VDD VSS sky130_fd_sc_hd__xor2_1_24/B sky130_fd_sc_hd__dfxtp_1_1332/CLK
+ sky130_fd_sc_hd__xnor2_1_100/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1343 VDD VSS sky130_fd_sc_hd__fa_2_1302/A sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__mux2_2_239/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1354 VDD VSS sky130_fd_sc_hd__fa_2_1276/A sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__and2_0_337/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1365 VDD VSS sky130_fd_sc_hd__fa_2_1287/A sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__mux2_2_233/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1376 VDD VSS sky130_fd_sc_hd__fa_2_1315/A sky130_fd_sc_hd__clkinv_8_102/Y
+ sky130_fd_sc_hd__mux2_2_263/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1387 VDD VSS sky130_fd_sc_hd__nor2_8_2/B sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__mux2_2_236/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1398 VDD VSS sky130_fd_sc_hd__mux2_2_249/A0 sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__o22ai_1_391/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_970 VDD VSS sky130_fd_sc_hd__nor2_2_14/A sky130_fd_sc_hd__clkinv_8_46/Y
+ sky130_fd_sc_hd__nor2b_1_108/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_981 VDD VSS sky130_fd_sc_hd__mux2_2_89/A0 sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__o22ai_1_214/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_992 VDD VSS sky130_fd_sc_hd__mux2_2_119/A0 sky130_fd_sc_hd__clkinv_8_63/Y
+ sky130_fd_sc_hd__dfxtp_1_992/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_590 VSS VDD sky130_fd_sc_hd__nand3_1_2/B sky130_fd_sc_hd__a22oi_1_4/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_820 sky130_fd_sc_hd__fa_2_819/B sky130_fd_sc_hd__fa_2_815/B
+ sky130_fd_sc_hd__fa_2_833/A sky130_fd_sc_hd__fa_2_820/B sky130_fd_sc_hd__fa_2_811/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_180 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_180/A sky130_fd_sc_hd__ha_2_179/A
+ sky130_fd_sc_hd__ha_2_180/SUM sky130_fd_sc_hd__ha_2_180/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_831 sky130_fd_sc_hd__fa_2_830/B sky130_fd_sc_hd__fa_2_828/B
+ sky130_fd_sc_hd__fa_2_835/B sky130_fd_sc_hd__ha_2_145/B sky130_fd_sc_hd__fa_2_793/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_191 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_191/A sky130_fd_sc_hd__ha_2_190/A
+ sky130_fd_sc_hd__ha_2_191/SUM sky130_fd_sc_hd__ha_2_191/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_842 sky130_fd_sc_hd__fa_2_841/CIN sky130_fd_sc_hd__fa_2_842/SUM
+ sky130_fd_sc_hd__fa_2_842/A sky130_fd_sc_hd__fa_2_842/B sky130_fd_sc_hd__fa_2_842/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_853 sky130_fd_sc_hd__fa_2_852/CIN sky130_fd_sc_hd__fa_2_853/SUM
+ sky130_fd_sc_hd__fa_2_853/A sky130_fd_sc_hd__fa_2_853/B sky130_fd_sc_hd__fa_2_853/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_864 sky130_fd_sc_hd__xor2_1_15/B sky130_fd_sc_hd__fa_2_864/SUM
+ sky130_fd_sc_hd__fa_2_864/A sky130_fd_sc_hd__fa_2_864/B sky130_fd_sc_hd__fa_2_864/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_875 sky130_fd_sc_hd__fa_2_874/CIN sky130_fd_sc_hd__fa_2_875/SUM
+ sky130_fd_sc_hd__fa_2_875/A sky130_fd_sc_hd__fa_2_875/B sky130_fd_sc_hd__fa_2_875/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_886 sky130_fd_sc_hd__fa_2_885/CIN sky130_fd_sc_hd__nand2_1_46/B
+ sky130_fd_sc_hd__ha_2_157/A sky130_fd_sc_hd__fa_2_886/B sky130_fd_sc_hd__fa_2_886/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_897 sky130_fd_sc_hd__fa_2_896/CIN sky130_fd_sc_hd__fa_2_897/SUM
+ sky130_fd_sc_hd__fa_2_897/A sky130_fd_sc_hd__fa_2_897/B sky130_fd_sc_hd__fa_2_897/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_6 sky130_fd_sc_hd__inv_2_6/A sky130_fd_sc_hd__inv_2_7/A VDD
+ VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__nor3_2_8 sky130_fd_sc_hd__nor3_2_8/C sky130_fd_sc_hd__nor3_2_8/Y
+ sky130_fd_sc_hd__nor3_2_8/A sky130_fd_sc_hd__nor3_2_9/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_2
Xsky130_fd_sc_hd__nor2_1_16 sky130_fd_sc_hd__nor3_1_27/B sky130_fd_sc_hd__nor2_1_16/Y
+ sky130_fd_sc_hd__nor3_1_26/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_120 VSS VDD sky130_fd_sc_hd__mux2_2_120/A1 sky130_fd_sc_hd__mux2_2_120/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_120/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_27 sky130_fd_sc_hd__nor2_1_27/B sky130_fd_sc_hd__nor2_1_27/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_131 VSS VDD sky130_fd_sc_hd__mux2_2_131/A1 sky130_fd_sc_hd__mux2_2_131/A0
+ sky130_fd_sc_hd__mux2_2_135/S sky130_fd_sc_hd__mux2_2_131/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_38 sky130_fd_sc_hd__fa_2_964/A sky130_fd_sc_hd__nor2_1_38/Y
+ sky130_fd_sc_hd__nor2_1_39/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_142 VSS VDD sky130_fd_sc_hd__mux2_2_142/A1 sky130_fd_sc_hd__mux2_2_142/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_142/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_49 sky130_fd_sc_hd__nor2_1_49/B sky130_fd_sc_hd__nor2_1_49/Y
+ sky130_fd_sc_hd__nor2_1_49/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_153 VSS VDD sky130_fd_sc_hd__mux2_2_153/A1 sky130_fd_sc_hd__mux2_2_153/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_153/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_164 VSS VDD sky130_fd_sc_hd__mux2_2_164/A1 sky130_fd_sc_hd__mux2_2_164/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_164/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_175 VSS VDD sky130_fd_sc_hd__mux2_2_175/A1 sky130_fd_sc_hd__mux2_2_175/A0
+ sky130_fd_sc_hd__nor2_8_1/A sky130_fd_sc_hd__mux2_2_175/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_186 VSS VDD sky130_fd_sc_hd__mux2_2_186/A1 sky130_fd_sc_hd__mux2_2_186/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_186/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_197 VSS VDD sky130_fd_sc_hd__mux2_2_197/A1 sky130_fd_sc_hd__mux2_2_197/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_197/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__maj3_1_102 sky130_fd_sc_hd__maj3_1_103/X sky130_fd_sc_hd__maj3_1_102/X
+ sky130_fd_sc_hd__maj3_1_102/B sky130_fd_sc_hd__maj3_1_102/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_113 sky130_fd_sc_hd__maj3_1_114/X sky130_fd_sc_hd__maj3_1_113/X
+ sky130_fd_sc_hd__maj3_1_113/B sky130_fd_sc_hd__maj3_1_113/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__and2_0_60 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_60/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_60/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_124 sky130_fd_sc_hd__maj3_1_125/X sky130_fd_sc_hd__maj3_1_124/X
+ sky130_fd_sc_hd__maj3_1_124/B sky130_fd_sc_hd__maj3_1_124/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_340 sky130_fd_sc_hd__nand2_1_464/Y sky130_fd_sc_hd__nand2_1_463/Y
+ sky130_fd_sc_hd__o22ai_1_340/Y sky130_fd_sc_hd__o22ai_1_340/A1 sky130_fd_sc_hd__a21o_2_19/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_71 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_74/A sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__ha_2_75/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_404 sky130_fd_sc_hd__o21a_1_39/B1 sky130_fd_sc_hd__fa_2_1201/A
+ sky130_fd_sc_hd__o21a_1_39/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_135 sky130_fd_sc_hd__maj3_1_136/X sky130_fd_sc_hd__maj3_1_135/X
+ sky130_fd_sc_hd__maj3_1_135/B sky130_fd_sc_hd__maj3_1_135/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_351 sky130_fd_sc_hd__o32ai_1_7/B2 sky130_fd_sc_hd__nor2_1_267/A
+ sky130_fd_sc_hd__o22ai_1_351/Y sky130_fd_sc_hd__o22ai_1_376/A1 sky130_fd_sc_hd__a222oi_1_24/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_82 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_82/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__and2_0_82/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_415 sky130_fd_sc_hd__nand2_1_415/Y sky130_fd_sc_hd__nand2_1_416/Y
+ sky130_fd_sc_hd__nand2_1_417/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_146 sky130_fd_sc_hd__maj3_1_147/X sky130_fd_sc_hd__maj3_1_146/X
+ sky130_fd_sc_hd__maj3_1_146/B sky130_fd_sc_hd__maj3_1_146/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_362 sky130_fd_sc_hd__o22ai_1_375/A2 sky130_fd_sc_hd__nor2_1_230/B
+ sky130_fd_sc_hd__o22ai_1_362/Y sky130_fd_sc_hd__nor2_1_231/B sky130_fd_sc_hd__o32ai_1_8/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_93 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_93/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_93/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_426 sky130_fd_sc_hd__nand2_1_426/Y sky130_fd_sc_hd__nand2_1_439/B
+ sky130_fd_sc_hd__o21ai_1_355/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_157 sky130_fd_sc_hd__maj3_1_158/X sky130_fd_sc_hd__maj3_1_157/X
+ sky130_fd_sc_hd__maj3_1_157/B sky130_fd_sc_hd__maj3_1_157/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_373 sky130_fd_sc_hd__o22ai_1_375/A2 sky130_fd_sc_hd__o22ai_1_373/B1
+ sky130_fd_sc_hd__o22ai_1_373/Y sky130_fd_sc_hd__nor2_1_235/B sky130_fd_sc_hd__o32ai_1_8/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_437 sky130_fd_sc_hd__nand2_1_437/Y sky130_fd_sc_hd__nand2_1_439/B
+ sky130_fd_sc_hd__o21ai_1_380/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_384 sky130_fd_sc_hd__nand2_1_514/Y sky130_fd_sc_hd__nand2_1_513/Y
+ sky130_fd_sc_hd__o22ai_1_384/Y sky130_fd_sc_hd__o22ai_1_397/A1 sky130_fd_sc_hd__a21o_2_25/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_448 sky130_fd_sc_hd__o21a_1_45/B1 sky130_fd_sc_hd__fa_2_1236/A
+ sky130_fd_sc_hd__o21a_1_45/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_395 sky130_fd_sc_hd__nand2_1_516/Y sky130_fd_sc_hd__nand2_1_515/Y
+ sky130_fd_sc_hd__o22ai_1_395/Y sky130_fd_sc_hd__o22ai_1_395/A1 sky130_fd_sc_hd__a21o_2_24/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_459 sky130_fd_sc_hd__nor2_1_242/A sky130_fd_sc_hd__fa_2_1244/A
+ sky130_fd_sc_hd__fa_2_1243/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_17 sky130_fd_sc_hd__ha_2_46/SUM sky130_fd_sc_hd__nor2b_1_17/Y
+ sky130_fd_sc_hd__or2_1_0/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_28 sky130_fd_sc_hd__ha_2_63/SUM sky130_fd_sc_hd__nor2b_1_28/Y
+ sky130_fd_sc_hd__or2_0_2/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_39 sky130_fd_sc_hd__xor2_1_8/X sky130_fd_sc_hd__nor2b_1_39/Y
+ sky130_fd_sc_hd__or2_0_3/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1006 sky130_fd_sc_hd__a21oi_1_404/A1 sky130_fd_sc_hd__a21boi_1_6/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1006/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1017 sky130_fd_sc_hd__nor2_1_266/A sky130_fd_sc_hd__fa_2_1258/A
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1028 sky130_fd_sc_hd__nor2_1_278/B sky130_fd_sc_hd__fa_2_1306/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1028/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_70 sky130_fd_sc_hd__buf_8_70/A sky130_fd_sc_hd__buf_8_70/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__clkinv_1_1039 sky130_fd_sc_hd__o32ai_1_9/A3 sky130_fd_sc_hd__fa_2_1276/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1039/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_81 sky130_fd_sc_hd__buf_8_81/A sky130_fd_sc_hd__buf_8_81/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_200 VDD VSS sky130_fd_sc_hd__nor3_2_6/A sky130_fd_sc_hd__clkinv_2_17/Y
+ sky130_fd_sc_hd__nand3_4_1/B VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_8_92 sky130_fd_sc_hd__ha_2_46/A sky130_fd_sc_hd__buf_8_92/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_211 VDD VSS sky130_fd_sc_hd__ha_2_70/A sky130_fd_sc_hd__dfxtp_1_212/CLK
+ sky130_fd_sc_hd__and2_0_82/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_222 VDD VSS sky130_fd_sc_hd__ha_2_81/A sky130_fd_sc_hd__dfxtp_1_223/CLK
+ sky130_fd_sc_hd__nor2b_1_41/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_233 VDD VSS sky130_fd_sc_hd__fa_2_876/A sky130_fd_sc_hd__dfxtp_1_462/CLK
+ sky130_fd_sc_hd__and2_0_180/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_244 VDD VSS sky130_fd_sc_hd__fa_2_865/A sky130_fd_sc_hd__dfxtp_1_266/CLK
+ sky130_fd_sc_hd__and2_0_174/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_255 VDD VSS sky130_fd_sc_hd__dfxtp_1_255/Q sky130_fd_sc_hd__dfxtp_1_258/CLK
+ sky130_fd_sc_hd__and2_0_218/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_266 VDD VSS sky130_fd_sc_hd__dfxtp_1_266/Q sky130_fd_sc_hd__dfxtp_1_266/CLK
+ sky130_fd_sc_hd__and2_0_229/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_277 VDD VSS sky130_fd_sc_hd__dfxtp_1_277/Q sky130_fd_sc_hd__dfxtp_1_277/CLK
+ sky130_fd_sc_hd__and2_0_207/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_288 VDD VSS sky130_fd_sc_hd__a22o_1_59/A1 sky130_fd_sc_hd__clkinv_4_31/Y
+ sky130_fd_sc_hd__nand2_1_133/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_299 VDD VSS sky130_fd_sc_hd__a22o_1_50/A1 sky130_fd_sc_hd__dfxtp_1_304/CLK
+ sky130_fd_sc_hd__and2_0_99/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o22ai_1_8 sky130_fd_sc_hd__fa_2_9/A sky130_fd_sc_hd__fa_2_80/B sky130_fd_sc_hd__fa_2_118/B
+ sky130_fd_sc_hd__fa_2_5/A sky130_fd_sc_hd__fa_2_2/A VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_105 sky130_fd_sc_hd__fa_2_102/B sky130_fd_sc_hd__fa_2_97/CIN
+ sky130_fd_sc_hd__ha_2_97/A sky130_fd_sc_hd__ha_2_97/B sky130_fd_sc_hd__ha_2_96/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_116 sky130_fd_sc_hd__fa_2_118/CIN sky130_fd_sc_hd__fa_2_113/A
+ sky130_fd_sc_hd__fa_2_76/B sky130_fd_sc_hd__fa_2_116/B sky130_fd_sc_hd__fa_2_116/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_127 sky130_fd_sc_hd__fa_2_126/B sky130_fd_sc_hd__fa_2_127/SUM
+ sky130_fd_sc_hd__fa_2_127/A sky130_fd_sc_hd__fa_2_127/B sky130_fd_sc_hd__fa_2_131/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_138 sky130_fd_sc_hd__fa_2_137/CIN sky130_fd_sc_hd__fa_2_138/SUM
+ sky130_fd_sc_hd__fa_2_91/A sky130_fd_sc_hd__fa_2_96/A sky130_fd_sc_hd__fa_2_66/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_149 sky130_fd_sc_hd__fa_2_146/CIN sky130_fd_sc_hd__nor2_1_252/A
+ sky130_fd_sc_hd__fa_2_149/A sky130_fd_sc_hd__fa_2_149/B sky130_fd_sc_hd__fa_2_149/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_100 VDD VSS sky130_fd_sc_hd__buf_2_100/X sky130_fd_sc_hd__buf_2_100/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_111 VDD VSS sky130_fd_sc_hd__buf_2_111/X sky130_fd_sc_hd__buf_2_111/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__fa_2_1310 sky130_fd_sc_hd__xor2_1_297/B sky130_fd_sc_hd__mux2_2_222/A0
+ sky130_fd_sc_hd__fa_2_1310/A sky130_fd_sc_hd__fa_2_1310/B sky130_fd_sc_hd__fa_2_1310/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_122 VDD VSS sky130_fd_sc_hd__buf_2_122/X sky130_fd_sc_hd__buf_2_122/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_15 sky130_fd_sc_hd__fa_2_31/A sky130_fd_sc_hd__fa_2_277/B
+ sky130_fd_sc_hd__fa_2_212/B sky130_fd_sc_hd__ha_2_99/A sky130_fd_sc_hd__fa_2_281/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_1321 sky130_fd_sc_hd__fa_2_1322/CIN sky130_fd_sc_hd__mux2_2_247/A1
+ sky130_fd_sc_hd__fa_2_1321/A sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1321/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_133 VDD VSS sky130_fd_sc_hd__buf_2_133/X sky130_fd_sc_hd__nand3_2_3/Y
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_26 sky130_fd_sc_hd__ha_2_110/B sky130_fd_sc_hd__fa_2_412/A
+ sky130_fd_sc_hd__fa_2_383/A sky130_fd_sc_hd__ha_2_108/B sky130_fd_sc_hd__fa_2_409/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_144 VDD VSS sky130_fd_sc_hd__buf_4_98/A sky130_fd_sc_hd__buf_2_144/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_37 sky130_fd_sc_hd__fa_2_546/A sky130_fd_sc_hd__fa_2_427/B
+ sky130_fd_sc_hd__o22ai_1_37/Y sky130_fd_sc_hd__ha_2_125/A sky130_fd_sc_hd__fa_2_566/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_155 VDD VSS sky130_fd_sc_hd__buf_4_104/A sky130_fd_sc_hd__buf_6_57/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_48 sky130_fd_sc_hd__fa_2_699/A sky130_fd_sc_hd__fa_2_700/B
+ sky130_fd_sc_hd__fa_2_569/B sky130_fd_sc_hd__fa_2_701/B sky130_fd_sc_hd__fa_2_698/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_166 VDD VSS sky130_fd_sc_hd__buf_2_166/X sky130_fd_sc_hd__nor3_1_19/Y
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_59 sky130_fd_sc_hd__o22ai_1_59/A2 sky130_fd_sc_hd__fa_2_956/A
+ sky130_fd_sc_hd__o22ai_1_59/Y sky130_fd_sc_hd__fa_2_955/A sky130_fd_sc_hd__o22ai_1_59/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_177 VDD VSS sky130_fd_sc_hd__buf_2_177/X sky130_fd_sc_hd__buf_2_177/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_188 VDD VSS sky130_fd_sc_hd__buf_2_188/X sky130_fd_sc_hd__buf_2_188/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_199 VDD VSS sky130_fd_sc_hd__buf_2_199/X sky130_fd_sc_hd__buf_2_199/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1140 VDD VSS sky130_fd_sc_hd__mux2_2_148/A0 sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__dfxtp_1_999/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1151 VDD VSS sky130_fd_sc_hd__mux2_2_141/A0 sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__o22ai_1_286/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1162 VDD VSS sky130_fd_sc_hd__fa_2_862/B sky130_fd_sc_hd__dfxtp_1_1179/CLK
+ sky130_fd_sc_hd__a21oi_1_375/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1173 VDD VSS sky130_fd_sc_hd__fa_2_851/B sky130_fd_sc_hd__dfxtp_1_1184/CLK
+ sky130_fd_sc_hd__a21oi_1_369/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1184 VDD VSS sky130_fd_sc_hd__fa_2_937/A sky130_fd_sc_hd__dfxtp_1_1184/CLK
+ sky130_fd_sc_hd__o21a_1_46/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1195 VDD VSS sky130_fd_sc_hd__fa_2_1244/A sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__mux2_2_212/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__ha_2_0 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_0/A sky130_fd_sc_hd__xor2_1_0/A
+ sky130_fd_sc_hd__ha_2_0/SUM sky130_fd_sc_hd__ha_2_0/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__buf_4_17 VDD VSS sky130_fd_sc_hd__buf_4_17/X sky130_fd_sc_hd__buf_8_25/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_28 VDD VSS sky130_fd_sc_hd__buf_4_28/X sky130_fd_sc_hd__buf_8_27/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_39 VDD VSS sky130_fd_sc_hd__buf_4_39/X sky130_fd_sc_hd__buf_4_39/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__clkbuf_1_11 VSS VDD sky130_fd_sc_hd__buf_4_9/A sky130_fd_sc_hd__clkbuf_4_3/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_22 VSS VDD sky130_fd_sc_hd__clkbuf_1_22/X sky130_fd_sc_hd__clkbuf_1_22/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_33 VSS VDD sky130_fd_sc_hd__clkbuf_1_33/X sky130_fd_sc_hd__clkbuf_1_33/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_44 VSS VDD sky130_fd_sc_hd__clkbuf_1_44/X sky130_fd_sc_hd__clkbuf_1_44/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_650 sky130_fd_sc_hd__fa_2_652/B sky130_fd_sc_hd__fa_2_650/SUM
+ sky130_fd_sc_hd__fa_2_650/A sky130_fd_sc_hd__fa_2_650/B sky130_fd_sc_hd__fa_2_654/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_55 VSS VDD sky130_fd_sc_hd__clkbuf_1_55/X sky130_fd_sc_hd__clkbuf_1_55/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_661 sky130_fd_sc_hd__fa_2_581/A sky130_fd_sc_hd__fa_2_582/B
+ sky130_fd_sc_hd__fa_2_661/A sky130_fd_sc_hd__fa_2_661/B sky130_fd_sc_hd__fa_2_666/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_66 VSS VDD sky130_fd_sc_hd__clkbuf_1_66/X sky130_fd_sc_hd__clkbuf_1_66/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_672 sky130_fd_sc_hd__fa_2_674/CIN sky130_fd_sc_hd__fa_2_666/B
+ sky130_fd_sc_hd__fa_2_672/A sky130_fd_sc_hd__fa_2_683/B sky130_fd_sc_hd__ha_2_130/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_77 VSS VDD sky130_fd_sc_hd__nand4_1_10/A sky130_fd_sc_hd__a22oi_2_11/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_683 sky130_fd_sc_hd__fa_2_680/A sky130_fd_sc_hd__fa_2_675/A
+ sky130_fd_sc_hd__fa_2_692/A sky130_fd_sc_hd__fa_2_683/B sky130_fd_sc_hd__fa_2_683/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_88 VSS VDD sky130_fd_sc_hd__clkbuf_1_88/X sky130_fd_sc_hd__nand3_2_0/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_694 sky130_fd_sc_hd__fa_2_573/A sky130_fd_sc_hd__fa_2_574/B
+ sky130_fd_sc_hd__fa_2_694/A sky130_fd_sc_hd__fa_2_694/B sky130_fd_sc_hd__fa_2_694/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_99 VSS VDD sky130_fd_sc_hd__clkbuf_1_99/X sky130_fd_sc_hd__nor3_1_7/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a21oi_1_207 sky130_fd_sc_hd__a21o_2_5/A2 sky130_fd_sc_hd__o22ai_1_175/Y
+ sky130_fd_sc_hd__a21oi_1_207/Y sky130_fd_sc_hd__fa_2_1051/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_218 sky130_fd_sc_hd__clkinv_1_729/Y sky130_fd_sc_hd__o21ai_1_252/Y
+ sky130_fd_sc_hd__a21oi_1_218/Y sky130_fd_sc_hd__nand2_1_331/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__or2_0_13 sky130_fd_sc_hd__or2_0_13/A sky130_fd_sc_hd__or2_0_13/X
+ sky130_fd_sc_hd__or2_0_13/B VSS VDD VSS VDD sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__a21oi_1_229 sky130_fd_sc_hd__a21o_2_5/X sky130_fd_sc_hd__o22ai_1_205/Y
+ sky130_fd_sc_hd__a21oi_1_229/Y sky130_fd_sc_hd__a211o_1_9/A1 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_2_14 sky130_fd_sc_hd__nor3_2_7/Y sky130_fd_sc_hd__a22oi_2_14/A2
+ sky130_fd_sc_hd__nor3_2_8/Y sky130_fd_sc_hd__a22oi_2_14/B2 sky130_fd_sc_hd__nand4_1_49/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__a22oi_2_25 sky130_fd_sc_hd__a22oi_2_25/A1 sky130_fd_sc_hd__a22oi_2_25/A2
+ sky130_fd_sc_hd__a22oi_2_25/B1 sky130_fd_sc_hd__a22oi_2_25/B2 sky130_fd_sc_hd__nand4_1_58/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__buf_12_0 sky130_fd_sc_hd__buf_6_8/X sky130_fd_sc_hd__buf_12_0/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__nand2_1_201 sky130_fd_sc_hd__nor2_1_20/B sky130_fd_sc_hd__nand2_1_201/B
+ sky130_fd_sc_hd__nor2_1_21/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_800 sky130_fd_sc_hd__o22ai_1_228/A1 sky130_fd_sc_hd__a21o_2_8/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_800/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_212 sky130_fd_sc_hd__xnor2_1_28/B sky130_fd_sc_hd__nand2_1_212/B
+ sky130_fd_sc_hd__nor2_1_30/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_811 sky130_fd_sc_hd__nor2_1_163/B sky130_fd_sc_hd__xor2_1_185/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_811/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_223 sky130_fd_sc_hd__o22ai_1_60/A2 sky130_fd_sc_hd__a31oi_1_2/A2
+ sky130_fd_sc_hd__nand2_1_223/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_822 sky130_fd_sc_hd__clkinv_1_822/Y sky130_fd_sc_hd__nor2_1_172/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_822/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_170 sky130_fd_sc_hd__a21oi_1_197/Y sky130_fd_sc_hd__a21oi_1_206/Y
+ sky130_fd_sc_hd__o22ai_1_170/Y sky130_fd_sc_hd__nor2_2_13/B sky130_fd_sc_hd__nor2_1_126/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_234 sky130_fd_sc_hd__xnor2_1_52/B sky130_fd_sc_hd__o21ai_1_76/B1
+ sky130_fd_sc_hd__o21ai_1_83/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_181 sky130_fd_sc_hd__nand4_1_86/A sky130_fd_sc_hd__o22ai_1_206/A1
+ sky130_fd_sc_hd__o22ai_1_181/Y sky130_fd_sc_hd__o22ai_1_206/B1 sky130_fd_sc_hd__nor2_1_120/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_833 sky130_fd_sc_hd__o22ai_1_252/B1 sky130_fd_sc_hd__fa_2_1134/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_833/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_245 sky130_fd_sc_hd__nand2_1_245/Y sky130_fd_sc_hd__nor2_1_54/B
+ sky130_fd_sc_hd__nor2_1_54/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_192 sky130_fd_sc_hd__nand4_1_86/A sky130_fd_sc_hd__o22ai_1_206/B1
+ sky130_fd_sc_hd__o22ai_1_192/Y sky130_fd_sc_hd__o22ai_1_206/A1 sky130_fd_sc_hd__nand4_1_86/C
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_844 sky130_fd_sc_hd__nor2_1_157/B sky130_fd_sc_hd__fa_2_1143/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_844/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_256 sky130_fd_sc_hd__o21a_1_6/B1 sky130_fd_sc_hd__fa_2_979/A
+ sky130_fd_sc_hd__o21a_1_6/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_855 sky130_fd_sc_hd__o22ai_1_265/B1 sky130_fd_sc_hd__fa_2_1152/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_855/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_267 sky130_fd_sc_hd__nand3_1_49/C sky130_fd_sc_hd__fa_2_986/A
+ sky130_fd_sc_hd__nor2_4_10/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand4_1_40 sky130_fd_sc_hd__nand4_1_40/C sky130_fd_sc_hd__nand4_1_40/B
+ sky130_fd_sc_hd__buf_2_290/A sky130_fd_sc_hd__nand4_1_40/D sky130_fd_sc_hd__nand4_1_40/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__clkinv_1_866 sky130_fd_sc_hd__nor3_1_39/B sky130_fd_sc_hd__o32ai_1_5/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_866/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_278 sky130_fd_sc_hd__nand2_1_278/Y sky130_fd_sc_hd__fa_2_1015/A
+ sky130_fd_sc_hd__nor2_4_10/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_877 sky130_fd_sc_hd__o31ai_1_7/B1 sky130_fd_sc_hd__a221oi_1_3/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_877/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand4_1_51 sky130_fd_sc_hd__nand4_1_51/C sky130_fd_sc_hd__nand4_1_51/B
+ sky130_fd_sc_hd__buf_2_270/A sky130_fd_sc_hd__nand4_1_51/D sky130_fd_sc_hd__nand4_1_51/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand2_1_289 sky130_fd_sc_hd__xnor2_1_73/B sky130_fd_sc_hd__nand2_1_289/B
+ sky130_fd_sc_hd__nand2_1_298/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_888 sky130_fd_sc_hd__nor2_1_205/A sky130_fd_sc_hd__or3_1_3/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_888/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand4_1_62 sky130_fd_sc_hd__nand4_1_62/C sky130_fd_sc_hd__nand4_1_62/B
+ sky130_fd_sc_hd__buf_2_265/A sky130_fd_sc_hd__buf_2_236/X sky130_fd_sc_hd__nand4_1_62/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__clkinv_1_899 sky130_fd_sc_hd__nand2_1_423/B sky130_fd_sc_hd__fa_2_300/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_899/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand4_1_73 sky130_fd_sc_hd__nand4_1_73/C sky130_fd_sc_hd__nand4_1_73/B
+ sky130_fd_sc_hd__nand2_1_6/B sky130_fd_sc_hd__nand4_1_73/D sky130_fd_sc_hd__nand4_1_73/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_84 sky130_fd_sc_hd__nand4_1_84/C sky130_fd_sc_hd__nand4_1_84/B
+ sky130_fd_sc_hd__nand4_1_84/Y sky130_fd_sc_hd__nand4_1_84/D sky130_fd_sc_hd__nand4_1_84/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__conb_1_11 sky130_fd_sc_hd__conb_1_11/LO sky130_fd_sc_hd__conb_1_11/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_22 sky130_fd_sc_hd__conb_1_22/LO sky130_fd_sc_hd__conb_1_22/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__mux2_2_6 VSS VDD sky130_fd_sc_hd__mux2_2_6/A1 sky130_fd_sc_hd__mux2_2_6/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_6/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1140 sky130_fd_sc_hd__fa_2_1141/CIN sky130_fd_sc_hd__and2_0_320/A
+ sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__fa_2_1140/B sky130_fd_sc_hd__xor2_1_182/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1151 sky130_fd_sc_hd__fa_2_1152/CIN sky130_fd_sc_hd__mux2_2_90/A1
+ sky130_fd_sc_hd__fa_2_1151/A sky130_fd_sc_hd__fa_2_1151/B sky130_fd_sc_hd__fa_2_1151/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1162 sky130_fd_sc_hd__fa_2_1163/CIN sky130_fd_sc_hd__mux2_2_119/A1
+ sky130_fd_sc_hd__fa_2_1162/A sky130_fd_sc_hd__fa_2_1172/B sky130_fd_sc_hd__fa_2_1162/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1173 sky130_fd_sc_hd__fa_2_1174/CIN sky130_fd_sc_hd__and2_0_324/A
+ sky130_fd_sc_hd__fa_2_1173/A sky130_fd_sc_hd__fa_2_1173/B sky130_fd_sc_hd__xor2_1_206/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1184 sky130_fd_sc_hd__fa_2_1185/CIN sky130_fd_sc_hd__mux2_2_139/A1
+ sky130_fd_sc_hd__fa_2_1184/A sky130_fd_sc_hd__fa_2_1184/B sky130_fd_sc_hd__fa_2_1184/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1195 sky130_fd_sc_hd__fa_2_1196/CIN sky130_fd_sc_hd__mux2_2_158/A1
+ sky130_fd_sc_hd__fa_2_1195/A sky130_fd_sc_hd__fa_2_1195/B sky130_fd_sc_hd__fa_2_1195/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o2bb2ai_1_2 sky130_fd_sc_hd__o2bb2ai_1_2/Y sky130_fd_sc_hd__nor2_1_18/Y
+ sky130_fd_sc_hd__ha_2_156/SUM sky130_fd_sc_hd__o21ai_1_31/A1 sky130_fd_sc_hd__maj3_1_3/C
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_480 sky130_fd_sc_hd__fa_2_482/B sky130_fd_sc_hd__fa_2_480/SUM
+ sky130_fd_sc_hd__fa_2_546/B sky130_fd_sc_hd__fa_2_480/B sky130_fd_sc_hd__fa_2_480/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_491 sky130_fd_sc_hd__fa_2_495/CIN sky130_fd_sc_hd__fa_2_489/B
+ sky130_fd_sc_hd__fa_2_491/A sky130_fd_sc_hd__fa_2_491/B sky130_fd_sc_hd__fa_2_500/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_1_107 sky130_fd_sc_hd__inv_2_69/A sky130_fd_sc_hd__inv_2_62/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_107/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_118 sky130_fd_sc_hd__clkinv_1_119/A sky130_fd_sc_hd__dfxtp_1_162/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_118/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_129 sky130_fd_sc_hd__buf_6_31/A sky130_fd_sc_hd__and2_4_0/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_129/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_7 VSS VDD sky130_fd_sc_hd__o21ai_1_7/A2 sky130_fd_sc_hd__or4_1_0/C
+ sky130_fd_sc_hd__a21oi_1_4/Y sky130_fd_sc_hd__o21ai_1_7/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__bufbuf_16_6 sky130_fd_sc_hd__inv_2_116/A sky130_fd_sc_hd__buf_6_74/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__nor2_1_201 sky130_fd_sc_hd__nor2_1_205/A sky130_fd_sc_hd__nor2_1_201/Y
+ sky130_fd_sc_hd__o31ai_1_7/A2 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_212 sky130_fd_sc_hd__nor2_1_212/B sky130_fd_sc_hd__nor2_1_212/Y
+ sky130_fd_sc_hd__nor2_1_212/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_223 sky130_fd_sc_hd__o21a_1_42/A1 sky130_fd_sc_hd__nor2_1_223/Y
+ sky130_fd_sc_hd__nor2_1_223/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_234 sky130_fd_sc_hd__nor2_1_234/B sky130_fd_sc_hd__nor2_1_234/Y
+ sky130_fd_sc_hd__nor2_1_234/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_245 sky130_fd_sc_hd__nor2_1_248/A sky130_fd_sc_hd__nor2_1_245/Y
+ sky130_fd_sc_hd__nor2_1_245/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_256 sky130_fd_sc_hd__or3_1_4/X sky130_fd_sc_hd__nor2_1_256/Y
+ sky130_fd_sc_hd__nor2_1_256/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_267 sky130_fd_sc_hd__o21a_1_55/A1 sky130_fd_sc_hd__nor2_1_267/Y
+ sky130_fd_sc_hd__nor2_1_267/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_278 sky130_fd_sc_hd__nor2_1_278/B sky130_fd_sc_hd__o21a_1_63/A1
+ sky130_fd_sc_hd__o21a_1_64/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_289 sky130_fd_sc_hd__or3_1_5/C sky130_fd_sc_hd__nor2_1_289/Y
+ sky130_fd_sc_hd__or3_1_5/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_430 sky130_fd_sc_hd__buf_8_189/X sky130_fd_sc_hd__buf_12_493/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_441 sky130_fd_sc_hd__buf_4_116/X sky130_fd_sc_hd__buf_12_485/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_300 sky130_fd_sc_hd__clkbuf_1_376/X sky130_fd_sc_hd__nor2_2_5/Y
+ sky130_fd_sc_hd__buf_2_207/X sky130_fd_sc_hd__clkbuf_1_463/X sky130_fd_sc_hd__nand4_1_74/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_452 sky130_fd_sc_hd__buf_6_76/X sky130_fd_sc_hd__buf_12_487/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_311 sky130_fd_sc_hd__nor2_2_4/Y sky130_fd_sc_hd__clkbuf_1_377/X
+ sky130_fd_sc_hd__a22oi_1_311/B2 sky130_fd_sc_hd__clkbuf_4_179/X sky130_fd_sc_hd__nand4_1_77/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_463 sky130_fd_sc_hd__buf_12_463/A sky130_fd_sc_hd__buf_12_479/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_322 sky130_fd_sc_hd__nor2b_1_88/A sky130_fd_sc_hd__nor2_1_39/A
+ sky130_fd_sc_hd__nor2_1_38/Y sky130_fd_sc_hd__nor2_1_39/B sky130_fd_sc_hd__o31ai_1_4/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_474 sky130_fd_sc_hd__buf_12_474/A sky130_fd_sc_hd__buf_12_474/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_333 sky130_fd_sc_hd__a21oi_1_96/A1 sky130_fd_sc_hd__a211o_1_8/A2
+ sky130_fd_sc_hd__nand2_1_264/A sky130_fd_sc_hd__o21ai_1_120/Y sky130_fd_sc_hd__a22oi_1_333/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_485 sky130_fd_sc_hd__buf_12_485/A sky130_fd_sc_hd__buf_12_485/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_344 sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__nor2_2_8/Y
+ sky130_fd_sc_hd__fa_2_1006/A sky130_fd_sc_hd__fa_2_1008/A sky130_fd_sc_hd__a22oi_1_344/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_496 sky130_fd_sc_hd__buf_12_496/A sky130_fd_sc_hd__buf_12_496/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_355 sky130_fd_sc_hd__clkinv_1_706/Y sky130_fd_sc_hd__o21ai_1_234/Y
+ sky130_fd_sc_hd__nand2_1_321/A sky130_fd_sc_hd__nand2_1_331/B sky130_fd_sc_hd__a22oi_1_355/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_366 sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__nor2_4_13/Y
+ sky130_fd_sc_hd__fa_2_1074/A sky130_fd_sc_hd__fa_2_1075/A sky130_fd_sc_hd__a22oi_1_366/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_377 sky130_fd_sc_hd__nor2_1_180/Y sky130_fd_sc_hd__nor2_1_182/Y
+ sky130_fd_sc_hd__fa_2_1149/A sky130_fd_sc_hd__fa_2_1145/A sky130_fd_sc_hd__a22oi_1_377/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_388 sky130_fd_sc_hd__clkinv_1_946/Y sky130_fd_sc_hd__nor3_1_40/B
+ sky130_fd_sc_hd__fa_2_1230/A sky130_fd_sc_hd__fa_2_1231/A sky130_fd_sc_hd__a22oi_1_388/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_630 sky130_fd_sc_hd__nand2_1_321/A sky130_fd_sc_hd__nor2_2_13/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_630/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22oi_1_399 sky130_fd_sc_hd__fa_2_1283/A sky130_fd_sc_hd__nor2_1_309/Y
+ sky130_fd_sc_hd__nor2_1_307/Y sky130_fd_sc_hd__fa_2_1279/A sky130_fd_sc_hd__a22oi_1_399/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_641 sky130_fd_sc_hd__o22ai_1_159/B2 sky130_fd_sc_hd__ha_2_190/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_641/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_652 sky130_fd_sc_hd__nor2_1_96/B sky130_fd_sc_hd__nand2_1_305/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_652/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_663 sky130_fd_sc_hd__clkinv_1_663/Y sky130_fd_sc_hd__nor2_1_93/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_663/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_674 sky130_fd_sc_hd__o21ai_1_192/A1 sky130_fd_sc_hd__nand2_1_294/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_674/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_685 sky130_fd_sc_hd__nor2_1_100/B sky130_fd_sc_hd__fa_2_1117/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_685/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_696 sky130_fd_sc_hd__nand2_1_318/A sky130_fd_sc_hd__a21oi_1_199/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_696/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand3_1_3 sky130_fd_sc_hd__nand3_1_3/Y sky130_fd_sc_hd__nand3_1_3/A
+ sky130_fd_sc_hd__nand3_1_3/C sky130_fd_sc_hd__nand3_1_3/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__xnor2_1_30 VSS VDD sky130_fd_sc_hd__nor2_1_34/B sky130_fd_sc_hd__xnor2_1_30/Y
+ sky130_fd_sc_hd__nor4_1_8/C VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_41 VSS VDD sky130_fd_sc_hd__xnor2_1_41/B sky130_fd_sc_hd__xnor2_1_41/Y
+ sky130_fd_sc_hd__nor2_1_44/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_52 VSS VDD sky130_fd_sc_hd__xnor2_1_52/B sky130_fd_sc_hd__xnor2_1_52/Y
+ sky130_fd_sc_hd__xnor2_1_52/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_63 VSS VDD sky130_fd_sc_hd__xnor2_1_63/B sky130_fd_sc_hd__xnor2_1_63/Y
+ sky130_fd_sc_hd__nor2_1_92/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_74 VSS VDD sky130_fd_sc_hd__xnor2_1_74/B sky130_fd_sc_hd__xnor2_1_74/Y
+ sky130_fd_sc_hd__nor2_1_95/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_85 VSS VDD sky130_fd_sc_hd__xnor2_1_85/B sky130_fd_sc_hd__xnor2_1_85/Y
+ sky130_fd_sc_hd__xnor2_1_85/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_96 VSS VDD sky130_fd_sc_hd__xor2_1_185/A sky130_fd_sc_hd__xnor2_1_96/Y
+ sky130_fd_sc_hd__xnor2_1_96/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkbuf_1_408 VSS VDD sky130_fd_sc_hd__clkbuf_1_408/X sky130_fd_sc_hd__clkbuf_1_408/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_419 VSS VDD sky130_fd_sc_hd__clkbuf_1_419/X sky130_fd_sc_hd__clkbuf_1_419/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o32ai_1_2 sky130_fd_sc_hd__nor3_1_38/C sky130_fd_sc_hd__o32ai_1_2/Y
+ sky130_fd_sc_hd__o32ai_1_2/A1 sky130_fd_sc_hd__o32ai_1_2/A3 sky130_fd_sc_hd__o32ai_1_2/B2
+ sky130_fd_sc_hd__o32ai_1_2/B1 VDD VSS VSS VDD sky130_fd_sc_hd__o32ai_1
Xsky130_fd_sc_hd__clkbuf_16_0 sky130_fd_sc_hd__clkbuf_16_5/A sky130_fd_sc_hd__buf_8_51/X
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__nor4_1_0 sky130_fd_sc_hd__inv_2_0/Y sky130_fd_sc_hd__inv_2_1/Y sky130_fd_sc_hd__nor4_1_0/Y
+ sky130_fd_sc_hd__nor4_1_0/A sky130_fd_sc_hd__nor4_1_0/B VDD VSS VSS VDD sky130_fd_sc_hd__nor4_1
Xsky130_fd_sc_hd__diode_2_160 sky130_fd_sc_hd__nand4_1_66/D VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_171 sky130_fd_sc_hd__clkbuf_4_179/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_182 sky130_fd_sc_hd__buf_2_246/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_193 sky130_fd_sc_hd__buf_2_249/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkinv_2_15 sky130_fd_sc_hd__inv_2_75/A sky130_fd_sc_hd__clkinv_2_15/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_15/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkbuf_4_202 sky130_fd_sc_hd__nand4_1_64/D sky130_fd_sc_hd__a22oi_1_257/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_2_26 sky130_fd_sc_hd__nand4_1_73/D sky130_fd_sc_hd__clkinv_2_26/A
+ VSS VDD VDD VSS VSS sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkbuf_4_213 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__nor2_1_140/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_2_37 sky130_fd_sc_hd__clkinv_4_26/A sky130_fd_sc_hd__clkinv_8_58/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_37/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkbuf_4_224 sky130_fd_sc_hd__nor3_2_0/A adc_bypass_en VSS VDD VDD
+ VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_2_48 sky130_fd_sc_hd__clkinv_4_57/A sky130_fd_sc_hd__clkinv_2_48/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_48/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__buf_12_260 sky130_fd_sc_hd__buf_12_260/A sky130_fd_sc_hd__buf_12_260/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_271 sky130_fd_sc_hd__inv_2_78/Y sky130_fd_sc_hd__buf_12_359/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_130 sky130_fd_sc_hd__clkbuf_4_72/X sky130_fd_sc_hd__clkbuf_4_73/X
+ sky130_fd_sc_hd__a22oi_1_130/B2 sky130_fd_sc_hd__buf_2_86/X sky130_fd_sc_hd__buf_2_104/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_282 sky130_fd_sc_hd__inv_2_91/Y sky130_fd_sc_hd__buf_12_282/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_141 sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__a22oi_2_12/A1
+ sky130_fd_sc_hd__buf_2_67/X sky130_fd_sc_hd__clkbuf_1_158/X sky130_fd_sc_hd__a22oi_1_141/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_293 sky130_fd_sc_hd__buf_8_145/X sky130_fd_sc_hd__buf_12_293/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_152 sky130_fd_sc_hd__clkbuf_1_351/X sky130_fd_sc_hd__clkbuf_1_353/X
+ sky130_fd_sc_hd__clkbuf_4_120/X sky130_fd_sc_hd__a22oi_1_152/A2 sky130_fd_sc_hd__nand4_1_33/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_163 sky130_fd_sc_hd__clkbuf_1_265/X sky130_fd_sc_hd__clkbuf_1_266/X
+ sky130_fd_sc_hd__clkbuf_1_278/X sky130_fd_sc_hd__a22oi_1_163/A2 sky130_fd_sc_hd__a22oi_1_163/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_174 sky130_fd_sc_hd__clkbuf_1_264/X sky130_fd_sc_hd__nor2_2_3/Y
+ sky130_fd_sc_hd__a22oi_1_174/B2 sky130_fd_sc_hd__clkbuf_4_131/X sky130_fd_sc_hd__nand4_1_38/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_185 sky130_fd_sc_hd__clkbuf_4_111/X sky130_fd_sc_hd__clkbuf_4_112/X
+ sky130_fd_sc_hd__a22oi_1_185/B2 sky130_fd_sc_hd__clkbuf_1_288/X sky130_fd_sc_hd__a22oi_1_185/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_196 sky130_fd_sc_hd__clkbuf_1_351/X sky130_fd_sc_hd__clkbuf_1_353/X
+ sky130_fd_sc_hd__clkinv_2_9/Y sky130_fd_sc_hd__a22oi_1_196/A2 sky130_fd_sc_hd__nand4_1_44/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_460 sky130_fd_sc_hd__a211o_1_6/A1 sky130_fd_sc_hd__nor2_1_77/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_460/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_471 sky130_fd_sc_hd__a211o_1_3/A1 sky130_fd_sc_hd__nor2_1_76/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_471/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_482 sky130_fd_sc_hd__o22ai_1_87/B2 sky130_fd_sc_hd__ha_2_172/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_482/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_493 sky130_fd_sc_hd__nor2_1_45/B sky130_fd_sc_hd__nand2_1_247/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_493/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_407 VSS VDD sky130_fd_sc_hd__a222oi_1_27/Y sky130_fd_sc_hd__nor2_1_267/A
+ sky130_fd_sc_hd__a22oi_1_389/Y sky130_fd_sc_hd__o21ai_1_407/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_418 VSS VDD sky130_fd_sc_hd__a222oi_1_30/Y sky130_fd_sc_hd__nor2_1_267/A
+ sky130_fd_sc_hd__nand2_1_486/Y sky130_fd_sc_hd__xor2_1_235/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_429 VSS VDD sky130_fd_sc_hd__a222oi_1_31/Y sky130_fd_sc_hd__nor2_1_267/A
+ sky130_fd_sc_hd__a22oi_1_393/Y sky130_fd_sc_hd__o21ai_1_429/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a21oi_1_390 sky130_fd_sc_hd__nor2_1_267/Y sky130_fd_sc_hd__nor2_1_258/Y
+ sky130_fd_sc_hd__a21oi_1_390/Y sky130_fd_sc_hd__fa_2_1232/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nor2_4_16 sky130_fd_sc_hd__nor3_1_39/A sky130_fd_sc_hd__nor2_4_16/A
+ sky130_fd_sc_hd__nor2_4_16/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__xor2_1_201 sky130_fd_sc_hd__fa_2_1173/A sky130_fd_sc_hd__fa_2_1178/B
+ sky130_fd_sc_hd__xor2_1_201/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_212 sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__fa_2_1206/B
+ sky130_fd_sc_hd__xor2_1_212/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_223 sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__fa_2_1195/B
+ sky130_fd_sc_hd__xor2_1_223/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_234 sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1241/B
+ sky130_fd_sc_hd__xor2_1_234/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_245 sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1230/B
+ sky130_fd_sc_hd__xor2_1_245/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_256 sky130_fd_sc_hd__xor2_1_267/B sky130_fd_sc_hd__fa_2_1258/B
+ sky130_fd_sc_hd__xor2_1_256/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_607 VDD VSS sky130_fd_sc_hd__and2_0_228/A sky130_fd_sc_hd__dfxtp_1_611/CLK
+ sky130_fd_sc_hd__fa_2_1027/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_267 sky130_fd_sc_hd__xor2_1_267/B sky130_fd_sc_hd__fa_2_1247/B
+ sky130_fd_sc_hd__xor2_1_267/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_618 VDD VSS sky130_fd_sc_hd__fa_2_820/B sky130_fd_sc_hd__dfxtp_1_626/CLK
+ sky130_fd_sc_hd__o21a_1_5/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_278 sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__xor2_1_278/X
+ sky130_fd_sc_hd__xor2_1_298/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_289 sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1282/B
+ sky130_fd_sc_hd__xor2_1_289/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_629 VDD VSS sky130_fd_sc_hd__fa_2_993/B sky130_fd_sc_hd__clkinv_8_41/Y
+ sky130_fd_sc_hd__and2_0_277/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_205 VSS VDD sky130_fd_sc_hd__buf_12_132/A sky130_fd_sc_hd__ha_2_43/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_216 VSS VDD sky130_fd_sc_hd__buf_8_106/A sky130_fd_sc_hd__buf_4_44/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_227 VSS VDD sky130_fd_sc_hd__clkbuf_1_228/A sky130_fd_sc_hd__buf_8_69/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_238 VSS VDD sky130_fd_sc_hd__buf_4_43/A sky130_fd_sc_hd__buf_8_83/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_249 VSS VDD sky130_fd_sc_hd__clkbuf_1_249/X sky130_fd_sc_hd__clkbuf_1_249/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_2_50 VDD VSS sky130_fd_sc_hd__buf_8_84/A sky130_fd_sc_hd__ha_2_45/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_61 VDD VSS sky130_fd_sc_hd__buf_2_61/X sky130_fd_sc_hd__buf_2_61/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_72 VDD VSS sky130_fd_sc_hd__buf_2_72/X sky130_fd_sc_hd__buf_2_72/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_83 VDD VSS sky130_fd_sc_hd__buf_2_83/X sky130_fd_sc_hd__buf_2_83/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_94 VDD VSS sky130_fd_sc_hd__buf_2_94/X sky130_fd_sc_hd__buf_2_94/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__diode_2_1 sky130_fd_sc_hd__buf_2_69/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__and2_0_203 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_203/X sky130_fd_sc_hd__and2_0_235/B
+ sky130_fd_sc_hd__and2_0_203/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_214 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_214/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_214/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_225 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_225/X sky130_fd_sc_hd__and2_0_235/B
+ sky130_fd_sc_hd__and2_0_225/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_236 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_236/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__fa_2_877/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_247 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_247/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__and2_0_247/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_258 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_258/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__fa_2_959/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_269 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_269/X sky130_fd_sc_hd__mux2_2_37/S
+ sky130_fd_sc_hd__and2_0_269/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__sdlclkp_2_8 sky130_fd_sc_hd__conb_1_18/LO sky130_fd_sc_hd__clkinv_8_104/A
+ sky130_fd_sc_hd__dfxtp_1_476/CLK sky130_fd_sc_hd__nand3_1_43/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__a22o_2_2 sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__ha_2_68/A
+ sky130_fd_sc_hd__a22o_2_2/X sky130_fd_sc_hd__dfxtp_1_3/Q sky130_fd_sc_hd__a22o_2_3/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_2
Xsky130_fd_sc_hd__o31ai_1_1 sky130_fd_sc_hd__o31ai_1_1/Y sky130_fd_sc_hd__xor2_1_9/A
+ sky130_fd_sc_hd__nor4_1_4/B sky130_fd_sc_hd__nor4_1_4/C sky130_fd_sc_hd__o31ai_1_1/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__o31ai_1
Xsky130_fd_sc_hd__clkinv_1_290 sky130_fd_sc_hd__fa_2_76/A sky130_fd_sc_hd__ha_2_91/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_290/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkbuf_4_11 sky130_fd_sc_hd__clkbuf_4_11/X sky130_fd_sc_hd__clkbuf_4_11/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_204 VSS VDD sky130_fd_sc_hd__xnor2_1_68/A sky130_fd_sc_hd__nor2_1_107/Y
+ sky130_fd_sc_hd__nand2_1_299/Y sky130_fd_sc_hd__xnor2_1_70/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_22 sky130_fd_sc_hd__clkbuf_4_22/X sky130_fd_sc_hd__clkbuf_4_22/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_215 VSS VDD sky130_fd_sc_hd__nand2_2_6/Y sky130_fd_sc_hd__o22ai_1_173/A2
+ sky130_fd_sc_hd__a21oi_1_191/Y sky130_fd_sc_hd__xor2_1_121/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_33 sky130_fd_sc_hd__a22oi_2_9/B2 sky130_fd_sc_hd__clkbuf_4_33/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_226 VSS VDD sky130_fd_sc_hd__nor2_1_127/A sky130_fd_sc_hd__nor2_1_130/Y
+ sky130_fd_sc_hd__a21oi_1_198/Y sky130_fd_sc_hd__xor2_1_127/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_44 sky130_fd_sc_hd__nand4_1_13/D sky130_fd_sc_hd__a22oi_1_72/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_237 VSS VDD sky130_fd_sc_hd__o22ai_1_204/B1 sky130_fd_sc_hd__nand4_1_86/C
+ sky130_fd_sc_hd__a21oi_1_211/Y sky130_fd_sc_hd__o21ai_1_237/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_55 sky130_fd_sc_hd__nand4_1_2/D sky130_fd_sc_hd__a22oi_1_35/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_248 VSS VDD sky130_fd_sc_hd__a21oi_1_234/Y sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__nand2b_1_16/Y sky130_fd_sc_hd__o21ai_1_248/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_66 sky130_fd_sc_hd__buf_2_40/A sky130_fd_sc_hd__dfxtp_1_260/Q
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_259 VSS VDD sky130_fd_sc_hd__a21oi_1_240/Y sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__a21oi_1_224/Y sky130_fd_sc_hd__xor2_1_103/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_77 sky130_fd_sc_hd__clkbuf_4_77/X sky130_fd_sc_hd__clkbuf_4_77/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_88 sky130_fd_sc_hd__clkbuf_4_88/X sky130_fd_sc_hd__clkbuf_4_88/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_99 sky130_fd_sc_hd__buf_12_153/A sky130_fd_sc_hd__buf_2_121/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__nor2_4_1 sky130_fd_sc_hd__nor2_4_1/Y sky130_fd_sc_hd__nor2_4_2/A
+ sky130_fd_sc_hd__inv_2_0/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__buf_8_150 sky130_fd_sc_hd__buf_8_150/A sky130_fd_sc_hd__buf_8_150/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_161 sky130_fd_sc_hd__buf_8_161/A sky130_fd_sc_hd__buf_8_161/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_172 sky130_fd_sc_hd__buf_8_172/A sky130_fd_sc_hd__buf_8_172/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_183 sky130_fd_sc_hd__inv_2_131/A sky130_fd_sc_hd__buf_8_183/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_194 sky130_fd_sc_hd__buf_6_59/X sky130_fd_sc_hd__buf_6_77/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_404 VDD VSS sky130_fd_sc_hd__nor2_1_60/A sky130_fd_sc_hd__dfxtp_1_425/CLK
+ sky130_fd_sc_hd__and2_0_128/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_415 VDD VSS sky130_fd_sc_hd__nor2_1_53/A sky130_fd_sc_hd__dfxtp_1_419/CLK
+ sky130_fd_sc_hd__and2_0_152/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_426 VDD VSS sky130_fd_sc_hd__dfxtp_1_426/Q sky130_fd_sc_hd__dfxtp_1_433/CLK
+ sky130_fd_sc_hd__nand2_1_112/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_437 VDD VSS sky130_fd_sc_hd__dfxtp_1_437/Q sky130_fd_sc_hd__dfxtp_1_452/CLK
+ sky130_fd_sc_hd__nand2_1_90/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_448 VDD VSS sky130_fd_sc_hd__dfxtp_1_994/D sky130_fd_sc_hd__dfxtp_1_448/CLK
+ sky130_fd_sc_hd__nand2_1_68/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_459 VDD VSS sky130_fd_sc_hd__dfxtp_1_459/Q sky130_fd_sc_hd__dfxtp_1_473/CLK
+ sky130_fd_sc_hd__and2_0_236/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2b_1_18 sky130_fd_sc_hd__nand2b_1_18/Y load_en sky130_fd_sc_hd__buf_6_86/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__fa_2_309 sky130_fd_sc_hd__fa_2_303/A sky130_fd_sc_hd__fa_2_306/B
+ sky130_fd_sc_hd__fa_2_309/A sky130_fd_sc_hd__fa_2_309/B sky130_fd_sc_hd__fa_2_309/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_8_14 sky130_fd_sc_hd__clkinv_8_14/Y sky130_fd_sc_hd__clkinv_8_14/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_25 sky130_fd_sc_hd__clkinv_8_26/A sky130_fd_sc_hd__clkinv_8_25/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_25/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_36 sky130_fd_sc_hd__clkinv_8_36/Y sky130_fd_sc_hd__clkinv_8_36/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_36/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_47 sky130_fd_sc_hd__clkinv_8_49/A sky130_fd_sc_hd__clkinv_8_47/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_47/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_58 sky130_fd_sc_hd__clkinv_8_59/A sky130_fd_sc_hd__clkinv_8_58/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_58/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_12 sky130_fd_sc_hd__inv_2_18/Y sky130_fd_sc_hd__buf_12_12/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__clkinv_8_69 sky130_fd_sc_hd__clkinv_8_70/A sky130_fd_sc_hd__clkinv_8_69/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_69/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_23 sky130_fd_sc_hd__buf_12_23/A sky130_fd_sc_hd__buf_12_23/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_34 sky130_fd_sc_hd__buf_8_45/X sky130_fd_sc_hd__buf_12_34/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_45 sky130_fd_sc_hd__buf_8_3/X sky130_fd_sc_hd__buf_12_45/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_56 sky130_fd_sc_hd__buf_8_40/X sky130_fd_sc_hd__buf_12_56/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_67 sky130_fd_sc_hd__buf_4_24/X sky130_fd_sc_hd__buf_12_67/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_78 sky130_fd_sc_hd__buf_4_22/X sky130_fd_sc_hd__buf_12_97/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_89 sky130_fd_sc_hd__buf_12_89/A sky130_fd_sc_hd__buf_12_89/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_2_7 VDD VSS sky130_fd_sc_hd__buf_2_7/X sky130_fd_sc_hd__buf_2_7/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1300 VDD VSS sky130_fd_sc_hd__mux2_2_172/A1 sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__a221oi_1_4/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1311 VDD VSS sky130_fd_sc_hd__fa_2_840/B sky130_fd_sc_hd__dfxtp_1_1326/CLK
+ sky130_fd_sc_hd__o21a_1_64/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1322 VDD VSS sky130_fd_sc_hd__fa_2_906/A sky130_fd_sc_hd__dfxtp_1_1322/CLK
+ sky130_fd_sc_hd__a21oi_1_425/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1333 VDD VSS sky130_fd_sc_hd__or2_0_12/A sky130_fd_sc_hd__clkinv_8_78/Y
+ sky130_fd_sc_hd__nor2b_1_127/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1344 VDD VSS sky130_fd_sc_hd__fa_2_1303/A sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__mux2_2_237/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1355 VDD VSS sky130_fd_sc_hd__fa_2_1277/A sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__mux2_2_261/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1366 VDD VSS sky130_fd_sc_hd__fa_2_1288/A sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__mux2_2_231/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1377 VDD VSS sky130_fd_sc_hd__fa_2_1316/A sky130_fd_sc_hd__clkinv_8_63/Y
+ sky130_fd_sc_hd__mux2_2_262/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1388 VDD VSS sky130_fd_sc_hd__nor2b_2_5/A sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__nor2b_1_132/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_960 VDD VSS sky130_fd_sc_hd__fa_2_1169/A sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__mux2_2_100/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1399 VDD VSS sky130_fd_sc_hd__mux2_2_246/A0 sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__o22ai_1_390/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_971 VDD VSS sky130_fd_sc_hd__mux2_2_117/A0 sky130_fd_sc_hd__clkinv_8_55/Y
+ sky130_fd_sc_hd__nor2_1_160/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_982 VDD VSS sky130_fd_sc_hd__mux2_2_87/A1 sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__o22ai_1_213/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_993 VDD VSS sky130_fd_sc_hd__mux2_2_118/A0 sky130_fd_sc_hd__clkinv_8_64/Y
+ sky130_fd_sc_hd__dfxtp_1_993/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_580 VSS VDD sky130_fd_sc_hd__nand3_1_10/B sky130_fd_sc_hd__a22oi_1_20/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_591 VSS VDD sky130_fd_sc_hd__nand3_1_1/B sky130_fd_sc_hd__a22oi_1_2/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_810 sky130_fd_sc_hd__fa_2_809/B sky130_fd_sc_hd__fa_2_810/SUM
+ sky130_fd_sc_hd__fa_2_810/A sky130_fd_sc_hd__fa_2_810/B sky130_fd_sc_hd__fa_2_810/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_170 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_170/A sky130_fd_sc_hd__nor2_1_91/A
+ sky130_fd_sc_hd__ha_2_170/SUM sky130_fd_sc_hd__ha_2_170/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_821 sky130_fd_sc_hd__fa_2_709/A sky130_fd_sc_hd__fa_2_710/B
+ sky130_fd_sc_hd__fa_2_821/A sky130_fd_sc_hd__fa_2_821/B sky130_fd_sc_hd__fa_2_826/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_181 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_181/A sky130_fd_sc_hd__ha_2_180/A
+ sky130_fd_sc_hd__ha_2_181/SUM sky130_fd_sc_hd__ha_2_181/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_832 sky130_fd_sc_hd__fa_2_705/A sky130_fd_sc_hd__fa_2_706/B
+ sky130_fd_sc_hd__fa_2_832/A sky130_fd_sc_hd__fa_2_832/B sky130_fd_sc_hd__fa_2_832/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_192 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_192/A sky130_fd_sc_hd__ha_2_191/A
+ sky130_fd_sc_hd__ha_2_192/SUM sky130_fd_sc_hd__ha_2_192/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_843 sky130_fd_sc_hd__fa_2_842/CIN sky130_fd_sc_hd__fa_2_843/SUM
+ sky130_fd_sc_hd__fa_2_843/A sky130_fd_sc_hd__fa_2_843/B sky130_fd_sc_hd__fa_2_843/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_854 sky130_fd_sc_hd__fa_2_853/CIN sky130_fd_sc_hd__fa_2_854/SUM
+ sky130_fd_sc_hd__fa_2_854/A sky130_fd_sc_hd__fa_2_854/B sky130_fd_sc_hd__fa_2_854/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_865 sky130_fd_sc_hd__fa_2_864/CIN sky130_fd_sc_hd__fa_2_865/SUM
+ sky130_fd_sc_hd__fa_2_865/A sky130_fd_sc_hd__fa_2_865/B sky130_fd_sc_hd__fa_2_865/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_876 sky130_fd_sc_hd__fa_2_875/CIN sky130_fd_sc_hd__fa_2_876/SUM
+ sky130_fd_sc_hd__fa_2_876/A sky130_fd_sc_hd__fa_2_876/B sky130_fd_sc_hd__fa_2_876/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_887 sky130_fd_sc_hd__fa_2_886/CIN sky130_fd_sc_hd__nand2_1_47/B
+ sky130_fd_sc_hd__ha_2_157/B sky130_fd_sc_hd__fa_2_887/B sky130_fd_sc_hd__o31ai_1_0/A3
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_898 sky130_fd_sc_hd__fa_2_897/CIN sky130_fd_sc_hd__fa_2_898/SUM
+ sky130_fd_sc_hd__fa_2_898/A sky130_fd_sc_hd__fa_2_898/B sky130_fd_sc_hd__fa_2_898/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_7 sky130_fd_sc_hd__inv_2_7/A sky130_fd_sc_hd__inv_2_7/Y VDD
+ VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__nor3_2_9 sky130_fd_sc_hd__nor3_2_9/C sky130_fd_sc_hd__nor3_2_9/Y
+ sky130_fd_sc_hd__nor3_2_9/A sky130_fd_sc_hd__nor3_2_9/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_2
Xsky130_fd_sc_hd__mux2_2_110 VSS VDD sky130_fd_sc_hd__mux2_2_110/A1 sky130_fd_sc_hd__mux2_2_110/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_110/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_17 sky130_fd_sc_hd__nor2_1_17/B sky130_fd_sc_hd__or2_0_4/B
+ sky130_fd_sc_hd__nor3_1_26/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_121 VSS VDD sky130_fd_sc_hd__mux2_2_121/A1 sky130_fd_sc_hd__mux2_2_121/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_121/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_28 sky130_fd_sc_hd__nor4_1_5/B sky130_fd_sc_hd__nor2_1_28/Y
+ sky130_fd_sc_hd__nor3_1_32/C VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_132 VSS VDD sky130_fd_sc_hd__mux2_2_132/A1 sky130_fd_sc_hd__mux2_2_132/A0
+ sky130_fd_sc_hd__mux2_2_135/S sky130_fd_sc_hd__mux2_2_132/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_39 sky130_fd_sc_hd__nor2_1_39/B sky130_fd_sc_hd__nor2_1_39/Y
+ sky130_fd_sc_hd__nor2_1_39/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_143 VSS VDD sky130_fd_sc_hd__mux2_2_143/A1 sky130_fd_sc_hd__mux2_2_143/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_143/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_154 VSS VDD sky130_fd_sc_hd__mux2_2_154/A1 sky130_fd_sc_hd__mux2_2_154/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_154/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_165 VSS VDD sky130_fd_sc_hd__mux2_2_165/A1 sky130_fd_sc_hd__mux2_2_165/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_165/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_176 VSS VDD sky130_fd_sc_hd__mux2_2_176/A1 sky130_fd_sc_hd__mux2_2_176/A0
+ sky130_fd_sc_hd__nor2_8_1/A sky130_fd_sc_hd__mux2_2_176/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_187 VSS VDD sky130_fd_sc_hd__mux2_2_187/A1 sky130_fd_sc_hd__mux2_2_187/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_187/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_198 VSS VDD sky130_fd_sc_hd__mux2_2_198/A1 sky130_fd_sc_hd__mux2_2_198/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_198/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__maj3_1_103 sky130_fd_sc_hd__maj3_1_104/X sky130_fd_sc_hd__maj3_1_103/X
+ sky130_fd_sc_hd__maj3_1_103/B sky130_fd_sc_hd__maj3_1_103/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__and2_0_50 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_50/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_50/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_114 sky130_fd_sc_hd__maj3_1_115/X sky130_fd_sc_hd__maj3_1_114/X
+ sky130_fd_sc_hd__maj3_1_114/B sky130_fd_sc_hd__maj3_1_114/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_330 sky130_fd_sc_hd__nand2_1_462/Y sky130_fd_sc_hd__nand2_1_461/Y
+ sky130_fd_sc_hd__o22ai_1_330/Y sky130_fd_sc_hd__nand2_1_474/B sky130_fd_sc_hd__o21ai_1_388/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_61 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_61/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_61/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_125 sky130_fd_sc_hd__maj3_1_126/X sky130_fd_sc_hd__maj3_1_125/X
+ sky130_fd_sc_hd__maj3_1_125/B sky130_fd_sc_hd__maj3_1_125/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_341 sky130_fd_sc_hd__nand2_1_464/Y sky130_fd_sc_hd__nand2_1_463/Y
+ sky130_fd_sc_hd__o22ai_1_341/Y sky130_fd_sc_hd__nand2_1_473/B sky130_fd_sc_hd__o21ai_1_387/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_72 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_73/A sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__ha_2_74/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_136 sky130_fd_sc_hd__maj3_1_137/X sky130_fd_sc_hd__maj3_1_136/X
+ sky130_fd_sc_hd__maj3_1_136/B sky130_fd_sc_hd__maj3_1_136/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_405 sky130_fd_sc_hd__o21a_1_40/B1 sky130_fd_sc_hd__fa_2_1199/A
+ sky130_fd_sc_hd__o21a_1_40/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_352 sky130_fd_sc_hd__nor2_1_257/A sky130_fd_sc_hd__nor2_1_268/A
+ sky130_fd_sc_hd__o22ai_1_352/Y sky130_fd_sc_hd__a21boi_1_6/Y sky130_fd_sc_hd__a222oi_1_30/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_83 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_83/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__and2_0_83/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_147 sky130_fd_sc_hd__maj3_1_148/X sky130_fd_sc_hd__maj3_1_147/X
+ sky130_fd_sc_hd__maj3_1_147/B sky130_fd_sc_hd__maj3_1_147/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_416 sky130_fd_sc_hd__nand2_1_416/Y sky130_fd_sc_hd__nand2_1_416/B
+ sky130_fd_sc_hd__nor2_8_0/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_363 sky130_fd_sc_hd__nor2_1_234/B sky130_fd_sc_hd__nor2_1_267/A
+ sky130_fd_sc_hd__o22ai_1_363/Y sky130_fd_sc_hd__o22ai_1_376/A1 sky130_fd_sc_hd__a222oi_1_29/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_94 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_94/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_94/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_427 sky130_fd_sc_hd__nand2_1_427/Y sky130_fd_sc_hd__nand2_1_439/B
+ sky130_fd_sc_hd__o21ai_1_359/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_158 sky130_fd_sc_hd__maj3_1_159/X sky130_fd_sc_hd__maj3_1_158/X
+ sky130_fd_sc_hd__maj3_1_158/B sky130_fd_sc_hd__maj3_1_158/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_374 sky130_fd_sc_hd__o32ai_1_8/A3 sky130_fd_sc_hd__o22ai_1_379/B1
+ sky130_fd_sc_hd__o22ai_1_374/Y sky130_fd_sc_hd__nor2_1_236/B sky130_fd_sc_hd__o21a_1_55/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_438 sky130_fd_sc_hd__nand2_1_438/Y sky130_fd_sc_hd__nor2b_2_3/A
+ sky130_fd_sc_hd__xor2_1_208/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_385 sky130_fd_sc_hd__nand2_1_514/Y sky130_fd_sc_hd__nand2_1_513/Y
+ sky130_fd_sc_hd__o22ai_1_385/Y sky130_fd_sc_hd__nand2_1_525/B sky130_fd_sc_hd__o21ai_1_441/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_449 sky130_fd_sc_hd__o21a_1_46/B1 sky130_fd_sc_hd__fa_2_1234/A
+ sky130_fd_sc_hd__o21a_1_46/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_396 sky130_fd_sc_hd__nand2_1_516/Y sky130_fd_sc_hd__nand2_1_515/Y
+ sky130_fd_sc_hd__o22ai_1_396/Y sky130_fd_sc_hd__nand2_1_524/B sky130_fd_sc_hd__o21ai_1_440/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2b_1_18 sky130_fd_sc_hd__ha_2_48/SUM sky130_fd_sc_hd__nor2b_1_18/Y
+ sky130_fd_sc_hd__or2_1_0/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__nor2b_1_29 sky130_fd_sc_hd__ha_2_61/SUM sky130_fd_sc_hd__nor2b_1_29/Y
+ sky130_fd_sc_hd__or2_0_2/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1007 sky130_fd_sc_hd__o21ai_1_425/B1 sky130_fd_sc_hd__nor2_1_262/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1007/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1018 sky130_fd_sc_hd__nor2_1_236/B sky130_fd_sc_hd__fa_2_1255/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1018/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_60 sky130_fd_sc_hd__buf_8_60/A sky130_fd_sc_hd__buf_8_60/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__clkinv_1_1029 sky130_fd_sc_hd__nor2_1_308/A sky130_fd_sc_hd__fa_2_1309/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1029/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_71 sky130_fd_sc_hd__inv_2_62/Y sky130_fd_sc_hd__buf_8_71/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_82 sky130_fd_sc_hd__inv_2_55/Y sky130_fd_sc_hd__buf_8_82/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_201 VDD VSS sky130_fd_sc_hd__ha_2_79/B sky130_fd_sc_hd__dfxtp_1_212/CLK
+ sky130_fd_sc_hd__and2_0_84/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_8_93 sky130_fd_sc_hd__buf_8_93/A sky130_fd_sc_hd__buf_8_93/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_212 VDD VSS sky130_fd_sc_hd__xor2_1_7/B sky130_fd_sc_hd__dfxtp_1_212/CLK
+ sky130_fd_sc_hd__and2_0_80/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_223 VDD VSS sky130_fd_sc_hd__ha_2_80/A sky130_fd_sc_hd__dfxtp_1_223/CLK
+ sky130_fd_sc_hd__nor2b_1_40/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_234 VDD VSS sky130_fd_sc_hd__fa_2_875/A sky130_fd_sc_hd__dfxtp_1_462/CLK
+ sky130_fd_sc_hd__and2_0_166/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_245 VDD VSS sky130_fd_sc_hd__fa_2_864/A sky130_fd_sc_hd__dfxtp_1_266/CLK
+ sky130_fd_sc_hd__and2_0_177/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_256 VDD VSS sky130_fd_sc_hd__dfxtp_1_256/Q sky130_fd_sc_hd__dfxtp_1_262/CLK
+ sky130_fd_sc_hd__and2_0_219/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_267 VDD VSS sky130_fd_sc_hd__dfxtp_1_267/Q sky130_fd_sc_hd__dfxtp_1_277/CLK
+ sky130_fd_sc_hd__and2_0_228/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_278 VDD VSS sky130_fd_sc_hd__xor2_1_14/B sky130_fd_sc_hd__dfxtp_1_463/CLK
+ sky130_fd_sc_hd__and2_0_206/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_289 VDD VSS sky130_fd_sc_hd__a22o_1_58/A1 sky130_fd_sc_hd__clkinv_4_31/Y
+ sky130_fd_sc_hd__nand2_1_131/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o22ai_1_9 sky130_fd_sc_hd__fa_2_9/A sky130_fd_sc_hd__fa_2_76/A sky130_fd_sc_hd__fa_2_126/A
+ sky130_fd_sc_hd__ha_2_91/A sky130_fd_sc_hd__fa_2_2/A VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_106 sky130_fd_sc_hd__fa_2_14/CIN sky130_fd_sc_hd__fa_2_99/B
+ sky130_fd_sc_hd__fa_2_5/A sky130_fd_sc_hd__ha_2_91/B sky130_fd_sc_hd__fa_2_2/B VSS
+ VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_117 sky130_fd_sc_hd__maj3_1_5/B sky130_fd_sc_hd__maj3_1_6/A
+ sky130_fd_sc_hd__fa_2_117/A sky130_fd_sc_hd__fa_2_117/B sky130_fd_sc_hd__fa_2_118/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_128 sky130_fd_sc_hd__fa_2_127/A sky130_fd_sc_hd__fa_2_122/B
+ sky130_fd_sc_hd__ha_2_97/B sky130_fd_sc_hd__ha_2_97/A sky130_fd_sc_hd__fa_2_76/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_139 sky130_fd_sc_hd__fa_2_141/CIN sky130_fd_sc_hd__fa_2_133/A
+ sky130_fd_sc_hd__fa_2_45/A sky130_fd_sc_hd__fa_2_139/B sky130_fd_sc_hd__fa_2_9/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_101 VDD VSS sky130_fd_sc_hd__buf_2_101/X sky130_fd_sc_hd__buf_2_101/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__fa_2_1300 sky130_fd_sc_hd__fa_2_1301/CIN sky130_fd_sc_hd__mux2_2_245/A1
+ sky130_fd_sc_hd__fa_2_1300/A sky130_fd_sc_hd__fa_2_1300/B sky130_fd_sc_hd__fa_2_1300/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_112 VDD VSS sky130_fd_sc_hd__buf_2_112/X sky130_fd_sc_hd__buf_2_112/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__fa_2_1311 sky130_fd_sc_hd__fa_2_1312/CIN sky130_fd_sc_hd__mux2_2_267/A1
+ sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1311/B sky130_fd_sc_hd__nor2_8_2/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_123 VDD VSS sky130_fd_sc_hd__buf_2_123/X sky130_fd_sc_hd__buf_2_123/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_16 sky130_fd_sc_hd__ha_2_91/B sky130_fd_sc_hd__fa_2_261/A
+ sky130_fd_sc_hd__fa_2_232/A sky130_fd_sc_hd__fa_2_5/A sky130_fd_sc_hd__fa_2_258/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_1322 sky130_fd_sc_hd__fa_2_1323/CIN sky130_fd_sc_hd__mux2_2_244/A1
+ sky130_fd_sc_hd__fa_2_1322/A sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1322/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_134 VDD VSS sky130_fd_sc_hd__buf_2_134/X sky130_fd_sc_hd__buf_8_133/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_27 sky130_fd_sc_hd__fa_2_404/A sky130_fd_sc_hd__fa_2_286/B
+ sky130_fd_sc_hd__o22ai_1_27/Y sky130_fd_sc_hd__ha_2_116/A sky130_fd_sc_hd__fa_2_424/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_145 VDD VSS sky130_fd_sc_hd__buf_2_145/X sky130_fd_sc_hd__buf_6_88/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_38 sky130_fd_sc_hd__fa_2_531/B sky130_fd_sc_hd__fa_2_554/A
+ sky130_fd_sc_hd__fa_2_553/B sky130_fd_sc_hd__ha_2_117/B sky130_fd_sc_hd__ha_2_124/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_156 VDD VSS sky130_fd_sc_hd__buf_4_105/A sky130_fd_sc_hd__buf_2_156/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_49 sky130_fd_sc_hd__fa_2_829/A sky130_fd_sc_hd__ha_2_140/A
+ sky130_fd_sc_hd__fa_2_741/A sky130_fd_sc_hd__fa_2_807/B sky130_fd_sc_hd__ha_2_145/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_167 VDD VSS sky130_fd_sc_hd__buf_2_167/X sky130_fd_sc_hd__nor3_1_20/Y
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_178 VDD VSS sky130_fd_sc_hd__buf_2_178/X sky130_fd_sc_hd__buf_2_178/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1130 VDD VSS sky130_fd_sc_hd__mux2_2_170/A0 sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__dfxtp_1_989/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_2_189 VDD VSS sky130_fd_sc_hd__buf_2_189/X sky130_fd_sc_hd__buf_2_189/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1141 VDD VSS sky130_fd_sc_hd__mux2_2_145/A0 sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__dfxtp_1_454/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1152 VDD VSS sky130_fd_sc_hd__mux2_2_138/A0 sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__o22ai_1_285/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1163 VDD VSS sky130_fd_sc_hd__fa_2_861/B sky130_fd_sc_hd__dfxtp_1_1180/CLK
+ sky130_fd_sc_hd__o21a_1_54/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1174 VDD VSS sky130_fd_sc_hd__fa_2_850/B sky130_fd_sc_hd__dfxtp_1_1180/CLK
+ sky130_fd_sc_hd__o21a_1_49/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1185 VDD VSS sky130_fd_sc_hd__fa_2_938/A sky130_fd_sc_hd__clkinv_4_24/Y
+ sky130_fd_sc_hd__a21oi_1_363/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1196 VDD VSS sky130_fd_sc_hd__fa_2_1245/A sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__mux2_2_209/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__ha_2_1 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_1/A sky130_fd_sc_hd__ha_2_0/B
+ sky130_fd_sc_hd__ha_2_1/SUM sky130_fd_sc_hd__ha_2_1/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__buf_4_18 VDD VSS sky130_fd_sc_hd__buf_6_17/A sky130_fd_sc_hd__buf_8_37/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_29 VDD VSS sky130_fd_sc_hd__buf_4_29/X sky130_fd_sc_hd__buf_8_17/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__dfxtp_1_790 VDD VSS sky130_fd_sc_hd__fa_2_1089/A sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__mux2_2_44/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_12 VSS VDD sky130_fd_sc_hd__clkbuf_4_5/A sky130_fd_sc_hd__clkbuf_4_4/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_23 VSS VDD sky130_fd_sc_hd__clkbuf_1_23/X sky130_fd_sc_hd__clkbuf_1_23/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_34 VSS VDD sky130_fd_sc_hd__clkbuf_1_34/X sky130_fd_sc_hd__clkbuf_1_34/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_640 sky130_fd_sc_hd__fa_2_639/A sky130_fd_sc_hd__fa_2_640/SUM
+ sky130_fd_sc_hd__fa_2_686/B sky130_fd_sc_hd__ha_2_134/A sky130_fd_sc_hd__ha_2_130/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_45 VSS VDD sky130_fd_sc_hd__clkbuf_1_45/X sky130_fd_sc_hd__clkbuf_1_45/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_651 sky130_fd_sc_hd__fa_2_650/A sky130_fd_sc_hd__fa_2_651/SUM
+ sky130_fd_sc_hd__ha_2_135/B sky130_fd_sc_hd__fa_2_659/A sky130_fd_sc_hd__ha_2_130/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_56 VSS VDD sky130_fd_sc_hd__clkbuf_1_56/X sky130_fd_sc_hd__clkbuf_1_56/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_662 sky130_fd_sc_hd__fa_2_661/B sky130_fd_sc_hd__fa_2_662/SUM
+ sky130_fd_sc_hd__fa_2_662/A sky130_fd_sc_hd__fa_2_662/B sky130_fd_sc_hd__fa_2_662/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_67 VSS VDD sky130_fd_sc_hd__clkbuf_1_67/X sky130_fd_sc_hd__clkbuf_1_67/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_673 sky130_fd_sc_hd__fa_2_674/B sky130_fd_sc_hd__fa_2_666/A
+ sky130_fd_sc_hd__fa_2_700/A sky130_fd_sc_hd__fa_2_673/B sky130_fd_sc_hd__fa_2_701/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_78 VSS VDD sky130_fd_sc_hd__nand4_1_9/A sky130_fd_sc_hd__a22oi_2_10/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_684 sky130_fd_sc_hd__fa_2_576/A sky130_fd_sc_hd__fa_2_577/B
+ sky130_fd_sc_hd__fa_2_684/A sky130_fd_sc_hd__fa_2_684/B sky130_fd_sc_hd__fa_2_688/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_89 VSS VDD sky130_fd_sc_hd__clkbuf_1_89/X sky130_fd_sc_hd__buf_2_25/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__and2_4_0 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__ha_2_59/B
+ sky130_fd_sc_hd__nor2_4_2/Y VSS VDD VSS VDD sky130_fd_sc_hd__and2_4
Xsky130_fd_sc_hd__fa_2_695 sky130_fd_sc_hd__fa_2_694/CIN sky130_fd_sc_hd__fa_2_695/SUM
+ sky130_fd_sc_hd__fa_2_695/A sky130_fd_sc_hd__fa_2_698/A sky130_fd_sc_hd__ha_2_134/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a21oi_1_208 sky130_fd_sc_hd__fa_2_1052/A sky130_fd_sc_hd__o22ai_1_180/Y
+ sky130_fd_sc_hd__a21oi_1_208/Y sky130_fd_sc_hd__nor2_4_12/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_219 sky130_fd_sc_hd__clkinv_1_731/Y sky130_fd_sc_hd__o22ai_1_196/Y
+ sky130_fd_sc_hd__a21oi_1_219/Y sky130_fd_sc_hd__nand2_1_331/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_2_15 sky130_fd_sc_hd__nor3_2_7/Y sky130_fd_sc_hd__a22oi_2_15/A2
+ sky130_fd_sc_hd__nor3_2_8/Y sky130_fd_sc_hd__a22oi_2_15/B2 sky130_fd_sc_hd__nand4_1_50/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__a22oi_2_26 sky130_fd_sc_hd__buf_2_165/X sky130_fd_sc_hd__a22oi_2_26/A2
+ sky130_fd_sc_hd__nor2_4_7/Y sky130_fd_sc_hd__a22oi_2_26/B2 sky130_fd_sc_hd__nand4_1_58/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__buf_12_1 sky130_fd_sc_hd__inv_2_22/Y sky130_fd_sc_hd__buf_12_1/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__nand2_1_202 sky130_fd_sc_hd__nor2_1_21/B sky130_fd_sc_hd__nand2_1_202/B
+ sky130_fd_sc_hd__nor2_1_22/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_801 sky130_fd_sc_hd__o22ai_1_230/A1 sky130_fd_sc_hd__a21o_2_9/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_801/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_213 sky130_fd_sc_hd__nor2_1_30/B sky130_fd_sc_hd__nand2_1_213/B
+ sky130_fd_sc_hd__nor2_1_31/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_160 sky130_fd_sc_hd__nand2_1_338/A sky130_fd_sc_hd__nand2_1_284/Y
+ sky130_fd_sc_hd__o22ai_1_160/Y sky130_fd_sc_hd__xnor2_1_84/Y sky130_fd_sc_hd__o22ai_1_160/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_812 sky130_fd_sc_hd__o31ai_1_6/A3 sky130_fd_sc_hd__xnor2_1_3/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_812/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_224 sky130_fd_sc_hd__a31oi_1_2/A2 sky130_fd_sc_hd__o22ai_1_60/B2
+ sky130_fd_sc_hd__fa_2_965/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_823 sky130_fd_sc_hd__o21ai_1_304/A2 sky130_fd_sc_hd__fa_2_1136/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_823/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_171 sky130_fd_sc_hd__a21oi_1_200/Y sky130_fd_sc_hd__a21oi_1_199/Y
+ sky130_fd_sc_hd__o22ai_1_171/Y sky130_fd_sc_hd__nor2_2_13/B sky130_fd_sc_hd__nor2_1_126/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_235 sky130_fd_sc_hd__xnor2_1_56/B sky130_fd_sc_hd__o21ai_1_75/B1
+ sky130_fd_sc_hd__o21ai_1_82/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_182 sky130_fd_sc_hd__o21a_1_16/A2 sky130_fd_sc_hd__nor2_1_116/B
+ sky130_fd_sc_hd__nor2_1_131/B sky130_fd_sc_hd__o22ai_1_191/A1 sky130_fd_sc_hd__o22ai_1_206/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_834 sky130_fd_sc_hd__nor2_1_145/B sky130_fd_sc_hd__fa_2_1131/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_834/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_246 sky130_fd_sc_hd__nand2_1_246/Y sky130_fd_sc_hd__nor2_1_53/B
+ sky130_fd_sc_hd__nor2_1_53/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_193 sky130_fd_sc_hd__o22ai_1_206/B1 sky130_fd_sc_hd__nor2_1_117/B
+ sky130_fd_sc_hd__o22ai_1_193/Y sky130_fd_sc_hd__o22ai_1_193/A1 sky130_fd_sc_hd__o22ai_1_206/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_845 sky130_fd_sc_hd__o22ai_1_262/A1 sky130_fd_sc_hd__nor2_1_182/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_845/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_257 sky130_fd_sc_hd__o21a_1_7/B1 sky130_fd_sc_hd__fa_2_977/A
+ sky130_fd_sc_hd__o21a_1_7/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand4_1_30 sky130_fd_sc_hd__nand4_1_30/C sky130_fd_sc_hd__nand4_1_30/B
+ sky130_fd_sc_hd__nand4_1_30/Y sky130_fd_sc_hd__nand4_1_30/D sky130_fd_sc_hd__buf_2_101/X
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__clkinv_1_856 sky130_fd_sc_hd__nor2_1_153/B sky130_fd_sc_hd__fa_2_1149/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_856/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_268 sky130_fd_sc_hd__nand3_1_49/A sky130_fd_sc_hd__fa_2_988/A
+ sky130_fd_sc_hd__a21o_2_3/A2 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand4_1_41 sky130_fd_sc_hd__nand4_1_41/C sky130_fd_sc_hd__nand4_1_41/B
+ sky130_fd_sc_hd__buf_2_289/A sky130_fd_sc_hd__nand4_1_41/D sky130_fd_sc_hd__nand4_1_41/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__clkinv_1_867 sky130_fd_sc_hd__nor2_1_214/A sky130_fd_sc_hd__nor2b_1_112/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_867/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_279 sky130_fd_sc_hd__nor2_1_76/A sky130_fd_sc_hd__nand2_1_282/B
+ sky130_fd_sc_hd__nand2_2_4/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_878 sky130_fd_sc_hd__o31ai_1_8/B1 sky130_fd_sc_hd__a21oi_1_322/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_878/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand4_1_52 sky130_fd_sc_hd__nand4_1_52/C sky130_fd_sc_hd__nand4_1_52/B
+ sky130_fd_sc_hd__buf_2_269/A sky130_fd_sc_hd__nand4_1_52/D sky130_fd_sc_hd__nand4_1_52/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__clkinv_1_889 sky130_fd_sc_hd__o32ai_1_4/B2 sky130_fd_sc_hd__fa_2_1193/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_889/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand4_1_63 sky130_fd_sc_hd__nand4_1_63/C sky130_fd_sc_hd__nand4_1_63/B
+ sky130_fd_sc_hd__nand4_1_63/Y sky130_fd_sc_hd__nand4_1_63/D sky130_fd_sc_hd__nand4_1_63/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_74 sky130_fd_sc_hd__nand4_1_74/C sky130_fd_sc_hd__nand4_1_74/B
+ sky130_fd_sc_hd__nand2_1_5/B sky130_fd_sc_hd__nand4_1_74/D sky130_fd_sc_hd__nand4_1_74/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_85 sky130_fd_sc_hd__nand4_1_85/C sky130_fd_sc_hd__nand4_1_85/B
+ sky130_fd_sc_hd__nand4_1_85/Y sky130_fd_sc_hd__nand4_1_85/D sky130_fd_sc_hd__nand4_1_85/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__conb_1_12 sky130_fd_sc_hd__conb_1_12/LO sky130_fd_sc_hd__conb_1_12/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_23 sky130_fd_sc_hd__conb_1_23/LO sky130_fd_sc_hd__conb_1_23/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__mux2_2_7 VSS VDD sky130_fd_sc_hd__mux2_2_7/A1 sky130_fd_sc_hd__mux2_2_7/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_7/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1130 sky130_fd_sc_hd__fa_2_1131/CIN sky130_fd_sc_hd__mux2_2_99/A1
+ sky130_fd_sc_hd__fa_2_1130/A sky130_fd_sc_hd__fa_2_1130/B sky130_fd_sc_hd__fa_2_1130/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1141 sky130_fd_sc_hd__fa_2_1142/CIN sky130_fd_sc_hd__and2_0_322/A
+ sky130_fd_sc_hd__fa_2_1141/A sky130_fd_sc_hd__fa_2_1141/B sky130_fd_sc_hd__fa_2_1141/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1152 sky130_fd_sc_hd__fa_2_1153/CIN sky130_fd_sc_hd__mux2_2_88/A1
+ sky130_fd_sc_hd__fa_2_1152/A sky130_fd_sc_hd__fa_2_1152/B sky130_fd_sc_hd__fa_2_1152/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1163 sky130_fd_sc_hd__fa_2_1164/CIN sky130_fd_sc_hd__mux2_2_118/A1
+ sky130_fd_sc_hd__fa_2_1163/A sky130_fd_sc_hd__fa_2_1172/B sky130_fd_sc_hd__fa_2_1163/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1174 sky130_fd_sc_hd__fa_2_1175/CIN sky130_fd_sc_hd__and2_0_327/A
+ sky130_fd_sc_hd__fa_2_1174/A sky130_fd_sc_hd__fa_2_1174/B sky130_fd_sc_hd__fa_2_1174/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1185 sky130_fd_sc_hd__fa_2_1186/CIN sky130_fd_sc_hd__mux2_2_137/A1
+ sky130_fd_sc_hd__fa_2_1185/A sky130_fd_sc_hd__fa_2_1185/B sky130_fd_sc_hd__fa_2_1185/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1196 sky130_fd_sc_hd__fa_2_1197/CIN sky130_fd_sc_hd__mux2_2_155/A1
+ sky130_fd_sc_hd__fa_2_1196/A sky130_fd_sc_hd__fa_2_1196/B sky130_fd_sc_hd__fa_2_1196/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o2bb2ai_1_3 sky130_fd_sc_hd__o2bb2ai_1_3/Y sky130_fd_sc_hd__nor2_1_18/Y
+ sky130_fd_sc_hd__ha_2_149/SUM sky130_fd_sc_hd__o21ai_1_31/A1 sky130_fd_sc_hd__maj3_1_1/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_470 sky130_fd_sc_hd__fa_2_471/A sky130_fd_sc_hd__fa_2_470/SUM
+ sky130_fd_sc_hd__ha_2_123/B sky130_fd_sc_hd__ha_2_122/B sky130_fd_sc_hd__fa_2_559/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_481 sky130_fd_sc_hd__fa_2_483/B sky130_fd_sc_hd__fa_2_479/A
+ sky130_fd_sc_hd__fa_2_546/A sky130_fd_sc_hd__ha_2_125/B sky130_fd_sc_hd__fa_2_564/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_492 sky130_fd_sc_hd__fa_2_491/A sky130_fd_sc_hd__fa_2_486/B
+ sky130_fd_sc_hd__ha_2_118/B sky130_fd_sc_hd__ha_2_125/A sky130_fd_sc_hd__fa_2_543/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_1_108 sky130_fd_sc_hd__inv_2_70/A sky130_fd_sc_hd__buf_8_68/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_108/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_119 sky130_fd_sc_hd__ha_2_47/A sky130_fd_sc_hd__clkinv_1_119/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_119/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_8 VSS VDD sky130_fd_sc_hd__nor4_1_2/A sky130_fd_sc_hd__o21ai_1_8/A1
+ sky130_fd_sc_hd__a21oi_1_5/Y sky130_fd_sc_hd__o21ai_1_8/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_1_202 sky130_fd_sc_hd__nor2_1_205/A sky130_fd_sc_hd__nor2_1_202/Y
+ sky130_fd_sc_hd__o31ai_1_8/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_213 sky130_fd_sc_hd__or3_1_3/X sky130_fd_sc_hd__nor2_1_213/Y
+ sky130_fd_sc_hd__nor2_1_213/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_224 sky130_fd_sc_hd__o21a_1_42/A1 sky130_fd_sc_hd__nor2_1_224/Y
+ sky130_fd_sc_hd__nor2_1_224/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_235 sky130_fd_sc_hd__nor2_1_235/B sky130_fd_sc_hd__o21a_1_49/A1
+ sky130_fd_sc_hd__o21a_1_50/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_246 sky130_fd_sc_hd__nor2_1_246/B sky130_fd_sc_hd__nor2_1_246/Y
+ sky130_fd_sc_hd__nor2_1_248/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_257 sky130_fd_sc_hd__nor2_1_257/B sky130_fd_sc_hd__nor2_1_257/Y
+ sky130_fd_sc_hd__nor2_1_257/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_268 sky130_fd_sc_hd__nor2_1_268/B sky130_fd_sc_hd__nor2_1_268/Y
+ sky130_fd_sc_hd__nor2_1_268/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_279 sky130_fd_sc_hd__o21a_1_68/A2 sky130_fd_sc_hd__o21a_1_64/A1
+ sky130_fd_sc_hd__o21a_1_65/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_420 sky130_fd_sc_hd__buf_8_183/X sky130_fd_sc_hd__buf_12_420/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_431 sky130_fd_sc_hd__buf_8_207/X sky130_fd_sc_hd__buf_12_495/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_442 sky130_fd_sc_hd__buf_4_115/X sky130_fd_sc_hd__buf_12_442/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_301 sky130_fd_sc_hd__clkbuf_4_165/X sky130_fd_sc_hd__clkinv_2_23/Y
+ sky130_fd_sc_hd__clkbuf_1_402/X sky130_fd_sc_hd__a22oi_1_301/A2 sky130_fd_sc_hd__a22oi_1_301/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_453 sky130_fd_sc_hd__buf_6_75/X sky130_fd_sc_hd__buf_12_476/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_312 sky130_fd_sc_hd__clkbuf_1_376/X sky130_fd_sc_hd__nor2_2_5/Y
+ sky130_fd_sc_hd__clkbuf_1_427/X sky130_fd_sc_hd__clkbuf_1_460/X sky130_fd_sc_hd__nand4_1_77/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_464 sky130_fd_sc_hd__buf_6_74/X sky130_fd_sc_hd__buf_12_492/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_323 sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_2_7/Y
+ sky130_fd_sc_hd__fa_2_995/A sky130_fd_sc_hd__fa_2_996/A sky130_fd_sc_hd__o21ai_1_91/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_475 sky130_fd_sc_hd__buf_12_475/A sky130_fd_sc_hd__buf_12_475/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_334 sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_2_8/Y
+ sky130_fd_sc_hd__fa_2_1011/A sky130_fd_sc_hd__fa_2_1014/A sky130_fd_sc_hd__a22oi_1_334/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_486 sky130_fd_sc_hd__buf_12_486/A sky130_fd_sc_hd__buf_12_486/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_345 sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_2_7/Y
+ sky130_fd_sc_hd__fa_2_997/A sky130_fd_sc_hd__fa_2_998/A sky130_fd_sc_hd__a22oi_1_345/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_497 sky130_fd_sc_hd__buf_12_497/A sky130_fd_sc_hd__buf_12_497/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_356 sky130_fd_sc_hd__clkinv_1_622/Y sky130_fd_sc_hd__o21ai_1_236/Y
+ sky130_fd_sc_hd__nand2_1_321/A sky130_fd_sc_hd__a211o_1_9/A1 sky130_fd_sc_hd__a22oi_1_356/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_367 sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__nor2_4_13/Y
+ sky130_fd_sc_hd__fa_2_1078/A sky130_fd_sc_hd__fa_2_1079/A sky130_fd_sc_hd__a22oi_1_367/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_378 sky130_fd_sc_hd__nor2_1_180/Y sky130_fd_sc_hd__nor2_1_182/Y
+ sky130_fd_sc_hd__fa_2_1148/A sky130_fd_sc_hd__fa_2_1144/A sky130_fd_sc_hd__a22oi_1_378/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_620 sky130_fd_sc_hd__o22ai_1_197/A2 sky130_fd_sc_hd__fa_2_1080/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_620/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22oi_1_389 sky130_fd_sc_hd__nor2_1_265/Y sky130_fd_sc_hd__nor2_1_267/Y
+ sky130_fd_sc_hd__fa_2_1233/A sky130_fd_sc_hd__fa_2_1229/A sky130_fd_sc_hd__a22oi_1_389/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_631 sky130_fd_sc_hd__o22ai_1_149/B2 sky130_fd_sc_hd__ha_2_200/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_631/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_642 sky130_fd_sc_hd__o22ai_1_160/B2 sky130_fd_sc_hd__ha_2_189/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_642/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_653 sky130_fd_sc_hd__nand2_1_290/B sky130_fd_sc_hd__nor2_1_109/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_653/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_664 sky130_fd_sc_hd__o21ai_1_197/A1 sky130_fd_sc_hd__nand2_1_299/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_664/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_675 sky130_fd_sc_hd__nor2_1_105/B sky130_fd_sc_hd__fa_2_1107/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_675/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_686 sky130_fd_sc_hd__nor2_1_111/B sky130_fd_sc_hd__fa_2_1118/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_686/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_697 sky130_fd_sc_hd__nand2_1_319/A sky130_fd_sc_hd__a222oi_1_2/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_697/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand3_1_4 sky130_fd_sc_hd__nand3_1_4/Y sky130_fd_sc_hd__nand3_1_4/A
+ sky130_fd_sc_hd__nand3_1_4/C sky130_fd_sc_hd__nand3_1_4/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__a222oi_1_40 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1310/A sky130_fd_sc_hd__nor2_2_18/Y
+ sky130_fd_sc_hd__nor3_1_41/A sky130_fd_sc_hd__xor2_1_298/A sky130_fd_sc_hd__nor2_4_19/B
+ sky130_fd_sc_hd__a222oi_1_40/Y sky130_fd_sc_hd__fa_2_1309/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_20 VSS VDD sky130_fd_sc_hd__nor2_1_23/B sky130_fd_sc_hd__xor2_1_18/B
+ sky130_fd_sc_hd__nor2_1_23/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_31 VSS VDD sky130_fd_sc_hd__nor2_1_33/B sky130_fd_sc_hd__xnor2_1_31/Y
+ sky130_fd_sc_hd__nor4_1_8/D VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_42 VSS VDD sky130_fd_sc_hd__xnor2_1_42/B sky130_fd_sc_hd__xnor2_1_42/Y
+ sky130_fd_sc_hd__nor2_1_44/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_53 VSS VDD sky130_fd_sc_hd__xnor2_1_53/B sky130_fd_sc_hd__xnor2_1_53/Y
+ sky130_fd_sc_hd__nor2_1_47/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_64 VSS VDD sky130_fd_sc_hd__xnor2_1_65/B sky130_fd_sc_hd__xnor2_1_64/Y
+ sky130_fd_sc_hd__xnor2_1_64/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_75 VSS VDD sky130_fd_sc_hd__xnor2_1_75/B sky130_fd_sc_hd__xnor2_1_75/Y
+ sky130_fd_sc_hd__nor2_1_95/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_86 VSS VDD sky130_fd_sc_hd__xnor2_1_86/B sky130_fd_sc_hd__xnor2_1_86/Y
+ sky130_fd_sc_hd__nor2_1_98/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_97 VSS VDD sky130_fd_sc_hd__xnor2_1_97/B sky130_fd_sc_hd__xnor2_1_97/Y
+ sky130_fd_sc_hd__fa_2_1241/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__a211oi_1_0 sky130_fd_sc_hd__nor2_1_8/A sky130_fd_sc_hd__nor2_1_8/Y
+ sky130_fd_sc_hd__nor2_1_23/A sky130_fd_sc_hd__a21oi_1_9/B1 sky130_fd_sc_hd__or4_1_1/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__clkbuf_1_409 VSS VDD sky130_fd_sc_hd__clkbuf_1_409/X sky130_fd_sc_hd__clkbuf_1_409/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o32ai_1_3 sky130_fd_sc_hd__o32ai_1_3/A2 sky130_fd_sc_hd__o32ai_1_3/Y
+ sky130_fd_sc_hd__fa_2_1175/A sky130_fd_sc_hd__o32ai_1_3/A3 sky130_fd_sc_hd__o32ai_1_3/B2
+ sky130_fd_sc_hd__fa_2_1174/A VDD VSS VSS VDD sky130_fd_sc_hd__o32ai_1
Xsky130_fd_sc_hd__clkbuf_16_1 sky130_fd_sc_hd__buf_12_112/A sky130_fd_sc_hd__buf_8_12/X
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__a22oi_1_0 sky130_fd_sc_hd__nor2_2_0/Y sky130_fd_sc_hd__clkinv_1_4/Y
+ sky130_fd_sc_hd__nand4_1_31/Y sky130_fd_sc_hd__nand4_1_15/Y sky130_fd_sc_hd__a22oi_1_0/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor4_1_1 sky130_fd_sc_hd__nor4_1_1/D sky130_fd_sc_hd__nor4_1_1/C
+ sky130_fd_sc_hd__nor4_1_1/Y sky130_fd_sc_hd__nor4_1_1/A sky130_fd_sc_hd__nor4_1_1/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__nor4_1
Xsky130_fd_sc_hd__diode_2_150 sky130_fd_sc_hd__buf_2_195/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_161 sky130_fd_sc_hd__nand4_1_73/D VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_172 sky130_fd_sc_hd__clkbuf_4_179/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_183 sky130_fd_sc_hd__dfxtp_1_92/D VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_194 sky130_fd_sc_hd__clkbuf_4_207/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkinv_2_16 sky130_fd_sc_hd__inv_2_83/A sky130_fd_sc_hd__a22o_1_14/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_16/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkbuf_4_203 sky130_fd_sc_hd__clkbuf_4_203/X sky130_fd_sc_hd__buf_8_185/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_214 sky130_fd_sc_hd__buf_6_50/A sky130_fd_sc_hd__dfxtp_1_1463/Q
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_2_27 sky130_fd_sc_hd__nand4_1_70/D sky130_fd_sc_hd__clkinv_2_27/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_27/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_2_38 sky130_fd_sc_hd__clkinv_4_27/A sky130_fd_sc_hd__clkinv_2_38/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_38/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkbuf_4_225 sky130_fd_sc_hd__nor2_1_2/A sky130_fd_sc_hd__dfxtp_1_282/Q
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_2_49 sky130_fd_sc_hd__clkinv_4_74/A sky130_fd_sc_hd__clkinv_4_73/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_49/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__buf_12_250 sky130_fd_sc_hd__buf_12_250/A sky130_fd_sc_hd__buf_12_250/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_261 sky130_fd_sc_hd__buf_12_261/A sky130_fd_sc_hd__buf_12_261/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_120 sky130_fd_sc_hd__a22oi_1_96/B1 sky130_fd_sc_hd__a22oi_1_96/A1
+ sky130_fd_sc_hd__clkbuf_1_145/X sky130_fd_sc_hd__a22oi_1_120/A2 sky130_fd_sc_hd__nand4_1_25/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_272 sky130_fd_sc_hd__inv_2_87/Y sky130_fd_sc_hd__buf_12_272/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_131 sky130_fd_sc_hd__a22oi_1_96/B1 sky130_fd_sc_hd__a22oi_1_96/A1
+ sky130_fd_sc_hd__clkbuf_1_142/X sky130_fd_sc_hd__a22oi_1_131/A2 sky130_fd_sc_hd__nand4_1_28/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_283 sky130_fd_sc_hd__inv_2_97/Y sky130_fd_sc_hd__buf_12_362/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_142 sky130_fd_sc_hd__clkbuf_4_72/X sky130_fd_sc_hd__clkbuf_4_73/X
+ sky130_fd_sc_hd__a22oi_1_142/B2 sky130_fd_sc_hd__buf_2_83/X sky130_fd_sc_hd__buf_2_101/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_294 sky130_fd_sc_hd__buf_8_144/X sky130_fd_sc_hd__buf_12_294/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_153 sky130_fd_sc_hd__clkbuf_4_111/X sky130_fd_sc_hd__clkbuf_4_112/X
+ sky130_fd_sc_hd__a22oi_1_153/B2 sky130_fd_sc_hd__clkbuf_1_296/X sky130_fd_sc_hd__a22oi_1_153/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_164 sky130_fd_sc_hd__clkbuf_1_351/X sky130_fd_sc_hd__clkbuf_1_353/X
+ sky130_fd_sc_hd__clkinv_2_13/Y sky130_fd_sc_hd__a22oi_1_164/A2 sky130_fd_sc_hd__nand4_1_36/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_175 sky130_fd_sc_hd__clkbuf_1_265/X sky130_fd_sc_hd__clkbuf_1_266/X
+ sky130_fd_sc_hd__clkbuf_1_275/X sky130_fd_sc_hd__a22oi_1_175/A2 sky130_fd_sc_hd__a22oi_1_175/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_186 sky130_fd_sc_hd__clkbuf_1_264/X sky130_fd_sc_hd__nor2_2_3/Y
+ sky130_fd_sc_hd__a22oi_1_186/B2 sky130_fd_sc_hd__clkbuf_4_128/X sky130_fd_sc_hd__nand4_1_41/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_197 sky130_fd_sc_hd__clkbuf_4_111/X sky130_fd_sc_hd__clkbuf_4_112/X
+ sky130_fd_sc_hd__a22oi_1_197/B2 sky130_fd_sc_hd__clkbuf_1_285/X sky130_fd_sc_hd__a22oi_1_197/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_450 sky130_fd_sc_hd__fa_2_951/B sky130_fd_sc_hd__nor2b_1_86/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_450/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_461 sky130_fd_sc_hd__clkinv_1_461/Y sky130_fd_sc_hd__a21oi_1_128/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_461/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_472 sky130_fd_sc_hd__nand2_1_264/A sky130_fd_sc_hd__nor2_2_9/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_472/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_483 sky130_fd_sc_hd__o22ai_1_88/B2 sky130_fd_sc_hd__ha_2_171/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_483/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_494 sky130_fd_sc_hd__o21ai_1_78/B1 sky130_fd_sc_hd__nor2_1_58/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_494/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_408 VSS VDD sky130_fd_sc_hd__o22ai_1_379/A2 sky130_fd_sc_hd__nor2_1_261/A
+ sky130_fd_sc_hd__a22oi_1_390/Y sky130_fd_sc_hd__o21ai_1_408/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_419 VSS VDD sky130_fd_sc_hd__o21ai_1_419/A2 sky130_fd_sc_hd__nor2_1_267/A
+ sky130_fd_sc_hd__nand2_1_486/Y sky130_fd_sc_hd__xor2_1_236/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a21oi_1_380 sky130_fd_sc_hd__nor2_2_17/Y sky130_fd_sc_hd__o21ai_1_393/Y
+ sky130_fd_sc_hd__nor2_1_249/B sky130_fd_sc_hd__fa_2_1247/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_391 sky130_fd_sc_hd__nand2_1_491/B sky130_fd_sc_hd__o22ai_1_358/Y
+ sky130_fd_sc_hd__a21oi_1_391/Y sky130_fd_sc_hd__o21ai_1_415/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nor2_4_17 sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__nor2_8_0/A
+ sky130_fd_sc_hd__nor2_4_17/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__xor2_1_202 sky130_fd_sc_hd__fa_2_1173/A sky130_fd_sc_hd__fa_2_1177/B
+ sky130_fd_sc_hd__xor2_1_202/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_213 sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__fa_2_1205/B
+ sky130_fd_sc_hd__xor2_1_213/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_224 sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__fa_2_1194/B
+ sky130_fd_sc_hd__xor2_1_224/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_235 sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1240/B
+ sky130_fd_sc_hd__xor2_1_235/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_246 sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1229/B
+ sky130_fd_sc_hd__xor2_1_246/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_257 sky130_fd_sc_hd__xor2_1_267/B sky130_fd_sc_hd__fa_2_1257/B
+ sky130_fd_sc_hd__xor2_1_257/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_608 VDD VSS sky130_fd_sc_hd__and2_0_229/A sky130_fd_sc_hd__dfxtp_1_611/CLK
+ sky130_fd_sc_hd__fa_2_1028/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_268 sky130_fd_sc_hd__fa_2_1242/A sky130_fd_sc_hd__fa_2_1246/B
+ sky130_fd_sc_hd__xor2_1_268/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_619 VDD VSS sky130_fd_sc_hd__ha_2_143/B sky130_fd_sc_hd__dfxtp_1_626/CLK
+ sky130_fd_sc_hd__a21oi_1_76/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_279 sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1292/B
+ sky130_fd_sc_hd__xor2_1_279/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_206 VSS VDD sky130_fd_sc_hd__bufbuf_16_3/A sky130_fd_sc_hd__clkinv_1_114/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_217 VSS VDD sky130_fd_sc_hd__buf_8_104/A sky130_fd_sc_hd__clkbuf_4_101/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_228 VSS VDD sky130_fd_sc_hd__clkbuf_1_228/X sky130_fd_sc_hd__clkbuf_1_228/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_239 VSS VDD sky130_fd_sc_hd__buf_4_44/A sky130_fd_sc_hd__buf_8_77/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_2_40 VDD VSS sky130_fd_sc_hd__buf_2_40/X sky130_fd_sc_hd__buf_2_40/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_51 VDD VSS sky130_fd_sc_hd__buf_8_74/A sky130_fd_sc_hd__ha_2_46/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_62 VDD VSS sky130_fd_sc_hd__buf_2_62/X sky130_fd_sc_hd__buf_2_62/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_73 VDD VSS sky130_fd_sc_hd__buf_2_73/X sky130_fd_sc_hd__buf_2_73/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_84 VDD VSS sky130_fd_sc_hd__buf_2_84/X sky130_fd_sc_hd__buf_2_84/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_95 VDD VSS sky130_fd_sc_hd__buf_2_95/X sky130_fd_sc_hd__buf_2_95/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__diode_2_2 sky130_fd_sc_hd__buf_2_122/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__and2_0_204 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_204/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__ha_2_166/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_215 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_215/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_215/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_226 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_226/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_226/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_237 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_237/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__fa_2_875/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_248 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_248/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__xnor2_1_27/Y sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_259 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_259/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__fa_2_960/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__sdlclkp_2_9 sky130_fd_sc_hd__conb_1_20/LO sky130_fd_sc_hd__clkinv_8_62/Y
+ sky130_fd_sc_hd__dfxtp_1_548/CLK sky130_fd_sc_hd__o21ai_1_32/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_2
Xsky130_fd_sc_hd__a22o_2_3 sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__ha_2_69/A
+ sky130_fd_sc_hd__a22o_2_3/X sky130_fd_sc_hd__dfxtp_1_2/Q sky130_fd_sc_hd__a22o_2_3/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_2
Xsky130_fd_sc_hd__o31ai_1_2 sky130_fd_sc_hd__o31ai_1_2/Y sky130_fd_sc_hd__nor3_1_31/C
+ sky130_fd_sc_hd__nor4_1_5/C sky130_fd_sc_hd__o31ai_1_2/A3 sky130_fd_sc_hd__o31ai_1_2/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__o31ai_1
Xsky130_fd_sc_hd__clkinv_1_280 sky130_fd_sc_hd__fa_2_86/A sky130_fd_sc_hd__ha_2_97/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_280/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_291 sky130_fd_sc_hd__fa_2_281/A sky130_fd_sc_hd__fa_2_31/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_291/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkbuf_4_12 sky130_fd_sc_hd__clkbuf_4_12/X sky130_fd_sc_hd__clkbuf_4_12/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_205 VSS VDD sky130_fd_sc_hd__xnor2_1_64/A sky130_fd_sc_hd__nor2_1_106/Y
+ sky130_fd_sc_hd__nand2_1_300/Y sky130_fd_sc_hd__xnor2_1_66/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_23 sky130_fd_sc_hd__clkbuf_4_23/X sky130_fd_sc_hd__clkbuf_4_23/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_216 VSS VDD sky130_fd_sc_hd__nand2_2_6/Y sky130_fd_sc_hd__a21oi_1_206/Y
+ sky130_fd_sc_hd__a21oi_1_192/Y sky130_fd_sc_hd__xor2_1_122/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_34 sky130_fd_sc_hd__a22oi_2_8/B2 sky130_fd_sc_hd__clkbuf_4_34/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_227 VSS VDD sky130_fd_sc_hd__nand2_2_6/Y sky130_fd_sc_hd__o21ai_1_227/A1
+ sky130_fd_sc_hd__a21oi_1_201/Y sky130_fd_sc_hd__xor2_1_128/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_45 sky130_fd_sc_hd__nand4_1_12/D sky130_fd_sc_hd__a22oi_1_68/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_238 VSS VDD sky130_fd_sc_hd__o22ai_1_204/B1 sky130_fd_sc_hd__nand4_1_86/D
+ sky130_fd_sc_hd__a21oi_1_212/Y sky130_fd_sc_hd__o21ai_1_238/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_56 sky130_fd_sc_hd__nand4_1_1/D sky130_fd_sc_hd__a22oi_1_31/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_249 VSS VDD sky130_fd_sc_hd__a211oi_1_9/Y sky130_fd_sc_hd__nor2_1_127/A
+ sky130_fd_sc_hd__a21oi_1_217/Y sky130_fd_sc_hd__xor2_1_99/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_67 sky130_fd_sc_hd__clkbuf_4_67/X sky130_fd_sc_hd__buf_2_40/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_78 sky130_fd_sc_hd__clkbuf_4_78/X sky130_fd_sc_hd__clkbuf_4_78/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_89 sky130_fd_sc_hd__clkbuf_4_89/X sky130_fd_sc_hd__clkbuf_4_89/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_8_140 sky130_fd_sc_hd__buf_8_140/A sky130_fd_sc_hd__buf_4_71/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_151 sky130_fd_sc_hd__buf_4_69/X sky130_fd_sc_hd__buf_8_171/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nor2_4_2 sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__nor2_4_2/A
+ sky130_fd_sc_hd__inv_2_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__buf_8_162 sky130_fd_sc_hd__buf_8_162/A sky130_fd_sc_hd__buf_6_43/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_173 sky130_fd_sc_hd__buf_8_173/A sky130_fd_sc_hd__buf_8_173/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_184 sky130_fd_sc_hd__buf_8_184/A sky130_fd_sc_hd__buf_8_184/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_195 sky130_fd_sc_hd__buf_8_213/A sky130_fd_sc_hd__buf_6_78/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_405 VDD VSS sky130_fd_sc_hd__fa_2_1041/A sky130_fd_sc_hd__dfxtp_1_425/CLK
+ sky130_fd_sc_hd__and2_0_123/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_416 VDD VSS sky130_fd_sc_hd__fa_2_1036/B sky130_fd_sc_hd__dfxtp_1_419/CLK
+ sky130_fd_sc_hd__and2_0_147/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_427 VDD VSS sky130_fd_sc_hd__dfxtp_1_427/Q sky130_fd_sc_hd__dfxtp_1_433/CLK
+ sky130_fd_sc_hd__nand2_1_110/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_438 VDD VSS sky130_fd_sc_hd__dfxtp_1_438/Q sky130_fd_sc_hd__dfxtp_1_452/CLK
+ sky130_fd_sc_hd__nand2_1_88/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_449 VDD VSS sky130_fd_sc_hd__dfxtp_1_995/D sky130_fd_sc_hd__dfxtp_1_454/CLK
+ sky130_fd_sc_hd__nand2_1_66/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkinv_8_15 sky130_fd_sc_hd__clkinv_8_15/Y sky130_fd_sc_hd__clkinv_8_15/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_26 sky130_fd_sc_hd__clkinv_8_33/A sky130_fd_sc_hd__clkinv_8_26/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_26/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_37 sky130_fd_sc_hd__clkinv_8_38/A sky130_fd_sc_hd__clkinv_8_37/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_37/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_48 sky130_fd_sc_hd__clkinv_8_48/Y sky130_fd_sc_hd__clkinv_8_49/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_48/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_59 sky130_fd_sc_hd__clkinv_8_59/Y sky130_fd_sc_hd__clkinv_8_59/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_59/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_13 sky130_fd_sc_hd__inv_2_35/Y sky130_fd_sc_hd__buf_12_94/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_24 sky130_fd_sc_hd__buf_8_34/A sky130_fd_sc_hd__buf_8_58/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_35 sky130_fd_sc_hd__buf_8_5/X sky130_fd_sc_hd__buf_12_35/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_90 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__xor2_1_90/X
+ sky130_fd_sc_hd__xor2_1_90/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_46 sky130_fd_sc_hd__buf_8_47/X sky130_fd_sc_hd__buf_12_46/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_57 sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__buf_12_57/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_68 sky130_fd_sc_hd__buf_4_26/X sky130_fd_sc_hd__buf_12_68/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_79 sky130_fd_sc_hd__buf_12_79/A sky130_fd_sc_hd__buf_12_79/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_2_8 VDD VSS sky130_fd_sc_hd__buf_2_8/X sky130_fd_sc_hd__buf_2_8/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1301 VDD VSS sky130_fd_sc_hd__ha_2_146/B sky130_fd_sc_hd__dfxtp_1_1329/CLK
+ sky130_fd_sc_hd__o32ai_1_10/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1312 VDD VSS sky130_fd_sc_hd__fa_2_839/B sky130_fd_sc_hd__dfxtp_1_1326/CLK
+ sky130_fd_sc_hd__a21oi_1_430/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1323 VDD VSS sky130_fd_sc_hd__fa_2_907/A sky130_fd_sc_hd__dfxtp_1_1326/CLK
+ sky130_fd_sc_hd__o21a_1_60/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1334 VDD VSS sky130_fd_sc_hd__fa_2_1293/B sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__and2_0_335/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1345 VDD VSS sky130_fd_sc_hd__fa_2_1304/A sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__mux2_2_234/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1356 VDD VSS sky130_fd_sc_hd__fa_2_1278/A sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__mux2_2_258/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1367 VDD VSS sky130_fd_sc_hd__fa_2_1289/A sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__mux2_2_229/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1378 VDD VSS sky130_fd_sc_hd__fa_2_1317/A sky130_fd_sc_hd__clkinv_8_63/Y
+ sky130_fd_sc_hd__mux2_2_259/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_950 VDD VSS sky130_fd_sc_hd__fa_2_1159/A sky130_fd_sc_hd__clkinv_8_64/Y
+ sky130_fd_sc_hd__mux2_2_122/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1389 VDD VSS sky130_fd_sc_hd__o32ai_1_11/A1 sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__nor2b_1_130/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_961 VDD VSS sky130_fd_sc_hd__fa_2_1170/A sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__mux2_2_97/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_972 VDD VSS sky130_fd_sc_hd__mux2_2_114/A0 sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__dfxtp_1_972/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_983 VDD VSS sky130_fd_sc_hd__mux2_2_85/A1 sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__o22ai_1_212/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_994 VDD VSS sky130_fd_sc_hd__mux2_2_115/A0 sky130_fd_sc_hd__clkinv_8_64/Y
+ sky130_fd_sc_hd__dfxtp_1_994/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_570 VSS VDD sky130_fd_sc_hd__nand2_1_9/A sky130_fd_sc_hd__nor3_2_0/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_581 VSS VDD sky130_fd_sc_hd__nand3_1_10/A sky130_fd_sc_hd__a22oi_1_21/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_592 VSS VDD sky130_fd_sc_hd__nand3_1_0/B sky130_fd_sc_hd__a22oi_1_0/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_800 sky130_fd_sc_hd__fa_2_799/B sky130_fd_sc_hd__fa_2_800/SUM
+ sky130_fd_sc_hd__fa_2_800/A sky130_fd_sc_hd__fa_2_800/B sky130_fd_sc_hd__fa_2_800/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_160 VSS VDD VSS VDD sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__ha_2_159/B
+ sky130_fd_sc_hd__ha_2_160/SUM sky130_fd_sc_hd__ha_2_160/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_811 sky130_fd_sc_hd__fa_2_813/CIN sky130_fd_sc_hd__fa_2_805/B
+ sky130_fd_sc_hd__fa_2_811/A sky130_fd_sc_hd__fa_2_823/B sky130_fd_sc_hd__fa_2_826/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_171 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_171/A sky130_fd_sc_hd__ha_2_170/A
+ sky130_fd_sc_hd__ha_2_171/SUM sky130_fd_sc_hd__ha_2_171/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_822 sky130_fd_sc_hd__fa_2_821/B sky130_fd_sc_hd__fa_2_822/SUM
+ sky130_fd_sc_hd__ha_2_140/B sky130_fd_sc_hd__fa_2_822/B sky130_fd_sc_hd__fa_2_822/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_182 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_182/A sky130_fd_sc_hd__ha_2_181/A
+ sky130_fd_sc_hd__ha_2_182/SUM sky130_fd_sc_hd__ha_2_182/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_833 sky130_fd_sc_hd__fa_2_832/CIN sky130_fd_sc_hd__fa_2_833/SUM
+ sky130_fd_sc_hd__fa_2_833/A sky130_fd_sc_hd__fa_2_834/A sky130_fd_sc_hd__ha_2_144/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_193 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_193/A sky130_fd_sc_hd__ha_2_192/A
+ sky130_fd_sc_hd__ha_2_193/SUM sky130_fd_sc_hd__ha_2_193/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_844 sky130_fd_sc_hd__fa_2_843/CIN sky130_fd_sc_hd__fa_2_844/SUM
+ sky130_fd_sc_hd__fa_2_844/A sky130_fd_sc_hd__fa_2_844/B sky130_fd_sc_hd__fa_2_844/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_855 sky130_fd_sc_hd__fa_2_854/CIN sky130_fd_sc_hd__fa_2_855/SUM
+ sky130_fd_sc_hd__fa_2_855/A sky130_fd_sc_hd__fa_2_855/B sky130_fd_sc_hd__fa_2_855/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_866 sky130_fd_sc_hd__fa_2_865/CIN sky130_fd_sc_hd__fa_2_866/SUM
+ sky130_fd_sc_hd__fa_2_866/A sky130_fd_sc_hd__fa_2_866/B sky130_fd_sc_hd__fa_2_866/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_877 sky130_fd_sc_hd__fa_2_876/CIN sky130_fd_sc_hd__fa_2_877/SUM
+ sky130_fd_sc_hd__fa_2_877/A sky130_fd_sc_hd__fa_2_877/B sky130_fd_sc_hd__nand2b_1_3/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_888 sky130_fd_sc_hd__xor2_1_24/A sky130_fd_sc_hd__fa_2_888/SUM
+ sky130_fd_sc_hd__fa_2_888/A sky130_fd_sc_hd__fa_2_888/B sky130_fd_sc_hd__fa_2_888/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_899 sky130_fd_sc_hd__fa_2_898/CIN sky130_fd_sc_hd__fa_2_899/SUM
+ sky130_fd_sc_hd__fa_2_899/A sky130_fd_sc_hd__fa_2_899/B sky130_fd_sc_hd__fa_2_899/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_8 sky130_fd_sc_hd__inv_2_8/A sky130_fd_sc_hd__inv_2_8/Y VDD
+ VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__mux2_2_100 VSS VDD sky130_fd_sc_hd__mux2_2_100/A1 sky130_fd_sc_hd__mux2_2_100/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_100/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_111 VSS VDD sky130_fd_sc_hd__mux2_2_111/A1 sky130_fd_sc_hd__mux2_2_111/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_111/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_18 sky130_fd_sc_hd__nor3_1_28/Y sky130_fd_sc_hd__nor2_1_18/Y
+ sky130_fd_sc_hd__inv_4_1/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_122 VSS VDD sky130_fd_sc_hd__mux2_2_122/A1 sky130_fd_sc_hd__mux2_2_122/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_122/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_29 sky130_fd_sc_hd__or4_1_2/C sky130_fd_sc_hd__nor2_1_29/Y
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_133 VSS VDD sky130_fd_sc_hd__mux2_2_133/A1 sky130_fd_sc_hd__mux2_2_133/A0
+ sky130_fd_sc_hd__mux2_2_135/S sky130_fd_sc_hd__mux2_2_133/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_144 VSS VDD sky130_fd_sc_hd__mux2_2_144/A1 sky130_fd_sc_hd__mux2_2_144/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_144/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_155 VSS VDD sky130_fd_sc_hd__mux2_2_155/A1 sky130_fd_sc_hd__mux2_2_155/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_155/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_166 VSS VDD sky130_fd_sc_hd__mux2_2_166/A1 sky130_fd_sc_hd__mux2_2_166/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_166/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_177 VSS VDD sky130_fd_sc_hd__mux2_2_177/A1 sky130_fd_sc_hd__mux2_2_177/A0
+ sky130_fd_sc_hd__nor2_8_1/A sky130_fd_sc_hd__mux2_2_177/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_188 VSS VDD sky130_fd_sc_hd__xor2_1_273/X sky130_fd_sc_hd__nand2_1_468/B
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_188/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_199 VSS VDD sky130_fd_sc_hd__mux2_2_199/A1 sky130_fd_sc_hd__mux2_2_199/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_199/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__and2_0_40 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_59/A sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__xor2_1_5/X sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_104 sky130_fd_sc_hd__maj3_1_105/X sky130_fd_sc_hd__maj3_1_104/X
+ sky130_fd_sc_hd__maj3_1_104/B sky130_fd_sc_hd__maj3_1_104/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_320 sky130_fd_sc_hd__o22ai_1_322/A2 sky130_fd_sc_hd__nor2_1_223/A
+ sky130_fd_sc_hd__o22ai_1_320/Y sky130_fd_sc_hd__nor2_1_193/B sky130_fd_sc_hd__o32ai_1_5/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_51 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_51/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_51/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_115 sky130_fd_sc_hd__maj3_1_116/X sky130_fd_sc_hd__maj3_1_115/X
+ sky130_fd_sc_hd__maj3_1_115/B sky130_fd_sc_hd__maj3_1_115/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_331 sky130_fd_sc_hd__nand2_1_462/Y sky130_fd_sc_hd__nand2_1_461/Y
+ sky130_fd_sc_hd__o22ai_1_331/Y sky130_fd_sc_hd__o22ai_1_344/A1 sky130_fd_sc_hd__a21o_2_21/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_62 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_83/A sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__ha_2_71/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_126 sky130_fd_sc_hd__maj3_1_127/X sky130_fd_sc_hd__maj3_1_126/X
+ sky130_fd_sc_hd__maj3_1_126/B sky130_fd_sc_hd__maj3_1_126/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_342 sky130_fd_sc_hd__nand2_1_464/Y sky130_fd_sc_hd__nand2_1_463/Y
+ sky130_fd_sc_hd__o22ai_1_342/Y sky130_fd_sc_hd__o22ai_1_342/A1 sky130_fd_sc_hd__a21o_2_20/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_73 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_73/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__and2_0_73/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_406 sky130_fd_sc_hd__o21a_1_41/B1 sky130_fd_sc_hd__fa_2_1196/A
+ sky130_fd_sc_hd__o21a_1_41/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_137 sky130_fd_sc_hd__maj3_1_138/X sky130_fd_sc_hd__maj3_1_137/X
+ sky130_fd_sc_hd__maj3_1_137/B sky130_fd_sc_hd__maj3_1_137/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_353 sky130_fd_sc_hd__nor2_1_268/A sky130_fd_sc_hd__nor2_1_265/A
+ sky130_fd_sc_hd__o22ai_1_353/Y sky130_fd_sc_hd__a21boi_1_5/Y sky130_fd_sc_hd__nor2_1_250/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_84 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_84/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__and2_0_84/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_417 sky130_fd_sc_hd__nand2_1_417/Y sky130_fd_sc_hd__mux2_2_171/S
+ sky130_fd_sc_hd__nand2_1_417/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_148 sky130_fd_sc_hd__maj3_1_149/X sky130_fd_sc_hd__maj3_1_148/X
+ sky130_fd_sc_hd__maj3_1_148/B sky130_fd_sc_hd__maj3_1_148/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_364 sky130_fd_sc_hd__o22ai_1_379/A2 sky130_fd_sc_hd__o22ai_1_364/B1
+ sky130_fd_sc_hd__o22ai_1_364/Y sky130_fd_sc_hd__nor2_1_228/B sky130_fd_sc_hd__o32ai_1_8/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_95 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_95/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_95/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_159 sky130_fd_sc_hd__maj3_1_160/X sky130_fd_sc_hd__maj3_1_159/X
+ sky130_fd_sc_hd__maj3_1_159/B sky130_fd_sc_hd__maj3_1_159/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_428 sky130_fd_sc_hd__nand2_1_428/Y sky130_fd_sc_hd__nor2b_2_3/A
+ sky130_fd_sc_hd__xor2_1_209/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_375 sky130_fd_sc_hd__o22ai_1_375/A2 sky130_fd_sc_hd__nor2_1_238/B
+ sky130_fd_sc_hd__o22ai_1_375/Y sky130_fd_sc_hd__nor2_1_239/B sky130_fd_sc_hd__o32ai_1_8/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_439 sky130_fd_sc_hd__nand2_1_439/Y sky130_fd_sc_hd__nand2_1_439/B
+ sky130_fd_sc_hd__o21ai_1_370/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_386 sky130_fd_sc_hd__nand2_1_514/Y sky130_fd_sc_hd__nand2_1_513/Y
+ sky130_fd_sc_hd__o22ai_1_386/Y sky130_fd_sc_hd__o22ai_1_399/A1 sky130_fd_sc_hd__a21o_2_26/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_397 sky130_fd_sc_hd__nand2_1_516/Y sky130_fd_sc_hd__nand2_1_515/Y
+ sky130_fd_sc_hd__o22ai_1_397/Y sky130_fd_sc_hd__o22ai_1_397/A1 sky130_fd_sc_hd__a21o_2_25/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2b_1_19 sky130_fd_sc_hd__ha_2_49/SUM sky130_fd_sc_hd__nor2b_1_19/Y
+ sky130_fd_sc_hd__or2_1_0/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1008 sky130_fd_sc_hd__nor2_1_263/A sky130_fd_sc_hd__xor2_1_253/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1008/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_50 sky130_fd_sc_hd__inv_2_36/Y sky130_fd_sc_hd__buf_8_50/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__clkinv_1_1019 sky130_fd_sc_hd__o21ai_1_436/A1 sky130_fd_sc_hd__fa_2_1256/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1019/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_61 sky130_fd_sc_hd__buf_8_61/A sky130_fd_sc_hd__buf_8_61/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_72 sky130_fd_sc_hd__buf_8_72/A sky130_fd_sc_hd__buf_8_72/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_83 sky130_fd_sc_hd__buf_8_83/A sky130_fd_sc_hd__buf_8_83/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_202 VDD VSS sky130_fd_sc_hd__ha_2_79/A sky130_fd_sc_hd__dfxtp_1_207/CLK
+ sky130_fd_sc_hd__and2_0_81/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_8_94 sky130_fd_sc_hd__buf_8_94/A sky130_fd_sc_hd__buf_8_94/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_213 VDD VSS sky130_fd_sc_hd__ha_2_89/B sky130_fd_sc_hd__dfxtp_1_224/CLK
+ sky130_fd_sc_hd__nor2b_1_38/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_224 VDD VSS sky130_fd_sc_hd__xor2_1_8/B sky130_fd_sc_hd__dfxtp_1_224/CLK
+ sky130_fd_sc_hd__nor2b_1_39/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_235 VDD VSS sky130_fd_sc_hd__fa_2_874/A sky130_fd_sc_hd__dfxtp_1_462/CLK
+ sky130_fd_sc_hd__and2_0_164/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_246 VDD VSS sky130_fd_sc_hd__xor2_1_15/A sky130_fd_sc_hd__dfxtp_1_266/CLK
+ sky130_fd_sc_hd__and2_0_184/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_257 VDD VSS sky130_fd_sc_hd__dfxtp_1_257/Q sky130_fd_sc_hd__dfxtp_1_258/CLK
+ sky130_fd_sc_hd__and2_0_220/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_268 VDD VSS sky130_fd_sc_hd__dfxtp_1_268/Q sky130_fd_sc_hd__dfxtp_1_277/CLK
+ sky130_fd_sc_hd__and2_0_226/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_279 VDD VSS sky130_fd_sc_hd__buf_2_262/A sky130_fd_sc_hd__dfxtp_1_282/CLK
+ sky130_fd_sc_hd__a211o_1_0/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_107 sky130_fd_sc_hd__fa_2_104/A sky130_fd_sc_hd__fa_2_99/A
+ sky130_fd_sc_hd__fa_2_82/A sky130_fd_sc_hd__ha_2_97/B sky130_fd_sc_hd__fa_2_96/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_118 sky130_fd_sc_hd__fa_2_121/B sky130_fd_sc_hd__fa_2_118/SUM
+ sky130_fd_sc_hd__fa_2_118/A sky130_fd_sc_hd__fa_2_118/B sky130_fd_sc_hd__fa_2_118/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_129 sky130_fd_sc_hd__fa_2_27/A sky130_fd_sc_hd__fa_2_29/B sky130_fd_sc_hd__fa_2_129/A
+ sky130_fd_sc_hd__fa_2_129/B sky130_fd_sc_hd__fa_2_134/SUM VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_102 VDD VSS sky130_fd_sc_hd__buf_2_102/X sky130_fd_sc_hd__buf_2_102/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__fa_2_1301 sky130_fd_sc_hd__fa_2_1302/CIN sky130_fd_sc_hd__mux2_2_242/A1
+ sky130_fd_sc_hd__fa_2_1301/A sky130_fd_sc_hd__fa_2_1301/B sky130_fd_sc_hd__fa_2_1301/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_113 VDD VSS sky130_fd_sc_hd__buf_4_38/A sky130_fd_sc_hd__buf_2_117/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__fa_2_1312 sky130_fd_sc_hd__fa_2_1313/CIN sky130_fd_sc_hd__mux2_2_266/A1
+ sky130_fd_sc_hd__fa_2_1312/A sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1312/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_124 VDD VSS sky130_fd_sc_hd__buf_2_124/X sky130_fd_sc_hd__buf_2_124/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_17 sky130_fd_sc_hd__fa_2_5/B sky130_fd_sc_hd__fa_2_144/B
+ sky130_fd_sc_hd__o22ai_1_17/Y sky130_fd_sc_hd__ha_2_97/A sky130_fd_sc_hd__fa_2_280/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_1323 sky130_fd_sc_hd__fa_2_1324/CIN sky130_fd_sc_hd__mux2_2_241/A1
+ sky130_fd_sc_hd__fa_2_1323/A sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1323/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_135 VDD VSS sky130_fd_sc_hd__buf_8_119/A sky130_fd_sc_hd__a22o_2_1/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_28 sky130_fd_sc_hd__fa_2_389/B sky130_fd_sc_hd__fa_2_412/A
+ sky130_fd_sc_hd__fa_2_411/B sky130_fd_sc_hd__ha_2_108/B sky130_fd_sc_hd__ha_2_115/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_146 VDD VSS sky130_fd_sc_hd__buf_2_146/X sky130_fd_sc_hd__buf_2_146/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_39 sky130_fd_sc_hd__fa_2_427/B sky130_fd_sc_hd__fa_2_559/B
+ sky130_fd_sc_hd__fa_2_463/A sky130_fd_sc_hd__ha_2_169/B sky130_fd_sc_hd__ha_2_125/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_157 VDD VSS sky130_fd_sc_hd__or2_1_2/B sky130_fd_sc_hd__nor2b_2_2/Y
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_168 VDD VSS sky130_fd_sc_hd__buf_2_168/X sky130_fd_sc_hd__buf_2_168/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_179 VDD VSS sky130_fd_sc_hd__buf_2_179/X sky130_fd_sc_hd__buf_2_179/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1120 VDD VSS sky130_fd_sc_hd__mux2_2_142/A0 sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__o22ai_1_273/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1131 VDD VSS sky130_fd_sc_hd__mux2_2_169/A0 sky130_fd_sc_hd__clkinv_8_64/Y
+ sky130_fd_sc_hd__dfxtp_1_990/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1142 VDD VSS sky130_fd_sc_hd__nand2_1_416/B sky130_fd_sc_hd__clkinv_8_78/Y
+ sky130_fd_sc_hd__xnor2_1_96/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1153 VDD VSS sky130_fd_sc_hd__mux2_2_136/A0 sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__o22ai_1_284/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1164 VDD VSS sky130_fd_sc_hd__fa_2_860/B sky130_fd_sc_hd__dfxtp_1_1180/CLK
+ sky130_fd_sc_hd__a21oi_1_374/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1175 VDD VSS sky130_fd_sc_hd__xnor2_1_9/A sky130_fd_sc_hd__dfxtp_1_1180/CLK
+ sky130_fd_sc_hd__xnor2_1_98/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1186 VDD VSS sky130_fd_sc_hd__fa_2_939/A sky130_fd_sc_hd__clkinv_4_24/Y
+ sky130_fd_sc_hd__o21a_1_45/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1197 VDD VSS sky130_fd_sc_hd__fa_2_1246/A sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__mux2_2_206/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__ha_2_2 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_2/A sky130_fd_sc_hd__ha_2_1/B
+ sky130_fd_sc_hd__ha_2_2/SUM sky130_fd_sc_hd__ha_2_2/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__buf_4_19 VDD VSS sky130_fd_sc_hd__buf_4_19/X sky130_fd_sc_hd__buf_8_26/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__dfxtp_1_780 VDD VSS sky130_fd_sc_hd__fa_2_1079/A sky130_fd_sc_hd__clkinv_8_55/Y
+ sky130_fd_sc_hd__mux2_2_64/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_791 VDD VSS sky130_fd_sc_hd__fa_2_1090/A sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__mux2_2_42/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_13 VSS VDD sky130_fd_sc_hd__clkbuf_4_6/A sky130_fd_sc_hd__buf_4_10/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_24 VSS VDD sky130_fd_sc_hd__clkbuf_1_24/X sky130_fd_sc_hd__clkbuf_1_24/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_630 sky130_fd_sc_hd__maj3_1_115/B sky130_fd_sc_hd__maj3_1_116/A
+ sky130_fd_sc_hd__fa_2_630/A sky130_fd_sc_hd__fa_2_630/B sky130_fd_sc_hd__fa_2_630/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_35 VSS VDD sky130_fd_sc_hd__clkbuf_1_35/X sky130_fd_sc_hd__clkbuf_1_35/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_641 sky130_fd_sc_hd__maj3_1_112/B sky130_fd_sc_hd__maj3_1_113/A
+ sky130_fd_sc_hd__fa_2_641/A sky130_fd_sc_hd__fa_2_641/B sky130_fd_sc_hd__fa_2_642/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_46 VSS VDD sky130_fd_sc_hd__clkbuf_1_46/X sky130_fd_sc_hd__clkbuf_1_46/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_652 sky130_fd_sc_hd__maj3_1_109/B sky130_fd_sc_hd__maj3_1_110/A
+ sky130_fd_sc_hd__fa_2_652/A sky130_fd_sc_hd__fa_2_652/B sky130_fd_sc_hd__fa_2_653/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_57 VSS VDD sky130_fd_sc_hd__clkbuf_1_57/X sky130_fd_sc_hd__clkbuf_1_57/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_663 sky130_fd_sc_hd__fa_2_664/CIN sky130_fd_sc_hd__fa_2_657/B
+ sky130_fd_sc_hd__fa_2_700/A sky130_fd_sc_hd__fa_2_689/B sky130_fd_sc_hd__fa_2_683/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_68 VSS VDD sky130_fd_sc_hd__clkbuf_1_68/X sky130_fd_sc_hd__clkbuf_1_68/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_674 sky130_fd_sc_hd__fa_2_676/CIN sky130_fd_sc_hd__fa_2_665/A
+ sky130_fd_sc_hd__ha_2_128/A sky130_fd_sc_hd__fa_2_674/B sky130_fd_sc_hd__fa_2_674/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_79 VSS VDD sky130_fd_sc_hd__nand4_1_8/A sky130_fd_sc_hd__a22oi_2_9/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_685 sky130_fd_sc_hd__fa_2_684/B sky130_fd_sc_hd__fa_2_685/SUM
+ sky130_fd_sc_hd__fa_2_685/A sky130_fd_sc_hd__fa_2_685/B sky130_fd_sc_hd__fa_2_689/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_696 sky130_fd_sc_hd__fa_2_572/A sky130_fd_sc_hd__fa_2_573/B
+ sky130_fd_sc_hd__fa_2_700/B sky130_fd_sc_hd__fa_2_696/B sky130_fd_sc_hd__fa_2_699/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a21oi_1_209 sky130_fd_sc_hd__a21o_2_5/A2 sky130_fd_sc_hd__o22ai_1_181/Y
+ sky130_fd_sc_hd__a21oi_1_209/Y sky130_fd_sc_hd__fa_2_1050/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_2_16 sky130_fd_sc_hd__buf_2_165/X sky130_fd_sc_hd__a22oi_2_16/A2
+ sky130_fd_sc_hd__nor2_4_7/Y sky130_fd_sc_hd__a22oi_2_16/B2 sky130_fd_sc_hd__nand4_1_50/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__a22oi_2_27 sky130_fd_sc_hd__buf_2_165/X sky130_fd_sc_hd__a22oi_2_27/A2
+ sky130_fd_sc_hd__nor2_4_7/Y sky130_fd_sc_hd__a22oi_2_27/B2 sky130_fd_sc_hd__nand4_1_59/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__buf_12_2 sky130_fd_sc_hd__inv_2_12/Y sky130_fd_sc_hd__buf_12_2/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__nand2_1_203 sky130_fd_sc_hd__nor2_1_22/B sky130_fd_sc_hd__nand2_1_203/B
+ sky130_fd_sc_hd__nor2_1_23/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_802 sky130_fd_sc_hd__o22ai_1_232/A1 sky130_fd_sc_hd__nor2_1_170/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_802/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_150 sky130_fd_sc_hd__nand2_1_338/A sky130_fd_sc_hd__nand2_1_284/Y
+ sky130_fd_sc_hd__o22ai_1_150/Y sky130_fd_sc_hd__xnor2_1_64/Y sky130_fd_sc_hd__o22ai_1_150/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_214 sky130_fd_sc_hd__nor2_1_31/B sky130_fd_sc_hd__nand2_1_214/B
+ sky130_fd_sc_hd__nor2_1_33/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_161 sky130_fd_sc_hd__nand2_1_338/A sky130_fd_sc_hd__nand2_1_284/Y
+ sky130_fd_sc_hd__o22ai_1_161/Y sky130_fd_sc_hd__xnor2_1_86/Y sky130_fd_sc_hd__o22ai_1_161/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_813 sky130_fd_sc_hd__nand2_1_368/B sky130_fd_sc_hd__fa_2_429/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_813/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_225 sky130_fd_sc_hd__o21ai_1_39/B1 sky130_fd_sc_hd__o22ai_1_59/A2
+ sky130_fd_sc_hd__fa_2_955/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_172 sky130_fd_sc_hd__nor2_1_126/A sky130_fd_sc_hd__nor2_2_13/B
+ sky130_fd_sc_hd__o22ai_1_172/Y sky130_fd_sc_hd__a21oi_1_202/Y sky130_fd_sc_hd__a222oi_1_2/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_824 sky130_fd_sc_hd__o22ai_1_247/A1 sky130_fd_sc_hd__fa_2_1132/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_824/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_236 sky130_fd_sc_hd__xnor2_1_60/B sky130_fd_sc_hd__o21ai_1_74/B1
+ sky130_fd_sc_hd__o21ai_1_81/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_183 sky130_fd_sc_hd__o22ai_1_204/B1 sky130_fd_sc_hd__nor2_1_117/B
+ sky130_fd_sc_hd__nor2_1_131/A sky130_fd_sc_hd__nor2_1_118/B sky130_fd_sc_hd__o22ai_1_206/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_835 sky130_fd_sc_hd__nor2_1_144/B sky130_fd_sc_hd__fa_2_1133/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_835/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_247 sky130_fd_sc_hd__nand2_1_247/Y sky130_fd_sc_hd__nor2_1_52/B
+ sky130_fd_sc_hd__nor2_1_52/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_194 sky130_fd_sc_hd__o21a_1_16/A2 sky130_fd_sc_hd__o22ai_1_194/B1
+ sky130_fd_sc_hd__nor2_1_135/B sky130_fd_sc_hd__nor2_1_120/B sky130_fd_sc_hd__o22ai_1_206/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand4_1_20 sky130_fd_sc_hd__nand4_1_20/C sky130_fd_sc_hd__nand4_1_20/B
+ sky130_fd_sc_hd__nand4_1_20/Y sky130_fd_sc_hd__nand4_1_20/D sky130_fd_sc_hd__buf_2_108/X
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__clkinv_1_846 sky130_fd_sc_hd__nand2_1_341/B sky130_fd_sc_hd__nor2b_1_104/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_846/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_258 sky130_fd_sc_hd__o21ai_1_89/B1 sky130_fd_sc_hd__nand2_1_282/B
+ sky130_fd_sc_hd__o21ai_1_90/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand4_1_31 sky130_fd_sc_hd__nand4_1_31/C sky130_fd_sc_hd__nand4_1_31/B
+ sky130_fd_sc_hd__nand4_1_31/Y sky130_fd_sc_hd__nand4_1_31/D sky130_fd_sc_hd__buf_2_100/X
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__clkinv_1_857 sky130_fd_sc_hd__o21a_1_29/A2 sky130_fd_sc_hd__fa_2_1151/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_857/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_269 sky130_fd_sc_hd__o211ai_1_7/C1 sky130_fd_sc_hd__a211o_1_6/A1
+ sky130_fd_sc_hd__a211o_1_8/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand4_1_42 sky130_fd_sc_hd__nand4_1_42/C sky130_fd_sc_hd__nand4_1_42/B
+ sky130_fd_sc_hd__buf_2_288/A sky130_fd_sc_hd__nand4_1_42/D sky130_fd_sc_hd__nand4_1_42/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__clkinv_1_868 sky130_fd_sc_hd__nor2_1_222/A sky130_fd_sc_hd__nor2b_2_3/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_868/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_879 sky130_fd_sc_hd__nor2_1_203/B sky130_fd_sc_hd__xor2_1_185/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_879/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand4_1_53 sky130_fd_sc_hd__nand4_1_53/C sky130_fd_sc_hd__nand4_1_53/B
+ sky130_fd_sc_hd__buf_2_268/A sky130_fd_sc_hd__nand4_1_53/D sky130_fd_sc_hd__nand4_1_53/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_64 sky130_fd_sc_hd__nand4_1_64/C sky130_fd_sc_hd__nand4_1_64/B
+ sky130_fd_sc_hd__nand4_1_64/Y sky130_fd_sc_hd__nand4_1_64/D sky130_fd_sc_hd__nand4_1_64/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_75 sky130_fd_sc_hd__nand4_1_75/C sky130_fd_sc_hd__nand4_1_75/B
+ sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__nand4_1_75/D sky130_fd_sc_hd__nand4_1_75/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_86 sky130_fd_sc_hd__nand4_1_86/C sky130_fd_sc_hd__nand4_1_86/B
+ sky130_fd_sc_hd__nand4_1_86/Y sky130_fd_sc_hd__nand4_1_86/D sky130_fd_sc_hd__nand4_1_86/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__conb_1_13 sky130_fd_sc_hd__conb_1_13/LO sky130_fd_sc_hd__conb_1_13/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_24 sky130_fd_sc_hd__conb_1_24/LO sky130_fd_sc_hd__conb_1_24/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__mux2_2_8 VSS VDD sky130_fd_sc_hd__mux2_2_8/A1 sky130_fd_sc_hd__mux2_2_8/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_8/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_90 VSS VDD sky130_fd_sc_hd__mux2_2_90/A1 sky130_fd_sc_hd__mux2_2_90/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_90/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1120 sky130_fd_sc_hd__fa_2_1121/CIN sky130_fd_sc_hd__fa_2_1120/SUM
+ sky130_fd_sc_hd__fa_2_1120/A sky130_fd_sc_hd__fa_2_1120/B sky130_fd_sc_hd__fa_2_1120/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1131 sky130_fd_sc_hd__fa_2_1132/CIN sky130_fd_sc_hd__mux2_2_96/A1
+ sky130_fd_sc_hd__fa_2_1131/A sky130_fd_sc_hd__fa_2_1131/B sky130_fd_sc_hd__fa_2_1131/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1142 sky130_fd_sc_hd__fa_2_1143/CIN sky130_fd_sc_hd__mux2_2_116/A1
+ sky130_fd_sc_hd__fa_2_1142/A sky130_fd_sc_hd__fa_2_1142/B sky130_fd_sc_hd__fa_2_1142/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1153 sky130_fd_sc_hd__fa_2_1154/CIN sky130_fd_sc_hd__mux2_2_86/A0
+ sky130_fd_sc_hd__fa_2_1153/A sky130_fd_sc_hd__fa_2_1153/B sky130_fd_sc_hd__fa_2_1153/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1164 sky130_fd_sc_hd__fa_2_1165/CIN sky130_fd_sc_hd__mux2_2_115/A1
+ sky130_fd_sc_hd__fa_2_1164/A sky130_fd_sc_hd__fa_2_1172/B sky130_fd_sc_hd__fa_2_1164/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1175 sky130_fd_sc_hd__fa_2_1176/CIN sky130_fd_sc_hd__mux2_2_165/A1
+ sky130_fd_sc_hd__fa_2_1175/A sky130_fd_sc_hd__fa_2_1175/B sky130_fd_sc_hd__fa_2_1175/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1186 sky130_fd_sc_hd__fa_2_1187/CIN sky130_fd_sc_hd__mux2_2_135/A0
+ sky130_fd_sc_hd__fa_2_1186/A sky130_fd_sc_hd__fa_2_1186/B sky130_fd_sc_hd__fa_2_1186/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1197 sky130_fd_sc_hd__fa_2_1198/CIN sky130_fd_sc_hd__mux2_2_152/A1
+ sky130_fd_sc_hd__fa_2_1197/A sky130_fd_sc_hd__fa_2_1197/B sky130_fd_sc_hd__fa_2_1197/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o2bb2ai_1_4 sky130_fd_sc_hd__o2bb2ai_1_4/Y sky130_fd_sc_hd__nor2_1_18/Y
+ sky130_fd_sc_hd__ha_2_154/SUM sky130_fd_sc_hd__o21ai_1_31/A1 sky130_fd_sc_hd__o21ai_1_29/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_460 sky130_fd_sc_hd__fa_2_456/CIN sky130_fd_sc_hd__or3_1_2/C
+ sky130_fd_sc_hd__fa_2_460/A sky130_fd_sc_hd__fa_2_460/B sky130_fd_sc_hd__fa_2_460/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_471 sky130_fd_sc_hd__maj3_1_102/B sky130_fd_sc_hd__maj3_1_103/A
+ sky130_fd_sc_hd__fa_2_471/A sky130_fd_sc_hd__fa_2_471/B sky130_fd_sc_hd__o22ai_1_33/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_482 sky130_fd_sc_hd__maj3_1_98/B sky130_fd_sc_hd__maj3_1_99/A
+ sky130_fd_sc_hd__fa_2_482/A sky130_fd_sc_hd__fa_2_482/B sky130_fd_sc_hd__fa_2_483/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_493 sky130_fd_sc_hd__fa_2_491/B sky130_fd_sc_hd__fa_2_486/A
+ sky130_fd_sc_hd__ha_2_124/A sky130_fd_sc_hd__ha_2_169/B sky130_fd_sc_hd__fa_2_546/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_1_109 sky130_fd_sc_hd__inv_2_71/A sky130_fd_sc_hd__buf_2_48/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_109/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_9 VSS VDD sky130_fd_sc_hd__o21ai_1_9/A2 sky130_fd_sc_hd__nor4_1_2/A
+ sky130_fd_sc_hd__nor2_1_22/A sky130_fd_sc_hd__o21ai_1_9/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__nor2_1_203 sky130_fd_sc_hd__nor2_1_203/B sky130_fd_sc_hd__nor2_1_203/Y
+ sky130_fd_sc_hd__nor2_1_205/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_214 sky130_fd_sc_hd__nor2_1_214/B sky130_fd_sc_hd__nor2_1_214/Y
+ sky130_fd_sc_hd__nor2_1_214/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_225 sky130_fd_sc_hd__nor2_1_225/B sky130_fd_sc_hd__nor2_1_225/Y
+ sky130_fd_sc_hd__nor2_1_225/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_236 sky130_fd_sc_hd__nor2_1_236/B sky130_fd_sc_hd__o21a_1_50/A1
+ sky130_fd_sc_hd__o21a_1_51/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_247 sky130_fd_sc_hd__or3_1_4/C sky130_fd_sc_hd__nor2_1_247/Y
+ sky130_fd_sc_hd__or3_1_4/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_258 sky130_fd_sc_hd__nor2_1_268/A sky130_fd_sc_hd__nor2_1_258/Y
+ sky130_fd_sc_hd__nor2_1_258/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_269 sky130_fd_sc_hd__nor2_1_303/A sky130_fd_sc_hd__o21a_1_56/A1
+ sky130_fd_sc_hd__o21a_1_57/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_410 sky130_fd_sc_hd__buf_6_69/X sky130_fd_sc_hd__buf_12_410/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_421 sky130_fd_sc_hd__buf_8_205/X sky130_fd_sc_hd__buf_12_421/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_432 sky130_fd_sc_hd__buf_8_212/X sky130_fd_sc_hd__buf_12_432/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_443 sky130_fd_sc_hd__buf_12_443/A sky130_fd_sc_hd__buf_12_443/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_302 sky130_fd_sc_hd__clkbuf_1_378/X sky130_fd_sc_hd__clkbuf_1_379/X
+ sky130_fd_sc_hd__clkbuf_4_167/X sky130_fd_sc_hd__buf_2_191/X sky130_fd_sc_hd__nand4_1_75/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_454 sky130_fd_sc_hd__buf_6_61/X sky130_fd_sc_hd__buf_12_454/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_313 sky130_fd_sc_hd__clkbuf_4_165/X sky130_fd_sc_hd__clkinv_2_23/Y
+ sky130_fd_sc_hd__clkbuf_1_399/X sky130_fd_sc_hd__a22oi_1_313/A2 sky130_fd_sc_hd__a22oi_1_313/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_465 sky130_fd_sc_hd__buf_12_465/A sky130_fd_sc_hd__buf_12_465/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_324 sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_2_7/Y
+ sky130_fd_sc_hd__fa_2_999/A sky130_fd_sc_hd__fa_2_1000/A sky130_fd_sc_hd__o21ai_1_92/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_476 sky130_fd_sc_hd__buf_12_476/A sky130_fd_sc_hd__buf_12_476/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_335 sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_2_7/Y
+ sky130_fd_sc_hd__fa_2_1007/A sky130_fd_sc_hd__fa_2_1008/A sky130_fd_sc_hd__a22oi_1_335/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_487 sky130_fd_sc_hd__buf_12_487/A sky130_fd_sc_hd__buf_12_487/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_346 sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_2_7/Y
+ sky130_fd_sc_hd__fa_2_1001/A sky130_fd_sc_hd__fa_2_1002/A sky130_fd_sc_hd__a22oi_1_346/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_498 sky130_fd_sc_hd__buf_12_498/A sky130_fd_sc_hd__buf_12_498/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_357 sky130_fd_sc_hd__clkinv_1_711/Y sky130_fd_sc_hd__nand2_1_333/B
+ sky130_fd_sc_hd__nand2_1_321/A sky130_fd_sc_hd__o21ai_1_238/Y sky130_fd_sc_hd__a22oi_1_357/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_368 sky130_fd_sc_hd__nor2_4_13/Y sky130_fd_sc_hd__nor2_2_12/Y
+ sky130_fd_sc_hd__fa_2_1082/A sky130_fd_sc_hd__fa_2_1084/A sky130_fd_sc_hd__a22oi_1_368/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_610 sky130_fd_sc_hd__nor2_1_91/B sky130_fd_sc_hd__fa_2_1045/COUT
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_610/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22oi_1_379 sky130_fd_sc_hd__clkinv_1_861/Y sky130_fd_sc_hd__nor3_1_39/B
+ sky130_fd_sc_hd__fa_2_1197/A sky130_fd_sc_hd__fa_2_1198/A sky130_fd_sc_hd__a22oi_1_379/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_621 sky130_fd_sc_hd__nand2_1_331/B sky130_fd_sc_hd__nor2_1_127/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_621/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_632 sky130_fd_sc_hd__o22ai_1_150/B2 sky130_fd_sc_hd__ha_2_199/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_632/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_643 sky130_fd_sc_hd__o22ai_1_161/B2 sky130_fd_sc_hd__ha_2_188/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_643/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_654 sky130_fd_sc_hd__nor2_1_95/B sky130_fd_sc_hd__nand2_1_304/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_654/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_665 sky130_fd_sc_hd__clkinv_1_665/Y sky130_fd_sc_hd__nor2_1_94/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_665/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_676 sky130_fd_sc_hd__nor2_1_106/B sky130_fd_sc_hd__fa_2_1108/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_676/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_687 sky130_fd_sc_hd__nor2_1_99/B sky130_fd_sc_hd__fa_2_1119/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_687/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_698 sky130_fd_sc_hd__clkinv_1_698/Y sky130_fd_sc_hd__a21oi_1_204/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_698/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand3_1_5 sky130_fd_sc_hd__nand3_1_5/Y sky130_fd_sc_hd__nand3_1_5/A
+ sky130_fd_sc_hd__nand3_1_5/C sky130_fd_sc_hd__nand3_1_5/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__a222oi_1_30 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1259/A sky130_fd_sc_hd__nor2_2_17/Y
+ sky130_fd_sc_hd__nor3_1_40/A sky130_fd_sc_hd__xor2_1_253/A sky130_fd_sc_hd__nor2_4_18/B
+ sky130_fd_sc_hd__a222oi_1_30/Y sky130_fd_sc_hd__fa_2_1258/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_41 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1297/A sky130_fd_sc_hd__nor2_2_18/Y
+ sky130_fd_sc_hd__nor3_1_41/A sky130_fd_sc_hd__fa_2_1299/A sky130_fd_sc_hd__nor3_1_41/B
+ sky130_fd_sc_hd__a222oi_1_41/Y sky130_fd_sc_hd__fa_2_1296/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_10 VSS VDD sky130_fd_sc_hd__xor2_1_15/X sky130_fd_sc_hd__xnor2_1_10/Y
+ sky130_fd_sc_hd__xnor2_1_10/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_21 VSS VDD sky130_fd_sc_hd__nor2_1_22/B sky130_fd_sc_hd__xor2_1_20/B
+ sky130_fd_sc_hd__nor2_1_22/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_32 VSS VDD sky130_fd_sc_hd__xor2_1_31/X sky130_fd_sc_hd__xnor2_1_32/Y
+ sky130_fd_sc_hd__xnor2_1_32/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_43 VSS VDD sky130_fd_sc_hd__xnor2_1_44/B sky130_fd_sc_hd__xnor2_1_43/Y
+ sky130_fd_sc_hd__xnor2_1_43/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_54 VSS VDD sky130_fd_sc_hd__xnor2_1_54/B sky130_fd_sc_hd__xnor2_1_54/Y
+ sky130_fd_sc_hd__nor2_1_47/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_65 VSS VDD sky130_fd_sc_hd__xnor2_1_65/B sky130_fd_sc_hd__xnor2_1_65/Y
+ sky130_fd_sc_hd__xnor2_1_65/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_76 VSS VDD sky130_fd_sc_hd__xnor2_1_77/B sky130_fd_sc_hd__xnor2_1_76/Y
+ sky130_fd_sc_hd__xnor2_1_76/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_87 VSS VDD sky130_fd_sc_hd__xnor2_1_87/B sky130_fd_sc_hd__xnor2_1_87/Y
+ sky130_fd_sc_hd__nor2_1_98/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_98 VSS VDD sky130_fd_sc_hd__xnor2_1_98/B sky130_fd_sc_hd__xnor2_1_98/Y
+ sky130_fd_sc_hd__fa_2_1259/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__a211oi_1_1 sky130_fd_sc_hd__fa_2_946/A sky130_fd_sc_hd__o21ai_1_35/Y
+ sky130_fd_sc_hd__nor3_1_34/C sky130_fd_sc_hd__nand4_1_84/B sky130_fd_sc_hd__nor3_1_34/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o32ai_1_4 sky130_fd_sc_hd__o32ai_1_4/A2 sky130_fd_sc_hd__o32ai_1_4/Y
+ sky130_fd_sc_hd__fa_2_1193/A sky130_fd_sc_hd__o32ai_1_4/A3 sky130_fd_sc_hd__o32ai_1_4/B2
+ sky130_fd_sc_hd__fa_2_1192/A VDD VSS VSS VDD sky130_fd_sc_hd__o32ai_1
Xsky130_fd_sc_hd__clkbuf_16_2 sky130_fd_sc_hd__buf_12_111/A sky130_fd_sc_hd__buf_8_14/X
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__fa_2_290 sky130_fd_sc_hd__fa_2_288/CIN sky130_fd_sc_hd__nor2_1_209/A
+ sky130_fd_sc_hd__fa_2_290/A sky130_fd_sc_hd__fa_2_290/B sky130_fd_sc_hd__fa_2_290/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor4_1_2 sky130_fd_sc_hd__or4_1_0/X sky130_fd_sc_hd__or4_1_1/X sky130_fd_sc_hd__nor4_1_2/Y
+ sky130_fd_sc_hd__nor4_1_2/A sky130_fd_sc_hd__nor4_1_2/B VDD VSS VSS VDD sky130_fd_sc_hd__nor4_1
Xsky130_fd_sc_hd__a22oi_1_1 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__a22oi_1_9/A1
+ sky130_fd_sc_hd__dfxtp_1_77/D sky130_fd_sc_hd__a22o_1_9/A1 sky130_fd_sc_hd__nand3_1_0/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__diode_2_140 sky130_fd_sc_hd__clkbuf_1_526/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_151 sky130_fd_sc_hd__buf_2_206/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_162 sky130_fd_sc_hd__nand4_1_67/D VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_173 sky130_fd_sc_hd__nand4_1_65/D VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_184 sky130_fd_sc_hd__buf_2_140/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_195 sky130_fd_sc_hd__clkbuf_1_527/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkinv_2_17 sky130_fd_sc_hd__clkinv_2_17/Y sky130_fd_sc_hd__clkinv_8_15/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_17/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkbuf_4_204 sky130_fd_sc_hd__buf_12_402/A sky130_fd_sc_hd__buf_6_58/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_2_28 sky130_fd_sc_hd__nand4_1_67/D sky130_fd_sc_hd__clkinv_2_28/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_28/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkbuf_4_215 sky130_fd_sc_hd__nand2_1_566/B sky130_fd_sc_hd__buf_4_66/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_2_39 sky130_fd_sc_hd__clkinv_4_29/A sky130_fd_sc_hd__clkinv_4_59/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_39/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkbuf_4_226 freq_eval_done sky130_fd_sc_hd__nor2_1_2/A VSS VDD
+ VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_12_240 sky130_fd_sc_hd__buf_12_240/A sky130_fd_sc_hd__buf_12_240/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_251 sky130_fd_sc_hd__buf_12_251/A sky130_fd_sc_hd__buf_12_251/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_110 sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__a22oi_2_12/A1
+ sky130_fd_sc_hd__buf_2_75/X sky130_fd_sc_hd__clkbuf_1_166/X sky130_fd_sc_hd__a22oi_1_110/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_262 sky130_fd_sc_hd__buf_12_262/A sky130_fd_sc_hd__buf_12_262/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_121 sky130_fd_sc_hd__a22oi_1_97/B1 sky130_fd_sc_hd__a22oi_1_97/A1
+ sky130_fd_sc_hd__buf_2_56/X sky130_fd_sc_hd__clkbuf_4_80/X sky130_fd_sc_hd__nand4_1_25/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_273 sky130_fd_sc_hd__inv_2_81/Y sky130_fd_sc_hd__buf_12_273/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_132 sky130_fd_sc_hd__a22oi_1_97/B1 sky130_fd_sc_hd__a22oi_1_97/A1
+ sky130_fd_sc_hd__buf_2_53/X sky130_fd_sc_hd__clkbuf_4_77/X sky130_fd_sc_hd__nand4_1_28/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_284 sky130_fd_sc_hd__inv_2_99/Y sky130_fd_sc_hd__buf_12_284/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_143 sky130_fd_sc_hd__a22oi_1_96/B1 sky130_fd_sc_hd__a22oi_1_96/A1
+ sky130_fd_sc_hd__clkbuf_1_139/X sky130_fd_sc_hd__a22oi_1_143/A2 sky130_fd_sc_hd__nand4_1_31/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_295 sky130_fd_sc_hd__buf_8_158/X sky130_fd_sc_hd__buf_12_367/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_154 sky130_fd_sc_hd__clkbuf_1_264/X sky130_fd_sc_hd__nor2_2_3/Y
+ sky130_fd_sc_hd__a22oi_1_154/B2 sky130_fd_sc_hd__clkbuf_4_136/X sky130_fd_sc_hd__nand4_1_33/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_165 sky130_fd_sc_hd__clkbuf_4_111/X sky130_fd_sc_hd__clkbuf_4_112/X
+ sky130_fd_sc_hd__a22oi_1_165/B2 sky130_fd_sc_hd__clkbuf_1_293/X sky130_fd_sc_hd__a22oi_1_165/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_176 sky130_fd_sc_hd__clkbuf_1_351/X sky130_fd_sc_hd__clkbuf_1_353/X
+ sky130_fd_sc_hd__clkinv_2_11/Y sky130_fd_sc_hd__a22oi_1_176/A2 sky130_fd_sc_hd__nand4_1_39/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_187 sky130_fd_sc_hd__clkbuf_1_265/X sky130_fd_sc_hd__clkbuf_1_266/X
+ sky130_fd_sc_hd__clkbuf_1_272/X sky130_fd_sc_hd__a22oi_1_187/A2 sky130_fd_sc_hd__a22oi_1_187/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_198 sky130_fd_sc_hd__clkbuf_1_264/X sky130_fd_sc_hd__nor2_2_3/Y
+ sky130_fd_sc_hd__a22oi_1_198/B2 sky130_fd_sc_hd__clkbuf_4_125/X sky130_fd_sc_hd__nand4_1_44/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_440 sky130_fd_sc_hd__fa_2_964/B sky130_fd_sc_hd__nor2b_1_88/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_440/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_2_10 sky130_fd_sc_hd__or2_1_1/B sky130_fd_sc_hd__ha_2_87/A
+ sky130_fd_sc_hd__buf_2_161/A sky130_fd_sc_hd__a22o_2_10/B2 sky130_fd_sc_hd__a22o_4_0/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_2
Xsky130_fd_sc_hd__clkinv_1_451 sky130_fd_sc_hd__fa_2_950/B sky130_fd_sc_hd__dfxtp_1_498/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_451/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_462 sky130_fd_sc_hd__a21oi_1_94/A1 sky130_fd_sc_hd__nor2_1_82/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_462/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_473 sky130_fd_sc_hd__o22ai_1_78/B2 sky130_fd_sc_hd__ha_2_181/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_473/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_484 sky130_fd_sc_hd__o21ai_1_71/A2 sky130_fd_sc_hd__ha_2_170/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_484/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_495 sky130_fd_sc_hd__nor2_1_44/B sky130_fd_sc_hd__nand2_1_246/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_495/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_409 VSS VDD sky130_fd_sc_hd__nor2_1_228/B sky130_fd_sc_hd__o21a_1_55/A1
+ sky130_fd_sc_hd__a21oi_1_394/Y sky130_fd_sc_hd__o21ai_1_409/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a21oi_1_370 sky130_fd_sc_hd__o21a_1_51/B1 sky130_fd_sc_hd__o21a_1_50/A1
+ sky130_fd_sc_hd__a21oi_1_370/Y sky130_fd_sc_hd__nor2_1_236/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_381 sky130_fd_sc_hd__nor2_2_17/Y sky130_fd_sc_hd__o21ai_1_394/Y
+ sky130_fd_sc_hd__nor2_1_250/B sky130_fd_sc_hd__fa_2_1229/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_392 sky130_fd_sc_hd__or2_0_11/B sky130_fd_sc_hd__o21ai_1_407/Y
+ sky130_fd_sc_hd__a21oi_1_392/Y sky130_fd_sc_hd__clkinv_1_990/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nor2_4_18 sky130_fd_sc_hd__nor3_1_40/A sky130_fd_sc_hd__nor2_4_18/A
+ sky130_fd_sc_hd__nor2_4_18/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__xor2_1_203 sky130_fd_sc_hd__fa_2_1173/A sky130_fd_sc_hd__fa_2_1176/B
+ sky130_fd_sc_hd__xor2_1_203/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_214 sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__fa_2_1204/B
+ sky130_fd_sc_hd__xor2_1_214/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_225 sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__fa_2_1193/B
+ sky130_fd_sc_hd__xor2_1_225/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_236 sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1239/B
+ sky130_fd_sc_hd__xor2_1_236/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_247 sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1228/B
+ sky130_fd_sc_hd__xor2_1_247/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_258 sky130_fd_sc_hd__xor2_1_267/B sky130_fd_sc_hd__fa_2_1256/B
+ sky130_fd_sc_hd__xor2_1_258/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_609 VDD VSS sky130_fd_sc_hd__and2_0_234/A sky130_fd_sc_hd__dfxtp_1_611/CLK
+ sky130_fd_sc_hd__fa_2_1029/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_269 sky130_fd_sc_hd__fa_2_1242/A sky130_fd_sc_hd__fa_2_1245/B
+ sky130_fd_sc_hd__xor2_1_269/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_207 VSS VDD sky130_fd_sc_hd__buf_8_109/A sky130_fd_sc_hd__clkbuf_1_230/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_218 VSS VDD sky130_fd_sc_hd__buf_8_93/A sky130_fd_sc_hd__buf_8_67/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_229 VSS VDD sky130_fd_sc_hd__clkbuf_1_230/A sky130_fd_sc_hd__buf_8_73/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_2_30 VDD VSS sky130_fd_sc_hd__inv_2_44/A sky130_fd_sc_hd__buf_8_56/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_41 VDD VSS sky130_fd_sc_hd__buf_2_41/X sky130_fd_sc_hd__buf_2_41/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_52 VDD VSS sky130_fd_sc_hd__buf_2_52/X sky130_fd_sc_hd__buf_2_52/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_63 VDD VSS sky130_fd_sc_hd__buf_2_63/X sky130_fd_sc_hd__buf_2_63/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_74 VDD VSS sky130_fd_sc_hd__buf_2_74/X sky130_fd_sc_hd__buf_2_74/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_85 VDD VSS sky130_fd_sc_hd__buf_2_85/X sky130_fd_sc_hd__buf_2_85/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_96 VDD VSS sky130_fd_sc_hd__buf_2_96/X sky130_fd_sc_hd__buf_2_96/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__diode_2_3 sky130_fd_sc_hd__clkbuf_1_247/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__and2_0_205 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_205/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__ha_2_167/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_216 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_216/X sky130_fd_sc_hd__and2_0_235/B
+ sky130_fd_sc_hd__and2_0_216/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_227 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_227/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_227/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_238 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_238/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__fa_2_876/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_249 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_249/X sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__xnor2_1_28/Y sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_270 sky130_fd_sc_hd__o22ai_1_0/A2 sky130_fd_sc_hd__ha_2_151/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_270/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_2_4 sky130_fd_sc_hd__nor2_4_4/Y sky130_fd_sc_hd__ha_2_71/A
+ sky130_fd_sc_hd__a22o_2_4/X sky130_fd_sc_hd__a22o_2_4/B2 sky130_fd_sc_hd__a22o_2_6/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_2
Xsky130_fd_sc_hd__clkinv_1_281 sky130_fd_sc_hd__fa_2_81/B sky130_fd_sc_hd__ha_2_96/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_281/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o31ai_1_3 sky130_fd_sc_hd__o31ai_1_3/Y sky130_fd_sc_hd__nor4_1_7/A
+ sky130_fd_sc_hd__nor4_1_7/B sky130_fd_sc_hd__xnor2_1_28/B sky130_fd_sc_hd__o31ai_1_3/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__o31ai_1
Xsky130_fd_sc_hd__clkinv_1_292 sky130_fd_sc_hd__fa_2_261/A sky130_fd_sc_hd__fa_2_5/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_292/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_0 sky130_fd_sc_hd__or2_0_0/A sky130_fd_sc_hd__o21ai_1_1/Y
+ sky130_fd_sc_hd__a21oi_1_0/Y sky130_fd_sc_hd__o21ai_1_1/A2 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkbuf_4_13 sky130_fd_sc_hd__clkbuf_4_13/X sky130_fd_sc_hd__clkbuf_4_13/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_206 VSS VDD sky130_fd_sc_hd__nand4_1_86/Y sky130_fd_sc_hd__fa_2_1050/A
+ sky130_fd_sc_hd__fa_2_1051/A sky130_fd_sc_hd__o21ai_1_206/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_24 sky130_fd_sc_hd__clkbuf_4_24/X sky130_fd_sc_hd__clkbuf_4_24/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_217 VSS VDD sky130_fd_sc_hd__nor2_1_130/Y sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__a21oi_1_193/Y sky130_fd_sc_hd__xor2_1_123/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_35 sky130_fd_sc_hd__a22oi_2_7/B2 sky130_fd_sc_hd__clkbuf_4_35/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_228 VSS VDD sky130_fd_sc_hd__o21a_1_16/A2 sky130_fd_sc_hd__nor2_1_113/B
+ sky130_fd_sc_hd__a22oi_1_350/Y sky130_fd_sc_hd__o21ai_1_228/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_46 sky130_fd_sc_hd__nand4_1_11/D sky130_fd_sc_hd__a22oi_1_64/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_239 VSS VDD sky130_fd_sc_hd__nor2_1_118/B sky130_fd_sc_hd__o21a_1_16/A2
+ sky130_fd_sc_hd__a21oi_1_213/Y sky130_fd_sc_hd__o21ai_1_239/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_57 sky130_fd_sc_hd__nand4_1_0/D sky130_fd_sc_hd__a22oi_1_28/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_68 sky130_fd_sc_hd__buf_2_41/A sky130_fd_sc_hd__dfxtp_1_261/Q
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_79 sky130_fd_sc_hd__clkbuf_4_79/X sky130_fd_sc_hd__clkbuf_4_79/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_8_130 sky130_fd_sc_hd__buf_8_130/A sky130_fd_sc_hd__buf_8_130/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_141 sky130_fd_sc_hd__buf_8_141/A sky130_fd_sc_hd__buf_4_80/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_152 sky130_fd_sc_hd__buf_8_152/A sky130_fd_sc_hd__buf_8_152/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nor2_4_3 sky130_fd_sc_hd__nor2_4_3/Y sky130_fd_sc_hd__nor2_4_3/A
+ sky130_fd_sc_hd__inv_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__buf_8_163 sky130_fd_sc_hd__buf_8_163/A sky130_fd_sc_hd__buf_8_163/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_174 sky130_fd_sc_hd__buf_8_174/A sky130_fd_sc_hd__buf_8_174/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_185 sky130_fd_sc_hd__buf_8_185/A sky130_fd_sc_hd__buf_8_185/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_196 sky130_fd_sc_hd__buf_8_196/A sky130_fd_sc_hd__buf_8_196/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_406 VDD VSS sky130_fd_sc_hd__nor2_1_61/A sky130_fd_sc_hd__dfxtp_1_425/CLK
+ sky130_fd_sc_hd__and2_0_118/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_417 VDD VSS sky130_fd_sc_hd__nor2_1_52/A sky130_fd_sc_hd__dfxtp_1_419/CLK
+ sky130_fd_sc_hd__and2_0_142/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_428 VDD VSS sky130_fd_sc_hd__dfxtp_1_428/Q sky130_fd_sc_hd__dfxtp_1_433/CLK
+ sky130_fd_sc_hd__nand2_1_108/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_439 VDD VSS sky130_fd_sc_hd__xnor2_1_99/A sky130_fd_sc_hd__dfxtp_1_452/CLK
+ sky130_fd_sc_hd__nand2_1_86/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a21o_2_20 sky130_fd_sc_hd__a21o_2_20/X sky130_fd_sc_hd__nor2_1_253/Y
+ sky130_fd_sc_hd__nor2_1_253/A sky130_fd_sc_hd__nor2_1_253/B VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__clkinv_8_16 sky130_fd_sc_hd__clkinv_8_16/Y sky130_fd_sc_hd__clkinv_4_9/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_27 sky130_fd_sc_hd__clkinv_8_28/A sky130_fd_sc_hd__clkinv_8_33/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_38 sky130_fd_sc_hd__clkinv_8_38/Y sky130_fd_sc_hd__clkinv_8_38/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_49 sky130_fd_sc_hd__clkinv_8_49/Y sky130_fd_sc_hd__clkinv_8_49/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_49/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_14 sky130_fd_sc_hd__inv_2_27/Y sky130_fd_sc_hd__buf_12_14/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_25 sky130_fd_sc_hd__buf_8_7/X sky130_fd_sc_hd__buf_12_95/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_80 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__fa_2_996/B
+ sky130_fd_sc_hd__xor2_1_80/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_36 sky130_fd_sc_hd__buf_8_36/X sky130_fd_sc_hd__buf_12_98/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_91 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__xor2_1_91/X
+ sky130_fd_sc_hd__xor2_1_91/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_47 sky130_fd_sc_hd__buf_8_6/X sky130_fd_sc_hd__buf_12_47/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_58 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__buf_8_60/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_69 sky130_fd_sc_hd__buf_4_20/X sky130_fd_sc_hd__buf_12_69/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_2_9 VDD VSS sky130_fd_sc_hd__buf_2_9/X sky130_fd_sc_hd__buf_2_9/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1302 VDD VSS sky130_fd_sc_hd__fa_2_849/B sky130_fd_sc_hd__dfxtp_1_1332/CLK
+ sky130_fd_sc_hd__a21oi_1_436/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1313 VDD VSS sky130_fd_sc_hd__fa_2_838/B sky130_fd_sc_hd__dfxtp_1_1329/CLK
+ sky130_fd_sc_hd__o21a_1_63/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1324 VDD VSS sky130_fd_sc_hd__fa_2_908/A sky130_fd_sc_hd__dfxtp_1_1326/CLK
+ sky130_fd_sc_hd__a21oi_1_424/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1335 VDD VSS sky130_fd_sc_hd__fa_2_1294/A sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__and2_0_336/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1346 VDD VSS sky130_fd_sc_hd__fa_2_1305/A sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__mux2_2_232/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1357 VDD VSS sky130_fd_sc_hd__fa_2_1279/A sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__mux2_2_255/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1368 VDD VSS sky130_fd_sc_hd__fa_2_1290/A sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__mux2_2_227/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_940 VDD VSS sky130_fd_sc_hd__fa_2_1132/A sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__mux2_2_94/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1379 VDD VSS sky130_fd_sc_hd__fa_2_1318/A sky130_fd_sc_hd__clkinv_8_63/Y
+ sky130_fd_sc_hd__mux2_2_256/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_951 VDD VSS sky130_fd_sc_hd__fa_2_1160/A sky130_fd_sc_hd__clkinv_8_63/Y
+ sky130_fd_sc_hd__mux2_2_121/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_962 VDD VSS sky130_fd_sc_hd__fa_2_1171/A sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__nand2_1_361/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_973 VDD VSS sky130_fd_sc_hd__mux2_2_111/A0 sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__o22ai_1_222/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_984 VDD VSS sky130_fd_sc_hd__mux2_2_83/A1 sky130_fd_sc_hd__clkinv_8_46/Y
+ sky130_fd_sc_hd__o22ai_1_211/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_995 VDD VSS sky130_fd_sc_hd__mux2_2_112/A0 sky130_fd_sc_hd__clkinv_8_64/Y
+ sky130_fd_sc_hd__dfxtp_1_995/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_560 VSS VDD sky130_fd_sc_hd__nand2_1_93/B sky130_fd_sc_hd__nand4_1_58/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_571 VSS VDD sky130_fd_sc_hd__dfxtp_1_77/D sky130_fd_sc_hd__nand4_1_47/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_582 VSS VDD sky130_fd_sc_hd__nand3_1_9/B sky130_fd_sc_hd__a22oi_1_18/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_150 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_150/A sky130_fd_sc_hd__ha_2_149/B
+ sky130_fd_sc_hd__ha_2_150/SUM sky130_fd_sc_hd__ha_2_150/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_593 VSS VDD sky130_fd_sc_hd__clkbuf_4_227/A sky130_fd_sc_hd__dfxtp_1_1456/Q
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_801 sky130_fd_sc_hd__fa_2_803/CIN sky130_fd_sc_hd__fa_2_796/B
+ sky130_fd_sc_hd__ha_2_145/A sky130_fd_sc_hd__fa_2_801/B sky130_fd_sc_hd__ha_2_141/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_161 VSS VDD VSS VDD sky130_fd_sc_hd__nor4_1_2/A sky130_fd_sc_hd__ha_2_160/B
+ sky130_fd_sc_hd__ha_2_161/SUM sky130_fd_sc_hd__ha_2_161/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_812 sky130_fd_sc_hd__fa_2_813/B sky130_fd_sc_hd__fa_2_805/A
+ sky130_fd_sc_hd__ha_2_145/A sky130_fd_sc_hd__fa_2_812/B sky130_fd_sc_hd__fa_2_833/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_172 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_172/A sky130_fd_sc_hd__ha_2_171/A
+ sky130_fd_sc_hd__ha_2_172/SUM sky130_fd_sc_hd__ha_2_172/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_823 sky130_fd_sc_hd__fa_2_822/CIN sky130_fd_sc_hd__fa_2_823/SUM
+ sky130_fd_sc_hd__fa_2_832/A sky130_fd_sc_hd__fa_2_823/B sky130_fd_sc_hd__fa_2_829/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_183 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_183/A sky130_fd_sc_hd__ha_2_182/A
+ sky130_fd_sc_hd__ha_2_183/SUM sky130_fd_sc_hd__ha_2_183/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_834 sky130_fd_sc_hd__fa_2_704/A sky130_fd_sc_hd__fa_2_705/B
+ sky130_fd_sc_hd__fa_2_834/A sky130_fd_sc_hd__fa_2_834/B sky130_fd_sc_hd__fa_2_834/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_194 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_194/A sky130_fd_sc_hd__ha_2_193/A
+ sky130_fd_sc_hd__ha_2_194/SUM sky130_fd_sc_hd__ha_2_194/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_845 sky130_fd_sc_hd__fa_2_844/CIN sky130_fd_sc_hd__fa_2_845/SUM
+ sky130_fd_sc_hd__fa_2_845/A sky130_fd_sc_hd__fa_2_845/B sky130_fd_sc_hd__fa_2_845/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_856 sky130_fd_sc_hd__fa_2_855/CIN sky130_fd_sc_hd__fa_2_856/SUM
+ sky130_fd_sc_hd__fa_2_856/A sky130_fd_sc_hd__fa_2_856/B sky130_fd_sc_hd__fa_2_856/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_867 sky130_fd_sc_hd__fa_2_866/CIN sky130_fd_sc_hd__fa_2_867/SUM
+ sky130_fd_sc_hd__fa_2_867/A sky130_fd_sc_hd__fa_2_867/B sky130_fd_sc_hd__fa_2_867/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_878 sky130_fd_sc_hd__xor2_1_16/B sky130_fd_sc_hd__nand2_1_38/B
+ sky130_fd_sc_hd__ha_2_149/A sky130_fd_sc_hd__fa_2_878/B sky130_fd_sc_hd__fa_2_878/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_889 sky130_fd_sc_hd__fa_2_888/CIN sky130_fd_sc_hd__fa_2_889/SUM
+ sky130_fd_sc_hd__fa_2_889/A sky130_fd_sc_hd__fa_2_889/B sky130_fd_sc_hd__fa_2_889/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__inv_2_9 sky130_fd_sc_hd__inv_2_9/A sky130_fd_sc_hd__inv_2_9/Y VDD
+ VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__mux2_2_101 VSS VDD sky130_fd_sc_hd__mux2_2_101/A1 sky130_fd_sc_hd__mux2_2_101/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_101/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_112 VSS VDD sky130_fd_sc_hd__mux2_2_112/A1 sky130_fd_sc_hd__mux2_2_112/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_112/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__nor2_1_19 sky130_fd_sc_hd__xor2_1_9/A sky130_fd_sc_hd__xor2_1_21/B
+ sky130_fd_sc_hd__nor4_1_4/C VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__mux2_2_123 VSS VDD sky130_fd_sc_hd__mux2_2_123/A1 sky130_fd_sc_hd__mux2_2_123/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_123/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_134 VSS VDD sky130_fd_sc_hd__mux2_2_134/A1 sky130_fd_sc_hd__mux2_2_134/A0
+ sky130_fd_sc_hd__mux2_2_135/S sky130_fd_sc_hd__mux2_2_134/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_145 VSS VDD sky130_fd_sc_hd__mux2_2_145/A1 sky130_fd_sc_hd__mux2_2_145/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_145/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_156 VSS VDD sky130_fd_sc_hd__mux2_2_156/A1 sky130_fd_sc_hd__mux2_2_156/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_156/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_167 VSS VDD sky130_fd_sc_hd__mux2_2_167/A1 sky130_fd_sc_hd__mux2_2_167/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_167/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_178 VSS VDD sky130_fd_sc_hd__mux2_2_178/A1 sky130_fd_sc_hd__mux2_2_178/A0
+ sky130_fd_sc_hd__nor2_8_1/A sky130_fd_sc_hd__mux2_2_178/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_189 VSS VDD sky130_fd_sc_hd__mux2_2_189/A1 sky130_fd_sc_hd__mux2_2_189/A0
+ sky130_fd_sc_hd__inv_2_139/Y sky130_fd_sc_hd__mux2_2_189/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__and2_0_30 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_30/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_31/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_310 sky130_fd_sc_hd__o22ai_1_318/A2 sky130_fd_sc_hd__o21a_1_42/A2
+ sky130_fd_sc_hd__o22ai_1_310/Y sky130_fd_sc_hd__nor2_1_195/B sky130_fd_sc_hd__o32ai_1_5/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_41 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_58/A sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__ha_2_56/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_105 sky130_fd_sc_hd__maj3_1_106/X sky130_fd_sc_hd__maj3_1_105/X
+ sky130_fd_sc_hd__o22ai_1_32/Y sky130_fd_sc_hd__maj3_1_105/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_321 sky130_fd_sc_hd__o32ai_1_5/A3 sky130_fd_sc_hd__nor2_1_196/B
+ sky130_fd_sc_hd__o22ai_1_321/Y sky130_fd_sc_hd__o22ai_1_321/A1 sky130_fd_sc_hd__o21a_1_42/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_52 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_52/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_52/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_116 sky130_fd_sc_hd__maj3_1_117/X sky130_fd_sc_hd__maj3_1_116/X
+ sky130_fd_sc_hd__maj3_1_116/B sky130_fd_sc_hd__maj3_1_116/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_332 sky130_fd_sc_hd__nand2_1_462/Y sky130_fd_sc_hd__nand2_1_461/Y
+ sky130_fd_sc_hd__o22ai_1_332/Y sky130_fd_sc_hd__nand2_1_475/B sky130_fd_sc_hd__o21ai_1_389/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_63 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_82/A sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__ha_2_70/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_127 sky130_fd_sc_hd__maj3_1_128/X sky130_fd_sc_hd__maj3_1_127/X
+ sky130_fd_sc_hd__maj3_1_127/B sky130_fd_sc_hd__maj3_1_127/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_343 sky130_fd_sc_hd__nand2_1_464/Y sky130_fd_sc_hd__nand2_1_463/Y
+ sky130_fd_sc_hd__o22ai_1_343/Y sky130_fd_sc_hd__nand2_1_474/B sky130_fd_sc_hd__o21ai_1_388/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_74 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_74/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__and2_0_74/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_138 sky130_fd_sc_hd__maj3_1_139/X sky130_fd_sc_hd__maj3_1_138/X
+ sky130_fd_sc_hd__maj3_1_138/B sky130_fd_sc_hd__maj3_1_138/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_407 sky130_fd_sc_hd__nor2_1_199/A sky130_fd_sc_hd__fa_2_1193/A
+ sky130_fd_sc_hd__fa_2_1192/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_354 sky130_fd_sc_hd__o32ai_1_6/B2 sky130_fd_sc_hd__nor2_1_267/A
+ sky130_fd_sc_hd__o22ai_1_354/Y sky130_fd_sc_hd__o22ai_1_376/A1 sky130_fd_sc_hd__a222oi_1_25/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_2_0 sky130_fd_sc_hd__nor2_2_0/B sky130_fd_sc_hd__nor2_2_0/Y
+ sky130_fd_sc_hd__nor4_1_0/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__and2_0_85 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_85/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__xnor2_1_4/Y sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_418 sky130_fd_sc_hd__nand2_1_418/Y sky130_fd_sc_hd__o31ai_1_8/A3
+ sky130_fd_sc_hd__o31ai_1_8/A2 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_149 sky130_fd_sc_hd__maj3_1_150/X sky130_fd_sc_hd__maj3_1_149/X
+ sky130_fd_sc_hd__maj3_1_149/B sky130_fd_sc_hd__maj3_1_149/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_365 sky130_fd_sc_hd__o32ai_1_8/A3 sky130_fd_sc_hd__nor2_1_231/B
+ sky130_fd_sc_hd__o22ai_1_365/Y sky130_fd_sc_hd__o22ai_1_365/A1 sky130_fd_sc_hd__o21a_1_55/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_96 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_96/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_96/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_429 sky130_fd_sc_hd__nand2_1_429/Y sky130_fd_sc_hd__nand2_1_439/B
+ sky130_fd_sc_hd__o21ai_1_362/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_376 sky130_fd_sc_hd__nor2_1_242/B sky130_fd_sc_hd__nor2_1_267/A
+ sky130_fd_sc_hd__o22ai_1_376/Y sky130_fd_sc_hd__o22ai_1_376/A1 sky130_fd_sc_hd__a222oi_1_33/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_387 sky130_fd_sc_hd__nand2_1_514/Y sky130_fd_sc_hd__nand2_1_513/Y
+ sky130_fd_sc_hd__o22ai_1_387/Y sky130_fd_sc_hd__nand2_1_526/B sky130_fd_sc_hd__o21ai_1_442/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_398 sky130_fd_sc_hd__nand2_1_516/Y sky130_fd_sc_hd__nand2_1_515/Y
+ sky130_fd_sc_hd__o22ai_1_398/Y sky130_fd_sc_hd__nand2_1_525/B sky130_fd_sc_hd__o21ai_1_441/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_8_40 sky130_fd_sc_hd__buf_8_40/A sky130_fd_sc_hd__buf_8_40/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__clkinv_1_1009 sky130_fd_sc_hd__o22ai_1_372/B1 sky130_fd_sc_hd__fa_2_1252/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1009/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_51 sky130_fd_sc_hd__ha_2_12/A sky130_fd_sc_hd__buf_8_51/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_62 sky130_fd_sc_hd__buf_8_62/A sky130_fd_sc_hd__buf_8_62/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_73 sky130_fd_sc_hd__ha_2_45/A sky130_fd_sc_hd__buf_8_73/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_84 sky130_fd_sc_hd__buf_8_84/A sky130_fd_sc_hd__buf_8_84/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_203 VDD VSS sky130_fd_sc_hd__ha_2_78/A sky130_fd_sc_hd__dfxtp_1_207/CLK
+ sky130_fd_sc_hd__and2_0_75/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_8_95 sky130_fd_sc_hd__buf_8_95/A sky130_fd_sc_hd__buf_8_95/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_214 VDD VSS sky130_fd_sc_hd__ha_2_89/A sky130_fd_sc_hd__dfxtp_1_224/CLK
+ sky130_fd_sc_hd__nor2b_1_42/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_225 VDD VSS sky130_fd_sc_hd__nor3_2_9/A sky130_fd_sc_hd__clkinv_4_20/Y
+ sky130_fd_sc_hd__buf_2_240/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_236 VDD VSS sky130_fd_sc_hd__fa_2_873/A sky130_fd_sc_hd__dfxtp_1_462/CLK
+ sky130_fd_sc_hd__and2_0_165/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_247 VDD VSS sky130_fd_sc_hd__buf_4_32/A sky130_fd_sc_hd__dfxtp_1_258/CLK
+ sky130_fd_sc_hd__and2_0_189/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_258 VDD VSS sky130_fd_sc_hd__dfxtp_1_258/Q sky130_fd_sc_hd__dfxtp_1_258/CLK
+ sky130_fd_sc_hd__and2_0_221/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_269 VDD VSS sky130_fd_sc_hd__dfxtp_1_269/Q sky130_fd_sc_hd__dfxtp_1_277/CLK
+ sky130_fd_sc_hd__and2_0_215/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_108 sky130_fd_sc_hd__fa_2_110/CIN sky130_fd_sc_hd__fa_2_103/A
+ sky130_fd_sc_hd__fa_2_66/B sky130_fd_sc_hd__fa_2_108/B sky130_fd_sc_hd__fa_2_14/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_119 sky130_fd_sc_hd__fa_2_120/CIN sky130_fd_sc_hd__fa_2_114/A
+ sky130_fd_sc_hd__fa_2_80/B sky130_fd_sc_hd__fa_2_87/B sky130_fd_sc_hd__fa_2_66/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_103 VDD VSS sky130_fd_sc_hd__buf_2_103/X sky130_fd_sc_hd__buf_2_103/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__fa_2_1302 sky130_fd_sc_hd__fa_2_1303/CIN sky130_fd_sc_hd__mux2_2_239/A1
+ sky130_fd_sc_hd__fa_2_1302/A sky130_fd_sc_hd__fa_2_1302/B sky130_fd_sc_hd__fa_2_1302/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_114 VDD VSS sky130_fd_sc_hd__buf_4_37/A sky130_fd_sc_hd__buf_2_116/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__fa_2_1313 sky130_fd_sc_hd__fa_2_1314/CIN sky130_fd_sc_hd__mux2_2_265/A1
+ sky130_fd_sc_hd__fa_2_1313/A sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1313/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_125 VDD VSS sky130_fd_sc_hd__buf_2_125/X sky130_fd_sc_hd__nand3_4_0/Y
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_18 sky130_fd_sc_hd__fa_2_238/B sky130_fd_sc_hd__fa_2_261/A
+ sky130_fd_sc_hd__fa_2_260/B sky130_fd_sc_hd__fa_2_5/A sky130_fd_sc_hd__fa_2_2/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_1324 sky130_fd_sc_hd__fa_2_1325/CIN sky130_fd_sc_hd__nand2_1_518/A
+ sky130_fd_sc_hd__fa_2_1324/A sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1324/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_136 VDD VSS sky130_fd_sc_hd__buf_8_124/A sky130_fd_sc_hd__a22o_2_2/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_29 sky130_fd_sc_hd__fa_2_286/B sky130_fd_sc_hd__fa_2_417/B
+ sky130_fd_sc_hd__fa_2_321/A sky130_fd_sc_hd__ha_2_112/A sky130_fd_sc_hd__ha_2_116/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_2_147 VDD VSS sky130_fd_sc_hd__buf_2_147/X sky130_fd_sc_hd__buf_2_147/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_158 VDD VSS sky130_fd_sc_hd__buf_2_246/A sky130_fd_sc_hd__buf_2_158/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1110 VDD VSS sky130_fd_sc_hd__nor3_1_39/C sky130_fd_sc_hd__clkinv_4_23/Y
+ sky130_fd_sc_hd__o21bai_1_3/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_2_169 VDD VSS sky130_fd_sc_hd__buf_2_169/X sky130_fd_sc_hd__buf_2_169/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1121 VDD VSS sky130_fd_sc_hd__mux2_2_139/A0 sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__o22ai_1_272/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1132 VDD VSS sky130_fd_sc_hd__mux2_2_168/A0 sky130_fd_sc_hd__clkinv_8_64/Y
+ sky130_fd_sc_hd__dfxtp_1_991/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1143 VDD VSS sky130_fd_sc_hd__mux2_2_164/A0 sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__nor2_1_201/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1154 VDD VSS sky130_fd_sc_hd__mux2_2_134/A1 sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__o22ai_1_283/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1165 VDD VSS sky130_fd_sc_hd__fa_2_859/B sky130_fd_sc_hd__dfxtp_1_1180/CLK
+ sky130_fd_sc_hd__a21oi_1_373/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1176 VDD VSS sky130_fd_sc_hd__fa_2_930/B sky130_fd_sc_hd__dfxtp_1_1179/CLK
+ sky130_fd_sc_hd__o32ai_1_6/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1187 VDD VSS sky130_fd_sc_hd__fa_2_940/A sky130_fd_sc_hd__clkinv_4_24/Y
+ sky130_fd_sc_hd__a21oi_1_362/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1198 VDD VSS sky130_fd_sc_hd__fa_2_1247/A sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__mux2_2_203/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_770 VDD VSS sky130_fd_sc_hd__fa_2_1069/B sky130_fd_sc_hd__clkinv_8_54/Y
+ sky130_fd_sc_hd__and2_0_302/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__ha_2_3 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_3/A sky130_fd_sc_hd__ha_2_2/B
+ sky130_fd_sc_hd__ha_2_3/SUM sky130_fd_sc_hd__ha_2_3/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__dfxtp_1_781 VDD VSS sky130_fd_sc_hd__fa_2_1080/A sky130_fd_sc_hd__clkinv_8_55/Y
+ sky130_fd_sc_hd__mux2_2_62/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_792 VDD VSS sky130_fd_sc_hd__fa_2_1091/A sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__mux2_2_39/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_390 VSS VDD sky130_fd_sc_hd__clkbuf_1_390/X sky130_fd_sc_hd__clkbuf_1_390/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_14 VSS VDD sky130_fd_sc_hd__buf_4_11/A sky130_fd_sc_hd__clkbuf_4_7/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_620 sky130_fd_sc_hd__fa_2_621/CIN sky130_fd_sc_hd__fa_2_615/B
+ sky130_fd_sc_hd__fa_2_698/A sky130_fd_sc_hd__fa_2_700/B sky130_fd_sc_hd__ha_2_128/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_25 VSS VDD sky130_fd_sc_hd__clkbuf_1_25/X sky130_fd_sc_hd__clkbuf_1_25/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_631 sky130_fd_sc_hd__fa_2_632/A sky130_fd_sc_hd__fa_2_627/B
+ sky130_fd_sc_hd__fa_2_686/B sky130_fd_sc_hd__fa_2_677/A sky130_fd_sc_hd__ha_2_131/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_36 VSS VDD sky130_fd_sc_hd__clkbuf_1_36/X sky130_fd_sc_hd__clkbuf_1_36/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_642 sky130_fd_sc_hd__fa_2_645/B sky130_fd_sc_hd__fa_2_642/SUM
+ sky130_fd_sc_hd__fa_2_642/A sky130_fd_sc_hd__fa_2_642/B sky130_fd_sc_hd__fa_2_647/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_47 VSS VDD sky130_fd_sc_hd__clkbuf_1_47/X sky130_fd_sc_hd__clkbuf_1_47/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_653 sky130_fd_sc_hd__fa_2_656/A sky130_fd_sc_hd__fa_2_653/SUM
+ sky130_fd_sc_hd__fa_2_653/A sky130_fd_sc_hd__fa_2_653/B sky130_fd_sc_hd__fa_2_659/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_58 VSS VDD sky130_fd_sc_hd__clkbuf_1_58/X sky130_fd_sc_hd__clkbuf_1_58/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_664 sky130_fd_sc_hd__fa_2_666/CIN sky130_fd_sc_hd__fa_2_660/A
+ sky130_fd_sc_hd__ha_2_129/B sky130_fd_sc_hd__fa_2_664/B sky130_fd_sc_hd__fa_2_664/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_69 VSS VDD sky130_fd_sc_hd__clkbuf_1_69/X sky130_fd_sc_hd__clkbuf_1_69/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_675 sky130_fd_sc_hd__fa_2_578/A sky130_fd_sc_hd__fa_2_579/B
+ sky130_fd_sc_hd__fa_2_675/A sky130_fd_sc_hd__fa_2_675/B sky130_fd_sc_hd__fa_2_681/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_686 sky130_fd_sc_hd__fa_2_685/B sky130_fd_sc_hd__fa_2_681/B
+ sky130_fd_sc_hd__fa_2_699/A sky130_fd_sc_hd__fa_2_686/B sky130_fd_sc_hd__fa_2_677/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_697 sky130_fd_sc_hd__fa_2_696/B sky130_fd_sc_hd__fa_2_694/B
+ sky130_fd_sc_hd__fa_2_701/B sky130_fd_sc_hd__ha_2_135/B sky130_fd_sc_hd__fa_2_659/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22oi_2_17 sky130_fd_sc_hd__nor3_2_7/Y sky130_fd_sc_hd__a22oi_2_17/A2
+ sky130_fd_sc_hd__nor3_2_8/Y sky130_fd_sc_hd__a22oi_2_17/B2 sky130_fd_sc_hd__nand4_1_51/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__a22oi_2_28 sky130_fd_sc_hd__buf_2_165/X sky130_fd_sc_hd__a22oi_2_28/A2
+ sky130_fd_sc_hd__nor2_4_7/Y sky130_fd_sc_hd__a22oi_2_28/B2 sky130_fd_sc_hd__nand4_1_60/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__buf_12_3 sky130_fd_sc_hd__inv_2_7/Y sky130_fd_sc_hd__buf_12_3/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__o22ai_1_140 sky130_fd_sc_hd__nand2_1_284/Y sky130_fd_sc_hd__nand2_2_5/Y
+ sky130_fd_sc_hd__o22ai_1_140/Y sky130_fd_sc_hd__xnor2_1_72/Y sky130_fd_sc_hd__o22ai_1_154/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_204 sky130_fd_sc_hd__nor2_1_23/B sky130_fd_sc_hd__nand2_1_204/B
+ sky130_fd_sc_hd__nor4_1_4/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_803 sky130_fd_sc_hd__o22ai_1_234/A1 sky130_fd_sc_hd__nor2_1_171/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_803/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_151 sky130_fd_sc_hd__nand2_1_338/A sky130_fd_sc_hd__nand2_1_284/Y
+ sky130_fd_sc_hd__o22ai_1_151/Y sky130_fd_sc_hd__xnor2_1_66/Y sky130_fd_sc_hd__o22ai_1_151/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_215 sky130_fd_sc_hd__nor2_1_33/B sky130_fd_sc_hd__nand2_1_215/B
+ sky130_fd_sc_hd__nor2_1_34/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_162 sky130_fd_sc_hd__nand2_1_338/A sky130_fd_sc_hd__nand2_1_284/Y
+ sky130_fd_sc_hd__o22ai_1_162/Y sky130_fd_sc_hd__xnor2_1_88/Y sky130_fd_sc_hd__o22ai_1_162/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_814 sky130_fd_sc_hd__nand2_1_369/B sky130_fd_sc_hd__fa_2_434/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_814/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_226 sky130_fd_sc_hd__nor2_1_77/A sky130_fd_sc_hd__o22ai_1_90/A1
+ sky130_fd_sc_hd__nand2_2_4/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_825 sky130_fd_sc_hd__nor2_1_149/B sky130_fd_sc_hd__fa_2_1125/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_825/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_173 sky130_fd_sc_hd__o22ai_1_173/A2 sky130_fd_sc_hd__a21oi_1_204/Y
+ sky130_fd_sc_hd__o22ai_1_173/Y sky130_fd_sc_hd__nor2_1_126/A sky130_fd_sc_hd__nor2_2_13/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_237 sky130_fd_sc_hd__o21ai_1_81/B1 sky130_fd_sc_hd__nor2_1_62/B
+ sky130_fd_sc_hd__nor2_1_62/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_184 sky130_fd_sc_hd__o21a_1_16/A2 sky130_fd_sc_hd__o22ai_1_184/B1
+ sky130_fd_sc_hd__nor2_1_132/B sky130_fd_sc_hd__nor2_1_115/B sky130_fd_sc_hd__o22ai_1_206/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand4_1_10 sky130_fd_sc_hd__nand4_1_10/C sky130_fd_sc_hd__nand4_1_10/B
+ sky130_fd_sc_hd__nand4_1_10/Y sky130_fd_sc_hd__nand4_1_10/D sky130_fd_sc_hd__nand4_1_10/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__clkinv_1_836 sky130_fd_sc_hd__clkinv_1_836/Y sky130_fd_sc_hd__nand2_1_386/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_836/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_248 sky130_fd_sc_hd__nand2_1_248/Y sky130_fd_sc_hd__nor2_1_51/B
+ sky130_fd_sc_hd__nor2_1_51/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand4_1_21 sky130_fd_sc_hd__nand4_1_21/C sky130_fd_sc_hd__nand4_1_21/B
+ sky130_fd_sc_hd__nand4_1_21/Y sky130_fd_sc_hd__nand4_1_21/D sky130_fd_sc_hd__buf_2_107/X
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__o22ai_1_195 sky130_fd_sc_hd__o22ai_1_206/B1 sky130_fd_sc_hd__o22ai_1_204/B1
+ sky130_fd_sc_hd__nor2_1_135/A sky130_fd_sc_hd__nor2_1_120/A sky130_fd_sc_hd__o22ai_1_195/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_847 sky130_fd_sc_hd__o32ai_1_2/B2 sky130_fd_sc_hd__o32ai_1_2/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_847/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_259 sky130_fd_sc_hd__o22ai_1_90/A2 sky130_fd_sc_hd__nor2_2_8/Y
+ sky130_fd_sc_hd__nor2_1_89/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand4_1_32 sky130_fd_sc_hd__nand4_1_32/C sky130_fd_sc_hd__nand4_1_32/B
+ sky130_fd_sc_hd__nand4_1_32/Y sky130_fd_sc_hd__nand4_1_32/D sky130_fd_sc_hd__nand4_1_32/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__clkinv_1_858 sky130_fd_sc_hd__nor2_2_15/B sky130_fd_sc_hd__nor2_2_14/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_858/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand4_1_43 sky130_fd_sc_hd__nand4_1_43/C sky130_fd_sc_hd__nand4_1_43/B
+ sky130_fd_sc_hd__buf_2_287/A sky130_fd_sc_hd__nand4_1_43/D sky130_fd_sc_hd__nand4_1_43/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__clkinv_1_869 sky130_fd_sc_hd__o32ai_1_3/A3 sky130_fd_sc_hd__fa_2_1174/A
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand4_1_54 sky130_fd_sc_hd__nand4_1_54/C sky130_fd_sc_hd__nand4_1_54/B
+ sky130_fd_sc_hd__nand4_1_54/Y sky130_fd_sc_hd__nand4_1_54/D sky130_fd_sc_hd__nand4_1_54/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_65 sky130_fd_sc_hd__nand4_1_65/C sky130_fd_sc_hd__nand4_1_65/B
+ sky130_fd_sc_hd__nand4_1_65/Y sky130_fd_sc_hd__nand4_1_65/D sky130_fd_sc_hd__nand4_1_65/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_76 sky130_fd_sc_hd__nand4_1_76/C sky130_fd_sc_hd__nand4_1_76/B
+ sky130_fd_sc_hd__nand2_1_3/B sky130_fd_sc_hd__nand4_1_76/D sky130_fd_sc_hd__nand4_1_76/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__conb_1_14 sky130_fd_sc_hd__conb_1_14/LO sky130_fd_sc_hd__conb_1_14/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_25 sky130_fd_sc_hd__conb_1_25/LO sky130_fd_sc_hd__conb_1_25/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__mux2_2_9 VSS VDD sky130_fd_sc_hd__mux2_2_9/A1 sky130_fd_sc_hd__mux2_2_9/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_9/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_80 VSS VDD sky130_fd_sc_hd__mux2_2_80/A1 sky130_fd_sc_hd__mux2_2_80/A0
+ sky130_fd_sc_hd__nor2_4_15/A sky130_fd_sc_hd__mux2_2_80/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_91 VSS VDD sky130_fd_sc_hd__mux2_2_91/A1 sky130_fd_sc_hd__mux2_2_91/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_91/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1110 sky130_fd_sc_hd__fa_2_1111/CIN sky130_fd_sc_hd__fa_2_1110/SUM
+ sky130_fd_sc_hd__fa_2_1110/A sky130_fd_sc_hd__fa_2_1110/B sky130_fd_sc_hd__fa_2_1110/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1121 sky130_fd_sc_hd__fa_2_1121/COUT sky130_fd_sc_hd__a22o_1_72/A2
+ sky130_fd_sc_hd__nor2_2_11/B sky130_fd_sc_hd__fa_2_1121/B sky130_fd_sc_hd__fa_2_1121/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1132 sky130_fd_sc_hd__fa_2_1133/CIN sky130_fd_sc_hd__mux2_2_94/A1
+ sky130_fd_sc_hd__fa_2_1132/A sky130_fd_sc_hd__fa_2_1132/B sky130_fd_sc_hd__fa_2_1132/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1143 sky130_fd_sc_hd__fa_2_1144/CIN sky130_fd_sc_hd__mux2_2_113/A1
+ sky130_fd_sc_hd__fa_2_1143/A sky130_fd_sc_hd__fa_2_1143/B sky130_fd_sc_hd__fa_2_1143/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1154 sky130_fd_sc_hd__fa_2_1155/CIN sky130_fd_sc_hd__mux2_2_84/A0
+ sky130_fd_sc_hd__fa_2_1154/A sky130_fd_sc_hd__fa_2_1154/B sky130_fd_sc_hd__fa_2_1154/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1165 sky130_fd_sc_hd__fa_2_1166/CIN sky130_fd_sc_hd__mux2_2_112/A1
+ sky130_fd_sc_hd__fa_2_1165/A sky130_fd_sc_hd__fa_2_1172/B sky130_fd_sc_hd__fa_2_1165/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1176 sky130_fd_sc_hd__fa_2_1177/CIN sky130_fd_sc_hd__mux2_2_162/A1
+ sky130_fd_sc_hd__fa_2_1176/A sky130_fd_sc_hd__fa_2_1176/B sky130_fd_sc_hd__fa_2_1176/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1187 sky130_fd_sc_hd__fa_2_1188/CIN sky130_fd_sc_hd__mux2_2_133/A0
+ sky130_fd_sc_hd__fa_2_1187/A sky130_fd_sc_hd__fa_2_1187/B sky130_fd_sc_hd__fa_2_1187/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1198 sky130_fd_sc_hd__fa_2_1199/CIN sky130_fd_sc_hd__mux2_2_149/A1
+ sky130_fd_sc_hd__fa_2_1198/A sky130_fd_sc_hd__fa_2_1198/B sky130_fd_sc_hd__fa_2_1198/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o2bb2ai_1_5 sky130_fd_sc_hd__o2bb2ai_1_5/Y sky130_fd_sc_hd__nor2_1_18/Y
+ sky130_fd_sc_hd__ha_2_150/SUM sky130_fd_sc_hd__o21ai_1_31/A1 sky130_fd_sc_hd__o22ai_1_0/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_450 sky130_fd_sc_hd__fa_2_446/A sky130_fd_sc_hd__fa_2_451/A
+ sky130_fd_sc_hd__fa_2_502/B sky130_fd_sc_hd__ha_2_117/B sky130_fd_sc_hd__fa_2_427/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_461 sky130_fd_sc_hd__fa_2_458/CIN sky130_fd_sc_hd__fa_2_462/CIN
+ sky130_fd_sc_hd__fa_2_566/B sky130_fd_sc_hd__fa_2_559/A sky130_fd_sc_hd__fa_2_543/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_472 sky130_fd_sc_hd__fa_2_473/A sky130_fd_sc_hd__fa_2_471/B
+ sky130_fd_sc_hd__ha_2_123/A sky130_fd_sc_hd__fa_2_567/A sky130_fd_sc_hd__fa_2_558/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_483 sky130_fd_sc_hd__fa_2_485/A sky130_fd_sc_hd__fa_2_483/SUM
+ sky130_fd_sc_hd__fa_2_483/A sky130_fd_sc_hd__fa_2_483/B sky130_fd_sc_hd__fa_2_488/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_494 sky130_fd_sc_hd__maj3_1_95/B sky130_fd_sc_hd__maj3_1_96/A
+ sky130_fd_sc_hd__fa_2_494/A sky130_fd_sc_hd__fa_2_494/B sky130_fd_sc_hd__fa_2_495/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor2_1_204 sky130_fd_sc_hd__or3_1_3/C sky130_fd_sc_hd__nor2_1_204/Y
+ sky130_fd_sc_hd__or3_1_3/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_215 sky130_fd_sc_hd__nor2_1_225/A sky130_fd_sc_hd__nor2_1_215/Y
+ sky130_fd_sc_hd__nor2_1_215/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_226 sky130_fd_sc_hd__nor2_1_226/B sky130_fd_sc_hd__fa_2_1242/A
+ sky130_fd_sc_hd__nor2_8_1/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_237 sky130_fd_sc_hd__o21a_1_55/A2 sky130_fd_sc_hd__o21a_1_51/A1
+ sky130_fd_sc_hd__o21a_1_52/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_248 sky130_fd_sc_hd__nor2_1_248/B sky130_fd_sc_hd__nor2_1_248/Y
+ sky130_fd_sc_hd__nor2_1_248/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_259 sky130_fd_sc_hd__nor2_1_259/B sky130_fd_sc_hd__nor2_1_259/Y
+ sky130_fd_sc_hd__nor2_1_268/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_400 sky130_fd_sc_hd__buf_6_61/A sky130_fd_sc_hd__buf_6_62/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_411 sky130_fd_sc_hd__bufbuf_8_7/X sky130_fd_sc_hd__buf_12_411/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_422 sky130_fd_sc_hd__buf_8_193/X sky130_fd_sc_hd__buf_12_494/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_433 sky130_fd_sc_hd__buf_8_212/X sky130_fd_sc_hd__buf_12_512/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_444 sky130_fd_sc_hd__buf_4_114/X sky130_fd_sc_hd__buf_12_499/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_303 sky130_fd_sc_hd__nor2_2_4/Y sky130_fd_sc_hd__clkbuf_1_377/X
+ sky130_fd_sc_hd__a22oi_1_303/B2 sky130_fd_sc_hd__clkbuf_4_181/X sky130_fd_sc_hd__nand4_1_75/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_455 sky130_fd_sc_hd__buf_12_455/A sky130_fd_sc_hd__buf_12_455/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_314 sky130_fd_sc_hd__clkbuf_1_378/X sky130_fd_sc_hd__clkbuf_1_379/X
+ sky130_fd_sc_hd__buf_2_219/X sky130_fd_sc_hd__buf_2_188/X sky130_fd_sc_hd__nand4_1_78/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_466 sky130_fd_sc_hd__buf_6_77/X sky130_fd_sc_hd__buf_12_466/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_325 sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__fa_2_989/A
+ sky130_fd_sc_hd__fa_2_992/A sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__a22oi_1_325/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_477 sky130_fd_sc_hd__buf_12_477/A sky130_fd_sc_hd__buf_12_477/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_336 sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_2_7/Y
+ sky130_fd_sc_hd__fa_2_1013/A sky130_fd_sc_hd__fa_2_1014/A sky130_fd_sc_hd__a22oi_1_336/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_488 sky130_fd_sc_hd__buf_12_488/A sky130_fd_sc_hd__buf_12_488/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_347 sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__nor2_4_13/Y
+ sky130_fd_sc_hd__fa_2_1071/A sky130_fd_sc_hd__fa_2_1072/A sky130_fd_sc_hd__a22oi_1_347/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_499 sky130_fd_sc_hd__buf_12_499/A sky130_fd_sc_hd__buf_12_499/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_358 sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__nor2_2_12/Y
+ sky130_fd_sc_hd__fa_2_1087/A sky130_fd_sc_hd__fa_2_1090/A sky130_fd_sc_hd__a22oi_1_358/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_600 sky130_fd_sc_hd__ha_2_175/B sky130_fd_sc_hd__fa_2_1040/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_600/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22oi_1_369 sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__nor2_4_13/Y
+ sky130_fd_sc_hd__fa_2_1073/A sky130_fd_sc_hd__fa_2_1074/A sky130_fd_sc_hd__a22oi_1_369/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_611 sky130_fd_sc_hd__fa_2_1045/B sky130_fd_sc_hd__nor2_2_6/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_611/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_622 sky130_fd_sc_hd__clkinv_1_622/Y sky130_fd_sc_hd__nor2_1_132/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_622/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_633 sky130_fd_sc_hd__o22ai_1_151/B2 sky130_fd_sc_hd__ha_2_198/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_633/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_644 sky130_fd_sc_hd__o22ai_1_162/B2 sky130_fd_sc_hd__ha_2_187/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_644/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_655 sky130_fd_sc_hd__nand2_1_289/B sky130_fd_sc_hd__nor2_1_108/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_655/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_666 sky130_fd_sc_hd__o21ai_1_196/A1 sky130_fd_sc_hd__nand2_1_298/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_666/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_677 sky130_fd_sc_hd__nor2_1_104/B sky130_fd_sc_hd__fa_2_1109/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_677/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_688 sky130_fd_sc_hd__nor2_1_112/B sky130_fd_sc_hd__fa_2_1120/B
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_699 sky130_fd_sc_hd__o21ai_1_225/A2 sky130_fd_sc_hd__o21a_1_9/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_699/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand3_1_6 sky130_fd_sc_hd__nand3_1_6/Y sky130_fd_sc_hd__nand3_1_6/A
+ sky130_fd_sc_hd__nand3_1_6/C sky130_fd_sc_hd__nand3_1_6/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__a222oi_1_20 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1208/A sky130_fd_sc_hd__nor2_2_16/Y
+ sky130_fd_sc_hd__nor3_1_39/A sky130_fd_sc_hd__xor2_1_208/A sky130_fd_sc_hd__nor2_4_16/B
+ sky130_fd_sc_hd__a222oi_1_20/Y sky130_fd_sc_hd__fa_2_1207/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_31 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1246/A sky130_fd_sc_hd__nor2_2_17/Y
+ sky130_fd_sc_hd__nor3_1_40/A sky130_fd_sc_hd__fa_2_1248/A sky130_fd_sc_hd__nor3_1_40/B
+ sky130_fd_sc_hd__a222oi_1_31/Y sky130_fd_sc_hd__fa_2_1245/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_42 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1296/A sky130_fd_sc_hd__nor2_2_18/Y
+ sky130_fd_sc_hd__nor3_1_41/A sky130_fd_sc_hd__fa_2_1298/A sky130_fd_sc_hd__nor3_1_41/B
+ sky130_fd_sc_hd__nor2_1_306/B sky130_fd_sc_hd__fa_2_1295/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_11 VSS VDD sky130_fd_sc_hd__xor2_1_16/X sky130_fd_sc_hd__xnor2_1_11/Y
+ sky130_fd_sc_hd__nor2_1_9/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_22 VSS VDD sky130_fd_sc_hd__xor2_1_24/X sky130_fd_sc_hd__xor2_1_23/B
+ sky130_fd_sc_hd__xnor2_1_23/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_33 VSS VDD sky130_fd_sc_hd__xnor2_1_33/B sky130_fd_sc_hd__xnor2_1_33/Y
+ sky130_fd_sc_hd__nor2_1_42/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_44 VSS VDD sky130_fd_sc_hd__xnor2_1_44/B sky130_fd_sc_hd__xnor2_1_44/Y
+ sky130_fd_sc_hd__xnor2_1_44/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_55 VSS VDD sky130_fd_sc_hd__xnor2_1_56/B sky130_fd_sc_hd__xnor2_1_55/Y
+ sky130_fd_sc_hd__xnor2_1_55/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_66 VSS VDD sky130_fd_sc_hd__xnor2_1_66/B sky130_fd_sc_hd__xnor2_1_66/Y
+ sky130_fd_sc_hd__nor2_1_93/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_77 VSS VDD sky130_fd_sc_hd__xnor2_1_77/B sky130_fd_sc_hd__xnor2_1_77/Y
+ sky130_fd_sc_hd__xnor2_1_77/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_88 VSS VDD sky130_fd_sc_hd__xnor2_1_89/B sky130_fd_sc_hd__xnor2_1_88/Y
+ sky130_fd_sc_hd__xnor2_1_88/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_99 VSS VDD sky130_fd_sc_hd__xor2_1_275/A sky130_fd_sc_hd__xnor2_1_99/Y
+ sky130_fd_sc_hd__xnor2_1_99/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__a211oi_1_2 sky130_fd_sc_hd__or3_1_0/B sky130_fd_sc_hd__o21ai_1_36/Y
+ sky130_fd_sc_hd__or3_1_0/A sky130_fd_sc_hd__nand4_1_84/A sky130_fd_sc_hd__or3_1_0/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o32ai_1_5 sky130_fd_sc_hd__nor3_1_39/C sky130_fd_sc_hd__o32ai_1_5/Y
+ sky130_fd_sc_hd__o32ai_1_5/A1 sky130_fd_sc_hd__o32ai_1_5/A3 sky130_fd_sc_hd__o32ai_1_5/B2
+ sky130_fd_sc_hd__o32ai_1_5/B1 VDD VSS VSS VDD sky130_fd_sc_hd__o32ai_1
Xsky130_fd_sc_hd__clkbuf_16_3 sky130_fd_sc_hd__buf_12_113/A sky130_fd_sc_hd__buf_6_16/X
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__fa_2_280 sky130_fd_sc_hd__fa_2_279/CIN sky130_fd_sc_hd__fa_2_280/SUM
+ sky130_fd_sc_hd__fa_2_280/A sky130_fd_sc_hd__fa_2_280/B sky130_fd_sc_hd__fa_2_250/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_291 sky130_fd_sc_hd__fa_2_288/A sky130_fd_sc_hd__fa_2_290/A
+ sky130_fd_sc_hd__ha_2_116/A sky130_fd_sc_hd__ha_2_116/B sky130_fd_sc_hd__fa_2_389/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22oi_1_2 sky130_fd_sc_hd__nor2_2_0/Y sky130_fd_sc_hd__clkinv_1_4/Y
+ sky130_fd_sc_hd__nand4_1_30/Y sky130_fd_sc_hd__nand4_1_14/Y sky130_fd_sc_hd__a22oi_1_2/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor4_1_3 sky130_fd_sc_hd__nor4_1_3/D sky130_fd_sc_hd__nor4_1_3/C
+ sky130_fd_sc_hd__nor4_1_3/Y sky130_fd_sc_hd__nor4_1_3/A sky130_fd_sc_hd__nor4_1_3/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__nor4_1
Xsky130_fd_sc_hd__diode_2_130 sky130_fd_sc_hd__buf_2_250/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_141 sky130_fd_sc_hd__buf_2_168/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_152 sky130_fd_sc_hd__a22o_1_18/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_163 sky130_fd_sc_hd__nand4_1_74/D VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_174 sky130_fd_sc_hd__nand4_1_65/D VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_185 sky130_fd_sc_hd__buf_2_140/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_196 sky130_fd_sc_hd__clkbuf_4_208/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkinv_2_18 sky130_fd_sc_hd__clkinv_4_13/A sky130_fd_sc_hd__clkinv_4_11/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_18/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkbuf_4_205 sky130_fd_sc_hd__buf_12_404/A sky130_fd_sc_hd__buf_8_188/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_216 sky130_fd_sc_hd__nand2_1_567/B sky130_fd_sc_hd__dfxtp_1_1450/Q
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_2_29 sky130_fd_sc_hd__nand4_1_66/D sky130_fd_sc_hd__clkinv_2_29/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_29/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkbuf_4_227 sky130_fd_sc_hd__clkbuf_4_227/X sky130_fd_sc_hd__clkbuf_4_227/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_12_230 sky130_fd_sc_hd__buf_12_230/A sky130_fd_sc_hd__buf_12_230/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_241 sky130_fd_sc_hd__buf_12_241/A sky130_fd_sc_hd__buf_12_241/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_100 sky130_fd_sc_hd__a22oi_1_96/B1 sky130_fd_sc_hd__a22oi_1_96/A1
+ sky130_fd_sc_hd__clkbuf_1_150/X sky130_fd_sc_hd__a22oi_1_100/A2 sky130_fd_sc_hd__nand4_1_20/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_252 sky130_fd_sc_hd__buf_12_252/A sky130_fd_sc_hd__buf_12_252/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_111 sky130_fd_sc_hd__clkbuf_4_72/X sky130_fd_sc_hd__clkbuf_4_73/X
+ sky130_fd_sc_hd__a22oi_1_111/B2 sky130_fd_sc_hd__buf_2_91/X sky130_fd_sc_hd__buf_2_106/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_263 sky130_fd_sc_hd__buf_12_263/A sky130_fd_sc_hd__buf_12_263/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_122 sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__a22oi_2_12/A1
+ sky130_fd_sc_hd__buf_2_72/X sky130_fd_sc_hd__clkbuf_1_163/X sky130_fd_sc_hd__a22oi_1_122/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_274 sky130_fd_sc_hd__inv_2_90/Y sky130_fd_sc_hd__buf_12_356/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_133 sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__a22oi_2_12/A1
+ sky130_fd_sc_hd__buf_2_69/X sky130_fd_sc_hd__clkbuf_1_160/X sky130_fd_sc_hd__a22oi_1_133/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_285 sky130_fd_sc_hd__buf_6_40/A sky130_fd_sc_hd__buf_12_285/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_144 sky130_fd_sc_hd__a22oi_1_97/B1 sky130_fd_sc_hd__a22oi_1_97/A1
+ sky130_fd_sc_hd__buf_2_52/X sky130_fd_sc_hd__clkbuf_4_74/X sky130_fd_sc_hd__nand4_1_31/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_296 sky130_fd_sc_hd__buf_8_159/X sky130_fd_sc_hd__buf_12_366/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_155 sky130_fd_sc_hd__clkbuf_1_265/X sky130_fd_sc_hd__clkbuf_1_266/X
+ sky130_fd_sc_hd__clkbuf_1_279/X sky130_fd_sc_hd__a22oi_1_155/A2 sky130_fd_sc_hd__a22oi_1_155/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_166 sky130_fd_sc_hd__clkbuf_1_264/X sky130_fd_sc_hd__nor2_2_3/Y
+ sky130_fd_sc_hd__a22oi_1_166/B2 sky130_fd_sc_hd__clkbuf_4_133/X sky130_fd_sc_hd__nand4_1_36/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_177 sky130_fd_sc_hd__clkbuf_4_111/X sky130_fd_sc_hd__clkbuf_4_112/X
+ sky130_fd_sc_hd__a22oi_1_177/B2 sky130_fd_sc_hd__clkbuf_1_290/X sky130_fd_sc_hd__a22oi_1_177/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_188 sky130_fd_sc_hd__clkbuf_1_351/X sky130_fd_sc_hd__clkbuf_1_353/X
+ sky130_fd_sc_hd__clkbuf_4_115/X sky130_fd_sc_hd__a22oi_1_188/A2 sky130_fd_sc_hd__nand4_1_42/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_430 sky130_fd_sc_hd__o21ai_1_39/A2 sky130_fd_sc_hd__fa_2_956/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_430/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22oi_1_199 sky130_fd_sc_hd__clkbuf_1_265/X sky130_fd_sc_hd__clkbuf_1_266/X
+ sky130_fd_sc_hd__clkbuf_1_269/X sky130_fd_sc_hd__a22oi_1_199/A2 sky130_fd_sc_hd__a22oi_1_199/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_441 sky130_fd_sc_hd__fa_2_962/B sky130_fd_sc_hd__dfxtp_1_486/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_441/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_2_11 sky130_fd_sc_hd__or2_1_1/B sky130_fd_sc_hd__ha_2_89/A
+ sky130_fd_sc_hd__buf_2_162/A sky130_fd_sc_hd__a22o_2_11/B2 sky130_fd_sc_hd__a22o_4_0/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_2
Xsky130_fd_sc_hd__clkinv_1_452 sky130_fd_sc_hd__fa_2_949/B sky130_fd_sc_hd__nor2b_1_87/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_452/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_463 sky130_fd_sc_hd__o21ai_1_112/A1 sky130_fd_sc_hd__fa_2_992/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_463/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_474 sky130_fd_sc_hd__o22ai_1_79/B2 sky130_fd_sc_hd__ha_2_180/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_474/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_485 sky130_fd_sc_hd__o21ai_1_72/A2 sky130_fd_sc_hd__o2bb2ai_1_31/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_485/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_496 sky130_fd_sc_hd__o21ai_1_79/B1 sky130_fd_sc_hd__nor2_1_57/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_496/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_360 sky130_fd_sc_hd__or2_0_10/B sky130_fd_sc_hd__nor3_1_39/C
+ sky130_fd_sc_hd__o21bai_1_3/A2 sky130_fd_sc_hd__nor3_1_39/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_371 sky130_fd_sc_hd__o21a_1_52/B1 sky130_fd_sc_hd__o21a_1_51/A1
+ sky130_fd_sc_hd__a21oi_1_371/Y sky130_fd_sc_hd__o21a_1_55/A2 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_382 sky130_fd_sc_hd__xor2_1_230/X sky130_fd_sc_hd__o21ai_1_395/Y
+ sky130_fd_sc_hd__a21oi_1_382/Y sky130_fd_sc_hd__nand2_1_470/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_393 sky130_fd_sc_hd__nor2_2_17/Y sky130_fd_sc_hd__o21ai_1_408/Y
+ sky130_fd_sc_hd__nor2_1_257/B sky130_fd_sc_hd__fa_2_1240/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nor2_4_19 sky130_fd_sc_hd__nor3_1_41/A sky130_fd_sc_hd__nor2_4_19/A
+ sky130_fd_sc_hd__nor2_4_19/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__xor2_1_204 sky130_fd_sc_hd__fa_2_1173/A sky130_fd_sc_hd__fa_2_1175/B
+ sky130_fd_sc_hd__xor2_1_204/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_215 sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__fa_2_1203/B
+ sky130_fd_sc_hd__xor2_1_215/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_226 sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__fa_2_1192/B
+ sky130_fd_sc_hd__xor2_1_226/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_237 sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1238/B
+ sky130_fd_sc_hd__xor2_1_237/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_248 sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1227/B
+ sky130_fd_sc_hd__xor2_1_248/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_259 sky130_fd_sc_hd__xor2_1_267/B sky130_fd_sc_hd__fa_2_1255/B
+ sky130_fd_sc_hd__xor2_1_259/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_208 VSS VDD sky130_fd_sc_hd__buf_12_126/A sky130_fd_sc_hd__buf_8_75/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_219 VSS VDD sky130_fd_sc_hd__buf_2_121/A sky130_fd_sc_hd__ha_2_47/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_2_20 VDD VSS sky130_fd_sc_hd__inv_2_6/A sky130_fd_sc_hd__ha_2_23/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_31 VDD VSS sky130_fd_sc_hd__buf_8_53/A sky130_fd_sc_hd__buf_8_1/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_42 VDD VSS sky130_fd_sc_hd__buf_2_42/X sky130_fd_sc_hd__buf_2_42/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_53 VDD VSS sky130_fd_sc_hd__buf_2_53/X sky130_fd_sc_hd__buf_2_53/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_64 VDD VSS sky130_fd_sc_hd__buf_2_64/X sky130_fd_sc_hd__buf_2_64/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_75 VDD VSS sky130_fd_sc_hd__buf_2_75/X sky130_fd_sc_hd__buf_2_75/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_86 VDD VSS sky130_fd_sc_hd__buf_2_86/X sky130_fd_sc_hd__buf_2_86/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_97 VDD VSS sky130_fd_sc_hd__buf_2_97/X sky130_fd_sc_hd__buf_2_97/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__diode_2_4 sky130_fd_sc_hd__clkbuf_1_247/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__and2_0_206 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_206/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_206/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_217 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_217/X sky130_fd_sc_hd__and2_0_235/B
+ sky130_fd_sc_hd__and2_0_217/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_228 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_228/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_228/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_239 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_239/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__fa_2_874/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_260 sky130_fd_sc_hd__o21ai_1_3/B1 sky130_fd_sc_hd__nor3_1_26/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_260/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_271 sky130_fd_sc_hd__maj3_1_0/C sky130_fd_sc_hd__ha_2_148/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_271/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_2_5 sky130_fd_sc_hd__nor2_4_4/Y sky130_fd_sc_hd__xor2_1_7/B
+ sky130_fd_sc_hd__nor2_1_7/B sky130_fd_sc_hd__a22o_2_5/B2 sky130_fd_sc_hd__a22o_2_6/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_2
Xsky130_fd_sc_hd__o31ai_1_4 sky130_fd_sc_hd__o31ai_1_4/Y sky130_fd_sc_hd__nor2_1_39/Y
+ sky130_fd_sc_hd__a31oi_1_2/Y sky130_fd_sc_hd__o31ai_1_4/A3 sky130_fd_sc_hd__o31ai_1_4/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__o31ai_1
Xsky130_fd_sc_hd__clkinv_1_282 sky130_fd_sc_hd__fa_2_76/B sky130_fd_sc_hd__ha_2_91/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_282/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_293 sky130_fd_sc_hd__fa_2_144/B sky130_fd_sc_hd__ha_2_97/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_293/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_1 sky130_fd_sc_hd__nand3_1_17/C sky130_fd_sc_hd__or2_0_0/B
+ sky130_fd_sc_hd__a21oi_1_1/Y sky130_fd_sc_hd__o21ai_1_2/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkbuf_4_14 sky130_fd_sc_hd__clkbuf_4_14/X sky130_fd_sc_hd__clkbuf_4_14/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_207 VSS VDD sky130_fd_sc_hd__nor2_1_127/A sky130_fd_sc_hd__nand2_1_316/Y
+ sky130_fd_sc_hd__nand2_1_315/Y sky130_fd_sc_hd__o21ai_1_207/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_25 sky130_fd_sc_hd__clkbuf_4_25/X sky130_fd_sc_hd__clkbuf_4_25/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_218 VSS VDD sky130_fd_sc_hd__a21oi_1_200/Y sky130_fd_sc_hd__nor2_1_126/A
+ sky130_fd_sc_hd__nand2_1_321/Y sky130_fd_sc_hd__o21ai_1_218/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_36 sky130_fd_sc_hd__a22oi_2_6/B2 sky130_fd_sc_hd__clkbuf_4_36/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_229 VSS VDD sky130_fd_sc_hd__o21ai_1_229/A2 sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__a21oi_1_203/Y sky130_fd_sc_hd__xor2_1_129/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_47 sky130_fd_sc_hd__nand4_1_10/D sky130_fd_sc_hd__a22oi_1_61/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_58 sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__clkinv_1_55/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_69 sky130_fd_sc_hd__clkbuf_4_69/X sky130_fd_sc_hd__buf_2_41/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__a21oi_1_190 sky130_fd_sc_hd__a21o_2_5/A2 sky130_fd_sc_hd__o21ai_1_210/Y
+ sky130_fd_sc_hd__a21oi_1_190/Y sky130_fd_sc_hd__fa_2_1077/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_120 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__buf_4_74/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_131 sky130_fd_sc_hd__buf_8_131/A sky130_fd_sc_hd__buf_8_131/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_142 sky130_fd_sc_hd__buf_8_142/A sky130_fd_sc_hd__buf_4_77/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_153 sky130_fd_sc_hd__buf_8_153/A sky130_fd_sc_hd__buf_4_88/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nor2_4_4 sky130_fd_sc_hd__nor2_4_4/Y sky130_fd_sc_hd__nor2_4_4/A
+ sky130_fd_sc_hd__inv_2_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__buf_8_164 sky130_fd_sc_hd__buf_8_164/A sky130_fd_sc_hd__buf_8_164/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_175 sky130_fd_sc_hd__buf_8_175/A sky130_fd_sc_hd__buf_8_175/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_186 sky130_fd_sc_hd__buf_8_186/A sky130_fd_sc_hd__buf_8_186/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_197 sky130_fd_sc_hd__inv_2_127/Y sky130_fd_sc_hd__buf_8_197/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_407 VDD VSS sky130_fd_sc_hd__fa_2_1043/A sky130_fd_sc_hd__dfxtp_1_425/CLK
+ sky130_fd_sc_hd__and2_0_114/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_418 VDD VSS sky130_fd_sc_hd__fa_2_1038/B sky130_fd_sc_hd__dfxtp_1_419/CLK
+ sky130_fd_sc_hd__and2_0_137/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_429 VDD VSS sky130_fd_sc_hd__dfxtp_1_429/Q sky130_fd_sc_hd__dfxtp_1_433/CLK
+ sky130_fd_sc_hd__nand2_1_106/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a21o_2_10 sky130_fd_sc_hd__a21o_2_10/X sky130_fd_sc_hd__nor2_1_170/Y
+ sky130_fd_sc_hd__nor2_1_170/A sky130_fd_sc_hd__nor2_1_170/B VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__a21o_2_21 sky130_fd_sc_hd__a21o_2_21/X sky130_fd_sc_hd__nor2_1_254/Y
+ sky130_fd_sc_hd__nor2_1_254/A sky130_fd_sc_hd__nor2_1_254/B VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__clkinv_8_17 sky130_fd_sc_hd__clkinv_8_17/Y sky130_fd_sc_hd__clkinv_8_17/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_17/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_28 sky130_fd_sc_hd__clkinv_8_29/A sky130_fd_sc_hd__clkinv_8_28/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_28/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_39 sky130_fd_sc_hd__clkinv_8_40/A sky130_fd_sc_hd__clkinv_8_62/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_39/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__buf_12_15 sky130_fd_sc_hd__buf_12_15/A sky130_fd_sc_hd__buf_12_15/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_70 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__xor2_1_70/X
+ sky130_fd_sc_hd__xor2_1_70/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_26 sky130_fd_sc_hd__buf_8_20/X sky130_fd_sc_hd__buf_12_92/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_81 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__fa_2_995/B
+ sky130_fd_sc_hd__xor2_1_81/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_37 sky130_fd_sc_hd__buf_8_16/X sky130_fd_sc_hd__buf_12_37/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_92 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__xor2_1_92/X
+ sky130_fd_sc_hd__xor2_1_92/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_48 sky130_fd_sc_hd__buf_8_0/X sky130_fd_sc_hd__buf_12_48/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_59 sky130_fd_sc_hd__buf_8_56/X sky130_fd_sc_hd__buf_12_88/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__dfxtp_1_1303 VDD VSS sky130_fd_sc_hd__fa_2_848/B sky130_fd_sc_hd__dfxtp_1_1322/CLK
+ sky130_fd_sc_hd__a21oi_1_435/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1314 VDD VSS sky130_fd_sc_hd__fa_2_837/B sky130_fd_sc_hd__dfxtp_1_1332/CLK
+ sky130_fd_sc_hd__a21oi_1_429/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1325 VDD VSS sky130_fd_sc_hd__fa_2_909/A sky130_fd_sc_hd__dfxtp_1_1326/CLK
+ sky130_fd_sc_hd__o21a_1_59/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1336 VDD VSS sky130_fd_sc_hd__fa_2_1295/A sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__mux2_2_260/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1347 VDD VSS sky130_fd_sc_hd__fa_2_1306/A sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__mux2_2_230/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1358 VDD VSS sky130_fd_sc_hd__fa_2_1280/A sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__mux2_2_252/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_930 VDD VSS sky130_fd_sc_hd__fa_2_1122/B sky130_fd_sc_hd__clkinv_8_55/Y
+ sky130_fd_sc_hd__and2_0_319/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1369 VDD VSS sky130_fd_sc_hd__fa_2_1291/A sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__mux2_2_225/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_941 VDD VSS sky130_fd_sc_hd__fa_2_1133/A sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__mux2_2_91/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_952 VDD VSS sky130_fd_sc_hd__fa_2_1161/A sky130_fd_sc_hd__clkinv_8_63/Y
+ sky130_fd_sc_hd__mux2_2_120/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_963 VDD VSS sky130_fd_sc_hd__fa_2_1172/A sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__nand2_1_363/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_974 VDD VSS sky130_fd_sc_hd__mux2_2_108/A0 sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__o22ai_1_221/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_985 VDD VSS sky130_fd_sc_hd__mux2_2_81/A1 sky130_fd_sc_hd__clkinv_8_46/Y
+ sky130_fd_sc_hd__o22ai_1_210/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_996 VDD VSS sky130_fd_sc_hd__mux2_2_109/A0 sky130_fd_sc_hd__clkinv_8_65/Y
+ sky130_fd_sc_hd__dfxtp_1_996/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_550 VSS VDD sky130_fd_sc_hd__nor2_8_0/A sky130_fd_sc_hd__mux2_2_135/S
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_561 VSS VDD sky130_fd_sc_hd__nand2_1_95/B sky130_fd_sc_hd__nand4_1_57/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_572 VSS VDD sky130_fd_sc_hd__dfxtp_1_60/D sky130_fd_sc_hd__nand4_1_46/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_140 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_140/A sky130_fd_sc_hd__fa_2_733/A
+ sky130_fd_sc_hd__fa_2_730/B sky130_fd_sc_hd__ha_2_140/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_583 VSS VDD sky130_fd_sc_hd__nand3_1_9/A sky130_fd_sc_hd__a22oi_1_19/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_151 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_151/A sky130_fd_sc_hd__ha_2_150/B
+ sky130_fd_sc_hd__ha_2_151/SUM sky130_fd_sc_hd__ha_2_151/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_594 VSS VDD sky130_fd_sc_hd__buf_2_285/A sky130_fd_sc_hd__dfxtp_1_1458/Q
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_802 sky130_fd_sc_hd__fa_2_803/B sky130_fd_sc_hd__fa_2_796/A
+ sky130_fd_sc_hd__ha_2_145/B sky130_fd_sc_hd__fa_2_812/B sky130_fd_sc_hd__fa_2_833/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_162 VSS VDD VSS VDD sky130_fd_sc_hd__or4_1_0/D sky130_fd_sc_hd__ha_2_161/B
+ sky130_fd_sc_hd__ha_2_162/SUM sky130_fd_sc_hd__ha_2_162/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_813 sky130_fd_sc_hd__fa_2_815/CIN sky130_fd_sc_hd__fa_2_804/A
+ sky130_fd_sc_hd__ha_2_140/B sky130_fd_sc_hd__fa_2_813/B sky130_fd_sc_hd__fa_2_813/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_173 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_173/A sky130_fd_sc_hd__ha_2_172/A
+ sky130_fd_sc_hd__ha_2_173/SUM sky130_fd_sc_hd__ha_2_173/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_824 sky130_fd_sc_hd__fa_2_826/CIN sky130_fd_sc_hd__fa_2_818/A
+ sky130_fd_sc_hd__fa_2_835/B sky130_fd_sc_hd__ha_2_144/A sky130_fd_sc_hd__fa_2_820/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_184 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_184/A sky130_fd_sc_hd__ha_2_183/A
+ sky130_fd_sc_hd__ha_2_184/SUM sky130_fd_sc_hd__ha_2_184/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_835 sky130_fd_sc_hd__fa_2_703/A sky130_fd_sc_hd__fa_2_704/B
+ sky130_fd_sc_hd__ha_2_145/A sky130_fd_sc_hd__fa_2_835/B sky130_fd_sc_hd__fa_2_832/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_195 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_195/A sky130_fd_sc_hd__ha_2_194/A
+ sky130_fd_sc_hd__ha_2_195/SUM sky130_fd_sc_hd__ha_2_195/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_846 sky130_fd_sc_hd__fa_2_845/CIN sky130_fd_sc_hd__fa_2_846/SUM
+ sky130_fd_sc_hd__fa_2_846/A sky130_fd_sc_hd__fa_2_846/B sky130_fd_sc_hd__fa_2_846/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_857 sky130_fd_sc_hd__fa_2_856/CIN sky130_fd_sc_hd__fa_2_857/SUM
+ sky130_fd_sc_hd__fa_2_857/A sky130_fd_sc_hd__fa_2_857/B sky130_fd_sc_hd__fa_2_857/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_868 sky130_fd_sc_hd__fa_2_867/CIN sky130_fd_sc_hd__fa_2_868/SUM
+ sky130_fd_sc_hd__fa_2_868/A sky130_fd_sc_hd__fa_2_868/B sky130_fd_sc_hd__fa_2_868/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__maj3_1_0 sky130_fd_sc_hd__maj3_1_0/C sky130_fd_sc_hd__maj3_1_0/X
+ sky130_fd_sc_hd__maj3_1_1/X sky130_fd_sc_hd__maj3_1_0/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__fa_2_879 sky130_fd_sc_hd__fa_2_878/CIN sky130_fd_sc_hd__nand2_1_39/B
+ sky130_fd_sc_hd__ha_2_150/A sky130_fd_sc_hd__fa_2_879/B sky130_fd_sc_hd__fa_2_879/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__mux2_2_102 VSS VDD sky130_fd_sc_hd__mux2_2_102/A1 sky130_fd_sc_hd__mux2_2_102/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_102/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_113 VSS VDD sky130_fd_sc_hd__mux2_2_113/A1 sky130_fd_sc_hd__mux2_2_113/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_113/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_124 VSS VDD sky130_fd_sc_hd__mux2_2_124/A1 sky130_fd_sc_hd__xor2_1_207/X
+ sky130_fd_sc_hd__mux2_2_135/S sky130_fd_sc_hd__mux2_2_124/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_135 VSS VDD sky130_fd_sc_hd__mux2_2_135/A1 sky130_fd_sc_hd__mux2_2_135/A0
+ sky130_fd_sc_hd__mux2_2_135/S sky130_fd_sc_hd__mux2_2_135/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_146 VSS VDD sky130_fd_sc_hd__mux2_2_146/A1 sky130_fd_sc_hd__mux2_2_146/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_146/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_157 VSS VDD sky130_fd_sc_hd__mux2_2_157/A1 sky130_fd_sc_hd__mux2_2_157/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_157/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_168 VSS VDD sky130_fd_sc_hd__mux2_2_168/A1 sky130_fd_sc_hd__mux2_2_168/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_168/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_179 VSS VDD sky130_fd_sc_hd__mux2_2_179/A1 sky130_fd_sc_hd__mux2_2_179/A0
+ sky130_fd_sc_hd__nor2_8_1/A sky130_fd_sc_hd__mux2_2_179/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__and2_0_20 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_20/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_18/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_300 sky130_fd_sc_hd__o22ai_1_322/A2 sky130_fd_sc_hd__nor2_1_218/A
+ sky130_fd_sc_hd__o22ai_1_300/Y sky130_fd_sc_hd__o22ai_1_309/B1 sky130_fd_sc_hd__o32ai_1_5/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_31 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_31/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_37/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_311 sky130_fd_sc_hd__o22ai_1_322/A2 sky130_fd_sc_hd__nor2_1_192/B
+ sky130_fd_sc_hd__o22ai_1_311/Y sky130_fd_sc_hd__o22ai_1_322/B1 sky130_fd_sc_hd__o32ai_1_5/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_42 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_57/A sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__ha_2_50/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_106 sky130_fd_sc_hd__maj3_1_107/X sky130_fd_sc_hd__maj3_1_106/X
+ sky130_fd_sc_hd__maj3_1_106/B sky130_fd_sc_hd__maj3_1_106/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_322 sky130_fd_sc_hd__o22ai_1_322/A2 sky130_fd_sc_hd__o22ai_1_322/B1
+ sky130_fd_sc_hd__o22ai_1_322/Y sky130_fd_sc_hd__nor2_1_195/B sky130_fd_sc_hd__o32ai_1_5/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_53 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_53/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_53/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_117 sky130_fd_sc_hd__maj3_1_118/X sky130_fd_sc_hd__maj3_1_117/X
+ sky130_fd_sc_hd__maj3_1_117/B sky130_fd_sc_hd__maj3_1_117/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_333 sky130_fd_sc_hd__nand2_1_462/Y sky130_fd_sc_hd__nand2_1_461/Y
+ sky130_fd_sc_hd__o22ai_1_333/Y sky130_fd_sc_hd__o22ai_1_346/A1 sky130_fd_sc_hd__a21o_2_22/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_64 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_81/A sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__ha_2_79/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_128 sky130_fd_sc_hd__maj3_1_129/X sky130_fd_sc_hd__maj3_1_128/X
+ sky130_fd_sc_hd__maj3_1_128/B sky130_fd_sc_hd__maj3_1_128/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_344 sky130_fd_sc_hd__nand2_1_464/Y sky130_fd_sc_hd__nand2_1_463/Y
+ sky130_fd_sc_hd__o22ai_1_344/Y sky130_fd_sc_hd__o22ai_1_344/A1 sky130_fd_sc_hd__a21o_2_21/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_75 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_75/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__and2_0_75/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_408 sky130_fd_sc_hd__o32ai_1_5/B1 sky130_fd_sc_hd__o32ai_1_5/A3
+ sky130_fd_sc_hd__o21bai_1_3/A2 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_139 sky130_fd_sc_hd__maj3_1_140/X sky130_fd_sc_hd__maj3_1_139/X
+ sky130_fd_sc_hd__maj3_1_139/B sky130_fd_sc_hd__maj3_1_139/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_355 sky130_fd_sc_hd__nor2_1_257/A sky130_fd_sc_hd__nor2_1_268/A
+ sky130_fd_sc_hd__o22ai_1_355/Y sky130_fd_sc_hd__a21boi_1_5/Y sky130_fd_sc_hd__a222oi_1_26/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_86 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_86/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_86/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nor2_2_1 sky130_fd_sc_hd__inv_2_2/Y sky130_fd_sc_hd__or2_1_1/B sky130_fd_sc_hd__nor2_4_4/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__nand2_1_419 sky130_fd_sc_hd__o31ai_1_8/A2 sky130_fd_sc_hd__nand2_1_419/B
+ sky130_fd_sc_hd__nor2_1_208/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_366 sky130_fd_sc_hd__o22ai_1_379/A2 sky130_fd_sc_hd__o22ai_1_366/B1
+ sky130_fd_sc_hd__o22ai_1_366/Y sky130_fd_sc_hd__nor2_1_230/B sky130_fd_sc_hd__o32ai_1_8/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_97 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_97/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_97/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_377 sky130_fd_sc_hd__o22ai_1_379/A2 sky130_fd_sc_hd__nor2_1_266/A
+ sky130_fd_sc_hd__o22ai_1_377/Y sky130_fd_sc_hd__nor2_1_236/B sky130_fd_sc_hd__o32ai_1_8/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_388 sky130_fd_sc_hd__nand2_1_514/Y sky130_fd_sc_hd__nand2_1_513/Y
+ sky130_fd_sc_hd__o22ai_1_388/Y sky130_fd_sc_hd__o22ai_1_401/A1 sky130_fd_sc_hd__a21o_2_27/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_399 sky130_fd_sc_hd__nand2_1_516/Y sky130_fd_sc_hd__nand2_1_515/Y
+ sky130_fd_sc_hd__o22ai_1_399/Y sky130_fd_sc_hd__o22ai_1_399/A1 sky130_fd_sc_hd__a21o_2_26/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_8_30 sky130_fd_sc_hd__inv_2_10/Y sky130_fd_sc_hd__buf_8_30/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_41 sky130_fd_sc_hd__buf_8_41/A sky130_fd_sc_hd__buf_8_41/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_52 sky130_fd_sc_hd__buf_8_53/A sky130_fd_sc_hd__buf_8_52/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_63 sky130_fd_sc_hd__buf_8_63/A sky130_fd_sc_hd__buf_8_63/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_74 sky130_fd_sc_hd__buf_8_74/A sky130_fd_sc_hd__buf_8_74/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_85 sky130_fd_sc_hd__buf_8_86/A sky130_fd_sc_hd__buf_8_85/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_204 VDD VSS sky130_fd_sc_hd__ha_2_77/A sky130_fd_sc_hd__dfxtp_1_207/CLK
+ sky130_fd_sc_hd__and2_0_77/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_8_96 sky130_fd_sc_hd__buf_8_96/A sky130_fd_sc_hd__buf_8_96/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_215 VDD VSS sky130_fd_sc_hd__ha_2_88/A sky130_fd_sc_hd__dfxtp_1_224/CLK
+ sky130_fd_sc_hd__nor2b_1_43/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_226 VDD VSS sky130_fd_sc_hd__nor3_2_9/B sky130_fd_sc_hd__clkinv_4_20/Y
+ sky130_fd_sc_hd__nor2_1_7/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_237 VDD VSS sky130_fd_sc_hd__fa_2_872/A sky130_fd_sc_hd__dfxtp_1_462/CLK
+ sky130_fd_sc_hd__and2_0_170/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_248 VDD VSS sky130_fd_sc_hd__buf_8_63/A sky130_fd_sc_hd__dfxtp_1_258/CLK
+ sky130_fd_sc_hd__and2_0_200/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_259 VDD VSS sky130_fd_sc_hd__dfxtp_1_259/Q sky130_fd_sc_hd__dfxtp_1_262/CLK
+ sky130_fd_sc_hd__and2_0_222/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_109 sky130_fd_sc_hd__maj3_1_7/B sky130_fd_sc_hd__maj3_1_8/A
+ sky130_fd_sc_hd__fa_2_109/A sky130_fd_sc_hd__fa_2_109/B sky130_fd_sc_hd__fa_2_110/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_104 VDD VSS sky130_fd_sc_hd__buf_2_104/X sky130_fd_sc_hd__buf_2_104/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__fa_2_1303 sky130_fd_sc_hd__fa_2_1304/CIN sky130_fd_sc_hd__mux2_2_237/A1
+ sky130_fd_sc_hd__fa_2_1303/A sky130_fd_sc_hd__fa_2_1303/B sky130_fd_sc_hd__fa_2_1303/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_115 VDD VSS sky130_fd_sc_hd__buf_8_67/A sky130_fd_sc_hd__ha_2_48/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__fa_2_1314 sky130_fd_sc_hd__fa_2_1315/CIN sky130_fd_sc_hd__mux2_2_264/A1
+ sky130_fd_sc_hd__fa_2_1314/A sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1314/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_126 VDD VSS sky130_fd_sc_hd__buf_2_126/X sky130_fd_sc_hd__buf_2_126/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o22ai_1_19 sky130_fd_sc_hd__fa_2_238/B sky130_fd_sc_hd__fa_2_265/B
+ sky130_fd_sc_hd__fa_2_268/A sky130_fd_sc_hd__ha_2_91/A sky130_fd_sc_hd__fa_2_2/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__fa_2_1325 sky130_fd_sc_hd__xor2_1_318/B sky130_fd_sc_hd__nand2_1_521/A
+ sky130_fd_sc_hd__fa_2_1325/A sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1325/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_137 VDD VSS sky130_fd_sc_hd__buf_4_97/A sky130_fd_sc_hd__inv_2_85/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_148 VDD VSS sky130_fd_sc_hd__buf_2_148/X sky130_fd_sc_hd__buf_2_148/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_159 VDD VSS sky130_fd_sc_hd__buf_2_159/X sky130_fd_sc_hd__buf_8_192/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1100 VDD VSS sky130_fd_sc_hd__fa_2_1219/A sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__mux2_2_151/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1111 VDD VSS sky130_fd_sc_hd__nor2_4_16/A sky130_fd_sc_hd__clkinv_4_23/Y
+ sky130_fd_sc_hd__nor2b_1_115/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1122 VDD VSS sky130_fd_sc_hd__mux2_2_137/A0 sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__o22ai_1_271/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1133 VDD VSS sky130_fd_sc_hd__mux2_2_167/A0 sky130_fd_sc_hd__clkinv_8_64/Y
+ sky130_fd_sc_hd__dfxtp_1_992/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1144 VDD VSS sky130_fd_sc_hd__mux2_2_161/A0 sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__a21oi_1_319/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1155 VDD VSS sky130_fd_sc_hd__mux2_2_132/A1 sky130_fd_sc_hd__clkinv_8_70/Y
+ sky130_fd_sc_hd__o22ai_1_282/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1166 VDD VSS sky130_fd_sc_hd__fa_2_858/B sky130_fd_sc_hd__dfxtp_1_1180/CLK
+ sky130_fd_sc_hd__o21a_1_53/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1177 VDD VSS sky130_fd_sc_hd__ha_2_169/A sky130_fd_sc_hd__dfxtp_1_1179/CLK
+ sky130_fd_sc_hd__a21oi_1_368/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1188 VDD VSS sky130_fd_sc_hd__fa_2_941/A sky130_fd_sc_hd__clkinv_4_24/Y
+ sky130_fd_sc_hd__o21a_1_44/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_760 VDD VSS sky130_fd_sc_hd__ha_2_133/B sky130_fd_sc_hd__dfxtp_1_764/CLK
+ sky130_fd_sc_hd__dfxtp_1_760/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1199 VDD VSS sky130_fd_sc_hd__fa_2_1248/A sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__mux2_2_200/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_771 VDD VSS sky130_fd_sc_hd__fa_2_1070/A sky130_fd_sc_hd__clkinv_8_54/Y
+ sky130_fd_sc_hd__and2_0_304/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__ha_2_4 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_4/A sky130_fd_sc_hd__ha_2_3/B
+ sky130_fd_sc_hd__ha_2_4/SUM sky130_fd_sc_hd__ha_2_4/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__dfxtp_1_782 VDD VSS sky130_fd_sc_hd__fa_2_1081/A sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__mux2_2_60/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_793 VDD VSS sky130_fd_sc_hd__xor2_1_88/A sky130_fd_sc_hd__clkinv_4_25/Y
+ sky130_fd_sc_hd__mux2_2_38/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_380 VSS VDD sky130_fd_sc_hd__a22oi_2_25/B1 sky130_fd_sc_hd__nor3_2_8/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_391 VSS VDD sky130_fd_sc_hd__a22oi_2_20/B2 sky130_fd_sc_hd__clkbuf_1_391/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_610 sky130_fd_sc_hd__maj3_1_120/B sky130_fd_sc_hd__maj3_1_121/A
+ sky130_fd_sc_hd__fa_2_610/A sky130_fd_sc_hd__fa_2_610/B sky130_fd_sc_hd__fa_2_611/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_15 VSS VDD sky130_fd_sc_hd__buf_6_8/A sky130_fd_sc_hd__dfxtp_1_459/Q
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_621 sky130_fd_sc_hd__fa_2_623/CIN sky130_fd_sc_hd__fa_2_618/A
+ sky130_fd_sc_hd__ha_2_130/B sky130_fd_sc_hd__fa_2_621/B sky130_fd_sc_hd__fa_2_621/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_26 VSS VDD sky130_fd_sc_hd__clkbuf_1_26/X sky130_fd_sc_hd__clkbuf_1_26/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_632 sky130_fd_sc_hd__fa_2_633/B sky130_fd_sc_hd__fa_2_630/B
+ sky130_fd_sc_hd__fa_2_632/A sky130_fd_sc_hd__fa_2_632/B sky130_fd_sc_hd__fa_2_635/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_37 VSS VDD sky130_fd_sc_hd__clkbuf_1_37/X sky130_fd_sc_hd__clkbuf_1_37/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_643 sky130_fd_sc_hd__fa_2_642/B sky130_fd_sc_hd__fa_2_643/SUM
+ sky130_fd_sc_hd__fa_2_695/A sky130_fd_sc_hd__ha_2_131/B sky130_fd_sc_hd__ha_2_131/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_48 VSS VDD sky130_fd_sc_hd__clkbuf_1_48/X sky130_fd_sc_hd__clkbuf_1_48/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_654 sky130_fd_sc_hd__fa_2_653/B sky130_fd_sc_hd__fa_2_654/SUM
+ sky130_fd_sc_hd__ha_2_129/B sky130_fd_sc_hd__ha_2_131/B sky130_fd_sc_hd__ha_2_131/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_59 VSS VDD sky130_fd_sc_hd__clkbuf_1_59/X sky130_fd_sc_hd__clkbuf_1_59/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_665 sky130_fd_sc_hd__fa_2_580/A sky130_fd_sc_hd__fa_2_581/B
+ sky130_fd_sc_hd__fa_2_665/A sky130_fd_sc_hd__fa_2_665/B sky130_fd_sc_hd__fa_2_671/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_676 sky130_fd_sc_hd__fa_2_675/B sky130_fd_sc_hd__fa_2_676/SUM
+ sky130_fd_sc_hd__fa_2_676/A sky130_fd_sc_hd__fa_2_676/B sky130_fd_sc_hd__fa_2_676/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_687 sky130_fd_sc_hd__fa_2_575/A sky130_fd_sc_hd__fa_2_576/B
+ sky130_fd_sc_hd__fa_2_687/A sky130_fd_sc_hd__fa_2_687/B sky130_fd_sc_hd__fa_2_692/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_698 sky130_fd_sc_hd__fa_2_571/A sky130_fd_sc_hd__fa_2_572/B
+ sky130_fd_sc_hd__fa_2_698/A sky130_fd_sc_hd__fa_2_698/B sky130_fd_sc_hd__fa_2_698/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22oi_2_18 sky130_fd_sc_hd__buf_2_165/X sky130_fd_sc_hd__a22oi_2_18/A2
+ sky130_fd_sc_hd__nor2_4_7/Y sky130_fd_sc_hd__a22oi_2_18/B2 sky130_fd_sc_hd__nand4_1_51/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__a22oi_2_29 sky130_fd_sc_hd__buf_2_165/X sky130_fd_sc_hd__a22oi_2_29/A2
+ sky130_fd_sc_hd__nor2_4_7/Y sky130_fd_sc_hd__a22oi_2_29/B2 sky130_fd_sc_hd__nand4_1_61/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__buf_12_4 sky130_fd_sc_hd__inv_2_20/Y sky130_fd_sc_hd__buf_12_4/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__o22ai_1_130 sky130_fd_sc_hd__nor2_1_88/A sky130_fd_sc_hd__o22ai_1_130/B1
+ sky130_fd_sc_hd__o22ai_1_130/Y sky130_fd_sc_hd__o22ai_1_132/B1 sky130_fd_sc_hd__o22ai_1_132/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_141 sky130_fd_sc_hd__nand2_1_284/Y sky130_fd_sc_hd__nand2_2_5/Y
+ sky130_fd_sc_hd__o22ai_1_141/Y sky130_fd_sc_hd__xnor2_1_74/Y sky130_fd_sc_hd__o22ai_1_155/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_205 sky130_fd_sc_hd__nor2_1_26/B sky130_fd_sc_hd__nor3_1_31/B
+ sky130_fd_sc_hd__or4_1_2/D VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_804 sky130_fd_sc_hd__o22ai_1_235/A1 sky130_fd_sc_hd__or3_1_2/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_804/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_152 sky130_fd_sc_hd__nand2_1_338/A sky130_fd_sc_hd__nand2_1_284/Y
+ sky130_fd_sc_hd__o22ai_1_152/Y sky130_fd_sc_hd__xnor2_1_68/Y sky130_fd_sc_hd__o22ai_1_152/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_216 sky130_fd_sc_hd__nor2_1_34/B sky130_fd_sc_hd__nand2_1_216/B
+ sky130_fd_sc_hd__nor2_1_35/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_815 sky130_fd_sc_hd__nand2_1_370/B sky130_fd_sc_hd__fa_2_426/SUM
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_163 sky130_fd_sc_hd__o21ai_1_199/Y sky130_fd_sc_hd__nand2_2_5/Y
+ sky130_fd_sc_hd__o22ai_1_163/Y sky130_fd_sc_hd__nand2_1_338/A sky130_fd_sc_hd__a22o_1_72/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_227 sky130_fd_sc_hd__o22ai_1_88/B1 sky130_fd_sc_hd__nor2_2_6/B
+ sky130_fd_sc_hd__nor2_2_6/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_174 sky130_fd_sc_hd__o22ai_1_204/B1 sky130_fd_sc_hd__nor2_1_118/B
+ sky130_fd_sc_hd__o22ai_1_174/Y sky130_fd_sc_hd__o22ai_1_194/B1 sky130_fd_sc_hd__o22ai_1_206/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_826 sky130_fd_sc_hd__nor2_1_176/A sky130_fd_sc_hd__fa_2_1137/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_826/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_238 sky130_fd_sc_hd__o21ai_1_82/B1 sky130_fd_sc_hd__nor2_1_61/B
+ sky130_fd_sc_hd__nor2_1_61/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_185 sky130_fd_sc_hd__o22ai_1_204/B1 sky130_fd_sc_hd__o22ai_1_190/A1
+ sky130_fd_sc_hd__nor2_1_132/A sky130_fd_sc_hd__nor2_1_116/B sky130_fd_sc_hd__o22ai_1_206/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand4_1_11 sky130_fd_sc_hd__nand4_1_11/C sky130_fd_sc_hd__nand4_1_11/B
+ sky130_fd_sc_hd__nand4_1_11/Y sky130_fd_sc_hd__nand4_1_11/D sky130_fd_sc_hd__nand4_1_11/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__clkinv_1_837 sky130_fd_sc_hd__o21ai_1_311/A2 sky130_fd_sc_hd__o21ai_1_322/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_837/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_249 sky130_fd_sc_hd__nand2_1_249/Y sky130_fd_sc_hd__nor2_1_50/B
+ sky130_fd_sc_hd__nor2_1_50/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_848 sky130_fd_sc_hd__nor2_1_183/B sky130_fd_sc_hd__o21ai_1_328/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_848/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_196 sky130_fd_sc_hd__a21oi_1_220/Y sky130_fd_sc_hd__o22ai_1_196/B1
+ sky130_fd_sc_hd__o22ai_1_196/Y sky130_fd_sc_hd__nor2_1_126/A sky130_fd_sc_hd__nor2_2_13/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand4_1_22 sky130_fd_sc_hd__nand4_1_22/C sky130_fd_sc_hd__nand4_1_22/B
+ sky130_fd_sc_hd__nand4_1_22/Y sky130_fd_sc_hd__nand4_1_22/D sky130_fd_sc_hd__buf_2_106/X
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_33 sky130_fd_sc_hd__nand4_1_33/C sky130_fd_sc_hd__nand4_1_33/B
+ sky130_fd_sc_hd__nand4_1_33/Y sky130_fd_sc_hd__nand4_1_33/D sky130_fd_sc_hd__nand4_1_33/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__clkinv_1_859 sky130_fd_sc_hd__nor2_1_158/B sky130_fd_sc_hd__o21bai_1_2/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_859/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand4_1_44 sky130_fd_sc_hd__nand4_1_44/C sky130_fd_sc_hd__nand4_1_44/B
+ sky130_fd_sc_hd__buf_2_286/A sky130_fd_sc_hd__nand4_1_44/D sky130_fd_sc_hd__nand4_1_44/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_55 sky130_fd_sc_hd__nand4_1_55/C sky130_fd_sc_hd__nand4_1_55/B
+ sky130_fd_sc_hd__buf_2_267/A sky130_fd_sc_hd__nand4_1_55/D sky130_fd_sc_hd__nand4_1_55/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_66 sky130_fd_sc_hd__nand4_1_66/C sky130_fd_sc_hd__nand4_1_66/B
+ sky130_fd_sc_hd__nand4_1_66/Y sky130_fd_sc_hd__nand4_1_66/D sky130_fd_sc_hd__nand4_1_66/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_77 sky130_fd_sc_hd__nand4_1_77/C sky130_fd_sc_hd__nand4_1_77/B
+ sky130_fd_sc_hd__nand2_1_2/B sky130_fd_sc_hd__nand4_1_77/D sky130_fd_sc_hd__nand4_1_77/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__conb_1_15 sky130_fd_sc_hd__conb_1_15/LO sky130_fd_sc_hd__conb_1_15/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_26 sky130_fd_sc_hd__conb_1_26/LO sky130_fd_sc_hd__conb_1_26/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__o21ai_1_390 VSS VDD sky130_fd_sc_hd__nand2_1_476/B sky130_fd_sc_hd__nor2_1_256/Y
+ sky130_fd_sc_hd__nor2_1_255/B sky130_fd_sc_hd__o21ai_1_390/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__mux2_2_70 VSS VDD sky130_fd_sc_hd__mux2_2_70/A1 sky130_fd_sc_hd__mux2_2_70/A0
+ sky130_fd_sc_hd__mux2_2_75/S sky130_fd_sc_hd__mux2_2_70/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_81 VSS VDD sky130_fd_sc_hd__mux2_2_81/A1 sky130_fd_sc_hd__mux2_2_81/A0
+ sky130_fd_sc_hd__nor2_4_15/A sky130_fd_sc_hd__mux2_2_81/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1100 sky130_fd_sc_hd__fa_2_1101/CIN sky130_fd_sc_hd__and2_0_306/A
+ sky130_fd_sc_hd__fa_2_1100/A sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1100/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__mux2_2_92 VSS VDD sky130_fd_sc_hd__xor2_1_183/X sky130_fd_sc_hd__mux2_2_92/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_92/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1111 sky130_fd_sc_hd__fa_2_1112/CIN sky130_fd_sc_hd__fa_2_1111/SUM
+ sky130_fd_sc_hd__fa_2_1111/A sky130_fd_sc_hd__fa_2_1111/B sky130_fd_sc_hd__fa_2_1111/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1122 sky130_fd_sc_hd__fa_2_1123/CIN sky130_fd_sc_hd__and2_0_319/A
+ sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__fa_2_1122/B sky130_fd_sc_hd__xor2_1_161/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1133 sky130_fd_sc_hd__fa_2_1134/CIN sky130_fd_sc_hd__mux2_2_91/A1
+ sky130_fd_sc_hd__fa_2_1133/A sky130_fd_sc_hd__fa_2_1133/B sky130_fd_sc_hd__fa_2_1133/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1144 sky130_fd_sc_hd__fa_2_1145/CIN sky130_fd_sc_hd__mux2_2_110/A1
+ sky130_fd_sc_hd__fa_2_1144/A sky130_fd_sc_hd__fa_2_1144/B sky130_fd_sc_hd__fa_2_1144/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1155 sky130_fd_sc_hd__fa_2_1156/CIN sky130_fd_sc_hd__mux2_2_82/A0
+ sky130_fd_sc_hd__fa_2_1155/A sky130_fd_sc_hd__fa_2_1155/B sky130_fd_sc_hd__fa_2_1155/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1166 sky130_fd_sc_hd__fa_2_1167/CIN sky130_fd_sc_hd__mux2_2_109/A1
+ sky130_fd_sc_hd__fa_2_1166/A sky130_fd_sc_hd__fa_2_1172/B sky130_fd_sc_hd__fa_2_1166/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1177 sky130_fd_sc_hd__fa_2_1178/CIN sky130_fd_sc_hd__mux2_2_159/A1
+ sky130_fd_sc_hd__fa_2_1177/A sky130_fd_sc_hd__fa_2_1177/B sky130_fd_sc_hd__fa_2_1177/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1188 sky130_fd_sc_hd__fa_2_1189/CIN sky130_fd_sc_hd__mux2_2_131/A0
+ sky130_fd_sc_hd__fa_2_1188/A sky130_fd_sc_hd__fa_2_1188/B sky130_fd_sc_hd__fa_2_1188/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1199 sky130_fd_sc_hd__fa_2_1200/CIN sky130_fd_sc_hd__mux2_2_146/A1
+ sky130_fd_sc_hd__fa_2_1199/A sky130_fd_sc_hd__fa_2_1199/B sky130_fd_sc_hd__fa_2_1199/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_590 VDD VSS sky130_fd_sc_hd__nor4_1_6/C sky130_fd_sc_hd__dfxtp_1_591/CLK
+ sky130_fd_sc_hd__a21o_2_0/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_440 sky130_fd_sc_hd__fa_2_436/B sky130_fd_sc_hd__fa_2_440/SUM
+ sky130_fd_sc_hd__ha_2_124/A sky130_fd_sc_hd__fa_2_535/A sky130_fd_sc_hd__fa_2_566/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o2bb2ai_1_6 sky130_fd_sc_hd__o2bb2ai_1_6/Y sky130_fd_sc_hd__nor2_1_18/Y
+ sky130_fd_sc_hd__ha_2_155/SUM sky130_fd_sc_hd__o21ai_1_31/A1 sky130_fd_sc_hd__maj3_1_2/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_451 sky130_fd_sc_hd__fa_2_445/A sky130_fd_sc_hd__fa_2_448/B
+ sky130_fd_sc_hd__fa_2_451/A sky130_fd_sc_hd__fa_2_451/B sky130_fd_sc_hd__fa_2_451/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_462 sky130_fd_sc_hd__fa_2_459/B sky130_fd_sc_hd__fa_2_463/CIN
+ sky130_fd_sc_hd__fa_2_462/A sky130_fd_sc_hd__fa_2_462/B sky130_fd_sc_hd__fa_2_462/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_473 sky130_fd_sc_hd__maj3_1_101/B sky130_fd_sc_hd__maj3_1_102/A
+ sky130_fd_sc_hd__fa_2_473/A sky130_fd_sc_hd__fa_2_473/B sky130_fd_sc_hd__fa_2_474/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_484 sky130_fd_sc_hd__fa_2_486/CIN sky130_fd_sc_hd__fa_2_482/A
+ sky130_fd_sc_hd__ha_2_124/B sky130_fd_sc_hd__fa_2_537/A sky130_fd_sc_hd__fa_2_484/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_2_0 VDD VSS sky130_fd_sc_hd__and2_2_0/A sky130_fd_sc_hd__and2_2_0/X
+ sky130_fd_sc_hd__inv_8_1/Y VDD VSS sky130_fd_sc_hd__and2_2
Xsky130_fd_sc_hd__fa_2_495 sky130_fd_sc_hd__fa_2_498/B sky130_fd_sc_hd__fa_2_495/SUM
+ sky130_fd_sc_hd__fa_2_495/A sky130_fd_sc_hd__fa_2_495/B sky130_fd_sc_hd__fa_2_495/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor2_1_205 sky130_fd_sc_hd__nor2_1_205/B sky130_fd_sc_hd__nor2_1_205/Y
+ sky130_fd_sc_hd__nor2_1_205/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_216 sky130_fd_sc_hd__nor2_1_216/B sky130_fd_sc_hd__nor2_1_216/Y
+ sky130_fd_sc_hd__nor2_1_225/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_227 sky130_fd_sc_hd__nor2_1_261/A sky130_fd_sc_hd__o21a_1_43/A1
+ sky130_fd_sc_hd__o21a_1_44/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_238 sky130_fd_sc_hd__nor2_1_238/B sky130_fd_sc_hd__o21a_1_52/A1
+ sky130_fd_sc_hd__o21a_1_53/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_249 sky130_fd_sc_hd__nor2_1_249/B sky130_fd_sc_hd__nor2_1_249/Y
+ sky130_fd_sc_hd__nor2_1_267/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_401 sky130_fd_sc_hd__buf_8_187/X sky130_fd_sc_hd__buf_12_451/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_412 sky130_fd_sc_hd__buf_8_190/X sky130_fd_sc_hd__buf_12_412/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_423 sky130_fd_sc_hd__buf_8_196/X sky130_fd_sc_hd__buf_12_478/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_434 sky130_fd_sc_hd__buf_8_198/X sky130_fd_sc_hd__buf_12_455/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_445 sky130_fd_sc_hd__buf_4_109/X sky130_fd_sc_hd__buf_12_445/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_304 sky130_fd_sc_hd__clkbuf_1_376/X sky130_fd_sc_hd__nor2_2_5/Y
+ sky130_fd_sc_hd__buf_2_206/X sky130_fd_sc_hd__clkbuf_1_462/X sky130_fd_sc_hd__nand4_1_75/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_456 sky130_fd_sc_hd__buf_6_65/X sky130_fd_sc_hd__buf_12_456/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_315 sky130_fd_sc_hd__nor2_2_4/Y sky130_fd_sc_hd__nor3_1_24/Y
+ sky130_fd_sc_hd__a22oi_1_315/B2 sky130_fd_sc_hd__clkbuf_4_178/X sky130_fd_sc_hd__nand4_1_78/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_467 sky130_fd_sc_hd__buf_6_64/X sky130_fd_sc_hd__buf_12_515/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_326 sky130_fd_sc_hd__fa_2_988/A sky130_fd_sc_hd__fa_2_990/A
+ sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__a22oi_1_326/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_478 sky130_fd_sc_hd__buf_12_478/A sky130_fd_sc_hd__buf_12_478/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_337 sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__nor2_2_8/Y
+ sky130_fd_sc_hd__fa_2_1013/A sky130_fd_sc_hd__fa_2_1015/A sky130_fd_sc_hd__a22oi_1_337/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_489 sky130_fd_sc_hd__buf_12_489/A sky130_fd_sc_hd__buf_12_489/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_348 sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__nor2_4_13/Y
+ sky130_fd_sc_hd__fa_2_1075/A sky130_fd_sc_hd__fa_2_1076/A sky130_fd_sc_hd__a22oi_1_348/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_359 sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__nor2_4_13/Y
+ sky130_fd_sc_hd__fa_2_1083/A sky130_fd_sc_hd__fa_2_1084/A sky130_fd_sc_hd__a22oi_1_359/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_601 sky130_fd_sc_hd__ha_2_176/B sky130_fd_sc_hd__fa_2_1039/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_601/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_612 sky130_fd_sc_hd__o21ai_1_92/A1 sky130_fd_sc_hd__nor2_2_8/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_612/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_623 sky130_fd_sc_hd__o21ai_1_230/A1 sky130_fd_sc_hd__fa_2_1068/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_623/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_634 sky130_fd_sc_hd__o22ai_1_152/B2 sky130_fd_sc_hd__ha_2_197/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_634/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_645 sky130_fd_sc_hd__o21ai_1_189/A2 sky130_fd_sc_hd__ha_2_186/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_645/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_656 sky130_fd_sc_hd__nor2_1_94/B sky130_fd_sc_hd__nand2_1_303/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_656/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_667 sky130_fd_sc_hd__clkinv_1_667/Y sky130_fd_sc_hd__nor2_1_95/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_667/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_678 sky130_fd_sc_hd__nor2_1_107/B sky130_fd_sc_hd__fa_2_1110/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_678/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_689 sky130_fd_sc_hd__o21ai_1_191/A2 sky130_fd_sc_hd__nor2_1_141/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_689/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand3_1_7 sky130_fd_sc_hd__nand3_1_7/Y sky130_fd_sc_hd__nand3_1_7/A
+ sky130_fd_sc_hd__nand3_1_7/C sky130_fd_sc_hd__nand3_1_7/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__a222oi_1_10 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1157/A sky130_fd_sc_hd__nor2_2_15/Y
+ sky130_fd_sc_hd__nor3_1_38/A sky130_fd_sc_hd__xor2_1_163/A sky130_fd_sc_hd__nor2_2_15/A
+ sky130_fd_sc_hd__a222oi_1_10/Y sky130_fd_sc_hd__fa_2_1156/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_21 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1195/A sky130_fd_sc_hd__nor2_2_16/Y
+ sky130_fd_sc_hd__nor3_1_39/A sky130_fd_sc_hd__fa_2_1197/A sky130_fd_sc_hd__nor3_1_39/B
+ sky130_fd_sc_hd__a222oi_1_21/Y sky130_fd_sc_hd__fa_2_1194/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_32 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1245/A sky130_fd_sc_hd__nor2_2_17/Y
+ sky130_fd_sc_hd__nor3_1_40/A sky130_fd_sc_hd__fa_2_1247/A sky130_fd_sc_hd__nor3_1_40/B
+ sky130_fd_sc_hd__nor2_1_264/B sky130_fd_sc_hd__fa_2_1244/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_43 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1295/A sky130_fd_sc_hd__nor2_2_18/Y
+ sky130_fd_sc_hd__nor3_1_41/A sky130_fd_sc_hd__fa_2_1297/A sky130_fd_sc_hd__nor3_1_41/B
+ sky130_fd_sc_hd__a222oi_1_43/Y sky130_fd_sc_hd__fa_2_1294/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_12 VSS VDD sky130_fd_sc_hd__xnor2_1_12/B sky130_fd_sc_hd__xnor2_1_12/Y
+ sky130_fd_sc_hd__ha_2_150/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_23 VSS VDD sky130_fd_sc_hd__xnor2_1_23/B sky130_fd_sc_hd__xnor2_1_23/Y
+ sky130_fd_sc_hd__xnor2_1_23/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_34 VSS VDD sky130_fd_sc_hd__xnor2_1_34/B sky130_fd_sc_hd__xnor2_1_34/Y
+ sky130_fd_sc_hd__nor2_1_42/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_45 VSS VDD sky130_fd_sc_hd__xnor2_1_45/B sky130_fd_sc_hd__xnor2_1_45/Y
+ sky130_fd_sc_hd__nor2_1_45/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_56 VSS VDD sky130_fd_sc_hd__xnor2_1_56/B sky130_fd_sc_hd__xnor2_1_56/Y
+ sky130_fd_sc_hd__xnor2_1_56/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_67 VSS VDD sky130_fd_sc_hd__xnor2_1_67/B sky130_fd_sc_hd__xnor2_1_67/Y
+ sky130_fd_sc_hd__nor2_1_93/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_78 VSS VDD sky130_fd_sc_hd__xnor2_1_78/B sky130_fd_sc_hd__xnor2_1_78/Y
+ sky130_fd_sc_hd__nor2_1_96/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_89 VSS VDD sky130_fd_sc_hd__xnor2_1_89/B sky130_fd_sc_hd__xnor2_1_89/Y
+ sky130_fd_sc_hd__xnor2_1_89/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__a211oi_1_3 sky130_fd_sc_hd__fa_2_962/A sky130_fd_sc_hd__o21ai_1_37/Y
+ sky130_fd_sc_hd__nor3_1_36/C sky130_fd_sc_hd__a31oi_1_1/A3 sky130_fd_sc_hd__nor3_1_36/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o32ai_1_6 sky130_fd_sc_hd__o32ai_1_6/A2 sky130_fd_sc_hd__o32ai_1_6/Y
+ sky130_fd_sc_hd__fa_2_1226/A sky130_fd_sc_hd__o32ai_1_6/A3 sky130_fd_sc_hd__o32ai_1_6/B2
+ sky130_fd_sc_hd__fa_2_1225/A VDD VSS VSS VDD sky130_fd_sc_hd__o32ai_1
Xsky130_fd_sc_hd__clkbuf_16_4 sky130_fd_sc_hd__buf_8_62/A sky130_fd_sc_hd__buf_12_66/X
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__fa_2_270 sky130_fd_sc_hd__fa_2_269/A sky130_fd_sc_hd__fa_2_264/B
+ sky130_fd_sc_hd__fa_2_15/B sky130_fd_sc_hd__ha_2_97/A sky130_fd_sc_hd__fa_2_258/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_281 sky130_fd_sc_hd__fa_2_283/CIN sky130_fd_sc_hd__fa_2_275/A
+ sky130_fd_sc_hd__fa_2_281/A sky130_fd_sc_hd__fa_2_281/B sky130_fd_sc_hd__fa_2_238/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_292 sky130_fd_sc_hd__fa_2_290/CIN sky130_fd_sc_hd__fa_2_292/SUM
+ sky130_fd_sc_hd__fa_2_292/A sky130_fd_sc_hd__fa_2_292/B sky130_fd_sc_hd__fa_2_292/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor4_1_4 sky130_fd_sc_hd__xor2_1_9/A sky130_fd_sc_hd__nor4_1_4/C
+ sky130_fd_sc_hd__nor4_1_4/Y sky130_fd_sc_hd__nor4_1_4/A sky130_fd_sc_hd__nor4_1_4/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__nor4_1
Xsky130_fd_sc_hd__a22oi_1_3 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__a22oi_1_9/A1
+ sky130_fd_sc_hd__dfxtp_1_60/D sky130_fd_sc_hd__a22o_1_8/A1 sky130_fd_sc_hd__nand3_1_1/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__diode_2_120 sky130_fd_sc_hd__clkbuf_4_189/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_131 sky130_fd_sc_hd__clkbuf_1_526/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_142 sky130_fd_sc_hd__buf_2_168/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_153 sky130_fd_sc_hd__buf_2_174/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_164 sky130_fd_sc_hd__nand4_1_75/D VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_175 sky130_fd_sc_hd__nand4_1_77/D VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_186 sky130_fd_sc_hd__buf_2_140/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_197 sky130_fd_sc_hd__buf_4_120/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkinv_2_19 sky130_fd_sc_hd__clkinv_2_19/Y sky130_fd_sc_hd__clkinv_4_78/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_2_19/w_94_21# sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkbuf_4_206 sky130_fd_sc_hd__buf_2_168/A sky130_fd_sc_hd__buf_2_249/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_217 sky130_fd_sc_hd__nor4_1_0/A sram_select[1] VSS VDD
+ VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_228 sky130_fd_sc_hd__a22oi_1_11/A2 sig_amplitude[2] VSS
+ VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_12_220 sky130_fd_sc_hd__buf_12_220/A sky130_fd_sc_hd__buf_12_252/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_231 sky130_fd_sc_hd__buf_12_231/A sky130_fd_sc_hd__buf_12_231/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_242 sky130_fd_sc_hd__buf_12_242/A sky130_fd_sc_hd__buf_12_242/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_101 sky130_fd_sc_hd__a22oi_1_97/B1 sky130_fd_sc_hd__a22oi_1_97/A1
+ sky130_fd_sc_hd__buf_2_61/X sky130_fd_sc_hd__clkbuf_4_85/X sky130_fd_sc_hd__nand4_1_20/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_253 sky130_fd_sc_hd__buf_12_253/A sky130_fd_sc_hd__buf_12_253/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_112 sky130_fd_sc_hd__a22oi_1_96/B1 sky130_fd_sc_hd__a22oi_1_96/A1
+ sky130_fd_sc_hd__clkbuf_1_147/X sky130_fd_sc_hd__a22oi_1_112/A2 sky130_fd_sc_hd__nand4_1_23/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_264 sky130_fd_sc_hd__buf_12_264/A sky130_fd_sc_hd__buf_12_264/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_123 sky130_fd_sc_hd__clkbuf_4_72/X sky130_fd_sc_hd__clkbuf_4_73/X
+ sky130_fd_sc_hd__a22oi_1_123/B2 sky130_fd_sc_hd__buf_2_88/X sky130_fd_sc_hd__clkbuf_4_90/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_275 sky130_fd_sc_hd__buf_12_275/A sky130_fd_sc_hd__buf_12_364/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_134 sky130_fd_sc_hd__clkbuf_4_72/X sky130_fd_sc_hd__clkbuf_4_73/X
+ sky130_fd_sc_hd__a22oi_1_134/B2 sky130_fd_sc_hd__buf_2_85/X sky130_fd_sc_hd__buf_2_103/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_286 sky130_fd_sc_hd__buf_12_286/A sky130_fd_sc_hd__buf_12_286/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_145 sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__a22oi_2_12/A1
+ sky130_fd_sc_hd__buf_2_66/X sky130_fd_sc_hd__clkbuf_1_157/X sky130_fd_sc_hd__a22oi_1_145/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_297 sky130_fd_sc_hd__buf_8_125/X sky130_fd_sc_hd__buf_12_353/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_156 sky130_fd_sc_hd__clkbuf_1_351/X sky130_fd_sc_hd__clkbuf_1_353/X
+ sky130_fd_sc_hd__clkbuf_4_119/X sky130_fd_sc_hd__a22oi_1_156/A2 sky130_fd_sc_hd__nand4_1_34/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_167 sky130_fd_sc_hd__clkbuf_1_265/X sky130_fd_sc_hd__clkbuf_1_266/X
+ sky130_fd_sc_hd__clkbuf_1_277/X sky130_fd_sc_hd__a22oi_1_167/A2 sky130_fd_sc_hd__a22oi_1_167/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_178 sky130_fd_sc_hd__clkbuf_1_264/X sky130_fd_sc_hd__nor2_2_3/Y
+ sky130_fd_sc_hd__a22oi_1_178/B2 sky130_fd_sc_hd__clkbuf_4_130/X sky130_fd_sc_hd__nand4_1_39/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_420 sky130_fd_sc_hd__o221ai_1_1/A2 sky130_fd_sc_hd__dfxtp_1_489/Q
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22oi_1_189 sky130_fd_sc_hd__clkbuf_4_111/X sky130_fd_sc_hd__clkbuf_4_112/X
+ sky130_fd_sc_hd__a22oi_1_189/B2 sky130_fd_sc_hd__clkbuf_1_287/X sky130_fd_sc_hd__a22oi_1_189/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_431 sky130_fd_sc_hd__or3_1_1/C sky130_fd_sc_hd__dfxtp_1_490/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_431/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_442 sky130_fd_sc_hd__fa_2_960/B sky130_fd_sc_hd__nand3_1_48/C
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_442/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_453 sky130_fd_sc_hd__fa_2_948/B sky130_fd_sc_hd__o21ai_1_36/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_453/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_464 sky130_fd_sc_hd__nor2_1_78/A sky130_fd_sc_hd__xor2_1_60/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_464/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_475 sky130_fd_sc_hd__o22ai_1_80/B2 sky130_fd_sc_hd__ha_2_179/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_475/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_486 sky130_fd_sc_hd__o21ai_1_74/B1 sky130_fd_sc_hd__nor2_1_62/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_486/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_497 sky130_fd_sc_hd__nor2_1_43/B sky130_fd_sc_hd__nand2_1_245/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_497/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_350 sky130_fd_sc_hd__fa_2_1208/A sky130_fd_sc_hd__nor2_1_220/Y
+ sky130_fd_sc_hd__a21oi_1_350/Y sky130_fd_sc_hd__nor3_1_39/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_361 sky130_fd_sc_hd__o21a_1_44/B1 sky130_fd_sc_hd__o21a_1_43/A1
+ sky130_fd_sc_hd__a21oi_1_361/Y sky130_fd_sc_hd__nor2_1_261/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_372 sky130_fd_sc_hd__o21a_1_53/B1 sky130_fd_sc_hd__o21a_1_52/A1
+ sky130_fd_sc_hd__a21oi_1_372/Y sky130_fd_sc_hd__nor2_1_238/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_383 sky130_fd_sc_hd__o21ai_1_406/Y sky130_fd_sc_hd__clkinv_1_986/Y
+ sky130_fd_sc_hd__a21oi_1_383/Y sky130_fd_sc_hd__nor2b_2_4/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_394 sky130_fd_sc_hd__fa_2_1238/A sky130_fd_sc_hd__o22ai_1_359/Y
+ sky130_fd_sc_hd__a21oi_1_394/Y sky130_fd_sc_hd__nor3_1_40/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__xor2_1_205 sky130_fd_sc_hd__fa_2_1173/A sky130_fd_sc_hd__fa_2_1174/B
+ sky130_fd_sc_hd__xor2_1_205/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_216 sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__fa_2_1202/B
+ sky130_fd_sc_hd__xor2_1_216/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_227 sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__xor2_1_227/X
+ sky130_fd_sc_hd__xor2_1_227/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_238 sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1237/B
+ sky130_fd_sc_hd__xor2_1_238/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_249 sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1226/B
+ sky130_fd_sc_hd__xor2_1_249/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__clkbuf_1_209 VSS VDD sky130_fd_sc_hd__buf_12_134/A sky130_fd_sc_hd__buf_8_67/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_2_10 VDD VSS sky130_fd_sc_hd__buf_2_10/X sky130_fd_sc_hd__buf_2_10/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_21 VDD VSS sky130_fd_sc_hd__buf_8_15/A sky130_fd_sc_hd__ha_2_26/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_32 VDD VSS sky130_fd_sc_hd__ha_2_12/A sky130_fd_sc_hd__buf_2_32/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_43 VDD VSS sky130_fd_sc_hd__buf_8_78/A sky130_fd_sc_hd__ha_2_32/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_54 VDD VSS sky130_fd_sc_hd__buf_2_54/X sky130_fd_sc_hd__buf_2_54/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_65 VDD VSS sky130_fd_sc_hd__buf_2_65/X sky130_fd_sc_hd__buf_2_65/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_76 VDD VSS sky130_fd_sc_hd__buf_2_76/X sky130_fd_sc_hd__buf_2_76/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_87 VDD VSS sky130_fd_sc_hd__buf_2_87/X sky130_fd_sc_hd__buf_2_87/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_98 VDD VSS sky130_fd_sc_hd__buf_8_77/A sky130_fd_sc_hd__buf_8_86/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__diode_2_5 sky130_fd_sc_hd__clkbuf_1_247/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__o211ai_1_70 sky130_fd_sc_hd__nor2_1_309/A sky130_fd_sc_hd__a21oi_1_474/Y
+ sky130_fd_sc_hd__xor2_1_289/A sky130_fd_sc_hd__nand2_1_544/Y sky130_fd_sc_hd__a21oi_1_466/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__and2_0_207 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_207/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_207/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_218 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_218/X sky130_fd_sc_hd__and2_0_235/B
+ sky130_fd_sc_hd__and2_0_218/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_229 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_229/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_229/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_250 sky130_fd_sc_hd__buf_12_396/A sky130_fd_sc_hd__clkinv_1_250/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_250/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_261 sky130_fd_sc_hd__nor2_1_13/B sky130_fd_sc_hd__ha_2_157/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_261/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_272 sky130_fd_sc_hd__a21oi_2_0/A2 sky130_fd_sc_hd__xor2_1_17/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_272/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_2_6 sky130_fd_sc_hd__nor2_4_4/Y sky130_fd_sc_hd__ha_2_70/A
+ sky130_fd_sc_hd__nor2_1_7/A sky130_fd_sc_hd__a22o_2_6/B2 sky130_fd_sc_hd__a22o_2_6/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22o_2
Xsky130_fd_sc_hd__o31ai_1_5 sky130_fd_sc_hd__o31ai_1_5/Y sky130_fd_sc_hd__xnor2_1_93/Y
+ sky130_fd_sc_hd__o31ai_1_6/A2 sky130_fd_sc_hd__o31ai_1_6/A3 sky130_fd_sc_hd__o31ai_1_5/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__o31ai_1
Xsky130_fd_sc_hd__clkinv_1_283 sky130_fd_sc_hd__fa_2_139/B sky130_fd_sc_hd__ha_2_95/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_283/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_294 sky130_fd_sc_hd__fa_2_238/B sky130_fd_sc_hd__fa_2_2/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_294/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_2 sky130_fd_sc_hd__or4_1_0/A sky130_fd_sc_hd__o21ai_1_5/Y
+ sky130_fd_sc_hd__a21oi_1_2/Y sky130_fd_sc_hd__o21ai_1_4/A2 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkbuf_4_15 sky130_fd_sc_hd__clkbuf_4_15/X sky130_fd_sc_hd__clkbuf_4_15/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_208 VSS VDD sky130_fd_sc_hd__nor2_1_139/A sky130_fd_sc_hd__nand2_1_339/A
+ sky130_fd_sc_hd__a21oi_1_188/Y sky130_fd_sc_hd__o21ai_1_208/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_26 sky130_fd_sc_hd__clkbuf_4_26/X sky130_fd_sc_hd__clkbuf_4_26/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_219 VSS VDD sky130_fd_sc_hd__nor2_1_132/Y sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__a21oi_1_194/Y sky130_fd_sc_hd__xor2_1_124/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_37 sky130_fd_sc_hd__a22oi_2_5/B2 sky130_fd_sc_hd__clkbuf_4_37/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_48 sky130_fd_sc_hd__nand4_1_9/D sky130_fd_sc_hd__a22oi_1_58/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_59 sky130_fd_sc_hd__buf_2_35/A sky130_fd_sc_hd__buf_2_119/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__a21oi_1_180 sky130_fd_sc_hd__o21a_1_10/B1 sky130_fd_sc_hd__o21a_1_9/A1
+ sky130_fd_sc_hd__dfxtp_1_766/D sky130_fd_sc_hd__nor2_1_113/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_191 sky130_fd_sc_hd__clkinv_1_698/Y sky130_fd_sc_hd__clkinv_1_694/Y
+ sky130_fd_sc_hd__a21oi_1_191/Y sky130_fd_sc_hd__nand2_1_331/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_110 sky130_fd_sc_hd__buf_8_110/A sky130_fd_sc_hd__buf_8_110/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_121 sky130_fd_sc_hd__inv_2_75/Y sky130_fd_sc_hd__buf_6_42/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_132 sky130_fd_sc_hd__buf_8_132/A sky130_fd_sc_hd__buf_8_132/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_143 sky130_fd_sc_hd__buf_8_143/A sky130_fd_sc_hd__buf_4_83/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_154 sky130_fd_sc_hd__buf_8_154/A sky130_fd_sc_hd__buf_4_92/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nor2_4_5 sky130_fd_sc_hd__nor2_4_5/Y sky130_fd_sc_hd__nor3_2_3/A
+ sky130_fd_sc_hd__nor2_4_5/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__buf_8_165 sky130_fd_sc_hd__buf_8_165/A sky130_fd_sc_hd__buf_8_165/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_176 sky130_fd_sc_hd__buf_8_176/A sky130_fd_sc_hd__buf_8_176/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_187 sky130_fd_sc_hd__buf_8_187/A sky130_fd_sc_hd__buf_8_187/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_198 sky130_fd_sc_hd__buf_8_198/A sky130_fd_sc_hd__buf_8_198/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_408 VDD VSS sky130_fd_sc_hd__nor2_1_62/A sky130_fd_sc_hd__dfxtp_1_425/CLK
+ sky130_fd_sc_hd__and2_0_108/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_419 VDD VSS sky130_fd_sc_hd__nor2_1_51/A sky130_fd_sc_hd__dfxtp_1_419/CLK
+ sky130_fd_sc_hd__and2_0_132/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a21o_2_11 sky130_fd_sc_hd__a21o_2_11/X sky130_fd_sc_hd__nor2_1_171/Y
+ sky130_fd_sc_hd__nor2_1_171/A sky130_fd_sc_hd__or3_1_2/X VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__a21o_2_22 sky130_fd_sc_hd__a21o_2_22/X sky130_fd_sc_hd__nor2_1_255/Y
+ sky130_fd_sc_hd__nor2_1_255/A sky130_fd_sc_hd__nor2_1_255/B VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__clkinv_8_18 sky130_fd_sc_hd__clkinv_2_7/A sky130_fd_sc_hd__clkinv_8_18/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_18/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__clkinv_8_29 sky130_fd_sc_hd__clkinv_8_30/A sky130_fd_sc_hd__clkinv_8_29/A
+ VSS VDD VSS VDD VSS sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__xor2_1_60 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__xor2_1_60/X
+ sky130_fd_sc_hd__xor2_1_60/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_16 sky130_fd_sc_hd__inv_2_38/Y sky130_fd_sc_hd__buf_12_16/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_71 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__xor2_1_71/X
+ sky130_fd_sc_hd__xor2_1_71/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_27 sky130_fd_sc_hd__buf_8_8/X sky130_fd_sc_hd__buf_12_27/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_82 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__fa_2_994/B
+ sky130_fd_sc_hd__xor2_1_82/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_38 sky130_fd_sc_hd__buf_8_30/X sky130_fd_sc_hd__buf_12_38/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_93 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__xor2_1_93/X
+ sky130_fd_sc_hd__xor2_1_93/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_49 sky130_fd_sc_hd__buf_8_32/X sky130_fd_sc_hd__buf_12_49/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__dfxtp_1_1304 VDD VSS sky130_fd_sc_hd__fa_2_847/B sky130_fd_sc_hd__dfxtp_1_1322/CLK
+ sky130_fd_sc_hd__o21a_1_67/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1315 VDD VSS sky130_fd_sc_hd__fa_2_836/B sky130_fd_sc_hd__dfxtp_1_1329/CLK
+ sky130_fd_sc_hd__o21a_1_62/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1326 VDD VSS sky130_fd_sc_hd__fa_2_910/A sky130_fd_sc_hd__dfxtp_1_1326/CLK
+ sky130_fd_sc_hd__a21oi_1_423/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1337 VDD VSS sky130_fd_sc_hd__fa_2_1296/A sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__mux2_2_257/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1348 VDD VSS sky130_fd_sc_hd__fa_2_1307/A sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__mux2_2_228/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_920 VDD VSS sky130_fd_sc_hd__fa_2_1149/A sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__mux2_2_95/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1359 VDD VSS sky130_fd_sc_hd__fa_2_1281/A sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__mux2_2_249/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_931 VDD VSS sky130_fd_sc_hd__fa_2_1123/A sky130_fd_sc_hd__clkinv_8_55/Y
+ sky130_fd_sc_hd__and2_0_321/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_942 VDD VSS sky130_fd_sc_hd__fa_2_1134/A sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__mux2_2_89/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_953 VDD VSS sky130_fd_sc_hd__fa_2_1162/A sky130_fd_sc_hd__clkinv_8_64/Y
+ sky130_fd_sc_hd__mux2_2_119/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_964 VDD VSS sky130_fd_sc_hd__nor2_4_14/B sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__mux2_2_92/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_975 VDD VSS sky130_fd_sc_hd__mux2_2_105/A0 sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__o22ai_1_220/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_986 VDD VSS sky130_fd_sc_hd__mux2_2_79/A1 sky130_fd_sc_hd__clkinv_8_46/Y
+ sky130_fd_sc_hd__o31ai_1_6/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_997 VDD VSS sky130_fd_sc_hd__mux2_2_106/A0 sky130_fd_sc_hd__clkinv_8_65/Y
+ sky130_fd_sc_hd__dfxtp_1_997/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_540 VSS VDD sky130_fd_sc_hd__clkbuf_1_540/X sky130_fd_sc_hd__clkbuf_1_540/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_551 VSS VDD sky130_fd_sc_hd__o31ai_1_7/A2 sky130_fd_sc_hd__xnor2_1_96/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_562 VSS VDD sky130_fd_sc_hd__nand2_1_101/B sky130_fd_sc_hd__nand4_1_54/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_130 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_130/A sky130_fd_sc_hd__fa_2_599/A
+ sky130_fd_sc_hd__fa_2_596/B sky130_fd_sc_hd__ha_2_130/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_573 VSS VDD sky130_fd_sc_hd__dfxtp_1_75/D sky130_fd_sc_hd__nand4_1_45/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_141 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_141/A sky130_fd_sc_hd__fa_2_736/A
+ sky130_fd_sc_hd__fa_2_733/B sky130_fd_sc_hd__ha_2_141/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_584 VSS VDD sky130_fd_sc_hd__nand3_1_8/B sky130_fd_sc_hd__a22oi_1_16/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_152 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_152/A sky130_fd_sc_hd__ha_2_151/B
+ sky130_fd_sc_hd__ha_2_152/SUM sky130_fd_sc_hd__ha_2_152/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_595 VSS VDD sky130_fd_sc_hd__buf_2_277/A sram_select[0]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_803 sky130_fd_sc_hd__fa_2_805/CIN sky130_fd_sc_hd__fa_2_795/A
+ sky130_fd_sc_hd__ha_2_142/A sky130_fd_sc_hd__fa_2_803/B sky130_fd_sc_hd__fa_2_803/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_163 VSS VDD VSS VDD sky130_fd_sc_hd__or4_1_1/C sky130_fd_sc_hd__ha_2_162/B
+ sky130_fd_sc_hd__ha_2_163/SUM sky130_fd_sc_hd__ha_2_163/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_814 sky130_fd_sc_hd__fa_2_711/A sky130_fd_sc_hd__fa_2_712/B
+ sky130_fd_sc_hd__fa_2_814/A sky130_fd_sc_hd__fa_2_814/B sky130_fd_sc_hd__fa_2_819/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_174 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_174/A sky130_fd_sc_hd__ha_2_173/A
+ sky130_fd_sc_hd__ha_2_174/SUM sky130_fd_sc_hd__ha_2_174/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_825 sky130_fd_sc_hd__fa_2_708/A sky130_fd_sc_hd__fa_2_709/B
+ sky130_fd_sc_hd__fa_2_825/A sky130_fd_sc_hd__fa_2_825/B sky130_fd_sc_hd__fa_2_829/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_185 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_185/A sky130_fd_sc_hd__ha_2_185/COUT
+ sky130_fd_sc_hd__ha_2_185/SUM sky130_fd_sc_hd__ha_2_185/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_836 sky130_fd_sc_hd__xnor2_1_7/B sky130_fd_sc_hd__fa_2_836/SUM
+ sky130_fd_sc_hd__fa_2_836/A sky130_fd_sc_hd__fa_2_836/B sky130_fd_sc_hd__fa_2_836/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_196 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_196/A sky130_fd_sc_hd__ha_2_195/A
+ sky130_fd_sc_hd__ha_2_196/SUM sky130_fd_sc_hd__ha_2_196/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_847 sky130_fd_sc_hd__fa_2_846/CIN sky130_fd_sc_hd__fa_2_847/SUM
+ sky130_fd_sc_hd__fa_2_847/A sky130_fd_sc_hd__fa_2_847/B sky130_fd_sc_hd__fa_2_847/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_858 sky130_fd_sc_hd__fa_2_857/CIN sky130_fd_sc_hd__fa_2_858/SUM
+ sky130_fd_sc_hd__fa_2_858/A sky130_fd_sc_hd__fa_2_858/B sky130_fd_sc_hd__fa_2_858/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_869 sky130_fd_sc_hd__fa_2_868/CIN sky130_fd_sc_hd__fa_2_869/SUM
+ sky130_fd_sc_hd__fa_2_869/A sky130_fd_sc_hd__fa_2_869/B sky130_fd_sc_hd__fa_2_869/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__maj3_1_1 sky130_fd_sc_hd__maj3_1_1/C sky130_fd_sc_hd__maj3_1_1/X
+ sky130_fd_sc_hd__maj3_1_1/B sky130_fd_sc_hd__maj3_1_1/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__mux2_2_103 VSS VDD sky130_fd_sc_hd__mux2_2_103/A1 sky130_fd_sc_hd__mux2_2_103/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_103/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_114 VSS VDD sky130_fd_sc_hd__mux2_2_114/A1 sky130_fd_sc_hd__mux2_2_114/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_114/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_125 VSS VDD sky130_fd_sc_hd__mux2_2_125/A1 sky130_fd_sc_hd__xor2_1_186/X
+ sky130_fd_sc_hd__mux2_2_135/S sky130_fd_sc_hd__mux2_2_125/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_136 VSS VDD sky130_fd_sc_hd__mux2_2_136/A1 sky130_fd_sc_hd__mux2_2_136/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_136/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_147 VSS VDD sky130_fd_sc_hd__mux2_2_147/A1 sky130_fd_sc_hd__mux2_2_147/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_147/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_158 VSS VDD sky130_fd_sc_hd__mux2_2_158/A1 sky130_fd_sc_hd__mux2_2_158/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_158/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_169 VSS VDD sky130_fd_sc_hd__mux2_2_169/A1 sky130_fd_sc_hd__mux2_2_169/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_169/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__and2_0_10 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_10/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_5/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_21 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_21/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__xor2_1_1/X sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_301 sky130_fd_sc_hd__nor2_1_225/A sky130_fd_sc_hd__nor2_1_214/A
+ sky130_fd_sc_hd__o22ai_1_301/Y sky130_fd_sc_hd__o22ai_1_301/A1 sky130_fd_sc_hd__nor2_1_217/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_32 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_32/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_38/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_312 sky130_fd_sc_hd__nor2_1_225/A sky130_fd_sc_hd__nor2_1_214/A
+ sky130_fd_sc_hd__o22ai_1_312/Y sky130_fd_sc_hd__a21oi_1_350/Y sky130_fd_sc_hd__nor2_1_225/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_43 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_56/A sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__ha_2_59/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_107 sky130_fd_sc_hd__maj3_1_107/C sky130_fd_sc_hd__maj3_1_107/X
+ sky130_fd_sc_hd__maj3_1_107/B sky130_fd_sc_hd__maj3_1_107/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_323 sky130_fd_sc_hd__a21oi_1_377/Y sky130_fd_sc_hd__nand2_1_445/B
+ sky130_fd_sc_hd__o22ai_1_323/Y sky130_fd_sc_hd__nor3_1_40/C sky130_fd_sc_hd__o32ai_1_8/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_54 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_54/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_54/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_118 sky130_fd_sc_hd__maj3_1_119/X sky130_fd_sc_hd__maj3_1_118/X
+ sky130_fd_sc_hd__maj3_1_118/B sky130_fd_sc_hd__maj3_1_118/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_334 sky130_fd_sc_hd__nand2_1_462/Y sky130_fd_sc_hd__nand2_1_461/Y
+ sky130_fd_sc_hd__o22ai_1_334/Y sky130_fd_sc_hd__nand2_1_476/B sky130_fd_sc_hd__o21ai_1_390/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_65 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_80/A sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__xor2_1_7/X sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_129 sky130_fd_sc_hd__maj3_1_130/X sky130_fd_sc_hd__maj3_1_129/X
+ sky130_fd_sc_hd__maj3_1_129/B sky130_fd_sc_hd__maj3_1_129/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_345 sky130_fd_sc_hd__nand2_1_464/Y sky130_fd_sc_hd__nand2_1_463/Y
+ sky130_fd_sc_hd__o22ai_1_345/Y sky130_fd_sc_hd__nand2_1_475/B sky130_fd_sc_hd__o21ai_1_389/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_76 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_76/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__and2_0_76/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_409 sky130_fd_sc_hd__nand2_1_409/Y sky130_fd_sc_hd__o31ai_1_7/A2
+ sky130_fd_sc_hd__xor2_1_185/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_356 sky130_fd_sc_hd__o22ai_1_375/A2 sky130_fd_sc_hd__nor2_1_229/B
+ sky130_fd_sc_hd__o22ai_1_356/Y sky130_fd_sc_hd__nor2_1_230/B sky130_fd_sc_hd__o32ai_1_8/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_2_2 sky130_fd_sc_hd__nor2_4_5/B sky130_fd_sc_hd__nor2_2_2/Y
+ sky130_fd_sc_hd__nor3_2_2/C VDD VSS VSS VDD sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__and2_0_87 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_87/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_87/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_367 sky130_fd_sc_hd__o22ai_1_375/A2 sky130_fd_sc_hd__o21a_1_55/A2
+ sky130_fd_sc_hd__o22ai_1_367/Y sky130_fd_sc_hd__nor2_1_238/B sky130_fd_sc_hd__o32ai_1_8/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_98 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_98/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_98/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_378 sky130_fd_sc_hd__o32ai_1_8/A3 sky130_fd_sc_hd__nor2_1_239/B
+ sky130_fd_sc_hd__o22ai_1_378/Y sky130_fd_sc_hd__o22ai_1_378/A1 sky130_fd_sc_hd__o21a_1_55/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_389 sky130_fd_sc_hd__nand2_1_514/Y sky130_fd_sc_hd__nand2_1_513/Y
+ sky130_fd_sc_hd__o22ai_1_389/Y sky130_fd_sc_hd__nand2_1_527/B sky130_fd_sc_hd__o21ai_1_443/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_8_20 sky130_fd_sc_hd__buf_8_20/A sky130_fd_sc_hd__buf_8_20/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_31 sky130_fd_sc_hd__buf_8_31/A sky130_fd_sc_hd__buf_8_31/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_42 sky130_fd_sc_hd__buf_8_42/A sky130_fd_sc_hd__buf_8_42/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_53 sky130_fd_sc_hd__buf_8_53/A sky130_fd_sc_hd__inv_2_43/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_64 sky130_fd_sc_hd__inv_2_60/Y sky130_fd_sc_hd__buf_8_64/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_75 sky130_fd_sc_hd__buf_8_75/A sky130_fd_sc_hd__buf_8_75/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_86 sky130_fd_sc_hd__buf_8_86/A sky130_fd_sc_hd__buf_8_86/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_205 VDD VSS sky130_fd_sc_hd__ha_2_76/A sky130_fd_sc_hd__dfxtp_1_207/CLK
+ sky130_fd_sc_hd__and2_0_76/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_8_97 sky130_fd_sc_hd__buf_8_97/A sky130_fd_sc_hd__buf_8_97/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_216 VDD VSS sky130_fd_sc_hd__ha_2_87/A sky130_fd_sc_hd__dfxtp_1_224/CLK
+ sky130_fd_sc_hd__nor2b_1_44/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_227 VDD VSS sky130_fd_sc_hd__nor3_2_8/A sky130_fd_sc_hd__clkinv_4_20/Y
+ sky130_fd_sc_hd__nor2_1_7/B VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_238 VDD VSS sky130_fd_sc_hd__fa_2_871/A sky130_fd_sc_hd__dfxtp_1_462/CLK
+ sky130_fd_sc_hd__and2_0_167/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_249 VDD VSS sky130_fd_sc_hd__buf_2_119/A sky130_fd_sc_hd__dfxtp_1_262/CLK
+ sky130_fd_sc_hd__and2_0_201/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_2_105 VDD VSS sky130_fd_sc_hd__buf_2_105/X sky130_fd_sc_hd__buf_2_105/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__fa_2_1304 sky130_fd_sc_hd__fa_2_1305/CIN sky130_fd_sc_hd__mux2_2_234/A1
+ sky130_fd_sc_hd__fa_2_1304/A sky130_fd_sc_hd__fa_2_1304/B sky130_fd_sc_hd__fa_2_1304/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_116 VDD VSS sky130_fd_sc_hd__buf_2_116/X sky130_fd_sc_hd__buf_2_116/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__fa_2_1315 sky130_fd_sc_hd__fa_2_1316/CIN sky130_fd_sc_hd__mux2_2_263/A1
+ sky130_fd_sc_hd__fa_2_1315/A sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1315/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_127 VDD VSS sky130_fd_sc_hd__inv_2_76/A sky130_fd_sc_hd__a22o_2_0/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_138 VDD VSS sky130_fd_sc_hd__buf_2_138/X sky130_fd_sc_hd__buf_6_49/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_149 VDD VSS sky130_fd_sc_hd__buf_4_99/A sky130_fd_sc_hd__buf_2_149/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1101 VDD VSS sky130_fd_sc_hd__fa_2_1220/A sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__mux2_2_148/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1112 VDD VSS sky130_fd_sc_hd__mux2_2_165/A0 sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__nor2_1_202/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1123 VDD VSS sky130_fd_sc_hd__mux2_2_135/A1 sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__o22ai_1_270/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1134 VDD VSS sky130_fd_sc_hd__mux2_2_166/A0 sky130_fd_sc_hd__clkinv_8_64/Y
+ sky130_fd_sc_hd__dfxtp_1_993/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1145 VDD VSS sky130_fd_sc_hd__mux2_2_158/A0 sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__o22ai_1_292/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1156 VDD VSS sky130_fd_sc_hd__mux2_2_130/A1 sky130_fd_sc_hd__clkinv_8_70/Y
+ sky130_fd_sc_hd__o22ai_1_281/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1167 VDD VSS sky130_fd_sc_hd__fa_2_857/B sky130_fd_sc_hd__dfxtp_1_1180/CLK
+ sky130_fd_sc_hd__a21oi_1_372/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1178 VDD VSS sky130_fd_sc_hd__fa_2_931/A sky130_fd_sc_hd__dfxtp_1_1179/CLK
+ sky130_fd_sc_hd__a21oi_1_367/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_750 VDD VSS sky130_fd_sc_hd__and2_0_174/A sky130_fd_sc_hd__dfxtp_1_768/CLK
+ sky130_fd_sc_hd__fa_2_1105/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1189 VDD VSS sky130_fd_sc_hd__fa_2_942/A sky130_fd_sc_hd__clkinv_4_24/Y
+ sky130_fd_sc_hd__a21oi_1_361/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_761 VDD VSS sky130_fd_sc_hd__ha_2_134/A sky130_fd_sc_hd__dfxtp_1_764/CLK
+ sky130_fd_sc_hd__o21a_1_12/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_772 VDD VSS sky130_fd_sc_hd__fa_2_1071/A sky130_fd_sc_hd__clkinv_8_54/Y
+ sky130_fd_sc_hd__and2_0_308/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__ha_2_5 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_5/A sky130_fd_sc_hd__ha_2_4/B
+ sky130_fd_sc_hd__ha_2_5/SUM sky130_fd_sc_hd__ha_2_5/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__dfxtp_1_783 VDD VSS sky130_fd_sc_hd__fa_2_1082/A sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__mux2_2_58/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_794 VDD VSS sky130_fd_sc_hd__fa_2_1046/B sky130_fd_sc_hd__clkinv_8_54/Y
+ sky130_fd_sc_hd__and2_0_301/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_370 VSS VDD sky130_fd_sc_hd__clkbuf_1_371/A sky130_fd_sc_hd__buf_6_43/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_381 VSS VDD sky130_fd_sc_hd__a22oi_2_25/A1 sky130_fd_sc_hd__nor3_2_7/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_600 sky130_fd_sc_hd__fa_2_602/CIN sky130_fd_sc_hd__fa_2_598/A
+ sky130_fd_sc_hd__ha_2_129/B sky130_fd_sc_hd__fa_2_689/B sky130_fd_sc_hd__fa_2_695/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_392 VSS VDD sky130_fd_sc_hd__clkbuf_1_392/X sky130_fd_sc_hd__clkbuf_1_392/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_611 sky130_fd_sc_hd__fa_2_614/A sky130_fd_sc_hd__fa_2_611/SUM
+ sky130_fd_sc_hd__fa_2_611/A sky130_fd_sc_hd__fa_2_611/B sky130_fd_sc_hd__fa_2_617/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_16 VSS VDD sky130_fd_sc_hd__buf_4_12/A sky130_fd_sc_hd__dfxtp_1_458/Q
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_622 sky130_fd_sc_hd__maj3_1_117/B sky130_fd_sc_hd__maj3_1_118/A
+ sky130_fd_sc_hd__fa_2_622/A sky130_fd_sc_hd__fa_2_622/B sky130_fd_sc_hd__fa_2_623/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_27 VSS VDD sky130_fd_sc_hd__clkbuf_1_27/X sky130_fd_sc_hd__clkbuf_1_27/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_633 sky130_fd_sc_hd__maj3_1_114/B sky130_fd_sc_hd__maj3_1_115/A
+ sky130_fd_sc_hd__fa_2_633/A sky130_fd_sc_hd__fa_2_633/B sky130_fd_sc_hd__fa_2_634/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_38 VSS VDD sky130_fd_sc_hd__clkbuf_1_38/X sky130_fd_sc_hd__clkbuf_1_38/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_644 sky130_fd_sc_hd__fa_2_646/B sky130_fd_sc_hd__fa_2_641/A
+ sky130_fd_sc_hd__fa_2_700/B sky130_fd_sc_hd__ha_2_132/B sky130_fd_sc_hd__ha_2_132/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_49 VSS VDD sky130_fd_sc_hd__clkbuf_1_49/X sky130_fd_sc_hd__clkbuf_1_49/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_655 sky130_fd_sc_hd__fa_2_657/A sky130_fd_sc_hd__fa_2_652/A
+ sky130_fd_sc_hd__ha_2_135/B sky130_fd_sc_hd__ha_2_132/A sky130_fd_sc_hd__ha_2_132/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_666 sky130_fd_sc_hd__fa_2_665/B sky130_fd_sc_hd__fa_2_666/SUM
+ sky130_fd_sc_hd__fa_2_666/A sky130_fd_sc_hd__fa_2_666/B sky130_fd_sc_hd__fa_2_666/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_677 sky130_fd_sc_hd__fa_2_679/CIN sky130_fd_sc_hd__fa_2_671/B
+ sky130_fd_sc_hd__fa_2_677/A sky130_fd_sc_hd__fa_2_689/B sky130_fd_sc_hd__fa_2_692/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_688 sky130_fd_sc_hd__fa_2_687/B sky130_fd_sc_hd__fa_2_688/SUM
+ sky130_fd_sc_hd__ha_2_130/B sky130_fd_sc_hd__fa_2_688/B sky130_fd_sc_hd__fa_2_688/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_699 sky130_fd_sc_hd__fa_2_698/CIN sky130_fd_sc_hd__fa_2_699/SUM
+ sky130_fd_sc_hd__fa_2_699/A sky130_fd_sc_hd__fa_2_700/A sky130_fd_sc_hd__ha_2_134/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22oi_2_19 sky130_fd_sc_hd__nor3_2_7/Y sky130_fd_sc_hd__a22oi_2_19/A2
+ sky130_fd_sc_hd__nor3_2_8/Y sky130_fd_sc_hd__a22oi_2_19/B2 sky130_fd_sc_hd__a22oi_2_19/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_2
Xsky130_fd_sc_hd__buf_12_5 sky130_fd_sc_hd__inv_2_21/Y sky130_fd_sc_hd__buf_12_5/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__o22ai_1_120 sky130_fd_sc_hd__o21a_1_8/A2 sky130_fd_sc_hd__o22ai_1_120/B1
+ sky130_fd_sc_hd__nor2_1_85/B sky130_fd_sc_hd__nor2_1_70/B sky130_fd_sc_hd__o21ai_1_92/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_131 sky130_fd_sc_hd__nor2_1_74/A sky130_fd_sc_hd__nor2_2_9/B
+ sky130_fd_sc_hd__o22ai_1_131/Y sky130_fd_sc_hd__a21oi_1_123/Y sky130_fd_sc_hd__a211oi_1_7/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_142 sky130_fd_sc_hd__nand2_1_284/Y sky130_fd_sc_hd__nand2_2_5/Y
+ sky130_fd_sc_hd__o22ai_1_142/Y sky130_fd_sc_hd__xnor2_1_76/Y sky130_fd_sc_hd__o22ai_1_156/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_206 sky130_fd_sc_hd__o31ai_1_2/B1 sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__nand2_1_206/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_153 sky130_fd_sc_hd__nand2_1_338/A sky130_fd_sc_hd__nand2_1_284/Y
+ sky130_fd_sc_hd__o22ai_1_153/Y sky130_fd_sc_hd__xnor2_1_70/Y sky130_fd_sc_hd__o22ai_1_153/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_805 sky130_fd_sc_hd__o31ai_1_6/A1 sky130_fd_sc_hd__xnor2_1_93/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_805/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_217 sky130_fd_sc_hd__o22a_1_0/A2 sky130_fd_sc_hd__o21ai_1_35/B1
+ sky130_fd_sc_hd__o21ai_1_35/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_816 sky130_fd_sc_hd__nand2_1_371/B sky130_fd_sc_hd__fa_2_442/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_816/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_164 sky130_fd_sc_hd__nand2_1_316/Y sky130_fd_sc_hd__nand2_2_6/A
+ sky130_fd_sc_hd__o22ai_1_164/Y sky130_fd_sc_hd__nand2_1_339/A sky130_fd_sc_hd__a21oi_1_188/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_228 sky130_fd_sc_hd__o21ai_1_56/B1 sky130_fd_sc_hd__nor2_1_91/B
+ sky130_fd_sc_hd__nor2_1_41/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_175 sky130_fd_sc_hd__o22ai_1_195/B2 sky130_fd_sc_hd__o22ai_1_206/A1
+ sky130_fd_sc_hd__o22ai_1_175/Y sky130_fd_sc_hd__o22ai_1_206/B1 sky130_fd_sc_hd__nor2_1_120/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_827 sky130_fd_sc_hd__o22ai_1_250/B1 sky130_fd_sc_hd__fa_2_1138/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_827/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_239 sky130_fd_sc_hd__o21ai_1_83/B1 sky130_fd_sc_hd__nor2_1_60/B
+ sky130_fd_sc_hd__nor2_1_60/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_186 sky130_fd_sc_hd__o22ai_1_204/B1 sky130_fd_sc_hd__nor2_1_118/B
+ sky130_fd_sc_hd__o22ai_1_186/Y sky130_fd_sc_hd__o22ai_1_193/A1 sky130_fd_sc_hd__o22ai_1_206/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand4_1_12 sky130_fd_sc_hd__nand4_1_12/C sky130_fd_sc_hd__nand4_1_12/B
+ sky130_fd_sc_hd__nand4_1_12/Y sky130_fd_sc_hd__nand4_1_12/D sky130_fd_sc_hd__nand4_1_12/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__clkinv_1_838 sky130_fd_sc_hd__clkinv_1_838/Y sky130_fd_sc_hd__a21boi_1_2/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_838/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand4_1_23 sky130_fd_sc_hd__nand4_1_23/C sky130_fd_sc_hd__nand4_1_23/B
+ sky130_fd_sc_hd__nand4_1_23/Y sky130_fd_sc_hd__nand4_1_23/D sky130_fd_sc_hd__nand4_1_23/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__o22ai_1_197 sky130_fd_sc_hd__o22ai_1_197/A2 sky130_fd_sc_hd__o22ai_1_204/B1
+ sky130_fd_sc_hd__o22ai_1_197/Y sky130_fd_sc_hd__o22ai_1_206/B1 sky130_fd_sc_hd__o22ai_1_197/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_849 sky130_fd_sc_hd__nor2_1_181/A sky130_fd_sc_hd__fa_2_1156/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_849/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand4_1_34 sky130_fd_sc_hd__nand4_1_34/C sky130_fd_sc_hd__nand4_1_34/B
+ sky130_fd_sc_hd__nand4_1_34/Y sky130_fd_sc_hd__nand4_1_34/D sky130_fd_sc_hd__nand4_1_34/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_45 sky130_fd_sc_hd__nand4_1_45/C sky130_fd_sc_hd__nand4_1_45/B
+ sky130_fd_sc_hd__nand4_1_45/Y sky130_fd_sc_hd__nand4_1_45/D sky130_fd_sc_hd__nand4_1_45/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_56 sky130_fd_sc_hd__nand4_1_56/C sky130_fd_sc_hd__nand4_1_56/B
+ sky130_fd_sc_hd__buf_2_266/A sky130_fd_sc_hd__nand4_1_56/D sky130_fd_sc_hd__nand4_1_56/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_67 sky130_fd_sc_hd__nand4_1_67/C sky130_fd_sc_hd__nand4_1_67/B
+ sky130_fd_sc_hd__nand4_1_67/Y sky130_fd_sc_hd__nand4_1_67/D sky130_fd_sc_hd__nand4_1_67/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_78 sky130_fd_sc_hd__nand4_1_78/C sky130_fd_sc_hd__nand4_1_78/B
+ sky130_fd_sc_hd__nand2_1_1/B sky130_fd_sc_hd__nand4_1_78/D sky130_fd_sc_hd__nand4_1_78/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__conb_1_16 sky130_fd_sc_hd__conb_1_16/LO sky130_fd_sc_hd__conb_1_16/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_27 sky130_fd_sc_hd__conb_1_27/LO sky130_fd_sc_hd__conb_1_27/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__a211oi_1_30 sky130_fd_sc_hd__nor3_1_40/A sky130_fd_sc_hd__nor2_1_266/Y
+ sky130_fd_sc_hd__o22ai_1_373/Y sky130_fd_sc_hd__a211oi_1_30/Y sky130_fd_sc_hd__fa_2_1256/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_380 VSS VDD sky130_fd_sc_hd__o22ai_1_318/A2 sky130_fd_sc_hd__o21a_1_42/A2
+ sky130_fd_sc_hd__a21oi_1_355/Y sky130_fd_sc_hd__o21ai_1_380/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_391 VSS VDD sky130_fd_sc_hd__o22ai_1_349/A1 sky130_fd_sc_hd__nor2_1_247/Y
+ sky130_fd_sc_hd__or3_1_4/X sky130_fd_sc_hd__o21ai_1_391/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__mux2_2_60 VSS VDD sky130_fd_sc_hd__mux2_2_60/A1 sky130_fd_sc_hd__mux2_2_60/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_60/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_71 VSS VDD sky130_fd_sc_hd__mux2_2_71/A1 sky130_fd_sc_hd__mux2_2_71/A0
+ sky130_fd_sc_hd__mux2_2_75/S sky130_fd_sc_hd__mux2_2_71/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_82 VSS VDD sky130_fd_sc_hd__mux2_2_82/A1 sky130_fd_sc_hd__mux2_2_82/A0
+ sky130_fd_sc_hd__nor2_4_15/A sky130_fd_sc_hd__mux2_2_82/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1101 sky130_fd_sc_hd__fa_2_1102/CIN sky130_fd_sc_hd__and2_0_310/A
+ sky130_fd_sc_hd__fa_2_1101/A sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1101/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__mux2_2_93 VSS VDD sky130_fd_sc_hd__mux2_2_93/A1 sky130_fd_sc_hd__mux2_2_93/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_93/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1112 sky130_fd_sc_hd__fa_2_1113/CIN sky130_fd_sc_hd__fa_2_1112/SUM
+ sky130_fd_sc_hd__fa_2_1112/A sky130_fd_sc_hd__fa_2_1112/B sky130_fd_sc_hd__fa_2_1112/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1123 sky130_fd_sc_hd__fa_2_1124/CIN sky130_fd_sc_hd__and2_0_321/A
+ sky130_fd_sc_hd__fa_2_1123/A sky130_fd_sc_hd__fa_2_1123/B sky130_fd_sc_hd__fa_2_1123/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1134 sky130_fd_sc_hd__fa_2_1135/CIN sky130_fd_sc_hd__mux2_2_89/A1
+ sky130_fd_sc_hd__fa_2_1134/A sky130_fd_sc_hd__fa_2_1134/B sky130_fd_sc_hd__fa_2_1134/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1145 sky130_fd_sc_hd__fa_2_1146/CIN sky130_fd_sc_hd__mux2_2_107/A1
+ sky130_fd_sc_hd__fa_2_1145/A sky130_fd_sc_hd__fa_2_1145/B sky130_fd_sc_hd__fa_2_1145/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1156 sky130_fd_sc_hd__fa_2_1157/CIN sky130_fd_sc_hd__mux2_2_80/A0
+ sky130_fd_sc_hd__fa_2_1156/A sky130_fd_sc_hd__fa_2_1156/B sky130_fd_sc_hd__fa_2_1156/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1167 sky130_fd_sc_hd__fa_2_1168/CIN sky130_fd_sc_hd__mux2_2_106/A1
+ sky130_fd_sc_hd__fa_2_1167/A sky130_fd_sc_hd__fa_2_1172/B sky130_fd_sc_hd__fa_2_1167/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1178 sky130_fd_sc_hd__fa_2_1179/CIN sky130_fd_sc_hd__mux2_2_156/A1
+ sky130_fd_sc_hd__fa_2_1178/A sky130_fd_sc_hd__fa_2_1178/B sky130_fd_sc_hd__fa_2_1178/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1189 sky130_fd_sc_hd__fa_2_1190/CIN sky130_fd_sc_hd__mux2_2_129/A0
+ sky130_fd_sc_hd__fa_2_1189/A sky130_fd_sc_hd__fa_2_1189/B sky130_fd_sc_hd__fa_2_1189/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_580 VDD VSS sky130_fd_sc_hd__nor4_1_7/B sky130_fd_sc_hd__dfxtp_1_591/CLK
+ sky130_fd_sc_hd__and2_0_249/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_591 VDD VSS sky130_fd_sc_hd__or4_1_2/A sky130_fd_sc_hd__dfxtp_1_591/CLK
+ sky130_fd_sc_hd__a21o_2_1/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_430 sky130_fd_sc_hd__fa_2_428/B sky130_fd_sc_hd__fa_2_429/B
+ sky130_fd_sc_hd__ha_2_117/B sky130_fd_sc_hd__fa_2_546/A sky130_fd_sc_hd__fa_2_427/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_441 sky130_fd_sc_hd__fa_2_431/B sky130_fd_sc_hd__fa_2_434/B
+ sky130_fd_sc_hd__ha_2_124/A sky130_fd_sc_hd__ha_2_124/B sky130_fd_sc_hd__fa_2_543/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o2bb2ai_1_7 sky130_fd_sc_hd__o2bb2ai_1_7/Y sky130_fd_sc_hd__nor2_1_18/Y
+ sky130_fd_sc_hd__ha_2_152/SUM sky130_fd_sc_hd__o21ai_1_31/A1 sky130_fd_sc_hd__nor2_1_11/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_452 sky130_fd_sc_hd__fa_2_448/CIN sky130_fd_sc_hd__nor2_1_171/A
+ sky130_fd_sc_hd__fa_2_452/A sky130_fd_sc_hd__fa_2_452/B sky130_fd_sc_hd__fa_2_452/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_463 sky130_fd_sc_hd__fa_2_456/A sky130_fd_sc_hd__fa_2_460/B
+ sky130_fd_sc_hd__fa_2_463/A sky130_fd_sc_hd__fa_2_463/B sky130_fd_sc_hd__fa_2_463/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_474 sky130_fd_sc_hd__fa_2_476/B sky130_fd_sc_hd__fa_2_474/SUM
+ sky130_fd_sc_hd__ha_2_119/B sky130_fd_sc_hd__fa_2_564/B sky130_fd_sc_hd__fa_2_474/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_485 sky130_fd_sc_hd__maj3_1_97/B sky130_fd_sc_hd__maj3_1_98/A
+ sky130_fd_sc_hd__fa_2_485/A sky130_fd_sc_hd__fa_2_485/B sky130_fd_sc_hd__fa_2_486/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_2_1 VDD VSS sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__and2_2_1/X
+ sky130_fd_sc_hd__ha_2_56/A VDD VSS sky130_fd_sc_hd__and2_2
Xsky130_fd_sc_hd__fa_2_496 sky130_fd_sc_hd__fa_2_497/CIN sky130_fd_sc_hd__fa_2_490/A
+ sky130_fd_sc_hd__ha_2_119/A sky130_fd_sc_hd__fa_2_554/A sky130_fd_sc_hd__fa_2_555/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor2_1_206 sky130_fd_sc_hd__nor2_1_206/B sky130_fd_sc_hd__nor2_1_206/Y
+ sky130_fd_sc_hd__nor2_1_224/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_217 sky130_fd_sc_hd__nor2_1_217/B sky130_fd_sc_hd__nor2_1_217/Y
+ sky130_fd_sc_hd__nor2_1_225/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_228 sky130_fd_sc_hd__nor2_1_228/B sky130_fd_sc_hd__o21a_1_44/A1
+ sky130_fd_sc_hd__o21a_1_45/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_239 sky130_fd_sc_hd__nor2_1_239/B sky130_fd_sc_hd__o21a_1_53/A1
+ sky130_fd_sc_hd__nor2_1_239/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_402 sky130_fd_sc_hd__buf_12_402/A sky130_fd_sc_hd__buf_12_500/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_413 sky130_fd_sc_hd__buf_8_220/X sky130_fd_sc_hd__buf_12_413/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_424 sky130_fd_sc_hd__buf_8_218/X sky130_fd_sc_hd__buf_12_424/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_435 sky130_fd_sc_hd__buf_8_213/X sky130_fd_sc_hd__buf_12_435/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_446 sky130_fd_sc_hd__buf_6_78/X sky130_fd_sc_hd__buf_12_446/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_305 sky130_fd_sc_hd__clkbuf_4_165/X sky130_fd_sc_hd__clkinv_2_23/Y
+ sky130_fd_sc_hd__clkbuf_1_401/X sky130_fd_sc_hd__a22oi_1_305/A2 sky130_fd_sc_hd__a22oi_1_305/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_457 sky130_fd_sc_hd__buf_6_62/X sky130_fd_sc_hd__buf_12_486/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_316 sky130_fd_sc_hd__clkbuf_1_376/X sky130_fd_sc_hd__nor2_2_5/Y
+ sky130_fd_sc_hd__buf_2_204/X sky130_fd_sc_hd__clkbuf_1_459/X sky130_fd_sc_hd__nand4_1_78/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_468 sky130_fd_sc_hd__buf_4_119/X sky130_fd_sc_hd__buf_12_468/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_327 sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__fa_2_991/A
+ sky130_fd_sc_hd__xor2_1_60/A sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__a22oi_1_327/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_479 sky130_fd_sc_hd__buf_12_479/A sky130_fd_sc_hd__buf_12_479/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_338 sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_2_7/Y
+ sky130_fd_sc_hd__fa_2_996/A sky130_fd_sc_hd__fa_2_997/A sky130_fd_sc_hd__a22oi_1_338/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_349 sky130_fd_sc_hd__nor2_2_12/Y sky130_fd_sc_hd__fa_2_1065/A
+ sky130_fd_sc_hd__fa_2_1068/A sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__a22oi_1_349/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_602 sky130_fd_sc_hd__ha_2_177/B sky130_fd_sc_hd__fa_2_1038/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_602/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_613 sky130_fd_sc_hd__o22ai_1_132/B1 sky130_fd_sc_hd__nor2_2_7/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_613/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_624 sky130_fd_sc_hd__nor2_1_128/A sky130_fd_sc_hd__xor2_1_87/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_624/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_635 sky130_fd_sc_hd__o22ai_1_153/B2 sky130_fd_sc_hd__ha_2_196/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_635/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_646 sky130_fd_sc_hd__o21ai_1_190/A2 sky130_fd_sc_hd__o2bb2ai_1_32/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_646/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_657 sky130_fd_sc_hd__nand2_1_288/B sky130_fd_sc_hd__nor2_1_107/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_657/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_668 sky130_fd_sc_hd__o21ai_1_195/A1 sky130_fd_sc_hd__nand2_1_297/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_668/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_679 sky130_fd_sc_hd__nor2_1_103/B sky130_fd_sc_hd__fa_2_1111/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_679/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand3_1_8 sky130_fd_sc_hd__nand3_1_8/Y sky130_fd_sc_hd__nand3_1_8/A
+ sky130_fd_sc_hd__nand3_1_8/C sky130_fd_sc_hd__nand3_1_8/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__a222oi_1_11 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1144/A sky130_fd_sc_hd__nor2_2_15/Y
+ sky130_fd_sc_hd__nor3_1_38/A sky130_fd_sc_hd__fa_2_1146/A sky130_fd_sc_hd__nor3_1_38/B
+ sky130_fd_sc_hd__a222oi_1_11/Y sky130_fd_sc_hd__fa_2_1143/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_22 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1194/A sky130_fd_sc_hd__nor2_2_16/Y
+ sky130_fd_sc_hd__nor3_1_39/A sky130_fd_sc_hd__fa_2_1196/A sky130_fd_sc_hd__nor3_1_39/B
+ sky130_fd_sc_hd__nor2_1_221/B sky130_fd_sc_hd__fa_2_1193/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_33 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1244/A sky130_fd_sc_hd__nor2_2_17/Y
+ sky130_fd_sc_hd__nor3_1_40/A sky130_fd_sc_hd__fa_2_1246/A sky130_fd_sc_hd__nor3_1_40/B
+ sky130_fd_sc_hd__a222oi_1_33/Y sky130_fd_sc_hd__fa_2_1243/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_13 VSS VDD sky130_fd_sc_hd__xnor2_1_19/Y sky130_fd_sc_hd__xnor2_1_13/Y
+ sky130_fd_sc_hd__ha_2_149/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_24 VSS VDD sky130_fd_sc_hd__xor2_1_26/X sky130_fd_sc_hd__xor2_1_25/B
+ sky130_fd_sc_hd__xnor2_1_25/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_35 VSS VDD sky130_fd_sc_hd__xnor2_1_36/B sky130_fd_sc_hd__xnor2_1_35/Y
+ sky130_fd_sc_hd__xnor2_1_35/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_46 VSS VDD sky130_fd_sc_hd__xnor2_1_46/B sky130_fd_sc_hd__xnor2_1_46/Y
+ sky130_fd_sc_hd__nor2_1_45/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_570 sky130_fd_sc_hd__nor2_1_321/B sky130_fd_sc_hd__nor2_1_323/A
+ sky130_fd_sc_hd__nor2_1_319/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_57 VSS VDD sky130_fd_sc_hd__xnor2_1_57/B sky130_fd_sc_hd__xnor2_1_57/Y
+ sky130_fd_sc_hd__nor2_1_48/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_68 VSS VDD sky130_fd_sc_hd__xnor2_1_69/B sky130_fd_sc_hd__xnor2_1_68/Y
+ sky130_fd_sc_hd__xnor2_1_68/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_79 VSS VDD sky130_fd_sc_hd__xnor2_1_79/B sky130_fd_sc_hd__xnor2_1_79/Y
+ sky130_fd_sc_hd__nor2_1_96/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__a211oi_1_4 sky130_fd_sc_hd__or3_1_1/B sky130_fd_sc_hd__o21ai_1_39/Y
+ sky130_fd_sc_hd__or3_1_1/A sky130_fd_sc_hd__a31oi_1_1/A1 sky130_fd_sc_hd__or3_1_1/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o32ai_1_7 sky130_fd_sc_hd__o32ai_1_7/A2 sky130_fd_sc_hd__o32ai_1_7/Y
+ sky130_fd_sc_hd__fa_2_1244/A sky130_fd_sc_hd__o32ai_1_7/A3 sky130_fd_sc_hd__o32ai_1_7/B2
+ sky130_fd_sc_hd__fa_2_1243/A VDD VSS VSS VDD sky130_fd_sc_hd__o32ai_1
Xsky130_fd_sc_hd__clkbuf_16_5 sky130_fd_sc_hd__buf_8_61/A sky130_fd_sc_hd__clkbuf_16_5/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__fa_2_260 sky130_fd_sc_hd__fa_2_263/B sky130_fd_sc_hd__fa_2_260/SUM
+ sky130_fd_sc_hd__fa_2_260/A sky130_fd_sc_hd__fa_2_260/B sky130_fd_sc_hd__fa_2_260/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_271 sky130_fd_sc_hd__fa_2_169/A sky130_fd_sc_hd__fa_2_171/B
+ sky130_fd_sc_hd__fa_2_271/A sky130_fd_sc_hd__fa_2_271/B sky130_fd_sc_hd__fa_2_276/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_282 sky130_fd_sc_hd__fa_2_165/CIN sky130_fd_sc_hd__fa_2_278/A
+ sky130_fd_sc_hd__ha_2_97/A sky130_fd_sc_hd__ha_2_99/A sky130_fd_sc_hd__fa_2_258/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_293 sky130_fd_sc_hd__fa_2_285/CIN sky130_fd_sc_hd__nor2_1_211/A
+ sky130_fd_sc_hd__fa_2_293/A sky130_fd_sc_hd__fa_2_293/B sky130_fd_sc_hd__fa_2_293/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor4_1_5 sky130_fd_sc_hd__nor4_1_5/D sky130_fd_sc_hd__nor4_1_5/C
+ sky130_fd_sc_hd__nor4_1_5/Y sky130_fd_sc_hd__or4_1_2/A sky130_fd_sc_hd__nor4_1_5/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__nor4_1
Xsky130_fd_sc_hd__a22oi_1_4 sky130_fd_sc_hd__nor2_2_0/Y sky130_fd_sc_hd__clkinv_1_4/Y
+ sky130_fd_sc_hd__nand4_1_29/Y sky130_fd_sc_hd__nand4_1_13/Y sky130_fd_sc_hd__a22oi_1_4/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__diode_2_110 sky130_fd_sc_hd__buf_2_225/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_121 sky130_fd_sc_hd__buf_2_250/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_132 sky130_fd_sc_hd__clkbuf_1_526/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_143 sky130_fd_sc_hd__buf_2_168/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_154 sky130_fd_sc_hd__clkbuf_4_172/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_165 sky130_fd_sc_hd__nand4_1_70/D VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_176 sky130_fd_sc_hd__nand4_1_77/D VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_187 sky130_fd_sc_hd__buf_6_53/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_198 sky130_fd_sc_hd__clkbuf_4_210/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkbuf_4_207 sky130_fd_sc_hd__buf_2_225/A sky130_fd_sc_hd__clkbuf_4_207/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_218 sky130_fd_sc_hd__nand3_1_16/A frequency_adc_done VSS
+ VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_12_210 sky130_fd_sc_hd__buf_6_22/X sky130_fd_sc_hd__buf_12_243/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_221 sky130_fd_sc_hd__buf_6_30/X sky130_fd_sc_hd__buf_12_229/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_232 sky130_fd_sc_hd__buf_12_232/A sky130_fd_sc_hd__buf_12_264/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_243 sky130_fd_sc_hd__buf_12_243/A sky130_fd_sc_hd__buf_12_260/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_90 sky130_fd_sc_hd__a21o_2_3/A2 sky130_fd_sc_hd__o21ai_1_107/Y
+ sky130_fd_sc_hd__a21oi_1_90/Y sky130_fd_sc_hd__fa_2_991/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_1_102 sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__a22oi_2_12/A1
+ sky130_fd_sc_hd__buf_2_77/X sky130_fd_sc_hd__clkbuf_1_168/X sky130_fd_sc_hd__a22oi_1_102/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_254 sky130_fd_sc_hd__buf_12_254/A sky130_fd_sc_hd__buf_12_254/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_113 sky130_fd_sc_hd__a22oi_1_97/B1 sky130_fd_sc_hd__a22oi_1_97/A1
+ sky130_fd_sc_hd__buf_2_58/X sky130_fd_sc_hd__clkbuf_4_82/X sky130_fd_sc_hd__nand4_1_23/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_265 sky130_fd_sc_hd__buf_12_265/A sky130_fd_sc_hd__buf_12_265/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_124 sky130_fd_sc_hd__a22oi_1_96/B1 sky130_fd_sc_hd__a22oi_1_96/A1
+ sky130_fd_sc_hd__clkbuf_1_144/X sky130_fd_sc_hd__a22oi_1_124/A2 sky130_fd_sc_hd__nand4_1_26/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_276 sky130_fd_sc_hd__buf_12_276/A sky130_fd_sc_hd__buf_6_41/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_135 sky130_fd_sc_hd__a22oi_1_96/B1 sky130_fd_sc_hd__a22oi_1_96/A1
+ sky130_fd_sc_hd__clkbuf_1_141/X sky130_fd_sc_hd__a22oi_1_135/A2 sky130_fd_sc_hd__nand4_1_29/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_287 sky130_fd_sc_hd__buf_8_129/X sky130_fd_sc_hd__buf_12_287/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_146 sky130_fd_sc_hd__clkbuf_4_72/X sky130_fd_sc_hd__clkbuf_4_73/X
+ sky130_fd_sc_hd__a22oi_1_146/B2 sky130_fd_sc_hd__buf_2_82/X sky130_fd_sc_hd__buf_2_100/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_298 sky130_fd_sc_hd__buf_8_122/X sky130_fd_sc_hd__buf_12_298/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_157 sky130_fd_sc_hd__clkbuf_4_111/X sky130_fd_sc_hd__clkbuf_4_112/X
+ sky130_fd_sc_hd__a22oi_1_157/B2 sky130_fd_sc_hd__clkbuf_1_295/X sky130_fd_sc_hd__a22oi_1_157/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_168 sky130_fd_sc_hd__clkbuf_1_351/X sky130_fd_sc_hd__clkbuf_1_353/X
+ sky130_fd_sc_hd__clkinv_2_12/Y sky130_fd_sc_hd__a22oi_1_168/A2 sky130_fd_sc_hd__nand4_1_37/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_410 sky130_fd_sc_hd__o221ai_1_0/B2 sky130_fd_sc_hd__nor2b_1_86/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_410/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22oi_1_179 sky130_fd_sc_hd__clkbuf_1_265/X sky130_fd_sc_hd__clkbuf_1_266/X
+ sky130_fd_sc_hd__clkbuf_1_274/X sky130_fd_sc_hd__a22oi_1_179/A2 sky130_fd_sc_hd__a22oi_1_179/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_421 sky130_fd_sc_hd__nand3_1_48/A sky130_fd_sc_hd__fa_2_960/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_421/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_432 sky130_fd_sc_hd__fa_2_968/B sky130_fd_sc_hd__dfxtp_1_480/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_432/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_443 sky130_fd_sc_hd__fa_2_959/B sky130_fd_sc_hd__dfxtp_1_489/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_443/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_454 sky130_fd_sc_hd__fa_2_947/B sky130_fd_sc_hd__dfxtp_1_501/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_454/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_465 sky130_fd_sc_hd__o22ai_1_77/B2 sky130_fd_sc_hd__ha_2_182/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_465/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_476 sky130_fd_sc_hd__o22ai_1_81/B2 sky130_fd_sc_hd__ha_2_178/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_476/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_487 sky130_fd_sc_hd__nor2_1_48/B sky130_fd_sc_hd__nand2_1_250/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_487/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_498 sky130_fd_sc_hd__o21ai_1_80/B1 sky130_fd_sc_hd__nor2_1_56/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_498/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_340 sky130_fd_sc_hd__fa_2_1183/A sky130_fd_sc_hd__o22ai_1_309/Y
+ sky130_fd_sc_hd__a21oi_1_340/Y sky130_fd_sc_hd__nor2_2_16/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_351 sky130_fd_sc_hd__or2_0_10/B sky130_fd_sc_hd__o21ai_1_375/Y
+ sky130_fd_sc_hd__a21oi_1_351/Y sky130_fd_sc_hd__o21ai_1_376/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_362 sky130_fd_sc_hd__o21a_1_45/B1 sky130_fd_sc_hd__o21a_1_44/A1
+ sky130_fd_sc_hd__a21oi_1_362/Y sky130_fd_sc_hd__nor2_1_228/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_373 sky130_fd_sc_hd__nor2_1_239/A sky130_fd_sc_hd__o21a_1_53/A1
+ sky130_fd_sc_hd__a21oi_1_373/Y sky130_fd_sc_hd__nor2_1_239/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_384 sky130_fd_sc_hd__clkinv_1_987/Y sky130_fd_sc_hd__clkinv_1_986/Y
+ sky130_fd_sc_hd__a21oi_1_384/Y sky130_fd_sc_hd__nand2_1_491/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_395 sky130_fd_sc_hd__fa_2_1232/A sky130_fd_sc_hd__o22ai_1_360/Y
+ sky130_fd_sc_hd__a21oi_1_395/Y sky130_fd_sc_hd__nor2_2_17/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__xor2_1_206 sky130_fd_sc_hd__fa_2_1173/A sky130_fd_sc_hd__xor2_1_206/X
+ sky130_fd_sc_hd__xor2_1_206/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_217 sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__fa_2_1201/B
+ sky130_fd_sc_hd__xor2_1_217/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_228 sky130_fd_sc_hd__xor2_1_228/B sky130_fd_sc_hd__xor2_1_228/X
+ sky130_fd_sc_hd__xor2_1_229/X VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_239 sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1236/B
+ sky130_fd_sc_hd__xor2_1_239/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_2_11 VDD VSS sky130_fd_sc_hd__buf_2_11/X sky130_fd_sc_hd__ha_2_13/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_22 VDD VSS sky130_fd_sc_hd__buf_2_22/X sky130_fd_sc_hd__buf_2_22/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_33 VDD VSS sky130_fd_sc_hd__ha_2_21/A sky130_fd_sc_hd__buf_2_33/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_44 VDD VSS sky130_fd_sc_hd__buf_2_44/X sky130_fd_sc_hd__ha_2_35/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_55 VDD VSS sky130_fd_sc_hd__buf_2_55/X sky130_fd_sc_hd__buf_2_55/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_66 VDD VSS sky130_fd_sc_hd__buf_2_66/X sky130_fd_sc_hd__buf_2_66/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_77 VDD VSS sky130_fd_sc_hd__buf_2_77/X sky130_fd_sc_hd__buf_2_77/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_88 VDD VSS sky130_fd_sc_hd__buf_2_88/X sky130_fd_sc_hd__buf_2_88/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_99 VDD VSS sky130_fd_sc_hd__buf_2_99/X sky130_fd_sc_hd__buf_2_99/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o211ai_1_60 sky130_fd_sc_hd__nor2_1_307/A sky130_fd_sc_hd__nor2_1_299/B
+ sky130_fd_sc_hd__xor2_1_306/A sky130_fd_sc_hd__nand2_1_530/Y sky130_fd_sc_hd__nand2_1_532/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__diode_2_6 sky130_fd_sc_hd__clkbuf_1_247/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__o211ai_1_71 sky130_fd_sc_hd__a21oi_1_474/Y sky130_fd_sc_hd__nor2_1_307/A
+ sky130_fd_sc_hd__xor2_1_293/A sky130_fd_sc_hd__a21oi_1_471/Y sky130_fd_sc_hd__nand2_1_545/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__and2_0_208 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_208/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_208/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_219 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_219/X sky130_fd_sc_hd__and2_0_235/B
+ sky130_fd_sc_hd__and2_0_219/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_240 sky130_fd_sc_hd__buf_8_211/A sky130_fd_sc_hd__clkinv_1_240/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_240/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_251 sky130_fd_sc_hd__inv_2_127/A sky130_fd_sc_hd__inv_2_117/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_251/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_262 sky130_fd_sc_hd__nor3_1_27/C sky130_fd_sc_hd__nor3_1_26/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_262/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_273 sky130_fd_sc_hd__nor3_1_26/C sky130_fd_sc_hd__nor3_1_27/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_273/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_2_7 sky130_fd_sc_hd__or2_1_1/B sky130_fd_sc_hd__ha_2_81/A sky130_fd_sc_hd__a22o_2_7/X
+ sky130_fd_sc_hd__a22o_2_7/B2 sky130_fd_sc_hd__a22o_4_0/B1 VDD VSS VDD VSS sky130_fd_sc_hd__a22o_2
Xsky130_fd_sc_hd__o31ai_1_6 sky130_fd_sc_hd__o31ai_1_6/Y sky130_fd_sc_hd__o31ai_1_6/A2
+ sky130_fd_sc_hd__o31ai_1_6/A1 sky130_fd_sc_hd__o31ai_1_6/A3 sky130_fd_sc_hd__o31ai_1_6/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__o31ai_1
Xsky130_fd_sc_hd__clkinv_1_284 sky130_fd_sc_hd__fa_2_66/B sky130_fd_sc_hd__fa_2_87/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_284/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_295 sky130_fd_sc_hd__fa_2_280/A sky130_fd_sc_hd__fa_2_5/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_295/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_3 sky130_fd_sc_hd__nor2_1_21/A sky130_fd_sc_hd__o21ai_1_6/Y
+ sky130_fd_sc_hd__a21oi_1_3/Y sky130_fd_sc_hd__xor2_1_11/X VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkbuf_4_16 sky130_fd_sc_hd__clkbuf_4_16/X sky130_fd_sc_hd__clkbuf_4_16/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__o21ai_1_209 VSS VDD sky130_fd_sc_hd__o21ai_1_209/A2 sky130_fd_sc_hd__o22ai_1_206/A1
+ sky130_fd_sc_hd__a22oi_1_347/Y sky130_fd_sc_hd__o21ai_1_209/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__clkbuf_4_27 sky130_fd_sc_hd__clkbuf_4_27/X sky130_fd_sc_hd__clkbuf_4_27/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_38 sky130_fd_sc_hd__clkbuf_4_38/X sky130_fd_sc_hd__clkbuf_4_38/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_49 sky130_fd_sc_hd__nand4_1_8/D sky130_fd_sc_hd__a22oi_1_55/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__a21oi_1_170 sky130_fd_sc_hd__clkinv_1_665/Y sky130_fd_sc_hd__nor2_1_94/B
+ sky130_fd_sc_hd__xnor2_1_73/A sky130_fd_sc_hd__xnor2_1_71/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_181 sky130_fd_sc_hd__o21a_1_11/B1 sky130_fd_sc_hd__o21a_1_10/A1
+ sky130_fd_sc_hd__dfxtp_1_764/D sky130_fd_sc_hd__nor2_1_114/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_192 sky130_fd_sc_hd__clkinv_1_695/Y sky130_fd_sc_hd__clkinv_1_694/Y
+ sky130_fd_sc_hd__a21oi_1_192/Y sky130_fd_sc_hd__nand2_1_331/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_100 sky130_fd_sc_hd__inv_2_63/Y sky130_fd_sc_hd__buf_8_100/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_111 sky130_fd_sc_hd__buf_8_111/A sky130_fd_sc_hd__buf_8_111/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_122 sky130_fd_sc_hd__buf_8_122/A sky130_fd_sc_hd__buf_8_122/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_133 sky130_fd_sc_hd__buf_8_133/A sky130_fd_sc_hd__buf_6_37/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_144 sky130_fd_sc_hd__inv_2_93/Y sky130_fd_sc_hd__buf_8_144/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nor2_4_6 sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__nor2_4_6/A
+ sky130_fd_sc_hd__nor2_4_6/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__buf_8_155 sky130_fd_sc_hd__buf_8_155/A sky130_fd_sc_hd__buf_8_155/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_166 sky130_fd_sc_hd__buf_8_166/A sky130_fd_sc_hd__buf_4_95/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_177 sky130_fd_sc_hd__buf_8_177/A sky130_fd_sc_hd__buf_8_177/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_188 sky130_fd_sc_hd__buf_8_188/A sky130_fd_sc_hd__buf_8_188/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_199 sky130_fd_sc_hd__buf_8_199/A sky130_fd_sc_hd__buf_8_199/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_409 VDD VSS sky130_fd_sc_hd__nor2_1_41/B sky130_fd_sc_hd__dfxtp_1_425/CLK
+ sky130_fd_sc_hd__and2_0_106/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a21o_2_12 sky130_fd_sc_hd__a21o_2_12/X sky130_fd_sc_hd__nor2_1_208/Y
+ sky130_fd_sc_hd__nor2_1_208/A sky130_fd_sc_hd__nor2_1_208/B VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__a21o_2_23 sky130_fd_sc_hd__a21o_2_23/X sky130_fd_sc_hd__nor2_1_256/Y
+ sky130_fd_sc_hd__nor2_1_256/A sky130_fd_sc_hd__or3_1_4/X VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__clkinv_8_19 sky130_fd_sc_hd__clkinv_8_19/Y sky130_fd_sc_hd__clkinv_8_0/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_19/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__xor2_1_50 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_977/B
+ sky130_fd_sc_hd__xor2_1_50/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_61 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__xor2_1_61/X
+ sky130_fd_sc_hd__xor2_1_61/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_17 sky130_fd_sc_hd__inv_2_41/Y sky130_fd_sc_hd__buf_12_17/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_72 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__xor2_1_72/X
+ sky130_fd_sc_hd__xor2_1_72/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_28 sky130_fd_sc_hd__buf_8_44/X sky130_fd_sc_hd__buf_12_28/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_83 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__xor2_1_83/X
+ sky130_fd_sc_hd__xor2_1_83/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_39 sky130_fd_sc_hd__buf_8_13/X sky130_fd_sc_hd__buf_12_39/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_94 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__xor2_1_94/X
+ sky130_fd_sc_hd__xor2_1_94/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2b_1_0 sky130_fd_sc_hd__nand2b_1_0/Y sky130_fd_sc_hd__nand3_2_2/A
+ sky130_fd_sc_hd__inv_8_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__dfxtp_1_1305 VDD VSS sky130_fd_sc_hd__fa_2_846/B sky130_fd_sc_hd__dfxtp_1_1322/CLK
+ sky130_fd_sc_hd__a21oi_1_434/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1316 VDD VSS sky130_fd_sc_hd__xnor2_1_7/A sky130_fd_sc_hd__dfxtp_1_1329/CLK
+ sky130_fd_sc_hd__xnor2_1_101/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1327 VDD VSS sky130_fd_sc_hd__fa_2_911/A sky130_fd_sc_hd__dfxtp_1_1329/CLK
+ sky130_fd_sc_hd__o21a_1_58/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1338 VDD VSS sky130_fd_sc_hd__fa_2_1297/A sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__mux2_2_254/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_910 VDD VSS sky130_fd_sc_hd__or2_0_9/A sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__nor2b_1_106/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1349 VDD VSS sky130_fd_sc_hd__fa_2_1308/A sky130_fd_sc_hd__clkinv_8_51/Y
+ sky130_fd_sc_hd__mux2_2_226/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_921 VDD VSS sky130_fd_sc_hd__fa_2_1150/A sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__mux2_2_93/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_932 VDD VSS sky130_fd_sc_hd__fa_2_1124/A sky130_fd_sc_hd__clkinv_8_55/Y
+ sky130_fd_sc_hd__mux2_2_117/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_943 VDD VSS sky130_fd_sc_hd__fa_2_1135/A sky130_fd_sc_hd__clkinv_8_46/Y
+ sky130_fd_sc_hd__mux2_2_87/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_954 VDD VSS sky130_fd_sc_hd__fa_2_1163/A sky130_fd_sc_hd__clkinv_8_64/Y
+ sky130_fd_sc_hd__mux2_2_118/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_965 VDD VSS sky130_fd_sc_hd__nor2b_1_104/A sky130_fd_sc_hd__clkinv_8_46/Y
+ sky130_fd_sc_hd__nor2b_1_111/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_976 VDD VSS sky130_fd_sc_hd__mux2_2_102/A0 sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__o22ai_1_219/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_987 VDD VSS sky130_fd_sc_hd__mux2_2_77/A1 sky130_fd_sc_hd__clkinv_8_46/Y
+ sky130_fd_sc_hd__dfxtp_1_987/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_998 VDD VSS sky130_fd_sc_hd__mux2_2_103/A0 sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__dfxtp_1_998/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_530 VSS VDD sky130_fd_sc_hd__buf_2_211/A sky130_fd_sc_hd__clkbuf_1_530/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_541 VSS VDD sky130_fd_sc_hd__clkbuf_1_541/X sky130_fd_sc_hd__clkbuf_1_541/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_552 VSS VDD sky130_fd_sc_hd__xor2_1_267/B sky130_fd_sc_hd__fa_2_1242/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_120 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_169/B sky130_fd_sc_hd__fa_2_487/B
+ sky130_fd_sc_hd__fa_2_483/A sky130_fd_sc_hd__ha_2_124/A sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_563 VSS VDD sky130_fd_sc_hd__nand2_1_111/B sky130_fd_sc_hd__nand4_1_49/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_131 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_131/A sky130_fd_sc_hd__fa_2_602/A
+ sky130_fd_sc_hd__fa_2_599/B sky130_fd_sc_hd__ha_2_131/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_574 VSS VDD sky130_fd_sc_hd__dfxtp_1_66/D sky130_fd_sc_hd__nand4_1_36/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_142 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_142/A sky130_fd_sc_hd__fa_2_739/A
+ sky130_fd_sc_hd__fa_2_736/B sky130_fd_sc_hd__ha_2_142/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_585 VSS VDD sky130_fd_sc_hd__nand3_1_7/B sky130_fd_sc_hd__a22oi_1_14/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_153 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_153/A sky130_fd_sc_hd__ha_2_152/B
+ sky130_fd_sc_hd__ha_2_153/SUM sky130_fd_sc_hd__ha_2_153/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_596 VSS VDD sky130_fd_sc_hd__dfxtp_1_63/D sky130_fd_sc_hd__nand4_1_33/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_804 sky130_fd_sc_hd__fa_2_713/A sky130_fd_sc_hd__fa_2_714/B
+ sky130_fd_sc_hd__fa_2_804/A sky130_fd_sc_hd__fa_2_804/B sky130_fd_sc_hd__fa_2_810/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_164 VSS VDD VSS VDD sky130_fd_sc_hd__or4_1_1/B sky130_fd_sc_hd__ha_2_163/B
+ sky130_fd_sc_hd__ha_2_164/SUM sky130_fd_sc_hd__ha_2_164/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_815 sky130_fd_sc_hd__fa_2_814/B sky130_fd_sc_hd__fa_2_815/SUM
+ sky130_fd_sc_hd__fa_2_815/A sky130_fd_sc_hd__fa_2_815/B sky130_fd_sc_hd__fa_2_815/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_175 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_175/A sky130_fd_sc_hd__ha_2_174/A
+ sky130_fd_sc_hd__ha_2_175/SUM sky130_fd_sc_hd__ha_2_175/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_826 sky130_fd_sc_hd__fa_2_825/B sky130_fd_sc_hd__fa_2_826/SUM
+ sky130_fd_sc_hd__fa_2_826/A sky130_fd_sc_hd__fa_2_834/B sky130_fd_sc_hd__fa_2_826/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_186 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_186/A sky130_fd_sc_hd__nor2_1_141/A
+ sky130_fd_sc_hd__ha_2_186/SUM sky130_fd_sc_hd__ha_2_186/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_837 sky130_fd_sc_hd__fa_2_836/CIN sky130_fd_sc_hd__fa_2_837/SUM
+ sky130_fd_sc_hd__fa_2_837/A sky130_fd_sc_hd__fa_2_837/B sky130_fd_sc_hd__fa_2_837/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_197 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_197/A sky130_fd_sc_hd__ha_2_196/A
+ sky130_fd_sc_hd__ha_2_197/SUM sky130_fd_sc_hd__ha_2_197/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_848 sky130_fd_sc_hd__fa_2_847/CIN sky130_fd_sc_hd__fa_2_848/SUM
+ sky130_fd_sc_hd__fa_2_848/A sky130_fd_sc_hd__fa_2_848/B sky130_fd_sc_hd__fa_2_848/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_859 sky130_fd_sc_hd__fa_2_858/CIN sky130_fd_sc_hd__fa_2_859/SUM
+ sky130_fd_sc_hd__fa_2_859/A sky130_fd_sc_hd__fa_2_859/B sky130_fd_sc_hd__fa_2_859/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__maj3_1_2 sky130_fd_sc_hd__maj3_1_3/X sky130_fd_sc_hd__maj3_1_2/X
+ sky130_fd_sc_hd__maj3_1_2/B sky130_fd_sc_hd__maj3_1_2/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__mux2_2_104 VSS VDD sky130_fd_sc_hd__mux2_2_104/A1 sky130_fd_sc_hd__mux2_2_104/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_104/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_115 VSS VDD sky130_fd_sc_hd__mux2_2_115/A1 sky130_fd_sc_hd__mux2_2_115/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_115/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_126 VSS VDD sky130_fd_sc_hd__mux2_2_126/A1 sky130_fd_sc_hd__mux2_2_126/A0
+ sky130_fd_sc_hd__mux2_2_135/S sky130_fd_sc_hd__mux2_2_126/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_137 VSS VDD sky130_fd_sc_hd__mux2_2_137/A1 sky130_fd_sc_hd__mux2_2_137/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_137/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_148 VSS VDD sky130_fd_sc_hd__mux2_2_148/A1 sky130_fd_sc_hd__mux2_2_148/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_148/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_159 VSS VDD sky130_fd_sc_hd__mux2_2_159/A1 sky130_fd_sc_hd__mux2_2_159/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_159/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__and2_0_11 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_11/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_6/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_22 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_22/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_17/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_302 sky130_fd_sc_hd__o22ai_1_322/A2 sky130_fd_sc_hd__o22ai_1_309/B1
+ sky130_fd_sc_hd__o22ai_1_302/Y sky130_fd_sc_hd__nor2_1_186/B sky130_fd_sc_hd__o22ai_1_318/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_33 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_33/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_39/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_313 sky130_fd_sc_hd__o32ai_1_5/A3 sky130_fd_sc_hd__o22ai_1_316/B1
+ sky130_fd_sc_hd__o22ai_1_313/Y sky130_fd_sc_hd__nor2_1_220/A sky130_fd_sc_hd__o21a_1_42/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_44 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_55/A sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__ha_2_53/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_108 sky130_fd_sc_hd__maj3_1_109/X sky130_fd_sc_hd__maj3_1_108/X
+ sky130_fd_sc_hd__maj3_1_108/B sky130_fd_sc_hd__maj3_1_108/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_324 sky130_fd_sc_hd__nand2_1_462/Y sky130_fd_sc_hd__o21ai_1_385/Y
+ sky130_fd_sc_hd__o22ai_1_324/Y sky130_fd_sc_hd__nand2_1_471/B sky130_fd_sc_hd__nand2_1_461/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_55 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_55/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_55/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_119 sky130_fd_sc_hd__maj3_1_120/X sky130_fd_sc_hd__maj3_1_119/X
+ sky130_fd_sc_hd__maj3_1_119/B sky130_fd_sc_hd__maj3_1_119/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_335 sky130_fd_sc_hd__nand2_1_462/Y sky130_fd_sc_hd__nand2_1_461/Y
+ sky130_fd_sc_hd__o22ai_1_335/Y sky130_fd_sc_hd__o22ai_1_348/A1 sky130_fd_sc_hd__a21o_2_23/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_66 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_79/A sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__ha_2_72/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_346 sky130_fd_sc_hd__nand2_1_464/Y sky130_fd_sc_hd__nand2_1_463/Y
+ sky130_fd_sc_hd__o22ai_1_346/Y sky130_fd_sc_hd__o22ai_1_346/A1 sky130_fd_sc_hd__a21o_2_22/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_77 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_77/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__and2_0_77/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_357 sky130_fd_sc_hd__o22ai_1_379/A2 sky130_fd_sc_hd__nor2_1_261/A
+ sky130_fd_sc_hd__o22ai_1_357/Y sky130_fd_sc_hd__o22ai_1_366/B1 sky130_fd_sc_hd__o32ai_1_8/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_2_3 sky130_fd_sc_hd__nor2_2_3/B sky130_fd_sc_hd__nor2_2_3/Y
+ sky130_fd_sc_hd__nor3_2_5/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__and2_0_88 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_88/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_88/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_368 sky130_fd_sc_hd__o22ai_1_379/A2 sky130_fd_sc_hd__nor2_1_235/B
+ sky130_fd_sc_hd__o22ai_1_368/Y sky130_fd_sc_hd__o22ai_1_379/B1 sky130_fd_sc_hd__o32ai_1_8/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_99 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_99/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_99/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_379 sky130_fd_sc_hd__o22ai_1_379/A2 sky130_fd_sc_hd__o22ai_1_379/B1
+ sky130_fd_sc_hd__o22ai_1_379/Y sky130_fd_sc_hd__nor2_1_238/B sky130_fd_sc_hd__o32ai_1_8/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_8_10 sky130_fd_sc_hd__buf_8_15/A sky130_fd_sc_hd__buf_8_10/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_21 sky130_fd_sc_hd__ha_2_26/A sky130_fd_sc_hd__buf_8_21/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_32 sky130_fd_sc_hd__buf_8_32/A sky130_fd_sc_hd__buf_8_32/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_43 sky130_fd_sc_hd__buf_8_43/A sky130_fd_sc_hd__buf_8_43/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_54 sky130_fd_sc_hd__buf_8_54/A sky130_fd_sc_hd__buf_8_54/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_65 sky130_fd_sc_hd__inv_2_68/A sky130_fd_sc_hd__buf_8_65/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_76 sky130_fd_sc_hd__buf_8_76/A sky130_fd_sc_hd__buf_8_83/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_87 sky130_fd_sc_hd__buf_8_87/A sky130_fd_sc_hd__buf_8_87/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_206 VDD VSS sky130_fd_sc_hd__ha_2_75/A sky130_fd_sc_hd__dfxtp_1_207/CLK
+ sky130_fd_sc_hd__and2_0_74/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_8_98 sky130_fd_sc_hd__inv_2_67/Y sky130_fd_sc_hd__buf_8_98/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_217 VDD VSS sky130_fd_sc_hd__ha_2_86/A sky130_fd_sc_hd__dfxtp_1_224/CLK
+ sky130_fd_sc_hd__nor2b_1_47/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_228 VDD VSS sky130_fd_sc_hd__nor2_2_5/A sky130_fd_sc_hd__clkinv_8_102/Y
+ sky130_fd_sc_hd__a22o_1_32/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_239 VDD VSS sky130_fd_sc_hd__fa_2_870/A sky130_fd_sc_hd__dfxtp_1_472/CLK
+ sky130_fd_sc_hd__and2_0_181/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_2_106 VDD VSS sky130_fd_sc_hd__buf_2_106/X sky130_fd_sc_hd__buf_2_106/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__fa_2_1305 sky130_fd_sc_hd__fa_2_1306/CIN sky130_fd_sc_hd__mux2_2_232/A1
+ sky130_fd_sc_hd__fa_2_1305/A sky130_fd_sc_hd__fa_2_1305/B sky130_fd_sc_hd__fa_2_1305/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_117 VDD VSS sky130_fd_sc_hd__buf_2_117/X sky130_fd_sc_hd__inv_2_46/Y
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__fa_2_1316 sky130_fd_sc_hd__fa_2_1317/CIN sky130_fd_sc_hd__mux2_2_262/A1
+ sky130_fd_sc_hd__fa_2_1316/A sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1316/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_128 VDD VSS sky130_fd_sc_hd__buf_8_135/A sky130_fd_sc_hd__a22o_2_3/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_139 VDD VSS sky130_fd_sc_hd__buf_2_139/X sky130_fd_sc_hd__buf_6_50/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1102 VDD VSS sky130_fd_sc_hd__fa_2_1221/A sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__mux2_2_145/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1113 VDD VSS sky130_fd_sc_hd__mux2_2_162/A0 sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__a21oi_1_318/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1124 VDD VSS sky130_fd_sc_hd__mux2_2_133/A1 sky130_fd_sc_hd__clkinv_8_70/Y
+ sky130_fd_sc_hd__o22ai_1_269/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1135 VDD VSS sky130_fd_sc_hd__mux2_2_163/A0 sky130_fd_sc_hd__clkinv_8_64/Y
+ sky130_fd_sc_hd__dfxtp_1_994/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1146 VDD VSS sky130_fd_sc_hd__mux2_2_155/A0 sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__o22ai_1_291/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1157 VDD VSS sky130_fd_sc_hd__mux2_2_128/A1 sky130_fd_sc_hd__clkinv_8_70/Y
+ sky130_fd_sc_hd__o22ai_1_280/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1168 VDD VSS sky130_fd_sc_hd__fa_2_856/B sky130_fd_sc_hd__dfxtp_1_1184/CLK
+ sky130_fd_sc_hd__o21a_1_52/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_740 VDD VSS sky130_fd_sc_hd__and2_0_166/A sky130_fd_sc_hd__dfxtp_1_744/CLK
+ sky130_fd_sc_hd__fa_2_1095/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1179 VDD VSS sky130_fd_sc_hd__fa_2_932/A sky130_fd_sc_hd__dfxtp_1_1179/CLK
+ sky130_fd_sc_hd__o21a_1_48/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_751 VDD VSS sky130_fd_sc_hd__and2_0_177/A sky130_fd_sc_hd__dfxtp_1_768/CLK
+ sky130_fd_sc_hd__fa_2_1106/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_762 VDD VSS sky130_fd_sc_hd__fa_2_659/A sky130_fd_sc_hd__dfxtp_1_764/CLK
+ sky130_fd_sc_hd__dfxtp_1_762/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_773 VDD VSS sky130_fd_sc_hd__fa_2_1072/A sky130_fd_sc_hd__clkinv_8_54/Y
+ sky130_fd_sc_hd__and2_0_311/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__ha_2_6 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_6/A sky130_fd_sc_hd__ha_2_5/B
+ sky130_fd_sc_hd__ha_2_6/SUM sky130_fd_sc_hd__ha_2_6/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__dfxtp_1_784 VDD VSS sky130_fd_sc_hd__fa_2_1083/A sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__mux2_2_56/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_795 VDD VSS sky130_fd_sc_hd__fa_2_1047/A sky130_fd_sc_hd__clkinv_8_54/Y
+ sky130_fd_sc_hd__and2_0_303/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_360 VSS VDD sky130_fd_sc_hd__clkbuf_1_361/A sky130_fd_sc_hd__buf_8_117/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_371 VSS VDD sky130_fd_sc_hd__buf_6_33/A sky130_fd_sc_hd__clkbuf_1_371/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_382 VSS VDD sky130_fd_sc_hd__clkbuf_1_382/X sky130_fd_sc_hd__clkbuf_1_541/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_393 VSS VDD sky130_fd_sc_hd__a22oi_2_19/B2 sky130_fd_sc_hd__clkbuf_1_393/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_601 sky130_fd_sc_hd__maj3_1_123/B sky130_fd_sc_hd__maj3_1_124/A
+ sky130_fd_sc_hd__fa_2_601/A sky130_fd_sc_hd__fa_2_601/B sky130_fd_sc_hd__fa_2_602/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_612 sky130_fd_sc_hd__fa_2_611/B sky130_fd_sc_hd__fa_2_612/SUM
+ sky130_fd_sc_hd__ha_2_130/B sky130_fd_sc_hd__ha_2_131/A sky130_fd_sc_hd__ha_2_129/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_17 VSS VDD sky130_fd_sc_hd__clkinv_1_21/A sky130_fd_sc_hd__ha_2_27/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_623 sky130_fd_sc_hd__fa_2_626/B sky130_fd_sc_hd__fa_2_623/SUM
+ sky130_fd_sc_hd__fa_2_623/A sky130_fd_sc_hd__fa_2_676/B sky130_fd_sc_hd__fa_2_623/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_28 VSS VDD sky130_fd_sc_hd__clkbuf_1_28/X sky130_fd_sc_hd__clkbuf_1_28/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_634 sky130_fd_sc_hd__fa_2_638/B sky130_fd_sc_hd__fa_2_634/SUM
+ sky130_fd_sc_hd__fa_2_634/A sky130_fd_sc_hd__fa_2_634/B sky130_fd_sc_hd__fa_2_640/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_39 VSS VDD sky130_fd_sc_hd__clkbuf_1_39/X sky130_fd_sc_hd__clkbuf_1_39/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_645 sky130_fd_sc_hd__maj3_1_111/B sky130_fd_sc_hd__maj3_1_112/A
+ sky130_fd_sc_hd__fa_2_645/A sky130_fd_sc_hd__fa_2_645/B sky130_fd_sc_hd__fa_2_646/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_656 sky130_fd_sc_hd__maj3_1_108/B sky130_fd_sc_hd__maj3_1_109/A
+ sky130_fd_sc_hd__fa_2_656/A sky130_fd_sc_hd__fa_2_656/B sky130_fd_sc_hd__fa_2_657/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_667 sky130_fd_sc_hd__fa_2_669/CIN sky130_fd_sc_hd__fa_2_662/B
+ sky130_fd_sc_hd__ha_2_135/A sky130_fd_sc_hd__fa_2_667/B sky130_fd_sc_hd__ha_2_131/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_678 sky130_fd_sc_hd__fa_2_679/B sky130_fd_sc_hd__fa_2_671/A
+ sky130_fd_sc_hd__ha_2_135/A sky130_fd_sc_hd__fa_2_678/B sky130_fd_sc_hd__fa_2_699/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_689 sky130_fd_sc_hd__fa_2_688/CIN sky130_fd_sc_hd__fa_2_689/SUM
+ sky130_fd_sc_hd__fa_2_698/A sky130_fd_sc_hd__fa_2_689/B sky130_fd_sc_hd__fa_2_695/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__conb_1_0 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__conb_1_0/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__buf_12_6 sky130_fd_sc_hd__inv_2_13/Y sky130_fd_sc_hd__buf_12_6/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__o22ai_1_110 sky130_fd_sc_hd__o21a_1_8/A2 sky130_fd_sc_hd__o22ai_1_110/B1
+ sky130_fd_sc_hd__nor2_1_82/B sky130_fd_sc_hd__nor2_1_65/B sky130_fd_sc_hd__o21ai_1_92/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_121 sky130_fd_sc_hd__o22ai_1_132/B1 sky130_fd_sc_hd__o22ai_1_130/B1
+ sky130_fd_sc_hd__nor2_1_85/A sky130_fd_sc_hd__nor2_1_70/A sky130_fd_sc_hd__o22ai_1_121/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_132 sky130_fd_sc_hd__nor2_1_87/A sky130_fd_sc_hd__o22ai_1_132/B1
+ sky130_fd_sc_hd__o22ai_1_132/Y sky130_fd_sc_hd__o21ai_1_92/A1 sky130_fd_sc_hd__o22ai_1_132/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_143 sky130_fd_sc_hd__nand2_1_284/Y sky130_fd_sc_hd__nand2_2_5/Y
+ sky130_fd_sc_hd__o22ai_1_143/Y sky130_fd_sc_hd__xnor2_1_78/Y sky130_fd_sc_hd__o22ai_1_157/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_207 sky130_fd_sc_hd__o31ai_1_2/A3 sky130_fd_sc_hd__or4_1_2/B
+ sky130_fd_sc_hd__or4_1_2/D VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2_2_10 sky130_fd_sc_hd__nor2_2_10/B sky130_fd_sc_hd__nor2_2_10/Y
+ sky130_fd_sc_hd__nor2_2_11/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__o22ai_1_154 sky130_fd_sc_hd__nand2_1_338/A sky130_fd_sc_hd__nand2_1_284/Y
+ sky130_fd_sc_hd__o22ai_1_154/Y sky130_fd_sc_hd__xnor2_1_72/Y sky130_fd_sc_hd__o22ai_1_154/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_806 sky130_fd_sc_hd__nor2_1_163/A sky130_fd_sc_hd__or3_1_2/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_806/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_218 sky130_fd_sc_hd__o22ai_1_58/B2 sky130_fd_sc_hd__o21ai_1_36/B1
+ sky130_fd_sc_hd__o21ai_1_36/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_817 sky130_fd_sc_hd__nand2_1_372/B sky130_fd_sc_hd__fa_2_448/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_817/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_165 sky130_fd_sc_hd__nand2_2_6/Y sky130_fd_sc_hd__nor2_1_127/A
+ sky130_fd_sc_hd__a211o_1_9/C1 sky130_fd_sc_hd__a21oi_1_189/Y sky130_fd_sc_hd__a21oi_1_190/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_229 sky130_fd_sc_hd__a22o_1_68/B2 sky130_fd_sc_hd__xnor2_1_34/B
+ sky130_fd_sc_hd__xnor2_1_33/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_176 sky130_fd_sc_hd__o21a_1_16/A2 sky130_fd_sc_hd__o22ai_1_190/A1
+ sky130_fd_sc_hd__nor2_1_129/B sky130_fd_sc_hd__nor2_1_116/B sky130_fd_sc_hd__o22ai_1_206/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_828 sky130_fd_sc_hd__nor2_1_143/B sky130_fd_sc_hd__fa_2_1135/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_828/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_187 sky130_fd_sc_hd__nand4_1_86/B sky130_fd_sc_hd__o22ai_1_206/A1
+ sky130_fd_sc_hd__o22ai_1_187/Y sky130_fd_sc_hd__o22ai_1_206/B1 sky130_fd_sc_hd__o22ai_1_195/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_839 sky130_fd_sc_hd__o21ai_1_317/B1 sky130_fd_sc_hd__nor2_1_177/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_839/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand4_1_13 sky130_fd_sc_hd__nand4_1_13/C sky130_fd_sc_hd__nand4_1_13/B
+ sky130_fd_sc_hd__nand4_1_13/Y sky130_fd_sc_hd__nand4_1_13/D sky130_fd_sc_hd__nand4_1_13/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__o211ai_1_0 sky130_fd_sc_hd__nor3_2_1/A sky130_fd_sc_hd__nor3_2_1/B
+ sky130_fd_sc_hd__o21a_1_0/A2 sky130_fd_sc_hd__nor3_1_2/C sky130_fd_sc_hd__nor3_1_4/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__nand4_1_24 sky130_fd_sc_hd__nand4_1_24/C sky130_fd_sc_hd__nand4_1_24/B
+ sky130_fd_sc_hd__nand4_1_24/Y sky130_fd_sc_hd__nand4_1_24/D sky130_fd_sc_hd__nand4_1_24/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__o22ai_1_198 sky130_fd_sc_hd__nor2_1_127/A sky130_fd_sc_hd__nor2_2_13/B
+ sky130_fd_sc_hd__o22ai_1_198/Y sky130_fd_sc_hd__a21oi_1_234/Y sky130_fd_sc_hd__a222oi_1_3/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand4_1_35 sky130_fd_sc_hd__nand4_1_35/C sky130_fd_sc_hd__nand4_1_35/B
+ sky130_fd_sc_hd__nand4_1_35/Y sky130_fd_sc_hd__nand4_1_35/D sky130_fd_sc_hd__nand4_1_35/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_46 sky130_fd_sc_hd__nand4_1_46/C sky130_fd_sc_hd__nand4_1_46/B
+ sky130_fd_sc_hd__nand4_1_46/Y sky130_fd_sc_hd__nand4_1_46/D sky130_fd_sc_hd__nand4_1_46/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_57 sky130_fd_sc_hd__nand4_1_57/C sky130_fd_sc_hd__nand4_1_57/B
+ sky130_fd_sc_hd__nand4_1_57/Y sky130_fd_sc_hd__nand4_1_57/D sky130_fd_sc_hd__nand4_1_57/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_68 sky130_fd_sc_hd__nand4_1_68/C sky130_fd_sc_hd__nand4_1_68/B
+ sky130_fd_sc_hd__nand4_1_68/Y sky130_fd_sc_hd__nand4_1_68/D sky130_fd_sc_hd__nand4_1_68/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_79 sky130_fd_sc_hd__nand4_1_79/C sky130_fd_sc_hd__nand4_1_79/B
+ sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__nand4_1_79/D sky130_fd_sc_hd__nand4_1_79/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__conb_1_17 sky130_fd_sc_hd__conb_1_17/LO sky130_fd_sc_hd__conb_1_17/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_28 sky130_fd_sc_hd__conb_1_28/LO sky130_fd_sc_hd__conb_1_28/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__a211oi_1_20 sky130_fd_sc_hd__nor2b_2_3/Y sky130_fd_sc_hd__o22ai_1_306/Y
+ sky130_fd_sc_hd__nor2_1_217/Y sky130_fd_sc_hd__a211oi_1_20/Y sky130_fd_sc_hd__o21ai_1_361/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_370 VSS VDD sky130_fd_sc_hd__o22ai_1_315/B1 sky130_fd_sc_hd__o21a_1_42/A1
+ sky130_fd_sc_hd__a21oi_1_343/Y sky130_fd_sc_hd__o21ai_1_370/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a211oi_1_31 sky130_fd_sc_hd__nor2b_2_4/Y sky130_fd_sc_hd__o22ai_1_376/Y
+ sky130_fd_sc_hd__nor2_1_268/Y sky130_fd_sc_hd__a211oi_1_31/Y sky130_fd_sc_hd__o21ai_1_437/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_381 VSS VDD sky130_fd_sc_hd__nor2_1_214/A sky130_fd_sc_hd__o21a_1_42/X
+ sky130_fd_sc_hd__a211oi_1_24/Y sky130_fd_sc_hd__xor2_1_205/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_392 VSS VDD sky130_fd_sc_hd__nor2_1_248/Y sky130_fd_sc_hd__or3_1_4/C
+ sky130_fd_sc_hd__nor2_1_245/A sky130_fd_sc_hd__o21ai_1_392/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__mux2_2_50 VSS VDD sky130_fd_sc_hd__mux2_2_50/A1 sky130_fd_sc_hd__mux2_2_50/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_50/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_61 VSS VDD sky130_fd_sc_hd__mux2_2_61/A1 sky130_fd_sc_hd__mux2_2_61/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_61/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_72 VSS VDD sky130_fd_sc_hd__mux2_2_72/A1 sky130_fd_sc_hd__mux2_2_72/A0
+ sky130_fd_sc_hd__mux2_2_75/S sky130_fd_sc_hd__mux2_2_72/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_83 VSS VDD sky130_fd_sc_hd__mux2_2_83/A1 sky130_fd_sc_hd__mux2_2_83/A0
+ sky130_fd_sc_hd__nor2_4_15/A sky130_fd_sc_hd__mux2_2_83/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1102 sky130_fd_sc_hd__fa_2_1103/CIN sky130_fd_sc_hd__and2_0_315/A
+ sky130_fd_sc_hd__fa_2_1102/A sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1102/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__mux2_2_94 VSS VDD sky130_fd_sc_hd__mux2_2_94/A1 sky130_fd_sc_hd__mux2_2_94/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_94/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1113 sky130_fd_sc_hd__fa_2_1114/CIN sky130_fd_sc_hd__fa_2_1113/SUM
+ sky130_fd_sc_hd__fa_2_1113/A sky130_fd_sc_hd__fa_2_1113/B sky130_fd_sc_hd__fa_2_1113/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1124 sky130_fd_sc_hd__fa_2_1125/CIN sky130_fd_sc_hd__mux2_2_117/A1
+ sky130_fd_sc_hd__fa_2_1124/A sky130_fd_sc_hd__fa_2_1124/B sky130_fd_sc_hd__fa_2_1124/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1135 sky130_fd_sc_hd__fa_2_1136/CIN sky130_fd_sc_hd__mux2_2_87/A0
+ sky130_fd_sc_hd__fa_2_1135/A sky130_fd_sc_hd__fa_2_1135/B sky130_fd_sc_hd__fa_2_1135/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1146 sky130_fd_sc_hd__fa_2_1147/CIN sky130_fd_sc_hd__mux2_2_104/A1
+ sky130_fd_sc_hd__fa_2_1146/A sky130_fd_sc_hd__fa_2_1146/B sky130_fd_sc_hd__fa_2_1146/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1157 sky130_fd_sc_hd__xor2_1_162/B sky130_fd_sc_hd__mux2_2_78/A0
+ sky130_fd_sc_hd__fa_2_1157/A sky130_fd_sc_hd__fa_2_1157/B sky130_fd_sc_hd__fa_2_1157/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1168 sky130_fd_sc_hd__fa_2_1169/CIN sky130_fd_sc_hd__mux2_2_103/A1
+ sky130_fd_sc_hd__fa_2_1168/A sky130_fd_sc_hd__fa_2_1172/B sky130_fd_sc_hd__fa_2_1168/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1179 sky130_fd_sc_hd__fa_2_1180/CIN sky130_fd_sc_hd__mux2_2_153/A1
+ sky130_fd_sc_hd__fa_2_1179/A sky130_fd_sc_hd__fa_2_1179/B sky130_fd_sc_hd__fa_2_1179/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_570 VDD VSS sky130_fd_sc_hd__a22o_1_35/B1 sky130_fd_sc_hd__dfxtp_1_576/CLK
+ sky130_fd_sc_hd__a22o_1_35/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_581 VDD VSS sky130_fd_sc_hd__nor4_1_6/A sky130_fd_sc_hd__dfxtp_1_594/CLK
+ sky130_fd_sc_hd__and2_0_245/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_592 VDD VSS sky130_fd_sc_hd__or4_1_2/B sky130_fd_sc_hd__dfxtp_1_595/CLK
+ sky130_fd_sc_hd__a21o_2_2/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_190 VSS VDD sky130_fd_sc_hd__clkbuf_1_190/X sky130_fd_sc_hd__nand3_1_29/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_420 sky130_fd_sc_hd__fa_2_419/B sky130_fd_sc_hd__fa_2_420/SUM
+ sky130_fd_sc_hd__fa_2_420/A sky130_fd_sc_hd__fa_2_420/B sky130_fd_sc_hd__fa_2_425/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_431 sky130_fd_sc_hd__fa_2_429/CIN sky130_fd_sc_hd__a21o_2_7/A1
+ sky130_fd_sc_hd__fa_2_431/A sky130_fd_sc_hd__fa_2_431/B sky130_fd_sc_hd__fa_2_431/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_442 sky130_fd_sc_hd__fa_2_435/CIN sky130_fd_sc_hd__fa_2_442/SUM
+ sky130_fd_sc_hd__fa_2_442/A sky130_fd_sc_hd__fa_2_442/B sky130_fd_sc_hd__fa_2_442/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o2bb2ai_1_8 sky130_fd_sc_hd__o2bb2ai_1_8/Y sky130_fd_sc_hd__nor2_1_18/Y
+ sky130_fd_sc_hd__ha_2_151/SUM sky130_fd_sc_hd__o21ai_1_31/A1 sky130_fd_sc_hd__o22ai_1_0/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_453 sky130_fd_sc_hd__fa_2_449/CIN sky130_fd_sc_hd__fa_2_455/A
+ sky130_fd_sc_hd__ha_2_125/A sky130_fd_sc_hd__ha_2_121/B sky130_fd_sc_hd__fa_2_551/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_464 sky130_fd_sc_hd__fa_2_460/CIN sky130_fd_sc_hd__or3_1_2/B
+ sky130_fd_sc_hd__fa_2_464/A sky130_fd_sc_hd__fa_2_464/B sky130_fd_sc_hd__maj3_1_82/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_475 sky130_fd_sc_hd__fa_2_477/CIN sky130_fd_sc_hd__fa_2_473/B
+ sky130_fd_sc_hd__ha_2_124/B sky130_fd_sc_hd__fa_2_535/A sky130_fd_sc_hd__fa_2_559/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_486 sky130_fd_sc_hd__fa_2_489/A sky130_fd_sc_hd__fa_2_486/SUM
+ sky130_fd_sc_hd__fa_2_486/A sky130_fd_sc_hd__fa_2_486/B sky130_fd_sc_hd__fa_2_486/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_497 sky130_fd_sc_hd__fa_2_499/CIN sky130_fd_sc_hd__fa_2_494/A
+ sky130_fd_sc_hd__fa_2_497/A sky130_fd_sc_hd__fa_2_497/B sky130_fd_sc_hd__fa_2_497/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor2_1_207 sky130_fd_sc_hd__nor2_1_207/B sky130_fd_sc_hd__nor2_1_207/Y
+ sky130_fd_sc_hd__nor2_1_224/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_218 sky130_fd_sc_hd__o21a_1_42/A1 sky130_fd_sc_hd__nor2_1_218/Y
+ sky130_fd_sc_hd__nor2_1_218/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_229 sky130_fd_sc_hd__nor2_1_229/B sky130_fd_sc_hd__o21a_1_45/A1
+ sky130_fd_sc_hd__o21a_1_46/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_403 sky130_fd_sc_hd__buf_8_197/X sky130_fd_sc_hd__buf_12_465/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_414 sky130_fd_sc_hd__buf_8_199/X sky130_fd_sc_hd__buf_12_463/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_425 sky130_fd_sc_hd__buf_8_210/X sky130_fd_sc_hd__buf_12_425/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_436 sky130_fd_sc_hd__buf_8_208/X sky130_fd_sc_hd__buf_12_443/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_447 sky130_fd_sc_hd__buf_4_118/X sky130_fd_sc_hd__buf_12_447/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_306 sky130_fd_sc_hd__clkbuf_1_378/X sky130_fd_sc_hd__clkbuf_1_379/X
+ sky130_fd_sc_hd__clkbuf_4_166/X sky130_fd_sc_hd__buf_2_190/X sky130_fd_sc_hd__nand4_1_76/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_458 sky130_fd_sc_hd__buf_6_72/X sky130_fd_sc_hd__buf_12_458/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_317 sky130_fd_sc_hd__clkbuf_4_165/X sky130_fd_sc_hd__clkinv_2_23/Y
+ sky130_fd_sc_hd__clkbuf_1_398/X sky130_fd_sc_hd__a22oi_1_317/A2 sky130_fd_sc_hd__a22oi_1_317/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_469 sky130_fd_sc_hd__buf_6_81/X sky130_fd_sc_hd__buf_12_469/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_328 sky130_fd_sc_hd__fa_2_989/A sky130_fd_sc_hd__fa_2_987/A
+ sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__nor2_2_7/Y sky130_fd_sc_hd__nand3_1_49/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_339 sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_2_8/Y
+ sky130_fd_sc_hd__fa_2_1004/A sky130_fd_sc_hd__fa_2_1007/A sky130_fd_sc_hd__a22oi_1_339/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_603 sky130_fd_sc_hd__ha_2_178/B sky130_fd_sc_hd__fa_2_1037/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_603/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_614 sky130_fd_sc_hd__a21o_2_3/A2 sky130_fd_sc_hd__o21a_1_8/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_614/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_625 sky130_fd_sc_hd__o21ai_1_251/A2 sky130_fd_sc_hd__a21o_2_5/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_625/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_636 sky130_fd_sc_hd__o22ai_1_154/B2 sky130_fd_sc_hd__ha_2_195/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_636/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_647 sky130_fd_sc_hd__nand2_1_293/B sky130_fd_sc_hd__nor2_1_112/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_647/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_658 sky130_fd_sc_hd__nor2_1_93/B sky130_fd_sc_hd__nand2_1_302/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_658/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_669 sky130_fd_sc_hd__clkinv_1_669/Y sky130_fd_sc_hd__nor2_1_96/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_669/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand3_1_9 sky130_fd_sc_hd__nand3_1_9/Y sky130_fd_sc_hd__nand3_1_9/A
+ sky130_fd_sc_hd__nand3_1_9/C sky130_fd_sc_hd__nand3_1_9/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__a21oi_1_500 sky130_fd_sc_hd__nor2_1_319/Y sky130_fd_sc_hd__or2_0_0/B
+ sky130_fd_sc_hd__nand2_1_568/A sky130_fd_sc_hd__nor2_1_318/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_12 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1143/A sky130_fd_sc_hd__nor2_2_15/Y
+ sky130_fd_sc_hd__nor3_1_38/A sky130_fd_sc_hd__fa_2_1145/A sky130_fd_sc_hd__nor3_1_38/B
+ sky130_fd_sc_hd__nor2_1_179/B sky130_fd_sc_hd__fa_2_1142/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_23 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1193/A sky130_fd_sc_hd__nor2_2_16/Y
+ sky130_fd_sc_hd__nor3_1_39/A sky130_fd_sc_hd__fa_2_1195/A sky130_fd_sc_hd__nor3_1_39/B
+ sky130_fd_sc_hd__a222oi_1_23/Y sky130_fd_sc_hd__fa_2_1192/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_34 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1294/A sky130_fd_sc_hd__nor2_2_18/Y
+ sky130_fd_sc_hd__nor3_1_41/A sky130_fd_sc_hd__fa_2_1296/A sky130_fd_sc_hd__nor3_1_41/B
+ sky130_fd_sc_hd__a222oi_1_34/Y sky130_fd_sc_hd__fa_2_1293/B sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_14 VSS VDD sky130_fd_sc_hd__maj3_1_1/A sky130_fd_sc_hd__xnor2_1_14/Y
+ sky130_fd_sc_hd__ha_2_148/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_25 VSS VDD sky130_fd_sc_hd__ha_2_117/B sky130_fd_sc_hd__xnor2_1_25/Y
+ sky130_fd_sc_hd__xnor2_1_25/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_36 VSS VDD sky130_fd_sc_hd__xnor2_1_36/B sky130_fd_sc_hd__xnor2_1_36/Y
+ sky130_fd_sc_hd__xnor2_1_36/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_560 sky130_fd_sc_hd__nand2_1_560/Y sky130_fd_sc_hd__buf_6_89/A
+ sky130_fd_sc_hd__nand2_1_560/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_47 VSS VDD sky130_fd_sc_hd__xnor2_1_48/B sky130_fd_sc_hd__xnor2_1_47/Y
+ sky130_fd_sc_hd__xnor2_1_47/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_571 sky130_fd_sc_hd__nor2b_1_142/A load_en sky130_fd_sc_hd__buf_6_86/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_58 VSS VDD sky130_fd_sc_hd__xnor2_1_58/B sky130_fd_sc_hd__xnor2_1_58/Y
+ sky130_fd_sc_hd__nor2_1_48/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_69 VSS VDD sky130_fd_sc_hd__xnor2_1_69/B sky130_fd_sc_hd__xnor2_1_69/Y
+ sky130_fd_sc_hd__xnor2_1_69/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__a211oi_1_5 sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__nor2_1_86/Y
+ sky130_fd_sc_hd__o22ai_1_128/Y sky130_fd_sc_hd__a211oi_1_5/Y sky130_fd_sc_hd__fa_2_1013/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__or4_1_0 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__or4_1_0/A sky130_fd_sc_hd__or4_1_0/X
+ sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__or4_1_0/D VDD VSS VDD VSS sky130_fd_sc_hd__or4_1
Xsky130_fd_sc_hd__o32ai_1_8 sky130_fd_sc_hd__nor3_1_40/C sky130_fd_sc_hd__o32ai_1_8/Y
+ sky130_fd_sc_hd__o32ai_1_8/A1 sky130_fd_sc_hd__o32ai_1_8/A3 sky130_fd_sc_hd__o32ai_1_8/B2
+ sky130_fd_sc_hd__o32ai_1_8/B1 VDD VSS VSS VDD sky130_fd_sc_hd__o32ai_1
Xsky130_fd_sc_hd__clkbuf_16_6 sky130_fd_sc_hd__buf_12_256/A sky130_fd_sc_hd__inv_2_57/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__fa_2_250 sky130_fd_sc_hd__fa_2_252/CIN sky130_fd_sc_hd__fa_2_245/A
+ sky130_fd_sc_hd__fa_2_250/A sky130_fd_sc_hd__fa_2_250/B sky130_fd_sc_hd__fa_2_250/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_261 sky130_fd_sc_hd__fa_2_262/CIN sky130_fd_sc_hd__fa_2_256/A
+ sky130_fd_sc_hd__fa_2_261/A sky130_fd_sc_hd__fa_2_273/A sky130_fd_sc_hd__fa_2_250/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_272 sky130_fd_sc_hd__fa_2_271/B sky130_fd_sc_hd__fa_2_272/SUM
+ sky130_fd_sc_hd__fa_2_272/A sky130_fd_sc_hd__fa_2_272/B sky130_fd_sc_hd__fa_2_277/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_283 sky130_fd_sc_hd__fa_2_167/B sky130_fd_sc_hd__fa_2_283/SUM
+ sky130_fd_sc_hd__fa_2_283/A sky130_fd_sc_hd__fa_2_283/B sky130_fd_sc_hd__fa_2_283/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_294 sky130_fd_sc_hd__fa_2_284/A sky130_fd_sc_hd__fa_2_285/B
+ sky130_fd_sc_hd__fa_2_389/B sky130_fd_sc_hd__fa_2_294/B sky130_fd_sc_hd__fa_2_297/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor4_1_6 sky130_fd_sc_hd__nor4_1_6/D sky130_fd_sc_hd__nor4_1_6/C
+ sky130_fd_sc_hd__nor4_1_6/Y sky130_fd_sc_hd__nor4_1_6/A sky130_fd_sc_hd__nor4_1_6/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__nor4_1
Xsky130_fd_sc_hd__a22oi_1_5 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__a22oi_1_9/A1
+ sky130_fd_sc_hd__dfxtp_1_75/D sky130_fd_sc_hd__a22o_1_7/A1 sky130_fd_sc_hd__nand3_1_2/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__diode_2_100 sky130_fd_sc_hd__inv_2_135/Y VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_111 sky130_fd_sc_hd__buf_2_225/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_122 sky130_fd_sc_hd__buf_2_250/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_133 sky130_fd_sc_hd__clkbuf_1_526/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_144 sky130_fd_sc_hd__buf_2_168/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_155 sky130_fd_sc_hd__clkbuf_4_172/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_166 sky130_fd_sc_hd__clkbuf_4_182/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_177 sky130_fd_sc_hd__nand4_1_79/D VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_188 sky130_fd_sc_hd__buf_6_49/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_199 sky130_fd_sc_hd__buf_2_266/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkbuf_4_208 sky130_fd_sc_hd__clkbuf_4_208/X sky130_fd_sc_hd__clkbuf_4_208/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_219 sky130_fd_sc_hd__a22o_1_9/A1 sig_amplitude[7] VSS VDD
+ VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_12_200 sky130_fd_sc_hd__buf_4_46/X sky130_fd_sc_hd__buf_12_200/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_211 sky130_fd_sc_hd__buf_12_211/A sky130_fd_sc_hd__buf_12_211/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_222 sky130_fd_sc_hd__buf_6_28/X sky130_fd_sc_hd__buf_12_231/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_233 sky130_fd_sc_hd__buf_12_233/A sky130_fd_sc_hd__buf_12_233/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_80 sky130_fd_sc_hd__nor2_1_70/B sky130_fd_sc_hd__o21a_1_7/A1
+ sky130_fd_sc_hd__a21oi_1_80/Y sky130_fd_sc_hd__o21ai_1_88/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_244 sky130_fd_sc_hd__buf_12_244/A sky130_fd_sc_hd__buf_12_244/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_103 sky130_fd_sc_hd__clkbuf_4_72/X sky130_fd_sc_hd__clkbuf_4_73/X
+ sky130_fd_sc_hd__clkbuf_1_255/X sky130_fd_sc_hd__buf_2_93/X sky130_fd_sc_hd__buf_2_108/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a21oi_1_91 sky130_fd_sc_hd__a21oi_1_91/A1 sky130_fd_sc_hd__o22ai_1_97/Y
+ sky130_fd_sc_hd__a21oi_1_91/Y sky130_fd_sc_hd__a211o_1_8/A2 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_255 sky130_fd_sc_hd__buf_12_255/A sky130_fd_sc_hd__buf_12_255/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_114 sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__a22oi_2_12/A1
+ sky130_fd_sc_hd__buf_2_74/X sky130_fd_sc_hd__clkbuf_1_165/X sky130_fd_sc_hd__a22oi_1_114/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_266 sky130_fd_sc_hd__inv_2_95/Y sky130_fd_sc_hd__buf_12_266/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_125 sky130_fd_sc_hd__a22oi_1_97/B1 sky130_fd_sc_hd__a22oi_1_97/A1
+ sky130_fd_sc_hd__buf_2_55/X sky130_fd_sc_hd__clkbuf_4_79/X sky130_fd_sc_hd__nand4_1_26/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_277 sky130_fd_sc_hd__buf_12_277/A sky130_fd_sc_hd__buf_12_358/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_136 sky130_fd_sc_hd__a22oi_1_97/B1 sky130_fd_sc_hd__a22oi_1_97/A1
+ sky130_fd_sc_hd__clkbuf_1_156/X sky130_fd_sc_hd__clkbuf_4_76/X sky130_fd_sc_hd__nand4_1_29/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_288 sky130_fd_sc_hd__buf_8_117/X sky130_fd_sc_hd__buf_12_288/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_147 sky130_fd_sc_hd__clkbuf_1_265/X sky130_fd_sc_hd__clkbuf_1_266/X
+ sky130_fd_sc_hd__clkbuf_1_281/X sky130_fd_sc_hd__a22oi_1_147/A2 sky130_fd_sc_hd__a22oi_1_147/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_299 sky130_fd_sc_hd__buf_8_160/X sky130_fd_sc_hd__buf_12_299/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_158 sky130_fd_sc_hd__clkbuf_1_264/X sky130_fd_sc_hd__nor2_2_3/Y
+ sky130_fd_sc_hd__a22oi_1_158/B2 sky130_fd_sc_hd__clkbuf_4_135/X sky130_fd_sc_hd__nand4_1_34/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_400 sky130_fd_sc_hd__nand3_1_45/C sky130_fd_sc_hd__or4_1_2/D
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_400/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22oi_1_169 sky130_fd_sc_hd__clkbuf_4_111/X sky130_fd_sc_hd__clkbuf_4_112/X
+ sky130_fd_sc_hd__a22oi_1_169/B2 sky130_fd_sc_hd__clkbuf_1_292/X sky130_fd_sc_hd__a22oi_1_169/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_411 sky130_fd_sc_hd__nor3_1_35/A sky130_fd_sc_hd__dfxtp_1_494/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_411/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_422 sky130_fd_sc_hd__nor2_1_37/A sky130_fd_sc_hd__fa_2_961/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_422/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_433 sky130_fd_sc_hd__fa_2_967/B sky130_fd_sc_hd__nor2_1_40/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_433/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_444 sky130_fd_sc_hd__fa_2_958/B sky130_fd_sc_hd__dfxtp_1_490/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_444/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_455 sky130_fd_sc_hd__fa_2_946/B sky130_fd_sc_hd__dfxtp_1_502/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_455/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_466 sky130_fd_sc_hd__o22ai_1_76/B2 sky130_fd_sc_hd__ha_2_183/SUM
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_477 sky130_fd_sc_hd__o22ai_1_82/B2 sky130_fd_sc_hd__ha_2_177/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_477/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_488 sky130_fd_sc_hd__o21ai_1_75/B1 sky130_fd_sc_hd__nor2_1_61/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_488/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_499 sky130_fd_sc_hd__nor2_1_42/B sky130_fd_sc_hd__nand2_1_244/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_499/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_330 sky130_fd_sc_hd__nor2_1_224/Y sky130_fd_sc_hd__nor2_1_215/Y
+ sky130_fd_sc_hd__a21oi_1_330/Y sky130_fd_sc_hd__fa_2_1181/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_341 sky130_fd_sc_hd__clkinv_1_921/Y sky130_fd_sc_hd__clkinv_1_919/Y
+ sky130_fd_sc_hd__a21oi_1_341/Y sky130_fd_sc_hd__nand2_1_439/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_352 sky130_fd_sc_hd__nor3_1_39/A sky130_fd_sc_hd__o22ai_1_313/Y
+ sky130_fd_sc_hd__a21oi_1_352/Y sky130_fd_sc_hd__fa_2_1206/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_363 sky130_fd_sc_hd__o21a_1_46/B1 sky130_fd_sc_hd__o21a_1_45/A1
+ sky130_fd_sc_hd__a21oi_1_363/Y sky130_fd_sc_hd__nor2_1_229/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_374 sky130_fd_sc_hd__o21a_1_54/B1 sky130_fd_sc_hd__nor2_1_240/Y
+ sky130_fd_sc_hd__a21oi_1_374/Y sky130_fd_sc_hd__nor2_1_240/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_385 sky130_fd_sc_hd__o21ai_1_406/Y sky130_fd_sc_hd__nor2_1_258/Y
+ sky130_fd_sc_hd__a21oi_1_385/Y sky130_fd_sc_hd__nor2b_1_119/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_396 sky130_fd_sc_hd__nor2_2_17/Y sky130_fd_sc_hd__o21ai_1_412/Y
+ sky130_fd_sc_hd__nor2_1_259/B sky130_fd_sc_hd__fa_2_1239/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_0 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_992/A sky130_fd_sc_hd__nor2_2_7/Y
+ sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__xor2_1_60/A sky130_fd_sc_hd__nor2_2_7/A
+ sky130_fd_sc_hd__a222oi_1_0/Y sky130_fd_sc_hd__fa_2_991/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xor2_1_207 sky130_fd_sc_hd__xor2_1_207/B sky130_fd_sc_hd__xor2_1_207/X
+ sky130_fd_sc_hd__xor2_1_208/X VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_390 sky130_fd_sc_hd__o21a_1_29/A1 sky130_fd_sc_hd__nor2_2_15/B
+ sky130_fd_sc_hd__nor2_2_15/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_218 sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__fa_2_1200/B
+ sky130_fd_sc_hd__xor2_1_218/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_229 sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__xor2_1_229/X
+ sky130_fd_sc_hd__nor2_8_0/B VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_2_12 VDD VSS sky130_fd_sc_hd__buf_2_12/X sky130_fd_sc_hd__ha_2_14/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_23 VDD VSS sky130_fd_sc_hd__buf_2_23/X sky130_fd_sc_hd__buf_2_23/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_34 VDD VSS sky130_fd_sc_hd__buf_4_33/A sky130_fd_sc_hd__buf_8_63/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_45 VDD VSS sky130_fd_sc_hd__buf_2_45/X sky130_fd_sc_hd__ha_2_38/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_56 VDD VSS sky130_fd_sc_hd__buf_2_56/X sky130_fd_sc_hd__buf_2_56/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_67 VDD VSS sky130_fd_sc_hd__buf_2_67/X sky130_fd_sc_hd__buf_2_67/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_78 VDD VSS sky130_fd_sc_hd__buf_2_78/X sky130_fd_sc_hd__buf_2_78/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_89 VDD VSS sky130_fd_sc_hd__buf_2_89/X sky130_fd_sc_hd__buf_2_89/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o211ai_1_50 sky130_fd_sc_hd__nor2_1_260/B sky130_fd_sc_hd__nor2_1_265/A
+ sky130_fd_sc_hd__xor2_1_263/A sky130_fd_sc_hd__nand2_1_481/Y sky130_fd_sc_hd__a21oi_1_385/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_61 sky130_fd_sc_hd__nor2_1_307/A sky130_fd_sc_hd__nor2_1_301/B
+ sky130_fd_sc_hd__xor2_1_307/A sky130_fd_sc_hd__nand2_1_531/Y sky130_fd_sc_hd__nand2_1_532/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__diode_2_7 sky130_fd_sc_hd__clkbuf_1_247/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__and2_0_209 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_209/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_209/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_230 sky130_fd_sc_hd__inv_2_122/A sky130_fd_sc_hd__a22o_2_9/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_230/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_241 sky130_fd_sc_hd__clkinv_1_242/A sky130_fd_sc_hd__inv_2_108/Y
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_252 sky130_fd_sc_hd__inv_2_128/A sky130_fd_sc_hd__buf_2_246/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_252/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_263 sky130_fd_sc_hd__nor2_1_12/B sky130_fd_sc_hd__ha_2_153/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_263/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_274 sky130_fd_sc_hd__o21ai_1_28/A1 sky130_fd_sc_hd__ha_2_157/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_274/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o31ai_1_7 sky130_fd_sc_hd__o31ai_1_7/Y sky130_fd_sc_hd__o31ai_1_7/A2
+ sky130_fd_sc_hd__o31ai_1_8/A2 sky130_fd_sc_hd__o31ai_1_8/A3 sky130_fd_sc_hd__o31ai_1_7/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__o31ai_1
Xsky130_fd_sc_hd__a22o_2_8 sky130_fd_sc_hd__or2_1_1/B sky130_fd_sc_hd__ha_2_84/A sky130_fd_sc_hd__a22o_2_8/X
+ sky130_fd_sc_hd__a22o_2_8/B2 sky130_fd_sc_hd__a22o_4_0/B1 VDD VSS VDD VSS sky130_fd_sc_hd__a22o_2
Xsky130_fd_sc_hd__clkinv_1_285 sky130_fd_sc_hd__fa_2_49/B sky130_fd_sc_hd__ha_2_95/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_285/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_296 sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__fa_2_15/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_296/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_4 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__a21oi_1_4/B1
+ sky130_fd_sc_hd__a21oi_1_4/Y sky130_fd_sc_hd__o21ai_1_7/A2 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkbuf_4_17 sky130_fd_sc_hd__clkbuf_4_17/X sky130_fd_sc_hd__clkbuf_4_17/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_28 sky130_fd_sc_hd__clkbuf_4_28/X sky130_fd_sc_hd__clkbuf_4_28/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_39 sky130_fd_sc_hd__clkbuf_4_39/X sky130_fd_sc_hd__clkbuf_4_39/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__a21oi_1_160 sky130_fd_sc_hd__nor2_2_11/Y sky130_fd_sc_hd__o22ai_1_159/Y
+ sky130_fd_sc_hd__a21oi_1_160/Y sky130_fd_sc_hd__fa_2_1117/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_171 sky130_fd_sc_hd__clkinv_1_663/Y sky130_fd_sc_hd__nor2_1_93/B
+ sky130_fd_sc_hd__xnor2_1_69/A sky130_fd_sc_hd__xnor2_1_67/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_182 sky130_fd_sc_hd__o21a_1_12/B1 sky130_fd_sc_hd__o21a_1_11/A1
+ sky130_fd_sc_hd__dfxtp_1_762/D sky130_fd_sc_hd__nor2_1_115/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_193 sky130_fd_sc_hd__nand2_1_331/B sky130_fd_sc_hd__o21ai_1_218/Y
+ sky130_fd_sc_hd__a21oi_1_193/Y sky130_fd_sc_hd__nand2_1_318/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_101 sky130_fd_sc_hd__inv_2_61/Y sky130_fd_sc_hd__buf_8_101/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_112 sky130_fd_sc_hd__buf_8_70/A sky130_fd_sc_hd__buf_4_51/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_123 sky130_fd_sc_hd__buf_8_123/A sky130_fd_sc_hd__buf_8_123/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_134 sky130_fd_sc_hd__and2_2_1/X sky130_fd_sc_hd__buf_8_170/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_145 sky130_fd_sc_hd__inv_2_94/Y sky130_fd_sc_hd__buf_8_145/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_156 sky130_fd_sc_hd__inv_2_92/Y sky130_fd_sc_hd__buf_8_156/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nor2_4_7 sky130_fd_sc_hd__nor2_4_7/Y sky130_fd_sc_hd__nor3_2_8/C
+ sky130_fd_sc_hd__nor2_4_8/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__buf_8_167 sky130_fd_sc_hd__buf_8_167/A sky130_fd_sc_hd__buf_6_36/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_178 sky130_fd_sc_hd__buf_8_178/A sky130_fd_sc_hd__buf_8_178/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_189 sky130_fd_sc_hd__inv_2_121/Y sky130_fd_sc_hd__buf_8_189/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__a21o_2_13 sky130_fd_sc_hd__a21o_2_13/X sky130_fd_sc_hd__nor2_1_209/Y
+ sky130_fd_sc_hd__nor2_1_209/A sky130_fd_sc_hd__nor2_1_209/B VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__a21o_2_24 sky130_fd_sc_hd__a21o_2_24/X sky130_fd_sc_hd__nor2_1_293/Y
+ sky130_fd_sc_hd__fa_2_3/SUM sky130_fd_sc_hd__nor2_1_293/B VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__xor2_1_40 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_987/B
+ sky130_fd_sc_hd__xor2_1_40/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_51 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_976/B
+ sky130_fd_sc_hd__xor2_1_51/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_62 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__xor2_1_62/X
+ sky130_fd_sc_hd__xor2_1_62/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_18 sky130_fd_sc_hd__inv_2_40/Y sky130_fd_sc_hd__buf_12_18/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_73 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__xor2_1_73/X
+ sky130_fd_sc_hd__xor2_1_73/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_29 sky130_fd_sc_hd__buf_8_9/X sky130_fd_sc_hd__buf_12_29/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_84 sky130_fd_sc_hd__xor2_1_84/B sky130_fd_sc_hd__xor2_1_84/X
+ sky130_fd_sc_hd__xor2_1_85/X VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_95 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__xor2_1_95/X
+ sky130_fd_sc_hd__xor2_1_95/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2b_1_1 sky130_fd_sc_hd__nand2b_1_1/Y sky130_fd_sc_hd__nand3_2_2/A
+ sky130_fd_sc_hd__inv_8_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__dfxtp_1_1306 VDD VSS sky130_fd_sc_hd__fa_2_845/B sky130_fd_sc_hd__dfxtp_1_1322/CLK
+ sky130_fd_sc_hd__a21oi_1_433/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1317 VDD VSS sky130_fd_sc_hd__fa_2_902/B sky130_fd_sc_hd__dfxtp_1_1329/CLK
+ sky130_fd_sc_hd__o32ai_1_9/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1328 VDD VSS sky130_fd_sc_hd__fa_2_912/A sky130_fd_sc_hd__dfxtp_1_1332/CLK
+ sky130_fd_sc_hd__a21oi_1_422/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_900 VDD VSS sky130_fd_sc_hd__fa_2_935/B sky130_fd_sc_hd__dfxtp_1_904/CLK
+ sky130_fd_sc_hd__o21a_1_21/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1339 VDD VSS sky130_fd_sc_hd__fa_2_1298/A sky130_fd_sc_hd__clkinv_8_70/Y
+ sky130_fd_sc_hd__mux2_2_251/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_911 VDD VSS sky130_fd_sc_hd__fa_2_1140/B sky130_fd_sc_hd__clkinv_8_55/Y
+ sky130_fd_sc_hd__and2_0_320/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_922 VDD VSS sky130_fd_sc_hd__fa_2_1151/A sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__mux2_2_90/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_933 VDD VSS sky130_fd_sc_hd__fa_2_1125/A sky130_fd_sc_hd__clkinv_8_55/Y
+ sky130_fd_sc_hd__mux2_2_114/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_944 VDD VSS sky130_fd_sc_hd__fa_2_1136/A sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__mux2_2_85/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_955 VDD VSS sky130_fd_sc_hd__fa_2_1164/A sky130_fd_sc_hd__clkinv_8_64/Y
+ sky130_fd_sc_hd__mux2_2_115/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_966 VDD VSS sky130_fd_sc_hd__o32ai_1_2/A1 sky130_fd_sc_hd__clkinv_8_46/Y
+ sky130_fd_sc_hd__nor2b_1_109/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_977 VDD VSS sky130_fd_sc_hd__mux2_2_99/A0 sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__o22ai_1_218/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_988 VDD VSS sky130_fd_sc_hd__mux2_2_123/A0 sky130_fd_sc_hd__clkinv_8_64/Y
+ sky130_fd_sc_hd__dfxtp_1_988/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_999 VDD VSS sky130_fd_sc_hd__mux2_2_100/A0 sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__dfxtp_1_999/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_520 VSS VDD sky130_fd_sc_hd__buf_2_233/A sky130_fd_sc_hd__clkbuf_1_533/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_531 VSS VDD sky130_fd_sc_hd__buf_2_172/A sky130_fd_sc_hd__clkbuf_1_531/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_542 VSS VDD sky130_fd_sc_hd__ha_2_95/B sky130_fd_sc_hd__ha_2_104/B
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_110 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_110/A sky130_fd_sc_hd__fa_2_342/CIN
+ sky130_fd_sc_hd__fa_2_338/B sky130_fd_sc_hd__ha_2_110/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_553 VSS VDD sky130_fd_sc_hd__and2_0_235/B sky130_fd_sc_hd__inv_4_1/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_121 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_169/B sky130_fd_sc_hd__fa_2_503/A
+ sky130_fd_sc_hd__ha_2_121/SUM sky130_fd_sc_hd__ha_2_121/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_564 VSS VDD sky130_fd_sc_hd__nand2_1_113/B sky130_fd_sc_hd__nand4_1_48/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_132 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_132/A sky130_fd_sc_hd__fa_2_605/A
+ sky130_fd_sc_hd__fa_2_602/B sky130_fd_sc_hd__ha_2_132/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_575 VSS VDD sky130_fd_sc_hd__nand3_1_15/C sky130_fd_sc_hd__a22oi_1_27/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_143 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_143/A sky130_fd_sc_hd__fa_2_822/B
+ sky130_fd_sc_hd__fa_2_819/A sky130_fd_sc_hd__ha_2_143/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_586 VSS VDD sky130_fd_sc_hd__nand3_1_6/B sky130_fd_sc_hd__a22oi_1_12/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_154 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_154/A sky130_fd_sc_hd__ha_2_153/B
+ sky130_fd_sc_hd__ha_2_154/SUM sky130_fd_sc_hd__ha_2_154/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_597 VSS VDD sky130_fd_sc_hd__clkbuf_1_598/A sig_frequency[4]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_805 sky130_fd_sc_hd__fa_2_804/B sky130_fd_sc_hd__fa_2_805/SUM
+ sky130_fd_sc_hd__fa_2_805/A sky130_fd_sc_hd__fa_2_805/B sky130_fd_sc_hd__fa_2_805/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_165 VSS VDD VSS VDD sky130_fd_sc_hd__nor4_1_2/B sky130_fd_sc_hd__ha_2_164/B
+ sky130_fd_sc_hd__ha_2_165/SUM sky130_fd_sc_hd__ha_2_165/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_816 sky130_fd_sc_hd__fa_2_815/A sky130_fd_sc_hd__fa_2_810/A
+ sky130_fd_sc_hd__fa_2_834/B sky130_fd_sc_hd__fa_2_829/A sky130_fd_sc_hd__ha_2_139/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_176 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_176/A sky130_fd_sc_hd__ha_2_175/A
+ sky130_fd_sc_hd__ha_2_176/SUM sky130_fd_sc_hd__ha_2_176/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_827 sky130_fd_sc_hd__fa_2_825/A sky130_fd_sc_hd__fa_2_821/A
+ sky130_fd_sc_hd__fa_2_833/A sky130_fd_sc_hd__ha_2_143/B sky130_fd_sc_hd__fa_2_793/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_187 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_187/A sky130_fd_sc_hd__ha_2_186/A
+ sky130_fd_sc_hd__ha_2_187/SUM sky130_fd_sc_hd__ha_2_187/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_838 sky130_fd_sc_hd__fa_2_837/CIN sky130_fd_sc_hd__fa_2_838/SUM
+ sky130_fd_sc_hd__fa_2_838/A sky130_fd_sc_hd__fa_2_838/B sky130_fd_sc_hd__fa_2_838/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_198 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_198/A sky130_fd_sc_hd__ha_2_197/A
+ sky130_fd_sc_hd__ha_2_198/SUM sky130_fd_sc_hd__ha_2_198/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_849 sky130_fd_sc_hd__fa_2_848/CIN sky130_fd_sc_hd__fa_2_849/SUM
+ sky130_fd_sc_hd__fa_2_849/A sky130_fd_sc_hd__fa_2_849/B sky130_fd_sc_hd__fa_2_849/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__maj3_1_3 sky130_fd_sc_hd__maj3_1_3/C sky130_fd_sc_hd__maj3_1_3/X
+ sky130_fd_sc_hd__maj3_1_3/B sky130_fd_sc_hd__maj3_1_3/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__mux2_2_105 VSS VDD sky130_fd_sc_hd__mux2_2_105/A1 sky130_fd_sc_hd__mux2_2_105/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_105/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_116 VSS VDD sky130_fd_sc_hd__mux2_2_116/A1 sky130_fd_sc_hd__mux2_2_116/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_116/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_127 VSS VDD sky130_fd_sc_hd__mux2_2_127/A1 sky130_fd_sc_hd__mux2_2_127/A0
+ sky130_fd_sc_hd__mux2_2_135/S sky130_fd_sc_hd__mux2_2_127/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_138 VSS VDD sky130_fd_sc_hd__mux2_2_138/A1 sky130_fd_sc_hd__mux2_2_138/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_138/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_149 VSS VDD sky130_fd_sc_hd__mux2_2_149/A1 sky130_fd_sc_hd__mux2_2_149/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_149/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__and2_0_12 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_12/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_7/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_23 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_23/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_11/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_303 sky130_fd_sc_hd__o22ai_1_322/A2 sky130_fd_sc_hd__o22ai_1_304/A1
+ sky130_fd_sc_hd__o22ai_1_303/Y sky130_fd_sc_hd__nor2_1_188/B sky130_fd_sc_hd__o32ai_1_5/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_34 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_34/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__and2_0_34/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_314 sky130_fd_sc_hd__o22ai_1_322/A2 sky130_fd_sc_hd__o22ai_1_322/B1
+ sky130_fd_sc_hd__o22ai_1_314/Y sky130_fd_sc_hd__o21a_1_42/A2 sky130_fd_sc_hd__o22ai_1_318/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_45 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_54/A sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__ha_2_51/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__maj3_1_109 sky130_fd_sc_hd__maj3_1_110/X sky130_fd_sc_hd__maj3_1_109/X
+ sky130_fd_sc_hd__maj3_1_109/B sky130_fd_sc_hd__maj3_1_109/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__o22ai_1_325 sky130_fd_sc_hd__nand2_1_462/Y sky130_fd_sc_hd__nand2_1_461/Y
+ sky130_fd_sc_hd__o22ai_1_325/Y sky130_fd_sc_hd__o22ai_1_338/A1 sky130_fd_sc_hd__a21o_2_18/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_56 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_56/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_56/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_336 sky130_fd_sc_hd__nand2_1_462/Y sky130_fd_sc_hd__nand2_1_461/Y
+ sky130_fd_sc_hd__o22ai_1_336/Y sky130_fd_sc_hd__o22ai_1_349/A1 sky130_fd_sc_hd__o21ai_1_391/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_67 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_78/A sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__ha_2_73/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_347 sky130_fd_sc_hd__nand2_1_464/Y sky130_fd_sc_hd__nand2_1_463/Y
+ sky130_fd_sc_hd__o22ai_1_347/Y sky130_fd_sc_hd__nand2_1_476/B sky130_fd_sc_hd__o21ai_1_390/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_78 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_78/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__and2_0_78/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_358 sky130_fd_sc_hd__nor2_1_268/A sky130_fd_sc_hd__nor2_1_257/A
+ sky130_fd_sc_hd__o22ai_1_358/Y sky130_fd_sc_hd__o22ai_1_358/A1 sky130_fd_sc_hd__nor2_1_260/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_2_4 sky130_fd_sc_hd__nor2_2_5/B sky130_fd_sc_hd__nor2_2_4/Y
+ sky130_fd_sc_hd__nor2_2_4/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__and2_0_89 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_89/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_89/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_369 sky130_fd_sc_hd__nor2_1_268/A sky130_fd_sc_hd__nor2_1_257/A
+ sky130_fd_sc_hd__o22ai_1_369/Y sky130_fd_sc_hd__a21oi_1_410/Y sky130_fd_sc_hd__nor2_1_268/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__buf_8_11 sky130_fd_sc_hd__ha_2_12/A sky130_fd_sc_hd__buf_8_11/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_22 sky130_fd_sc_hd__inv_2_24/Y sky130_fd_sc_hd__buf_8_22/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_33 sky130_fd_sc_hd__buf_8_33/A sky130_fd_sc_hd__buf_8_33/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_44 sky130_fd_sc_hd__buf_8_44/A sky130_fd_sc_hd__buf_8_44/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_55 sky130_fd_sc_hd__inv_2_15/Y sky130_fd_sc_hd__buf_8_55/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_66 sky130_fd_sc_hd__buf_8_66/A sky130_fd_sc_hd__buf_8_66/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_77 sky130_fd_sc_hd__buf_8_77/A sky130_fd_sc_hd__buf_8_77/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_88 sky130_fd_sc_hd__buf_8_88/A sky130_fd_sc_hd__buf_8_88/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_207 VDD VSS sky130_fd_sc_hd__ha_2_74/A sky130_fd_sc_hd__dfxtp_1_207/CLK
+ sky130_fd_sc_hd__and2_0_73/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_8_99 sky130_fd_sc_hd__ha_2_39/A sky130_fd_sc_hd__buf_8_99/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_218 VDD VSS sky130_fd_sc_hd__ha_2_85/A sky130_fd_sc_hd__dfxtp_1_224/CLK
+ sky130_fd_sc_hd__nor2b_1_48/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_229 VDD VSS sky130_fd_sc_hd__nor3_2_10/B sky130_fd_sc_hd__clkinv_8_102/Y
+ sky130_fd_sc_hd__a22o_1_28/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_2_107 VDD VSS sky130_fd_sc_hd__buf_2_107/X sky130_fd_sc_hd__buf_2_107/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__fa_2_1306 sky130_fd_sc_hd__fa_2_1307/CIN sky130_fd_sc_hd__mux2_2_230/A0
+ sky130_fd_sc_hd__fa_2_1306/A sky130_fd_sc_hd__fa_2_1306/B sky130_fd_sc_hd__fa_2_1306/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_118 VDD VSS sky130_fd_sc_hd__buf_4_36/A sky130_fd_sc_hd__buf_2_118/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__fa_2_1317 sky130_fd_sc_hd__fa_2_1318/CIN sky130_fd_sc_hd__mux2_2_259/A1
+ sky130_fd_sc_hd__fa_2_1317/A sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1317/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_129 VDD VSS sky130_fd_sc_hd__buf_8_155/A sky130_fd_sc_hd__and2_1_3/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1103 VDD VSS sky130_fd_sc_hd__fa_2_1222/A sky130_fd_sc_hd__clkinv_8_78/Y
+ sky130_fd_sc_hd__nand2_1_413/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1114 VDD VSS sky130_fd_sc_hd__mux2_2_159/A0 sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__o22ai_1_279/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1125 VDD VSS sky130_fd_sc_hd__mux2_2_131/A1 sky130_fd_sc_hd__clkinv_8_70/Y
+ sky130_fd_sc_hd__o22ai_1_268/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1136 VDD VSS sky130_fd_sc_hd__mux2_2_160/A0 sky130_fd_sc_hd__clkinv_8_64/Y
+ sky130_fd_sc_hd__dfxtp_1_995/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1147 VDD VSS sky130_fd_sc_hd__mux2_2_152/A0 sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__o22ai_1_290/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1158 VDD VSS sky130_fd_sc_hd__mux2_2_126/A1 sky130_fd_sc_hd__clkinv_8_70/Y
+ sky130_fd_sc_hd__o31ai_1_7/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_730 VDD VSS sky130_fd_sc_hd__mux2_2_12/A1 sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__o21ai_1_67/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1169 VDD VSS sky130_fd_sc_hd__fa_2_855/B sky130_fd_sc_hd__dfxtp_1_1184/CLK
+ sky130_fd_sc_hd__a21oi_1_371/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_741 VDD VSS sky130_fd_sc_hd__and2_0_164/A sky130_fd_sc_hd__dfxtp_1_744/CLK
+ sky130_fd_sc_hd__fa_2_1096/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_752 VDD VSS sky130_fd_sc_hd__and2_0_184/A sky130_fd_sc_hd__dfxtp_1_768/CLK
+ sky130_fd_sc_hd__xor2_1_139/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_763 VDD VSS sky130_fd_sc_hd__ha_2_134/B sky130_fd_sc_hd__dfxtp_1_768/CLK
+ sky130_fd_sc_hd__o21a_1_11/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_774 VDD VSS sky130_fd_sc_hd__fa_2_1073/A sky130_fd_sc_hd__clkinv_8_54/Y
+ sky130_fd_sc_hd__and2_0_312/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__ha_2_7 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_7/A sky130_fd_sc_hd__ha_2_6/B
+ sky130_fd_sc_hd__ha_2_7/SUM sky130_fd_sc_hd__ha_2_7/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__dfxtp_1_785 VDD VSS sky130_fd_sc_hd__fa_2_1084/A sky130_fd_sc_hd__clkinv_8_56/Y
+ sky130_fd_sc_hd__mux2_2_54/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_796 VDD VSS sky130_fd_sc_hd__fa_2_1048/A sky130_fd_sc_hd__clkinv_8_54/Y
+ sky130_fd_sc_hd__and2_0_307/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_350 VSS VDD sky130_fd_sc_hd__buf_8_164/A sky130_fd_sc_hd__clkbuf_1_363/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_361 VSS VDD sky130_fd_sc_hd__buf_8_139/A sky130_fd_sc_hd__clkbuf_1_361/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_372 VSS VDD sky130_fd_sc_hd__buf_4_91/A sky130_fd_sc_hd__buf_4_90/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_383 VSS VDD sky130_fd_sc_hd__clkbuf_1_383/X sky130_fd_sc_hd__clkbuf_1_383/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_602 sky130_fd_sc_hd__fa_2_604/B sky130_fd_sc_hd__fa_2_602/SUM
+ sky130_fd_sc_hd__fa_2_602/A sky130_fd_sc_hd__fa_2_602/B sky130_fd_sc_hd__fa_2_602/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_394 VSS VDD sky130_fd_sc_hd__a22oi_2_17/B2 sky130_fd_sc_hd__clkbuf_1_394/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_613 sky130_fd_sc_hd__fa_2_615/A sky130_fd_sc_hd__fa_2_610/A
+ sky130_fd_sc_hd__fa_2_692/A sky130_fd_sc_hd__ha_2_132/A sky130_fd_sc_hd__fa_2_683/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_18 VSS VDD sky130_fd_sc_hd__a22oi_2_9/B1 sky130_fd_sc_hd__nor3_2_3/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_624 sky130_fd_sc_hd__fa_2_625/CIN sky130_fd_sc_hd__fa_2_619/A
+ sky130_fd_sc_hd__fa_2_700/B sky130_fd_sc_hd__fa_2_624/B sky130_fd_sc_hd__ha_2_129/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_29 VSS VDD sky130_fd_sc_hd__clkbuf_1_29/X sky130_fd_sc_hd__clkbuf_1_29/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_635 sky130_fd_sc_hd__fa_2_634/B sky130_fd_sc_hd__fa_2_635/SUM
+ sky130_fd_sc_hd__ha_2_132/B sky130_fd_sc_hd__ha_2_130/B sky130_fd_sc_hd__fa_2_700/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_646 sky130_fd_sc_hd__fa_2_649/B sky130_fd_sc_hd__fa_2_646/SUM
+ sky130_fd_sc_hd__fa_2_646/A sky130_fd_sc_hd__fa_2_646/B sky130_fd_sc_hd__fa_2_651/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_657 sky130_fd_sc_hd__fa_2_660/B sky130_fd_sc_hd__fa_2_657/SUM
+ sky130_fd_sc_hd__fa_2_657/A sky130_fd_sc_hd__fa_2_657/B sky130_fd_sc_hd__o22ai_1_46/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_668 sky130_fd_sc_hd__fa_2_669/B sky130_fd_sc_hd__fa_2_662/A
+ sky130_fd_sc_hd__ha_2_135/B sky130_fd_sc_hd__fa_2_678/B sky130_fd_sc_hd__fa_2_699/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_679 sky130_fd_sc_hd__fa_2_681/CIN sky130_fd_sc_hd__fa_2_670/A
+ sky130_fd_sc_hd__ha_2_130/B sky130_fd_sc_hd__fa_2_679/B sky130_fd_sc_hd__fa_2_679/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__conb_1_1 sky130_fd_sc_hd__conb_1_1/LO sky130_fd_sc_hd__conb_1_1/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__buf_12_7 sky130_fd_sc_hd__inv_2_11/Y sky130_fd_sc_hd__buf_12_7/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__o22ai_1_100 sky130_fd_sc_hd__o22ai_1_130/B1 sky130_fd_sc_hd__nor2_1_68/B
+ sky130_fd_sc_hd__o22ai_1_100/Y sky130_fd_sc_hd__o22ai_1_120/B1 sky130_fd_sc_hd__o21ai_1_92/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_111 sky130_fd_sc_hd__o22ai_1_130/B1 sky130_fd_sc_hd__o22ai_1_116/A1
+ sky130_fd_sc_hd__nor2_1_82/A sky130_fd_sc_hd__nor2_1_66/B sky130_fd_sc_hd__o22ai_1_132/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_122 sky130_fd_sc_hd__o22ai_1_92/A1 sky130_fd_sc_hd__o22ai_1_122/B1
+ sky130_fd_sc_hd__o22ai_1_122/Y sky130_fd_sc_hd__nor2_1_76/A sky130_fd_sc_hd__nor2_2_9/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_133 sky130_fd_sc_hd__nor2_2_9/B sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__o22ai_1_133/Y sky130_fd_sc_hd__a21oi_1_127/Y sky130_fd_sc_hd__a21boi_0_1/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_144 sky130_fd_sc_hd__nand2_1_284/Y sky130_fd_sc_hd__nand2_2_5/Y
+ sky130_fd_sc_hd__o22ai_1_144/Y sky130_fd_sc_hd__xnor2_1_80/Y sky130_fd_sc_hd__o22ai_1_158/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_208 sky130_fd_sc_hd__nor3_1_31/C sky130_fd_sc_hd__nor2_1_28/Y
+ sky130_fd_sc_hd__or4_1_2/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_155 sky130_fd_sc_hd__nand2_1_338/A sky130_fd_sc_hd__nand2_1_284/Y
+ sky130_fd_sc_hd__o22ai_1_155/Y sky130_fd_sc_hd__xnor2_1_74/Y sky130_fd_sc_hd__o22ai_1_155/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_807 sky130_fd_sc_hd__o32ai_1_1/B2 sky130_fd_sc_hd__fa_2_1142/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_807/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_2_11 sky130_fd_sc_hd__nor2_2_11/B sky130_fd_sc_hd__nor2_2_11/Y
+ sky130_fd_sc_hd__nor2_2_11/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__nand2_1_219 sky130_fd_sc_hd__o21ai_1_35/B1 sky130_fd_sc_hd__o22a_1_0/B2
+ sky130_fd_sc_hd__xor2_1_31/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_818 sky130_fd_sc_hd__clkinv_1_818/Y sky130_fd_sc_hd__nand2_1_376/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_818/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_166 sky130_fd_sc_hd__nor2_2_13/B sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__o22ai_1_166/Y sky130_fd_sc_hd__a21oi_1_220/Y sky130_fd_sc_hd__a21oi_1_190/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_177 sky130_fd_sc_hd__o22ai_1_204/B1 sky130_fd_sc_hd__o22ai_1_191/A1
+ sky130_fd_sc_hd__nor2_1_129/A sky130_fd_sc_hd__nor2_1_117/B sky130_fd_sc_hd__o22ai_1_206/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_829 sky130_fd_sc_hd__nor2_1_146/B sky130_fd_sc_hd__fa_2_1129/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_829/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_188 sky130_fd_sc_hd__o21a_1_16/A2 sky130_fd_sc_hd__nor2_1_119/B
+ sky130_fd_sc_hd__nor2_1_133/B sky130_fd_sc_hd__o22ai_1_194/B1 sky130_fd_sc_hd__o22ai_1_206/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand4_1_14 sky130_fd_sc_hd__nand4_1_14/C sky130_fd_sc_hd__nand4_1_14/B
+ sky130_fd_sc_hd__nand4_1_14/Y sky130_fd_sc_hd__nand4_1_14/D sky130_fd_sc_hd__nand4_1_14/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__o211ai_1_1 sky130_fd_sc_hd__nand4_1_81/Y sky130_fd_sc_hd__nand4_1_80/Y
+ sky130_fd_sc_hd__o211ai_1_1/Y sky130_fd_sc_hd__o21ai_1_3/B1 sky130_fd_sc_hd__o211ai_1_1/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__nand4_1_25 sky130_fd_sc_hd__nand4_1_25/C sky130_fd_sc_hd__nand4_1_25/B
+ sky130_fd_sc_hd__nand4_1_25/Y sky130_fd_sc_hd__nand4_1_25/D sky130_fd_sc_hd__nand4_1_25/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__o22ai_1_199 sky130_fd_sc_hd__nor2_2_13/B sky130_fd_sc_hd__nor2_1_127/A
+ sky130_fd_sc_hd__o22ai_1_199/Y sky130_fd_sc_hd__o21a_1_16/X sky130_fd_sc_hd__a21oi_1_238/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand4_1_36 sky130_fd_sc_hd__nand4_1_36/C sky130_fd_sc_hd__nand4_1_36/B
+ sky130_fd_sc_hd__nand4_1_36/Y sky130_fd_sc_hd__nand4_1_36/D sky130_fd_sc_hd__nand4_1_36/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_47 sky130_fd_sc_hd__nand4_1_47/C sky130_fd_sc_hd__nand4_1_47/B
+ sky130_fd_sc_hd__nand4_1_47/Y sky130_fd_sc_hd__nand4_1_47/D sky130_fd_sc_hd__nand4_1_47/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_58 sky130_fd_sc_hd__nand4_1_58/C sky130_fd_sc_hd__nand4_1_58/B
+ sky130_fd_sc_hd__nand4_1_58/Y sky130_fd_sc_hd__nand4_1_58/D sky130_fd_sc_hd__nand4_1_58/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_69 sky130_fd_sc_hd__nand4_1_69/C sky130_fd_sc_hd__nand4_1_69/B
+ sky130_fd_sc_hd__nand4_1_69/Y sky130_fd_sc_hd__nand4_1_69/D sky130_fd_sc_hd__nand4_1_69/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__conb_1_18 sky130_fd_sc_hd__conb_1_18/LO sky130_fd_sc_hd__conb_1_18/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_29 sky130_fd_sc_hd__conb_1_29/LO sky130_fd_sc_hd__conb_1_29/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__a211oi_1_10 sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__nor2_1_138/Y
+ sky130_fd_sc_hd__o22ai_1_206/Y sky130_fd_sc_hd__a211oi_1_10/Y sky130_fd_sc_hd__fa_2_1084/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_360 VSS VDD sky130_fd_sc_hd__nor2_1_214/A sky130_fd_sc_hd__o21ai_1_360/A1
+ sky130_fd_sc_hd__a211oi_1_20/Y sky130_fd_sc_hd__xor2_1_226/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a211oi_1_21 sky130_fd_sc_hd__nor2_2_16/Y sky130_fd_sc_hd__nor2_1_218/Y
+ sky130_fd_sc_hd__o22ai_1_307/Y sky130_fd_sc_hd__nor2_1_217/B sky130_fd_sc_hd__fa_2_1187/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_371 VSS VDD sky130_fd_sc_hd__o22ai_1_319/A1 sky130_fd_sc_hd__nor2_1_195/B
+ sky130_fd_sc_hd__o21ai_1_371/B1 sky130_fd_sc_hd__o21ai_1_371/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a211oi_1_32 sky130_fd_sc_hd__nor2_1_309/Y sky130_fd_sc_hd__nor2_1_299/Y
+ sky130_fd_sc_hd__nor2_1_300/Y sky130_fd_sc_hd__a211oi_1_32/Y sky130_fd_sc_hd__fa_2_1284/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_382 VSS VDD sky130_fd_sc_hd__o22ai_1_318/A2 sky130_fd_sc_hd__o21ai_1_382/A1
+ sky130_fd_sc_hd__a21oi_1_357/Y sky130_fd_sc_hd__o21ai_1_382/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_393 VSS VDD sky130_fd_sc_hd__nor2_1_241/B sky130_fd_sc_hd__o22ai_1_379/A2
+ sky130_fd_sc_hd__a22oi_1_387/Y sky130_fd_sc_hd__o21ai_1_393/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__mux2_2_40 VSS VDD sky130_fd_sc_hd__mux2_2_40/A1 sky130_fd_sc_hd__xor2_1_86/X
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_40/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_51 VSS VDD sky130_fd_sc_hd__mux2_2_51/A1 sky130_fd_sc_hd__mux2_2_51/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_51/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_62 VSS VDD sky130_fd_sc_hd__mux2_2_62/A1 sky130_fd_sc_hd__mux2_2_62/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_62/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_73 VSS VDD sky130_fd_sc_hd__mux2_2_73/A1 sky130_fd_sc_hd__mux2_2_73/A0
+ sky130_fd_sc_hd__mux2_2_75/S sky130_fd_sc_hd__mux2_2_73/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_84 VSS VDD sky130_fd_sc_hd__mux2_2_84/A1 sky130_fd_sc_hd__mux2_2_84/A0
+ sky130_fd_sc_hd__nor2_4_15/A sky130_fd_sc_hd__mux2_2_84/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1103 sky130_fd_sc_hd__fa_2_1104/CIN sky130_fd_sc_hd__and2_0_316/A
+ sky130_fd_sc_hd__fa_2_1103/A sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1103/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__mux2_2_95 VSS VDD sky130_fd_sc_hd__mux2_2_95/A1 sky130_fd_sc_hd__mux2_2_95/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_95/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1114 sky130_fd_sc_hd__fa_2_1115/CIN sky130_fd_sc_hd__fa_2_1114/SUM
+ sky130_fd_sc_hd__fa_2_1114/A sky130_fd_sc_hd__fa_2_1114/B sky130_fd_sc_hd__fa_2_1114/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1125 sky130_fd_sc_hd__fa_2_1126/CIN sky130_fd_sc_hd__mux2_2_114/A1
+ sky130_fd_sc_hd__fa_2_1125/A sky130_fd_sc_hd__fa_2_1125/B sky130_fd_sc_hd__fa_2_1125/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1136 sky130_fd_sc_hd__fa_2_1137/CIN sky130_fd_sc_hd__mux2_2_85/A0
+ sky130_fd_sc_hd__fa_2_1136/A sky130_fd_sc_hd__fa_2_1136/B sky130_fd_sc_hd__fa_2_1136/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1147 sky130_fd_sc_hd__fa_2_1148/CIN sky130_fd_sc_hd__mux2_2_101/A1
+ sky130_fd_sc_hd__fa_2_1147/A sky130_fd_sc_hd__fa_2_1147/B sky130_fd_sc_hd__fa_2_1147/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1158 sky130_fd_sc_hd__fa_2_1159/CIN sky130_fd_sc_hd__mux2_2_123/A1
+ sky130_fd_sc_hd__fa_2_1172/B sky130_fd_sc_hd__fa_2_1158/B sky130_fd_sc_hd__fa_2_1172/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1169 sky130_fd_sc_hd__fa_2_1170/CIN sky130_fd_sc_hd__mux2_2_100/A1
+ sky130_fd_sc_hd__fa_2_1169/A sky130_fd_sc_hd__fa_2_1172/B sky130_fd_sc_hd__fa_2_1169/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_560 VDD VSS sky130_fd_sc_hd__dfxtp_1_560/Q sky130_fd_sc_hd__dfxtp_1_576/CLK
+ sky130_fd_sc_hd__dfxtp_1_560/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_571 VDD VSS sky130_fd_sc_hd__and2_0_203/A sky130_fd_sc_hd__dfxtp_1_571/CLK
+ sky130_fd_sc_hd__dfxtp_1_572/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_582 VDD VSS sky130_fd_sc_hd__nor4_1_7/C sky130_fd_sc_hd__dfxtp_1_591/CLK
+ sky130_fd_sc_hd__and2_0_248/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_593 VDD VSS sky130_fd_sc_hd__or4_1_2/D sky130_fd_sc_hd__dfxtp_1_595/CLK
+ sky130_fd_sc_hd__and2_0_247/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_180 VSS VDD sky130_fd_sc_hd__nand4_1_26/B sky130_fd_sc_hd__a22oi_1_126/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_191 VSS VDD sky130_fd_sc_hd__clkbuf_1_192/A sky130_fd_sc_hd__nand3_1_27/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_410 sky130_fd_sc_hd__maj3_1_57/B sky130_fd_sc_hd__maj3_1_58/A
+ sky130_fd_sc_hd__fa_2_410/A sky130_fd_sc_hd__fa_2_410/B sky130_fd_sc_hd__fa_2_411/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_421 sky130_fd_sc_hd__fa_2_420/A sky130_fd_sc_hd__fa_2_415/B
+ sky130_fd_sc_hd__ha_2_116/B sky130_fd_sc_hd__ha_2_116/A sky130_fd_sc_hd__fa_2_409/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_432 sky130_fd_sc_hd__fa_2_429/A sky130_fd_sc_hd__fa_2_431/A
+ sky130_fd_sc_hd__ha_2_125/A sky130_fd_sc_hd__ha_2_125/B sky130_fd_sc_hd__fa_2_531/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o2bb2ai_1_9 sky130_fd_sc_hd__o2bb2ai_1_9/Y sky130_fd_sc_hd__nor2_1_18/Y
+ sky130_fd_sc_hd__ha_2_148/SUM sky130_fd_sc_hd__o21ai_1_31/A1 sky130_fd_sc_hd__maj3_1_0/C
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_443 sky130_fd_sc_hd__fa_2_437/B sky130_fd_sc_hd__fa_2_444/CIN
+ sky130_fd_sc_hd__fa_2_546/A sky130_fd_sc_hd__ha_2_123/A sky130_fd_sc_hd__fa_2_551/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_454 sky130_fd_sc_hd__fa_2_451/B sky130_fd_sc_hd__fa_2_455/CIN
+ sky130_fd_sc_hd__fa_2_537/A sky130_fd_sc_hd__fa_2_454/B sky130_fd_sc_hd__fa_2_454/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_465 sky130_fd_sc_hd__maj3_1_107/B sky130_fd_sc_hd__fa_2_465/SUM
+ sky130_fd_sc_hd__fa_2_502/B sky130_fd_sc_hd__ha_2_169/B sky130_fd_sc_hd__ha_2_121/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_476 sky130_fd_sc_hd__maj3_1_100/B sky130_fd_sc_hd__maj3_1_101/A
+ sky130_fd_sc_hd__fa_2_476/A sky130_fd_sc_hd__fa_2_476/B sky130_fd_sc_hd__fa_2_477/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_487 sky130_fd_sc_hd__fa_2_490/CIN sky130_fd_sc_hd__fa_2_485/B
+ sky130_fd_sc_hd__ha_2_125/B sky130_fd_sc_hd__fa_2_487/B sky130_fd_sc_hd__fa_2_487/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_498 sky130_fd_sc_hd__maj3_1_94/B sky130_fd_sc_hd__maj3_1_95/A
+ sky130_fd_sc_hd__fa_2_498/A sky130_fd_sc_hd__fa_2_498/B sky130_fd_sc_hd__fa_2_499/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor2_1_208 sky130_fd_sc_hd__nor2_1_208/B sky130_fd_sc_hd__nor2_1_208/Y
+ sky130_fd_sc_hd__nor2_1_208/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_219 sky130_fd_sc_hd__nor2_1_225/A sky130_fd_sc_hd__nor2_1_219/Y
+ sky130_fd_sc_hd__nor2_1_220/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__buf_12_404 sky130_fd_sc_hd__buf_12_404/A sky130_fd_sc_hd__buf_12_404/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_415 sky130_fd_sc_hd__buf_8_221/X sky130_fd_sc_hd__buf_12_415/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_426 sky130_fd_sc_hd__buf_8_211/X sky130_fd_sc_hd__buf_12_482/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_437 sky130_fd_sc_hd__buf_12_437/A sky130_fd_sc_hd__buf_12_474/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_448 sky130_fd_sc_hd__buf_4_111/X sky130_fd_sc_hd__buf_12_448/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_307 sky130_fd_sc_hd__nor2_2_4/Y sky130_fd_sc_hd__clkbuf_1_377/X
+ sky130_fd_sc_hd__a22oi_1_307/B2 sky130_fd_sc_hd__clkbuf_4_180/X sky130_fd_sc_hd__nand4_1_76/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_459 sky130_fd_sc_hd__buf_6_68/X sky130_fd_sc_hd__buf_12_459/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_318 sky130_fd_sc_hd__nor3_1_22/Y sky130_fd_sc_hd__nor3_1_23/Y
+ sky130_fd_sc_hd__buf_2_218/X sky130_fd_sc_hd__buf_2_187/X sky130_fd_sc_hd__nand4_1_79/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_329 sky130_fd_sc_hd__a21oi_1_89/A1 sky130_fd_sc_hd__a211o_1_8/A2
+ sky130_fd_sc_hd__nand2_1_264/A sky130_fd_sc_hd__o21ai_1_115/Y sky130_fd_sc_hd__o211ai_1_7/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_604 sky130_fd_sc_hd__ha_2_179/B sky130_fd_sc_hd__fa_2_1036/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_604/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_615 sky130_fd_sc_hd__a211o_1_8/A2 sky130_fd_sc_hd__nor2_1_74/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_615/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_626 sky130_fd_sc_hd__clkinv_1_626/Y sky130_fd_sc_hd__nand2_1_284/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_626/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_637 sky130_fd_sc_hd__o22ai_1_155/B2 sky130_fd_sc_hd__ha_2_194/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_637/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_648 sky130_fd_sc_hd__nor2_1_98/B sky130_fd_sc_hd__nand2_1_307/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_648/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_659 sky130_fd_sc_hd__nand2_1_287/B sky130_fd_sc_hd__nor2_1_106/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_659/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_501 sky130_fd_sc_hd__nor2_1_322/A sky130_fd_sc_hd__nor2_1_321/Y
+ sky130_fd_sc_hd__a21oi_1_501/Y sky130_fd_sc_hd__nor2_1_321/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__o21ai_1_190 VSS VDD sky130_fd_sc_hd__o21ai_1_190/A2 sky130_fd_sc_hd__nand2_1_284/Y
+ sky130_fd_sc_hd__a21oi_1_165/Y sky130_fd_sc_hd__o21ai_1_190/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_13 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1142/A sky130_fd_sc_hd__nor2_2_15/Y
+ sky130_fd_sc_hd__nor3_1_38/A sky130_fd_sc_hd__fa_2_1144/A sky130_fd_sc_hd__nor3_1_38/B
+ sky130_fd_sc_hd__a222oi_1_13/Y sky130_fd_sc_hd__fa_2_1141/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_24 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1243/A sky130_fd_sc_hd__nor2_2_17/Y
+ sky130_fd_sc_hd__nor3_1_40/A sky130_fd_sc_hd__fa_2_1245/A sky130_fd_sc_hd__nor3_1_40/B
+ sky130_fd_sc_hd__a222oi_1_24/Y sky130_fd_sc_hd__fa_2_1242/B sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_35 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1276/A sky130_fd_sc_hd__nor2_2_18/Y
+ sky130_fd_sc_hd__nor3_1_41/A sky130_fd_sc_hd__fa_2_1278/A sky130_fd_sc_hd__nor3_1_41/B
+ sky130_fd_sc_hd__a222oi_1_35/Y sky130_fd_sc_hd__fa_2_1275/B sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_15 VSS VDD sky130_fd_sc_hd__xor2_1_21/X sky130_fd_sc_hd__xnor2_1_15/Y
+ sky130_fd_sc_hd__ha_2_156/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_26 VSS VDD sky130_fd_sc_hd__nor2_1_31/B sky130_fd_sc_hd__xnor2_1_26/Y
+ sky130_fd_sc_hd__nor4_1_6/B VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_550 sky130_fd_sc_hd__nand3_1_52/A sky130_fd_sc_hd__nand3_1_9/Y
+ sky130_fd_sc_hd__nor2_1_314/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_37 VSS VDD sky130_fd_sc_hd__xnor2_1_37/B sky130_fd_sc_hd__xnor2_1_37/Y
+ sky130_fd_sc_hd__nor2_1_43/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_561 sky130_fd_sc_hd__nand2_1_561/Y sky130_fd_sc_hd__buf_4_62/A
+ sky130_fd_sc_hd__nand2_1_561/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_48 VSS VDD sky130_fd_sc_hd__xnor2_1_48/B sky130_fd_sc_hd__xnor2_1_48/Y
+ sky130_fd_sc_hd__xnor2_1_48/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__xnor2_1_59 VSS VDD sky130_fd_sc_hd__xnor2_1_60/B sky130_fd_sc_hd__xnor2_1_59/Y
+ sky130_fd_sc_hd__xnor2_1_59/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_1130 sky130_fd_sc_hd__clkinv_4_39/A sky130_fd_sc_hd__buf_6_85/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1130/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a211oi_1_6 sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__nor2_1_87/Y
+ sky130_fd_sc_hd__o22ai_1_130/Y sky130_fd_sc_hd__a211oi_1_6/Y sky130_fd_sc_hd__fa_2_1012/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__dfxtp_1_390 VDD VSS sky130_fd_sc_hd__fa_2_1118/B sky130_fd_sc_hd__dfxtp_1_391/CLK
+ sky130_fd_sc_hd__and2_0_115/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__or4_1_1 sky130_fd_sc_hd__or4_1_1/C sky130_fd_sc_hd__or4_1_1/A sky130_fd_sc_hd__or4_1_1/X
+ sky130_fd_sc_hd__or4_1_1/B sky130_fd_sc_hd__or4_1_1/D VDD VSS VDD VSS sky130_fd_sc_hd__or4_1
Xsky130_fd_sc_hd__o32ai_1_9 sky130_fd_sc_hd__o32ai_1_9/A2 sky130_fd_sc_hd__o32ai_1_9/Y
+ sky130_fd_sc_hd__fa_2_1277/A sky130_fd_sc_hd__o32ai_1_9/A3 sky130_fd_sc_hd__o32ai_1_9/B2
+ sky130_fd_sc_hd__fa_2_1276/A VDD VSS VSS VDD sky130_fd_sc_hd__o32ai_1
Xsky130_fd_sc_hd__clkbuf_16_7 sky130_fd_sc_hd__buf_12_255/A sky130_fd_sc_hd__buf_4_53/X
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__fa_2_240 sky130_fd_sc_hd__maj3_1_35/B sky130_fd_sc_hd__maj3_1_36/A
+ sky130_fd_sc_hd__fa_2_240/A sky130_fd_sc_hd__fa_2_240/B sky130_fd_sc_hd__fa_2_241/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_251 sky130_fd_sc_hd__maj3_1_33/B sky130_fd_sc_hd__maj3_1_34/A
+ sky130_fd_sc_hd__fa_2_251/A sky130_fd_sc_hd__fa_2_251/B sky130_fd_sc_hd__fa_2_252/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_262 sky130_fd_sc_hd__fa_2_264/CIN sky130_fd_sc_hd__fa_2_259/A
+ sky130_fd_sc_hd__fa_2_281/B sky130_fd_sc_hd__fa_2_262/B sky130_fd_sc_hd__fa_2_262/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_273 sky130_fd_sc_hd__fa_2_272/A sky130_fd_sc_hd__fa_2_273/SUM
+ sky130_fd_sc_hd__fa_2_273/A sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__fa_2_281/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_284 sky130_fd_sc_hd__fa_2_292/CIN sky130_fd_sc_hd__nor2_1_210/A
+ sky130_fd_sc_hd__fa_2_284/A sky130_fd_sc_hd__fa_2_284/B sky130_fd_sc_hd__fa_2_284/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_0 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_0/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__or2_0_0/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__fa_2_295 sky130_fd_sc_hd__fa_2_285/A sky130_fd_sc_hd__fa_2_293/B
+ sky130_fd_sc_hd__fa_2_424/B sky130_fd_sc_hd__fa_2_295/B sky130_fd_sc_hd__fa_2_298/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor4_1_7 sky130_fd_sc_hd__nor4_1_7/D sky130_fd_sc_hd__nor4_1_7/C
+ sky130_fd_sc_hd__nor4_1_7/Y sky130_fd_sc_hd__nor4_1_7/A sky130_fd_sc_hd__nor4_1_7/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__nor4_1
Xsky130_fd_sc_hd__a22oi_1_6 sky130_fd_sc_hd__nor2_2_0/Y sky130_fd_sc_hd__clkinv_1_4/Y
+ sky130_fd_sc_hd__nand4_1_28/Y sky130_fd_sc_hd__nand4_1_12/Y sky130_fd_sc_hd__a22oi_1_6/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__diode_2_101 sky130_fd_sc_hd__inv_2_135/Y VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_112 sky130_fd_sc_hd__buf_2_225/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_123 sky130_fd_sc_hd__buf_2_250/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_134 sky130_fd_sc_hd__clkbuf_1_526/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_145 sky130_fd_sc_hd__buf_2_168/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_156 sky130_fd_sc_hd__clkbuf_4_174/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_167 sky130_fd_sc_hd__clkbuf_4_182/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_178 sky130_fd_sc_hd__nand4_1_79/D VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_189 sky130_fd_sc_hd__buf_2_153/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__buf_2_290 VDD VSS sky130_fd_sc_hd__buf_2_290/X sky130_fd_sc_hd__buf_2_290/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__clkbuf_4_209 sky130_fd_sc_hd__buf_2_250/A sky130_fd_sc_hd__buf_2_251/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_12_201 sky130_fd_sc_hd__buf_12_201/A sky130_fd_sc_hd__buf_12_201/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_212 sky130_fd_sc_hd__buf_12_212/A sky130_fd_sc_hd__buf_12_212/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_223 sky130_fd_sc_hd__buf_6_29/X sky130_fd_sc_hd__buf_12_223/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_70 sky130_fd_sc_hd__nand2_1_246/Y sky130_fd_sc_hd__nor2_1_53/Y
+ sky130_fd_sc_hd__xnor2_1_43/A sky130_fd_sc_hd__xnor2_1_41/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_234 sky130_fd_sc_hd__buf_12_234/A sky130_fd_sc_hd__buf_12_234/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_81 sky130_fd_sc_hd__nor2_2_9/A sky130_fd_sc_hd__nor2_1_71/Y
+ sky130_fd_sc_hd__a21oi_1_81/Y sky130_fd_sc_hd__a32o_1_0/A3 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_245 sky130_fd_sc_hd__buf_12_245/A sky130_fd_sc_hd__buf_12_245/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_92 sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__o211ai_1_6/Y
+ sky130_fd_sc_hd__a21oi_1_92/Y sky130_fd_sc_hd__fa_2_991/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_1_104 sky130_fd_sc_hd__a22oi_1_96/B1 sky130_fd_sc_hd__a22oi_1_96/A1
+ sky130_fd_sc_hd__clkbuf_1_149/X sky130_fd_sc_hd__a22oi_1_104/A2 sky130_fd_sc_hd__nand4_1_21/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_256 sky130_fd_sc_hd__buf_12_256/A sky130_fd_sc_hd__buf_12_256/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_115 sky130_fd_sc_hd__clkbuf_4_72/X sky130_fd_sc_hd__clkbuf_4_73/X
+ sky130_fd_sc_hd__a22oi_1_115/B2 sky130_fd_sc_hd__buf_2_90/X sky130_fd_sc_hd__clkbuf_4_92/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_267 sky130_fd_sc_hd__buf_12_267/A sky130_fd_sc_hd__buf_12_267/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_126 sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__a22oi_2_12/A1
+ sky130_fd_sc_hd__buf_2_71/X sky130_fd_sc_hd__clkbuf_1_162/X sky130_fd_sc_hd__a22oi_1_126/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_278 sky130_fd_sc_hd__inv_2_102/Y sky130_fd_sc_hd__buf_12_278/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_137 sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__a22oi_2_12/A1
+ sky130_fd_sc_hd__buf_2_68/X sky130_fd_sc_hd__clkbuf_1_159/X sky130_fd_sc_hd__a22oi_1_137/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_289 sky130_fd_sc_hd__buf_6_39/X sky130_fd_sc_hd__buf_12_289/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_148 sky130_fd_sc_hd__clkbuf_1_351/X sky130_fd_sc_hd__clkbuf_1_353/X
+ sky130_fd_sc_hd__clkbuf_4_121/X sky130_fd_sc_hd__a22oi_1_148/A2 sky130_fd_sc_hd__nand4_1_32/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_159 sky130_fd_sc_hd__clkbuf_1_265/X sky130_fd_sc_hd__clkbuf_1_266/X
+ sky130_fd_sc_hd__clkbuf_1_336/X sky130_fd_sc_hd__a22oi_1_159/A2 sky130_fd_sc_hd__a22oi_1_159/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_401 sky130_fd_sc_hd__nor4_1_5/C sky130_fd_sc_hd__nor2_1_29/Y
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_412 sky130_fd_sc_hd__a21oi_1_24/A2 sky130_fd_sc_hd__nand2b_1_7/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_412/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_423 sky130_fd_sc_hd__nor3_1_36/A sky130_fd_sc_hd__dfxtp_1_486/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_423/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_434 sky130_fd_sc_hd__fa_2_966/B sky130_fd_sc_hd__nand2_1_223/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_434/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_445 sky130_fd_sc_hd__fa_2_957/B sky130_fd_sc_hd__nor2b_1_89/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_445/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_456 sky130_fd_sc_hd__fa_2_945/B sky130_fd_sc_hd__nor2_1_36/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_456/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_467 sky130_fd_sc_hd__o22ai_1_75/B2 sky130_fd_sc_hd__ha_2_184/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_467/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_478 sky130_fd_sc_hd__o22ai_1_83/B2 sky130_fd_sc_hd__ha_2_176/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_478/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_489 sky130_fd_sc_hd__nor2_1_47/B sky130_fd_sc_hd__nand2_1_249/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_489/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_320 sky130_fd_sc_hd__nor2_2_16/Y sky130_fd_sc_hd__o21ai_1_339/Y
+ sky130_fd_sc_hd__nor2_1_206/B sky130_fd_sc_hd__fa_2_1196/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_331 sky130_fd_sc_hd__nand2_1_439/B sky130_fd_sc_hd__o22ai_1_301/Y
+ sky130_fd_sc_hd__a21oi_1_331/Y sky130_fd_sc_hd__o21ai_1_361/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_342 sky130_fd_sc_hd__nor2b_2_3/Y sky130_fd_sc_hd__o21ai_1_369/Y
+ sky130_fd_sc_hd__a21oi_1_342/Y sky130_fd_sc_hd__o21ai_1_382/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_353 sky130_fd_sc_hd__fa_2_1205/A sky130_fd_sc_hd__o22ai_1_314/Y
+ sky130_fd_sc_hd__a21oi_1_353/Y sky130_fd_sc_hd__nor3_1_39/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_364 sky130_fd_sc_hd__o21a_1_47/B1 sky130_fd_sc_hd__o21a_1_46/A1
+ sky130_fd_sc_hd__a21oi_1_364/Y sky130_fd_sc_hd__nor2_1_230/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_90 sky130_fd_sc_hd__clkbuf_4_208/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_375 sky130_fd_sc_hd__nor2_1_241/A sky130_fd_sc_hd__o21a_1_54/A1
+ sky130_fd_sc_hd__a21oi_1_375/Y sky130_fd_sc_hd__nor2_1_241/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_386 sky130_fd_sc_hd__fa_2_1232/A sky130_fd_sc_hd__o22ai_1_356/Y
+ sky130_fd_sc_hd__a21oi_1_386/Y sky130_fd_sc_hd__nor3_1_40/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_397 sky130_fd_sc_hd__fa_2_1235/A sky130_fd_sc_hd__o22ai_1_361/Y
+ sky130_fd_sc_hd__a21oi_1_397/Y sky130_fd_sc_hd__nor2_2_17/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_1 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1015/A sky130_fd_sc_hd__nor2_2_7/Y
+ sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_4_9/B sky130_fd_sc_hd__nor2_2_7/A
+ sky130_fd_sc_hd__a222oi_1_1/Y sky130_fd_sc_hd__fa_2_1014/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2_1_380 sky130_fd_sc_hd__nand2_1_380/Y sky130_fd_sc_hd__fa_2_1139/A
+ sky130_fd_sc_hd__nor3_1_38/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xor2_1_208 sky130_fd_sc_hd__xor2_1_209/X sky130_fd_sc_hd__xor2_1_208/X
+ sky130_fd_sc_hd__xor2_1_208/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_391 sky130_fd_sc_hd__nor2_1_183/A sky130_fd_sc_hd__nor2b_1_104/A
+ sky130_fd_sc_hd__o32ai_1_2/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_990 sky130_fd_sc_hd__clkinv_1_990/Y sky130_fd_sc_hd__nor2_1_257/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_990/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor2_1_219 sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__fa_2_1199/B
+ sky130_fd_sc_hd__xor2_1_219/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_2_13 VDD VSS sky130_fd_sc_hd__buf_2_13/X sky130_fd_sc_hd__ha_2_15/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_24 VDD VSS sky130_fd_sc_hd__buf_2_24/X sky130_fd_sc_hd__buf_2_24/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_35 VDD VSS sky130_fd_sc_hd__buf_2_35/X sky130_fd_sc_hd__buf_2_35/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_46 VDD VSS sky130_fd_sc_hd__buf_8_76/A sky130_fd_sc_hd__ha_2_39/B
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_57 VDD VSS sky130_fd_sc_hd__buf_2_57/X sky130_fd_sc_hd__buf_2_57/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_68 VDD VSS sky130_fd_sc_hd__buf_2_68/X sky130_fd_sc_hd__buf_2_68/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_79 VDD VSS sky130_fd_sc_hd__buf_2_79/X sky130_fd_sc_hd__buf_2_79/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o211ai_1_40 sky130_fd_sc_hd__a21oi_1_335/Y sky130_fd_sc_hd__nor2_1_224/A
+ sky130_fd_sc_hd__xor2_1_220/A sky130_fd_sc_hd__a211oi_1_18/Y sky130_fd_sc_hd__nand2_1_431/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_51 sky130_fd_sc_hd__nor2_1_257/A sky130_fd_sc_hd__a222oi_1_26/Y
+ sky130_fd_sc_hd__xor2_1_264/A sky130_fd_sc_hd__nand2_1_482/Y sky130_fd_sc_hd__a21oi_1_387/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_62 sky130_fd_sc_hd__nor2_1_302/B sky130_fd_sc_hd__nor2_1_307/A
+ sky130_fd_sc_hd__xor2_1_308/A sky130_fd_sc_hd__nand2_1_533/Y sky130_fd_sc_hd__a21oi_1_445/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__diode_2_8 sky130_fd_sc_hd__clkbuf_1_247/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__nor4_1_10 sky130_fd_sc_hd__nor4_1_10/D sky130_fd_sc_hd__nor4_1_10/C
+ sky130_fd_sc_hd__nor4_1_10/Y sky130_fd_sc_hd__nor4_1_10/A sky130_fd_sc_hd__nor4_1_10/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__nor4_1
Xsky130_fd_sc_hd__clkinv_1_220 sky130_fd_sc_hd__clkinv_2_30/A sky130_fd_sc_hd__a22o_1_24/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_220/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_231 sky130_fd_sc_hd__inv_2_123/A sky130_fd_sc_hd__buf_8_202/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_231/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_242 sky130_fd_sc_hd__buf_8_184/A sky130_fd_sc_hd__clkinv_1_242/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_242/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_253 sky130_fd_sc_hd__inv_2_129/A sky130_fd_sc_hd__inv_2_125/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_253/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_264 sky130_fd_sc_hd__maj3_1_3/C sky130_fd_sc_hd__ha_2_156/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_264/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_275 sky130_fd_sc_hd__fa_2_45/A sky130_fd_sc_hd__ha_2_94/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_275/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_2_9 sky130_fd_sc_hd__or2_1_1/B sky130_fd_sc_hd__ha_2_86/A sky130_fd_sc_hd__a22o_2_9/X
+ sky130_fd_sc_hd__a22o_2_9/B2 sky130_fd_sc_hd__a22o_4_0/B1 VDD VSS VDD VSS sky130_fd_sc_hd__a22o_2
Xsky130_fd_sc_hd__o31ai_1_8 sky130_fd_sc_hd__o31ai_1_8/Y sky130_fd_sc_hd__o31ai_1_8/A2
+ sky130_fd_sc_hd__o31ai_1_8/A1 sky130_fd_sc_hd__o31ai_1_8/A3 sky130_fd_sc_hd__o31ai_1_8/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__o31ai_1
Xsky130_fd_sc_hd__clkinv_1_286 sky130_fd_sc_hd__fa_2_96/A sky130_fd_sc_hd__fa_2_67/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_286/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_297 sky130_fd_sc_hd__fa_2_274/A sky130_fd_sc_hd__fa_2_242/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_297/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_5 sky130_fd_sc_hd__o21ai_1_8/A1 sky130_fd_sc_hd__nor2_1_22/A
+ sky130_fd_sc_hd__a21oi_1_5/Y sky130_fd_sc_hd__nor4_1_2/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkbuf_4_18 sky130_fd_sc_hd__clkbuf_4_18/X sky130_fd_sc_hd__clkbuf_4_18/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_29 sky130_fd_sc_hd__clkbuf_4_29/X sky130_fd_sc_hd__clkbuf_4_29/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__a21oi_1_150 sky130_fd_sc_hd__nor2_2_11/Y sky130_fd_sc_hd__o22ai_1_149/Y
+ sky130_fd_sc_hd__a21oi_1_150/Y sky130_fd_sc_hd__fa_2_1107/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_161 sky130_fd_sc_hd__nor2_2_11/Y sky130_fd_sc_hd__o22ai_1_160/Y
+ sky130_fd_sc_hd__a21oi_1_161/Y sky130_fd_sc_hd__fa_2_1118/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_172 sky130_fd_sc_hd__clkinv_1_661/Y sky130_fd_sc_hd__nor2_1_92/B
+ sky130_fd_sc_hd__xnor2_1_65/A sky130_fd_sc_hd__xnor2_1_63/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_183 sky130_fd_sc_hd__o21a_1_13/B1 sky130_fd_sc_hd__o21a_1_12/A1
+ sky130_fd_sc_hd__dfxtp_1_760/D sky130_fd_sc_hd__nor2_1_116/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_194 sky130_fd_sc_hd__nand2_1_319/A sky130_fd_sc_hd__o21ai_1_220/Y
+ sky130_fd_sc_hd__a21oi_1_194/Y sky130_fd_sc_hd__a211o_1_9/A1 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_102 sky130_fd_sc_hd__inv_2_69/Y sky130_fd_sc_hd__buf_8_102/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_113 sky130_fd_sc_hd__buf_8_113/A sky130_fd_sc_hd__buf_6_24/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_124 sky130_fd_sc_hd__buf_8_124/A sky130_fd_sc_hd__buf_6_38/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_135 sky130_fd_sc_hd__buf_8_135/A sky130_fd_sc_hd__buf_4_79/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_146 sky130_fd_sc_hd__buf_8_146/A sky130_fd_sc_hd__buf_4_87/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nor2_4_8 sky130_fd_sc_hd__nor2_4_8/Y sky130_fd_sc_hd__nor3_2_9/A
+ sky130_fd_sc_hd__nor2_4_8/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__buf_8_157 sky130_fd_sc_hd__inv_2_76/A sky130_fd_sc_hd__buf_8_169/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_168 sky130_fd_sc_hd__buf_4_68/X sky130_fd_sc_hd__buf_8_168/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_179 sky130_fd_sc_hd__buf_8_179/A sky130_fd_sc_hd__buf_8_179/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__a21o_2_14 sky130_fd_sc_hd__a21o_2_14/X sky130_fd_sc_hd__nor2_1_210/Y
+ sky130_fd_sc_hd__nor2_1_210/A sky130_fd_sc_hd__nor2_1_210/B VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__a21o_2_25 sky130_fd_sc_hd__a21o_2_25/X sky130_fd_sc_hd__nor2_1_294/Y
+ sky130_fd_sc_hd__fa_2_7/SUM sky130_fd_sc_hd__nor2_1_294/B VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__xor2_1_30 sky130_fd_sc_hd__xor2_1_30/B sky130_fd_sc_hd__xor2_1_30/X
+ sky130_fd_sc_hd__xor2_1_30/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_41 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_986/B
+ sky130_fd_sc_hd__xor2_1_41/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_52 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_975/B
+ sky130_fd_sc_hd__xor2_1_52/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_63 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__xor2_1_63/X
+ sky130_fd_sc_hd__xor2_1_63/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__buf_12_19 sky130_fd_sc_hd__inv_2_39/Y sky130_fd_sc_hd__buf_12_19/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__xor2_1_74 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__xor2_1_74/X
+ sky130_fd_sc_hd__xor2_1_74/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_85 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__xor2_1_85/X
+ sky130_fd_sc_hd__xor2_1_85/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_96 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__xor2_1_96/X
+ sky130_fd_sc_hd__xor2_1_96/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2b_1_2 sky130_fd_sc_hd__nand3_4_1/A sky130_fd_sc_hd__dfxtp_1_81/Q
+ sky130_fd_sc_hd__a22o_2_3/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__dfxtp_1_1307 VDD VSS sky130_fd_sc_hd__fa_2_844/B sky130_fd_sc_hd__dfxtp_1_1322/CLK
+ sky130_fd_sc_hd__o21a_1_66/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1318 VDD VSS sky130_fd_sc_hd__ha_2_168/A sky130_fd_sc_hd__dfxtp_1_1332/CLK
+ sky130_fd_sc_hd__a21oi_1_428/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1329 VDD VSS sky130_fd_sc_hd__fa_2_913/A sky130_fd_sc_hd__dfxtp_1_1329/CLK
+ sky130_fd_sc_hd__o21a_1_57/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_901 VDD VSS sky130_fd_sc_hd__fa_2_936/B sky130_fd_sc_hd__dfxtp_1_902/CLK
+ sky130_fd_sc_hd__dfxtp_1_901/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_912 VDD VSS sky130_fd_sc_hd__fa_2_1141/A sky130_fd_sc_hd__clkinv_8_55/Y
+ sky130_fd_sc_hd__and2_0_322/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_923 VDD VSS sky130_fd_sc_hd__fa_2_1152/A sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__mux2_2_88/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_934 VDD VSS sky130_fd_sc_hd__fa_2_1126/A sky130_fd_sc_hd__clkinv_8_55/Y
+ sky130_fd_sc_hd__mux2_2_111/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_945 VDD VSS sky130_fd_sc_hd__fa_2_1137/A sky130_fd_sc_hd__clkinv_8_46/Y
+ sky130_fd_sc_hd__mux2_2_83/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_956 VDD VSS sky130_fd_sc_hd__fa_2_1165/A sky130_fd_sc_hd__clkinv_8_65/Y
+ sky130_fd_sc_hd__mux2_2_112/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a221oi_1_0 sky130_fd_sc_hd__o21ai_1_6/B1 sky130_fd_sc_hd__o21ai_1_7/Y
+ sky130_fd_sc_hd__nor2_1_9/B sky130_fd_sc_hd__nor2_1_9/A sky130_fd_sc_hd__nor2_1_9/Y
+ sky130_fd_sc_hd__or4_1_1/A VSS VDD VDD VSS sky130_fd_sc_hd__a221oi_1
Xsky130_fd_sc_hd__dfxtp_1_967 VDD VSS sky130_fd_sc_hd__nor2_2_15/A sky130_fd_sc_hd__clkinv_8_46/Y
+ sky130_fd_sc_hd__nor2b_1_107/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_978 VDD VSS sky130_fd_sc_hd__mux2_2_96/A0 sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__o22ai_1_217/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_989 VDD VSS sky130_fd_sc_hd__mux2_2_122/A0 sky130_fd_sc_hd__clkinv_8_64/Y
+ sky130_fd_sc_hd__dfxtp_1_989/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_510 VSS VDD sky130_fd_sc_hd__buf_8_216/A sky130_fd_sc_hd__buf_2_240/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_521 VSS VDD sky130_fd_sc_hd__clkbuf_1_521/X sky130_fd_sc_hd__clkbuf_1_521/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_532 VSS VDD sky130_fd_sc_hd__clkbuf_1_532/X sky130_fd_sc_hd__clkbuf_1_532/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_100 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_91/A sky130_fd_sc_hd__fa_2_191/CIN
+ sky130_fd_sc_hd__fa_2_187/B sky130_fd_sc_hd__ha_2_91/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_543 VSS VDD sky130_fd_sc_hd__fa_2_57/A sky130_fd_sc_hd__ha_2_99/B
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_111 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_112/A sky130_fd_sc_hd__fa_2_345/B
+ sky130_fd_sc_hd__fa_2_341/A sky130_fd_sc_hd__ha_2_115/A sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_554 VSS VDD sky130_fd_sc_hd__fa_2_32/A sky130_fd_sc_hd__ha_2_95/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_122 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_123/B sky130_fd_sc_hd__fa_2_526/CIN
+ sky130_fd_sc_hd__fa_2_518/A sky130_fd_sc_hd__ha_2_122/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_565 VSS VDD sky130_fd_sc_hd__buf_4_60/A sky130_fd_sc_hd__dfxtp_1_1458/Q
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_133 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_133/A sky130_fd_sc_hd__fa_2_688/B
+ sky130_fd_sc_hd__fa_2_685/A sky130_fd_sc_hd__ha_2_133/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_576 VSS VDD sky130_fd_sc_hd__nand3_1_14/B sky130_fd_sc_hd__a22oi_1_26/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_144 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_144/A sky130_fd_sc_hd__fa_2_828/A
+ sky130_fd_sc_hd__ha_2_144/SUM sky130_fd_sc_hd__ha_2_144/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_587 VSS VDD sky130_fd_sc_hd__nand3_1_5/B sky130_fd_sc_hd__a22oi_1_10/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_155 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_155/A sky130_fd_sc_hd__ha_2_154/B
+ sky130_fd_sc_hd__ha_2_155/SUM sky130_fd_sc_hd__ha_2_155/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_598 VSS VDD sky130_fd_sc_hd__a22o_1_3/A1 sky130_fd_sc_hd__clkbuf_1_598/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_806 sky130_fd_sc_hd__fa_2_808/CIN sky130_fd_sc_hd__fa_2_800/B
+ sky130_fd_sc_hd__fa_2_806/A sky130_fd_sc_hd__fa_2_817/B sky130_fd_sc_hd__ha_2_140/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_166 VSS VDD VSS VDD sky130_fd_sc_hd__or4_1_1/D sky130_fd_sc_hd__ha_2_165/B
+ sky130_fd_sc_hd__ha_2_166/SUM sky130_fd_sc_hd__ha_2_166/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_817 sky130_fd_sc_hd__fa_2_814/A sky130_fd_sc_hd__fa_2_809/A
+ sky130_fd_sc_hd__fa_2_826/A sky130_fd_sc_hd__fa_2_817/B sky130_fd_sc_hd__fa_2_817/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_177 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_177/A sky130_fd_sc_hd__ha_2_176/A
+ sky130_fd_sc_hd__ha_2_177/SUM sky130_fd_sc_hd__ha_2_177/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_828 sky130_fd_sc_hd__fa_2_707/A sky130_fd_sc_hd__fa_2_708/B
+ sky130_fd_sc_hd__fa_2_828/A sky130_fd_sc_hd__fa_2_828/B sky130_fd_sc_hd__fa_2_828/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_188 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_188/A sky130_fd_sc_hd__ha_2_187/A
+ sky130_fd_sc_hd__ha_2_188/SUM sky130_fd_sc_hd__ha_2_188/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_839 sky130_fd_sc_hd__fa_2_838/CIN sky130_fd_sc_hd__fa_2_839/SUM
+ sky130_fd_sc_hd__fa_2_839/A sky130_fd_sc_hd__fa_2_839/B sky130_fd_sc_hd__fa_2_839/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_199 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_199/A sky130_fd_sc_hd__ha_2_198/A
+ sky130_fd_sc_hd__ha_2_199/SUM sky130_fd_sc_hd__ha_2_199/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__maj3_1_4 sky130_fd_sc_hd__maj3_1_5/X sky130_fd_sc_hd__maj3_1_4/X
+ sky130_fd_sc_hd__maj3_1_4/B sky130_fd_sc_hd__maj3_1_4/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__ha_2_90 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_99/A sky130_fd_sc_hd__maj3_1_29/C
+ sky130_fd_sc_hd__ha_2_90/SUM sky130_fd_sc_hd__ha_2_99/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__mux2_2_106 VSS VDD sky130_fd_sc_hd__mux2_2_106/A1 sky130_fd_sc_hd__mux2_2_106/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_106/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_117 VSS VDD sky130_fd_sc_hd__mux2_2_117/A1 sky130_fd_sc_hd__mux2_2_117/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_117/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_128 VSS VDD sky130_fd_sc_hd__mux2_2_128/A1 sky130_fd_sc_hd__mux2_2_128/A0
+ sky130_fd_sc_hd__mux2_2_135/S sky130_fd_sc_hd__mux2_2_128/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_139 VSS VDD sky130_fd_sc_hd__mux2_2_139/A1 sky130_fd_sc_hd__mux2_2_139/A0
+ sky130_fd_sc_hd__mux2_2_171/S sky130_fd_sc_hd__mux2_2_139/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__and2_0_13 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_13/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_9/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_24 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_24/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_32/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_304 sky130_fd_sc_hd__o22ai_1_322/A2 sky130_fd_sc_hd__nor2_1_185/B
+ sky130_fd_sc_hd__o22ai_1_304/Y sky130_fd_sc_hd__o22ai_1_304/A1 sky130_fd_sc_hd__o32ai_1_5/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_35 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_35/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_33/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_315 sky130_fd_sc_hd__o22ai_1_322/A2 sky130_fd_sc_hd__o22ai_1_315/B1
+ sky130_fd_sc_hd__o22ai_1_315/Y sky130_fd_sc_hd__nor2_1_196/B sky130_fd_sc_hd__o32ai_1_5/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_46 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_53/A sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__ha_2_55/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_326 sky130_fd_sc_hd__nand2_1_462/Y sky130_fd_sc_hd__nand2_1_461/Y
+ sky130_fd_sc_hd__o22ai_1_326/Y sky130_fd_sc_hd__nand2_1_472/B sky130_fd_sc_hd__o21ai_1_386/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_57 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_57/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_57/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_337 sky130_fd_sc_hd__nand2_1_464/Y sky130_fd_sc_hd__o21ai_1_385/Y
+ sky130_fd_sc_hd__o22ai_1_337/Y sky130_fd_sc_hd__nand2_1_471/B sky130_fd_sc_hd__nand2_1_463/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_68 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_77/A sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__ha_2_77/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_348 sky130_fd_sc_hd__nand2_1_464/Y sky130_fd_sc_hd__nand2_1_463/Y
+ sky130_fd_sc_hd__o22ai_1_348/Y sky130_fd_sc_hd__o22ai_1_348/A1 sky130_fd_sc_hd__a21o_2_23/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_79 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_79/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__and2_0_79/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_359 sky130_fd_sc_hd__o22ai_1_379/A2 sky130_fd_sc_hd__o22ai_1_366/B1
+ sky130_fd_sc_hd__o22ai_1_359/Y sky130_fd_sc_hd__nor2_1_229/B sky130_fd_sc_hd__o22ai_1_375/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_2_5 sky130_fd_sc_hd__nor2_2_5/B sky130_fd_sc_hd__nor2_2_5/Y
+ sky130_fd_sc_hd__nor2_2_5/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__buf_8_12 sky130_fd_sc_hd__buf_8_49/A sky130_fd_sc_hd__buf_8_12/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_23 sky130_fd_sc_hd__buf_8_23/A sky130_fd_sc_hd__buf_8_23/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_34 sky130_fd_sc_hd__buf_8_34/A sky130_fd_sc_hd__buf_8_34/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_45 sky130_fd_sc_hd__buf_8_45/A sky130_fd_sc_hd__buf_8_45/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_56 sky130_fd_sc_hd__buf_8_56/A sky130_fd_sc_hd__buf_8_56/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_67 sky130_fd_sc_hd__buf_8_67/A sky130_fd_sc_hd__buf_8_67/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_78 sky130_fd_sc_hd__buf_8_78/A sky130_fd_sc_hd__buf_8_78/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_89 sky130_fd_sc_hd__buf_8_89/A sky130_fd_sc_hd__buf_8_89/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_208 VDD VSS sky130_fd_sc_hd__ha_2_73/A sky130_fd_sc_hd__dfxtp_1_212/CLK
+ sky130_fd_sc_hd__and2_0_78/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_219 VDD VSS sky130_fd_sc_hd__ha_2_84/A sky130_fd_sc_hd__dfxtp_1_224/CLK
+ sky130_fd_sc_hd__nor2b_1_49/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_2_108 VDD VSS sky130_fd_sc_hd__buf_2_108/X sky130_fd_sc_hd__buf_2_108/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__fa_2_1307 sky130_fd_sc_hd__fa_2_1308/CIN sky130_fd_sc_hd__mux2_2_228/A0
+ sky130_fd_sc_hd__fa_2_1307/A sky130_fd_sc_hd__fa_2_1307/B sky130_fd_sc_hd__fa_2_1307/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_119 VDD VSS sky130_fd_sc_hd__buf_2_119/X sky130_fd_sc_hd__buf_2_119/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__fa_2_1318 sky130_fd_sc_hd__fa_2_1319/CIN sky130_fd_sc_hd__mux2_2_256/A1
+ sky130_fd_sc_hd__fa_2_1318/A sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1318/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1104 VDD VSS sky130_fd_sc_hd__fa_2_1223/A sky130_fd_sc_hd__clkinv_8_78/Y
+ sky130_fd_sc_hd__nand2_1_415/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1115 VDD VSS sky130_fd_sc_hd__mux2_2_156/A0 sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__o22ai_1_278/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1126 VDD VSS sky130_fd_sc_hd__mux2_2_129/A1 sky130_fd_sc_hd__clkinv_8_70/Y
+ sky130_fd_sc_hd__o22ai_1_267/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1137 VDD VSS sky130_fd_sc_hd__mux2_2_157/A0 sky130_fd_sc_hd__clkinv_8_64/Y
+ sky130_fd_sc_hd__dfxtp_1_996/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1148 VDD VSS sky130_fd_sc_hd__mux2_2_149/A0 sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__o22ai_1_289/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_720 VDD VSS sky130_fd_sc_hd__mux2_2_34/A0 sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__o21ai_1_57/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1159 VDD VSS sky130_fd_sc_hd__mux2_2_124/A1 sky130_fd_sc_hd__clkinv_8_70/Y
+ sky130_fd_sc_hd__a221oi_1_3/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_731 VDD VSS sky130_fd_sc_hd__mux2_2_10/A1 sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__o21ai_1_68/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_742 VDD VSS sky130_fd_sc_hd__and2_0_165/A sky130_fd_sc_hd__dfxtp_1_744/CLK
+ sky130_fd_sc_hd__fa_2_1097/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_753 VDD VSS sky130_fd_sc_hd__fa_2_667/B sky130_fd_sc_hd__dfxtp_1_755/CLK
+ sky130_fd_sc_hd__dfxtp_1_753/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_764 VDD VSS sky130_fd_sc_hd__ha_2_135/B sky130_fd_sc_hd__dfxtp_1_764/CLK
+ sky130_fd_sc_hd__dfxtp_1_764/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_775 VDD VSS sky130_fd_sc_hd__fa_2_1074/A sky130_fd_sc_hd__clkinv_8_54/Y
+ sky130_fd_sc_hd__and2_0_318/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__ha_2_8 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_8/A sky130_fd_sc_hd__ha_2_7/B
+ sky130_fd_sc_hd__ha_2_8/SUM sky130_fd_sc_hd__ha_2_8/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__dfxtp_1_786 VDD VSS sky130_fd_sc_hd__fa_2_1085/A sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__mux2_2_52/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_797 VDD VSS sky130_fd_sc_hd__fa_2_1049/A sky130_fd_sc_hd__clkinv_8_54/Y
+ sky130_fd_sc_hd__and2_0_309/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_340 VSS VDD sky130_fd_sc_hd__buf_8_148/A sky130_fd_sc_hd__buf_6_34/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_351 VSS VDD sky130_fd_sc_hd__clkbuf_1_351/X sky130_fd_sc_hd__nor3_1_14/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_362 VSS VDD sky130_fd_sc_hd__clkbuf_1_362/X sky130_fd_sc_hd__buf_6_39/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_373 VSS VDD sky130_fd_sc_hd__buf_8_192/A sky130_fd_sc_hd__buf_2_158/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_384 VSS VDD sky130_fd_sc_hd__clkbuf_1_384/X sky130_fd_sc_hd__clkbuf_1_384/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_395 VSS VDD sky130_fd_sc_hd__a22oi_2_15/B2 sky130_fd_sc_hd__clkbuf_1_395/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_603 sky130_fd_sc_hd__fa_2_605/B sky130_fd_sc_hd__fa_2_601/A
+ sky130_fd_sc_hd__fa_2_683/B sky130_fd_sc_hd__ha_2_130/B sky130_fd_sc_hd__fa_2_700/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_614 sky130_fd_sc_hd__maj3_1_119/B sky130_fd_sc_hd__maj3_1_120/A
+ sky130_fd_sc_hd__fa_2_614/A sky130_fd_sc_hd__fa_2_614/B sky130_fd_sc_hd__fa_2_615/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_19 VSS VDD sky130_fd_sc_hd__clkbuf_1_19/X sky130_fd_sc_hd__clkbuf_1_19/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_625 sky130_fd_sc_hd__fa_2_627/CIN sky130_fd_sc_hd__fa_2_622/A
+ sky130_fd_sc_hd__fa_2_692/A sky130_fd_sc_hd__fa_2_625/B sky130_fd_sc_hd__fa_2_625/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_636 sky130_fd_sc_hd__fa_2_634/A sky130_fd_sc_hd__fa_2_632/B
+ sky130_fd_sc_hd__ha_2_133/A sky130_fd_sc_hd__ha_2_133/B sky130_fd_sc_hd__fa_2_624/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_647 sky130_fd_sc_hd__fa_2_646/A sky130_fd_sc_hd__fa_2_647/SUM
+ sky130_fd_sc_hd__ha_2_134/B sky130_fd_sc_hd__ha_2_134/A sky130_fd_sc_hd__fa_2_624/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_658 sky130_fd_sc_hd__fa_2_662/CIN sky130_fd_sc_hd__fa_2_656/B
+ sky130_fd_sc_hd__ha_2_128/A sky130_fd_sc_hd__ha_2_126/A sky130_fd_sc_hd__fa_2_658/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_669 sky130_fd_sc_hd__fa_2_671/CIN sky130_fd_sc_hd__fa_2_661/A
+ sky130_fd_sc_hd__ha_2_132/A sky130_fd_sc_hd__fa_2_669/B sky130_fd_sc_hd__fa_2_669/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__conb_1_2 sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__conb_1_2/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__buf_12_8 sky130_fd_sc_hd__inv_2_16/Y sky130_fd_sc_hd__buf_12_8/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__o22ai_1_101 sky130_fd_sc_hd__o22ai_1_121/B2 sky130_fd_sc_hd__o21ai_1_92/A1
+ sky130_fd_sc_hd__o22ai_1_101/Y sky130_fd_sc_hd__o22ai_1_132/B1 sky130_fd_sc_hd__nor2_1_70/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_112 sky130_fd_sc_hd__o22ai_1_130/B1 sky130_fd_sc_hd__nor2_1_68/B
+ sky130_fd_sc_hd__o22ai_1_112/Y sky130_fd_sc_hd__o22ai_1_119/A1 sky130_fd_sc_hd__o22ai_1_132/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_123 sky130_fd_sc_hd__o22ai_1_123/A2 sky130_fd_sc_hd__o22ai_1_130/B1
+ sky130_fd_sc_hd__o22ai_1_123/Y sky130_fd_sc_hd__o22ai_1_132/B1 sky130_fd_sc_hd__o22ai_1_123/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_134 sky130_fd_sc_hd__nor2_2_9/B sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__o22ai_1_134/Y sky130_fd_sc_hd__a21oi_1_132/Y sky130_fd_sc_hd__a21boi_1_0/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_145 sky130_fd_sc_hd__nand2_1_284/Y sky130_fd_sc_hd__nand2_2_5/Y
+ sky130_fd_sc_hd__o22ai_1_145/Y sky130_fd_sc_hd__xnor2_1_82/Y sky130_fd_sc_hd__o22ai_1_159/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_209 sky130_fd_sc_hd__o21ai_1_32/B1 sky130_fd_sc_hd__buf_2_263/X
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_156 sky130_fd_sc_hd__nand2_1_338/A sky130_fd_sc_hd__nand2_1_284/Y
+ sky130_fd_sc_hd__o22ai_1_156/Y sky130_fd_sc_hd__xnor2_1_76/Y sky130_fd_sc_hd__o22ai_1_156/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_808 sky130_fd_sc_hd__nor2_1_156/B sky130_fd_sc_hd__fa_2_1144/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_808/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_2_12 sky130_fd_sc_hd__nor2_4_13/B sky130_fd_sc_hd__nor2_2_12/Y
+ sky130_fd_sc_hd__nor2_2_13/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__clkinv_1_819 sky130_fd_sc_hd__clkinv_1_819/Y sky130_fd_sc_hd__a21boi_1_1/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_819/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_167 sky130_fd_sc_hd__nor2_2_13/B sky130_fd_sc_hd__nor2_1_126/A
+ sky130_fd_sc_hd__o22ai_1_167/Y sky130_fd_sc_hd__o22ai_1_173/A2 sky130_fd_sc_hd__nor2_1_134/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_178 sky130_fd_sc_hd__o21a_1_16/A2 sky130_fd_sc_hd__nor2_1_114/B
+ sky130_fd_sc_hd__nor2_1_130/B sky130_fd_sc_hd__o22ai_1_184/B1 sky130_fd_sc_hd__o22ai_1_206/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_189 sky130_fd_sc_hd__o22ai_1_204/B1 sky130_fd_sc_hd__nor2_1_120/B
+ sky130_fd_sc_hd__nor2_1_133/A sky130_fd_sc_hd__nor2_1_120/A sky130_fd_sc_hd__o22ai_1_206/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand4_1_15 sky130_fd_sc_hd__nand4_1_15/C sky130_fd_sc_hd__nand4_1_15/B
+ sky130_fd_sc_hd__nand4_1_15/Y sky130_fd_sc_hd__nand4_1_15/D sky130_fd_sc_hd__nand4_1_15/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__o211ai_1_2 sky130_fd_sc_hd__o31ai_1_1/B1 sky130_fd_sc_hd__xor2_1_10/X
+ sky130_fd_sc_hd__nor4_1_1/B sky130_fd_sc_hd__nand2_1_32/Y sky130_fd_sc_hd__a21oi_1_8/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__nand4_1_26 sky130_fd_sc_hd__nand4_1_26/C sky130_fd_sc_hd__nand4_1_26/B
+ sky130_fd_sc_hd__nand4_1_26/Y sky130_fd_sc_hd__nand4_1_26/D sky130_fd_sc_hd__buf_2_105/X
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_37 sky130_fd_sc_hd__nand4_1_37/C sky130_fd_sc_hd__nand4_1_37/B
+ sky130_fd_sc_hd__nand4_1_37/Y sky130_fd_sc_hd__nand4_1_37/D sky130_fd_sc_hd__nand4_1_37/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_48 sky130_fd_sc_hd__nand4_1_48/C sky130_fd_sc_hd__nand4_1_48/B
+ sky130_fd_sc_hd__nand4_1_48/Y sky130_fd_sc_hd__nand4_1_48/D sky130_fd_sc_hd__nand4_1_48/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_59 sky130_fd_sc_hd__nand4_1_59/C sky130_fd_sc_hd__nand4_1_59/B
+ sky130_fd_sc_hd__nand4_1_59/Y sky130_fd_sc_hd__nand4_1_59/D sky130_fd_sc_hd__nand4_1_59/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__conb_1_19 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__conb_1_19/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__o21ai_1_350 VSS VDD sky130_fd_sc_hd__nor2_1_216/B sky130_fd_sc_hd__nor2_1_214/A
+ sky130_fd_sc_hd__a21oi_1_330/Y sky130_fd_sc_hd__o21ai_1_350/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a211oi_1_11 sky130_fd_sc_hd__nor2_1_182/Y sky130_fd_sc_hd__nor2_1_172/Y
+ sky130_fd_sc_hd__nor2_1_173/Y sky130_fd_sc_hd__a211oi_1_11/Y sky130_fd_sc_hd__fa_2_1131/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__a211oi_1_22 sky130_fd_sc_hd__nor2b_1_112/Y sky130_fd_sc_hd__nor2_1_221/Y
+ sky130_fd_sc_hd__o21ai_1_379/Y sky130_fd_sc_hd__a211oi_1_22/Y sky130_fd_sc_hd__o21ai_1_380/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_361 VSS VDD sky130_fd_sc_hd__o22ai_1_318/A2 sky130_fd_sc_hd__nor2_1_189/B
+ sky130_fd_sc_hd__a21oi_1_339/Y sky130_fd_sc_hd__o21ai_1_361/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_372 VSS VDD sky130_fd_sc_hd__a21oi_1_356/Y sky130_fd_sc_hd__nor2_1_224/A
+ sky130_fd_sc_hd__a21oi_1_347/Y sky130_fd_sc_hd__xor2_1_200/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a211oi_1_33 sky130_fd_sc_hd__nor2b_1_126/Y sky130_fd_sc_hd__o21ai_1_465/Y
+ sky130_fd_sc_hd__nor2_1_301/Y sky130_fd_sc_hd__a211oi_1_33/Y sky130_fd_sc_hd__o21ai_1_467/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_383 VSS VDD sky130_fd_sc_hd__o22ai_1_318/A2 sky130_fd_sc_hd__nor2_1_197/B
+ sky130_fd_sc_hd__a21oi_1_358/Y sky130_fd_sc_hd__o21ai_1_383/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_394 VSS VDD sky130_fd_sc_hd__nor2_1_233/B sky130_fd_sc_hd__o22ai_1_379/A2
+ sky130_fd_sc_hd__a22oi_1_388/Y sky130_fd_sc_hd__o21ai_1_394/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__mux2_2_30 VSS VDD sky130_fd_sc_hd__mux2_2_30/A1 sky130_fd_sc_hd__mux2_2_30/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_30/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_41 VSS VDD sky130_fd_sc_hd__mux2_2_41/A1 sky130_fd_sc_hd__mux2_2_41/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_41/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_52 VSS VDD sky130_fd_sc_hd__mux2_2_52/A1 sky130_fd_sc_hd__mux2_2_52/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_52/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_63 VSS VDD sky130_fd_sc_hd__mux2_2_63/A1 sky130_fd_sc_hd__mux2_2_63/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_63/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_74 VSS VDD sky130_fd_sc_hd__mux2_2_74/A1 sky130_fd_sc_hd__mux2_2_74/A0
+ sky130_fd_sc_hd__mux2_2_75/S sky130_fd_sc_hd__mux2_2_74/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_85 VSS VDD sky130_fd_sc_hd__mux2_2_85/A1 sky130_fd_sc_hd__mux2_2_85/A0
+ sky130_fd_sc_hd__nor2_4_15/A sky130_fd_sc_hd__mux2_2_85/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1104 sky130_fd_sc_hd__fa_2_1105/CIN sky130_fd_sc_hd__and2_0_317/A
+ sky130_fd_sc_hd__fa_2_1104/A sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1104/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__mux2_2_96 VSS VDD sky130_fd_sc_hd__mux2_2_96/A1 sky130_fd_sc_hd__mux2_2_96/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_96/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1115 sky130_fd_sc_hd__fa_2_1116/CIN sky130_fd_sc_hd__fa_2_1115/SUM
+ sky130_fd_sc_hd__fa_2_1115/A sky130_fd_sc_hd__fa_2_1115/B sky130_fd_sc_hd__fa_2_1115/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1126 sky130_fd_sc_hd__fa_2_1127/CIN sky130_fd_sc_hd__mux2_2_111/A1
+ sky130_fd_sc_hd__fa_2_1126/A sky130_fd_sc_hd__fa_2_1126/B sky130_fd_sc_hd__fa_2_1126/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1137 sky130_fd_sc_hd__fa_2_1138/CIN sky130_fd_sc_hd__mux2_2_83/A0
+ sky130_fd_sc_hd__fa_2_1137/A sky130_fd_sc_hd__fa_2_1137/B sky130_fd_sc_hd__fa_2_1137/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1148 sky130_fd_sc_hd__fa_2_1149/CIN sky130_fd_sc_hd__mux2_2_98/A1
+ sky130_fd_sc_hd__fa_2_1148/A sky130_fd_sc_hd__fa_2_1148/B sky130_fd_sc_hd__fa_2_1148/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1159 sky130_fd_sc_hd__fa_2_1160/CIN sky130_fd_sc_hd__mux2_2_122/A1
+ sky130_fd_sc_hd__fa_2_1159/A sky130_fd_sc_hd__fa_2_1172/B sky130_fd_sc_hd__fa_2_1159/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_550 VDD VSS sky130_fd_sc_hd__a22o_1_33/B1 sky130_fd_sc_hd__dfxtp_1_595/CLK
+ sky130_fd_sc_hd__a22o_1_33/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_561 VDD VSS sky130_fd_sc_hd__and2_0_219/A sky130_fd_sc_hd__dfxtp_1_577/CLK
+ sky130_fd_sc_hd__dfxtp_1_562/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_572 VDD VSS sky130_fd_sc_hd__dfxtp_1_572/Q sky130_fd_sc_hd__dfxtp_1_595/CLK
+ sky130_fd_sc_hd__nor2_1_25/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_583 VDD VSS sky130_fd_sc_hd__nor4_1_7/D sky130_fd_sc_hd__dfxtp_1_591/CLK
+ sky130_fd_sc_hd__and2_0_250/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_594 VDD VSS sky130_fd_sc_hd__buf_2_252/A sky130_fd_sc_hd__dfxtp_1_594/CLK
+ sky130_fd_sc_hd__nor4_1_5/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_170 VSS VDD sky130_fd_sc_hd__a22oi_1_94/A2 sky130_fd_sc_hd__clkbuf_1_170/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_181 VSS VDD sky130_fd_sc_hd__nand4_1_25/B sky130_fd_sc_hd__clkbuf_1_243/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_192 VSS VDD sky130_fd_sc_hd__clkbuf_1_192/X sky130_fd_sc_hd__clkbuf_1_192/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_400 sky130_fd_sc_hd__fa_2_397/A sky130_fd_sc_hd__fa_2_392/A
+ sky130_fd_sc_hd__fa_2_404/A sky130_fd_sc_hd__ha_2_116/B sky130_fd_sc_hd__fa_2_417/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_411 sky130_fd_sc_hd__fa_2_414/B sky130_fd_sc_hd__fa_2_411/SUM
+ sky130_fd_sc_hd__fa_2_411/A sky130_fd_sc_hd__fa_2_411/B sky130_fd_sc_hd__fa_2_411/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_422 sky130_fd_sc_hd__fa_2_320/B sky130_fd_sc_hd__fa_2_423/CIN
+ sky130_fd_sc_hd__fa_2_425/B sky130_fd_sc_hd__fa_2_422/B sky130_fd_sc_hd__fa_2_395/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_433 sky130_fd_sc_hd__fa_2_434/CIN sky130_fd_sc_hd__a21o_2_8/A1
+ sky130_fd_sc_hd__fa_2_433/A sky130_fd_sc_hd__fa_2_433/B sky130_fd_sc_hd__fa_2_433/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_444 sky130_fd_sc_hd__fa_2_435/A sky130_fd_sc_hd__fa_2_442/A
+ sky130_fd_sc_hd__fa_2_567/B sky130_fd_sc_hd__fa_2_444/B sky130_fd_sc_hd__fa_2_444/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_455 sky130_fd_sc_hd__fa_2_448/A sky130_fd_sc_hd__fa_2_452/B
+ sky130_fd_sc_hd__fa_2_455/A sky130_fd_sc_hd__fa_2_455/B sky130_fd_sc_hd__fa_2_455/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_466 sky130_fd_sc_hd__maj3_1_106/B sky130_fd_sc_hd__maj3_1_107/A
+ sky130_fd_sc_hd__ha_2_122/B sky130_fd_sc_hd__ha_2_118/B sky130_fd_sc_hd__fa_2_502/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_477 sky130_fd_sc_hd__fa_2_479/B sky130_fd_sc_hd__fa_2_477/SUM
+ sky130_fd_sc_hd__ha_2_124/B sky130_fd_sc_hd__fa_2_559/A sky130_fd_sc_hd__fa_2_477/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_488 sky130_fd_sc_hd__fa_2_487/CIN sky130_fd_sc_hd__fa_2_488/SUM
+ sky130_fd_sc_hd__fa_2_546/A sky130_fd_sc_hd__ha_2_119/A sky130_fd_sc_hd__fa_2_559/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_499 sky130_fd_sc_hd__fa_2_504/B sky130_fd_sc_hd__fa_2_499/SUM
+ sky130_fd_sc_hd__fa_2_499/A sky130_fd_sc_hd__fa_2_499/B sky130_fd_sc_hd__fa_2_499/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor2_1_209 sky130_fd_sc_hd__nor2_1_209/B sky130_fd_sc_hd__nor2_1_209/Y
+ sky130_fd_sc_hd__nor2_1_209/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__and2_0_190 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_190/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__ha_2_160/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_405 sky130_fd_sc_hd__buf_6_59/X sky130_fd_sc_hd__bufbuf_8_9/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_416 sky130_fd_sc_hd__buf_12_416/A sky130_fd_sc_hd__buf_12_416/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_427 sky130_fd_sc_hd__buf_12_427/A sky130_fd_sc_hd__buf_12_427/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_438 sky130_fd_sc_hd__buf_2_245/X sky130_fd_sc_hd__buf_12_473/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_449 sky130_fd_sc_hd__buf_6_71/X sky130_fd_sc_hd__buf_12_449/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_308 sky130_fd_sc_hd__clkbuf_1_376/X sky130_fd_sc_hd__nor2_2_5/Y
+ sky130_fd_sc_hd__buf_2_205/X sky130_fd_sc_hd__clkbuf_1_461/X sky130_fd_sc_hd__nand4_1_76/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_319 sky130_fd_sc_hd__nor2_2_4/Y sky130_fd_sc_hd__nor3_1_24/Y
+ sky130_fd_sc_hd__a22oi_1_319/B2 sky130_fd_sc_hd__clkbuf_4_177/X sky130_fd_sc_hd__nand4_1_79/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_605 sky130_fd_sc_hd__ha_2_180/B sky130_fd_sc_hd__fa_2_1035/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_605/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_616 sky130_fd_sc_hd__o22ai_1_130/B1 sky130_fd_sc_hd__nor2_4_10/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_616/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_627 sky130_fd_sc_hd__o21ai_1_171/A2 sky130_fd_sc_hd__nor2_2_11/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_627/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_638 sky130_fd_sc_hd__o22ai_1_156/B2 sky130_fd_sc_hd__ha_2_193/SUM
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_649 sky130_fd_sc_hd__nand2_1_292/B sky130_fd_sc_hd__nor2_1_111/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_649/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_180 VSS VDD sky130_fd_sc_hd__nand2_2_5/Y sky130_fd_sc_hd__xnor2_1_73/Y
+ sky130_fd_sc_hd__a21oi_1_155/Y sky130_fd_sc_hd__o21ai_1_180/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_191 VSS VDD sky130_fd_sc_hd__o21ai_1_191/A2 sky130_fd_sc_hd__nand2_1_284/Y
+ sky130_fd_sc_hd__a21oi_1_165/Y sky130_fd_sc_hd__o21ai_1_191/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_14 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1192/A sky130_fd_sc_hd__nor2_2_16/Y
+ sky130_fd_sc_hd__nor3_1_39/A sky130_fd_sc_hd__fa_2_1194/A sky130_fd_sc_hd__nor3_1_39/B
+ sky130_fd_sc_hd__a222oi_1_14/Y sky130_fd_sc_hd__fa_2_1191/B sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_25 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1225/A sky130_fd_sc_hd__nor2_2_17/Y
+ sky130_fd_sc_hd__nor3_1_40/A sky130_fd_sc_hd__fa_2_1227/A sky130_fd_sc_hd__nor3_1_40/B
+ sky130_fd_sc_hd__a222oi_1_25/Y sky130_fd_sc_hd__fa_2_1224/B sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_36 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1292/A sky130_fd_sc_hd__nor2_2_18/Y
+ sky130_fd_sc_hd__nor3_1_41/A sky130_fd_sc_hd__nor2_4_19/B sky130_fd_sc_hd__xor2_1_299/A
+ sky130_fd_sc_hd__a222oi_1_36/Y sky130_fd_sc_hd__fa_2_1291/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__xnor2_1_16 VSS VDD sky130_fd_sc_hd__maj3_1_3/B sky130_fd_sc_hd__xnor2_1_16/Y
+ sky130_fd_sc_hd__ha_2_155/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_540 sky130_fd_sc_hd__nand2_1_540/Y sky130_fd_sc_hd__nand2_1_543/B
+ sky130_fd_sc_hd__o21ai_1_485/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_27 VSS VDD sky130_fd_sc_hd__nor2_1_30/B sky130_fd_sc_hd__xnor2_1_27/Y
+ sky130_fd_sc_hd__nor4_1_7/C VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_551 sky130_fd_sc_hd__a31oi_1_4/A3 sky130_fd_sc_hd__nand3_1_12/Y
+ sky130_fd_sc_hd__nor2_1_312/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_38 VSS VDD sky130_fd_sc_hd__xnor2_1_38/B sky130_fd_sc_hd__xnor2_1_38/Y
+ sky130_fd_sc_hd__nor2_1_43/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_562 sky130_fd_sc_hd__nand2_1_562/Y sky130_fd_sc_hd__buf_6_84/X
+ sky130_fd_sc_hd__nand2_1_562/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_49 VSS VDD sky130_fd_sc_hd__xnor2_1_49/B sky130_fd_sc_hd__xnor2_1_49/Y
+ sky130_fd_sc_hd__nor2_1_46/Y VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_1120 sky130_fd_sc_hd__nor2_1_322/B sky130_fd_sc_hd__nor2_1_320/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1120/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1131 sky130_fd_sc_hd__clkinv_4_40/A sky130_fd_sc_hd__nand2_1_566/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1131/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a211oi_1_7 sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__nor2_1_88/Y
+ sky130_fd_sc_hd__o22ai_1_132/Y sky130_fd_sc_hd__a211oi_1_7/Y sky130_fd_sc_hd__fa_2_1008/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__dfxtp_1_380 VDD VSS sky130_fd_sc_hd__fa_2_1108/B sky130_fd_sc_hd__dfxtp_1_380/CLK
+ sky130_fd_sc_hd__and2_0_187/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_0 sky130_fd_sc_hd__nand3_1_0/C sky130_fd_sc_hd__nand2_1_0/B
+ sky130_fd_sc_hd__nand2_1_9/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_391 VDD VSS sky130_fd_sc_hd__nor2_1_99/A sky130_fd_sc_hd__dfxtp_1_391/CLK
+ sky130_fd_sc_hd__and2_0_110/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__or4_1_2 sky130_fd_sc_hd__or4_1_2/C sky130_fd_sc_hd__or4_1_2/A sky130_fd_sc_hd__or4_1_2/X
+ sky130_fd_sc_hd__or4_1_2/B sky130_fd_sc_hd__or4_1_2/D VDD VSS VDD VSS sky130_fd_sc_hd__or4_1
Xsky130_fd_sc_hd__clkbuf_16_8 sky130_fd_sc_hd__buf_12_370/A sky130_fd_sc_hd__inv_2_86/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__fa_2_230 sky130_fd_sc_hd__fa_2_232/CIN sky130_fd_sc_hd__fa_2_226/A
+ sky130_fd_sc_hd__fa_2_230/A sky130_fd_sc_hd__fa_2_230/B sky130_fd_sc_hd__fa_2_230/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_241 sky130_fd_sc_hd__fa_2_245/B sky130_fd_sc_hd__fa_2_241/SUM
+ sky130_fd_sc_hd__fa_2_241/A sky130_fd_sc_hd__fa_2_241/B sky130_fd_sc_hd__fa_2_241/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_252 sky130_fd_sc_hd__fa_2_255/B sky130_fd_sc_hd__fa_2_252/SUM
+ sky130_fd_sc_hd__fa_2_252/A sky130_fd_sc_hd__fa_2_252/B sky130_fd_sc_hd__fa_2_252/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_263 sky130_fd_sc_hd__maj3_1_30/B sky130_fd_sc_hd__maj3_1_31/A
+ sky130_fd_sc_hd__fa_2_263/A sky130_fd_sc_hd__fa_2_263/B sky130_fd_sc_hd__fa_2_264/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_274 sky130_fd_sc_hd__fa_2_272/B sky130_fd_sc_hd__fa_2_269/B
+ sky130_fd_sc_hd__fa_2_274/A sky130_fd_sc_hd__fa_2_280/A sky130_fd_sc_hd__fa_2_261/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_285 sky130_fd_sc_hd__fa_2_284/CIN sky130_fd_sc_hd__fa_2_285/SUM
+ sky130_fd_sc_hd__fa_2_285/A sky130_fd_sc_hd__fa_2_285/B sky130_fd_sc_hd__fa_2_285/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_1 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_1/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__and2_0_1/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__fa_2_296 sky130_fd_sc_hd__fa_2_292/A sky130_fd_sc_hd__fa_2_284/B
+ sky130_fd_sc_hd__fa_2_424/B sky130_fd_sc_hd__fa_2_296/B sky130_fd_sc_hd__fa_2_392/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor4_1_8 sky130_fd_sc_hd__nor4_1_8/D sky130_fd_sc_hd__nor4_1_8/C
+ sky130_fd_sc_hd__nor4_1_8/Y sky130_fd_sc_hd__nor4_1_8/A sky130_fd_sc_hd__nor4_1_8/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__nor4_1
Xsky130_fd_sc_hd__a22oi_1_7 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__a22oi_1_9/A1
+ sky130_fd_sc_hd__buf_2_286/X sky130_fd_sc_hd__a22oi_1_7/A2 sky130_fd_sc_hd__nand3_1_3/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__diode_2_102 sky130_fd_sc_hd__inv_2_135/Y VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_113 sky130_fd_sc_hd__buf_2_225/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_124 sky130_fd_sc_hd__buf_2_250/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_135 sky130_fd_sc_hd__clkbuf_1_526/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_146 sky130_fd_sc_hd__buf_2_168/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_157 sky130_fd_sc_hd__clkbuf_4_174/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_168 sky130_fd_sc_hd__clkbuf_4_187/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_179 sky130_fd_sc_hd__a22o_4_0/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__buf_2_280 VDD VSS sky130_fd_sc_hd__buf_2_280/X sig_frequency[1]
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_291 VDD VSS sky130_fd_sc_hd__buf_2_291/X sig_frequency[7]
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_12_202 sky130_fd_sc_hd__buf_4_54/X sky130_fd_sc_hd__buf_12_202/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_213 sky130_fd_sc_hd__buf_12_213/A sky130_fd_sc_hd__buf_12_213/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_60 sky130_fd_sc_hd__a21oi_1_60/A1 sky130_fd_sc_hd__nor2_1_47/B
+ sky130_fd_sc_hd__xnor2_1_56/A sky130_fd_sc_hd__xnor2_1_54/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_224 sky130_fd_sc_hd__buf_12_224/A sky130_fd_sc_hd__buf_12_224/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_71 sky130_fd_sc_hd__nand2_1_245/Y sky130_fd_sc_hd__nor2_1_54/Y
+ sky130_fd_sc_hd__xnor2_1_39/A sky130_fd_sc_hd__xnor2_1_37/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_235 sky130_fd_sc_hd__buf_12_235/A sky130_fd_sc_hd__buf_12_235/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_82 sky130_fd_sc_hd__a21o_2_3/A2 sky130_fd_sc_hd__o21ai_1_91/Y
+ sky130_fd_sc_hd__a21oi_1_82/Y sky130_fd_sc_hd__fa_2_997/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_246 sky130_fd_sc_hd__buf_12_246/A sky130_fd_sc_hd__buf_12_246/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_93 sky130_fd_sc_hd__fa_2_992/A sky130_fd_sc_hd__nor2_1_78/Y
+ sky130_fd_sc_hd__a21oi_1_93/Y sky130_fd_sc_hd__nor2_4_10/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_1_105 sky130_fd_sc_hd__a22oi_1_97/B1 sky130_fd_sc_hd__a22oi_1_97/A1
+ sky130_fd_sc_hd__buf_2_60/X sky130_fd_sc_hd__clkbuf_4_84/X sky130_fd_sc_hd__nand4_1_21/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_257 sky130_fd_sc_hd__buf_12_257/A sky130_fd_sc_hd__buf_12_257/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_116 sky130_fd_sc_hd__a22oi_1_96/B1 sky130_fd_sc_hd__a22oi_1_96/A1
+ sky130_fd_sc_hd__clkbuf_1_146/X sky130_fd_sc_hd__a22oi_1_116/A2 sky130_fd_sc_hd__nand4_1_24/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_268 sky130_fd_sc_hd__buf_12_268/A sky130_fd_sc_hd__buf_12_365/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_127 sky130_fd_sc_hd__clkbuf_4_72/X sky130_fd_sc_hd__clkbuf_4_73/X
+ sky130_fd_sc_hd__a22oi_1_127/B2 sky130_fd_sc_hd__buf_2_87/X sky130_fd_sc_hd__buf_2_105/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_279 sky130_fd_sc_hd__inv_2_100/Y sky130_fd_sc_hd__buf_12_357/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_138 sky130_fd_sc_hd__clkbuf_4_72/X sky130_fd_sc_hd__clkbuf_4_73/X
+ sky130_fd_sc_hd__a22oi_1_138/B2 sky130_fd_sc_hd__buf_2_84/X sky130_fd_sc_hd__buf_2_102/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_149 sky130_fd_sc_hd__clkbuf_4_111/X sky130_fd_sc_hd__clkbuf_4_112/X
+ sky130_fd_sc_hd__a22oi_1_149/B2 sky130_fd_sc_hd__clkbuf_1_297/X sky130_fd_sc_hd__a22oi_1_149/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_402 sky130_fd_sc_hd__a21o_2_2/B1 sky130_fd_sc_hd__o21ai_1_32/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_402/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_413 sky130_fd_sc_hd__o22a_1_0/B2 sky130_fd_sc_hd__xnor2_1_32/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_413/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_424 sky130_fd_sc_hd__nor2_1_39/B sky130_fd_sc_hd__fa_2_963/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_424/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_435 sky130_fd_sc_hd__fa_2_963/B sky130_fd_sc_hd__nor2_1_39/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_435/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_446 sky130_fd_sc_hd__fa_2_956/B sky130_fd_sc_hd__o21ai_1_39/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_446/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_457 sky130_fd_sc_hd__fa_2_944/B sky130_fd_sc_hd__o21ai_1_35/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_457/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_468 sky130_fd_sc_hd__o22ai_1_89/A1 sky130_fd_sc_hd__nor2_1_41/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_468/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_479 sky130_fd_sc_hd__o22ai_1_84/B2 sky130_fd_sc_hd__ha_2_175/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_479/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_310 sky130_fd_sc_hd__o21a_1_38/B1 sky130_fd_sc_hd__o21a_1_37/A1
+ sky130_fd_sc_hd__a21oi_1_310/Y sky130_fd_sc_hd__nor2_1_193/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_321 sky130_fd_sc_hd__nor2_2_16/Y sky130_fd_sc_hd__o21ai_1_340/Y
+ sky130_fd_sc_hd__nor2_1_207/B sky130_fd_sc_hd__fa_2_1178/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_332 sky130_fd_sc_hd__or2_0_10/B sky130_fd_sc_hd__o21ai_1_353/Y
+ sky130_fd_sc_hd__a21oi_1_332/Y sky130_fd_sc_hd__clkinv_1_905/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_343 sky130_fd_sc_hd__fa_2_1199/A sky130_fd_sc_hd__o22ai_1_310/Y
+ sky130_fd_sc_hd__a21oi_1_343/Y sky130_fd_sc_hd__nor3_1_39/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_354 sky130_fd_sc_hd__fa_2_1199/A sky130_fd_sc_hd__o22ai_1_315/Y
+ sky130_fd_sc_hd__a21oi_1_354/Y sky130_fd_sc_hd__nor2_2_16/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_80 sky130_fd_sc_hd__inv_12_0/Y VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_365 sky130_fd_sc_hd__nor2_1_231/A sky130_fd_sc_hd__o21a_1_47/A1
+ sky130_fd_sc_hd__a21oi_1_365/Y sky130_fd_sc_hd__nor2_1_231/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_91 sky130_fd_sc_hd__clkbuf_1_535/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_376 sky130_fd_sc_hd__nor2_1_242/A sky130_fd_sc_hd__nor2_1_242/Y
+ sky130_fd_sc_hd__a21oi_1_376/Y sky130_fd_sc_hd__nor2_1_242/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_387 sky130_fd_sc_hd__clkinv_1_987/Y sky130_fd_sc_hd__nor2_1_258/Y
+ sky130_fd_sc_hd__a21oi_1_387/Y sky130_fd_sc_hd__nor2b_2_4/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_398 sky130_fd_sc_hd__fa_2_1230/A sky130_fd_sc_hd__o22ai_1_362/Y
+ sky130_fd_sc_hd__a21oi_1_398/Y sky130_fd_sc_hd__nor3_1_40/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_2 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1068/A sky130_fd_sc_hd__nor2_4_13/Y
+ sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__xor2_1_87/A sky130_fd_sc_hd__nor2_4_13/A
+ sky130_fd_sc_hd__a222oi_1_2/Y sky130_fd_sc_hd__fa_2_1067/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2_1_370 sky130_fd_sc_hd__a21o_2_8/A2 sky130_fd_sc_hd__nand2_1_370/B
+ sky130_fd_sc_hd__a21o_2_9/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_381 sky130_fd_sc_hd__nand2_1_381/Y sky130_fd_sc_hd__nor2b_1_105/Y
+ sky130_fd_sc_hd__o21ai_1_301/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_980 sky130_fd_sc_hd__nand2_1_471/B sky130_fd_sc_hd__fa_2_144/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_980/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor2_1_209 sky130_fd_sc_hd__nor2_4_17/Y sky130_fd_sc_hd__xor2_1_209/X
+ sky130_fd_sc_hd__xor2_1_209/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2_1_392 sky130_fd_sc_hd__o32ai_1_5/A3 sky130_fd_sc_hd__nor2_4_16/B
+ sky130_fd_sc_hd__nor2_4_16/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_991 sky130_fd_sc_hd__o21ai_1_412/A2 sky130_fd_sc_hd__fa_2_1238/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_991/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_2_14 VDD VSS sky130_fd_sc_hd__buf_2_14/X sky130_fd_sc_hd__ha_2_16/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_25 VDD VSS sky130_fd_sc_hd__buf_2_25/X sky130_fd_sc_hd__buf_2_25/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_36 VDD VSS sky130_fd_sc_hd__buf_4_35/A sky130_fd_sc_hd__buf_2_36/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_47 VDD VSS sky130_fd_sc_hd__buf_2_47/X sky130_fd_sc_hd__buf_2_47/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_58 VDD VSS sky130_fd_sc_hd__buf_2_58/X sky130_fd_sc_hd__buf_2_58/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_69 VDD VSS sky130_fd_sc_hd__buf_2_69/X sky130_fd_sc_hd__buf_2_69/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o211ai_1_30 sky130_fd_sc_hd__nor2_1_180/A sky130_fd_sc_hd__a21oi_1_290/Y
+ sky130_fd_sc_hd__xor2_1_148/A sky130_fd_sc_hd__nand2_1_383/Y sky130_fd_sc_hd__nand2_1_386/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_41 sky130_fd_sc_hd__a21oi_1_335/Y sky130_fd_sc_hd__nor2_1_222/A
+ sky130_fd_sc_hd__xor2_1_224/A sky130_fd_sc_hd__a21oi_1_332/Y sky130_fd_sc_hd__nand2_1_433/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_52 sky130_fd_sc_hd__a21oi_1_395/Y sky130_fd_sc_hd__nor2_1_267/A
+ sky130_fd_sc_hd__xor2_1_265/A sky130_fd_sc_hd__a211oi_1_25/Y sky130_fd_sc_hd__nand2_1_483/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__diode_2_9 sky130_fd_sc_hd__clkbuf_1_247/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__o211ai_1_63 sky130_fd_sc_hd__nor2_1_299/A sky130_fd_sc_hd__a222oi_1_36/Y
+ sky130_fd_sc_hd__xor2_1_309/A sky130_fd_sc_hd__nand2_1_534/Y sky130_fd_sc_hd__a21oi_1_447/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__nor4_1_11 sky130_fd_sc_hd__nor4_1_11/D sky130_fd_sc_hd__nor4_1_11/C
+ sky130_fd_sc_hd__nor4_1_11/Y sky130_fd_sc_hd__nor4_1_11/A sky130_fd_sc_hd__nor4_1_11/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__nor4_1
Xsky130_fd_sc_hd__clkinv_1_210 sky130_fd_sc_hd__clkinv_2_24/A sky130_fd_sc_hd__a22oi_1_301/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_210/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_221 sky130_fd_sc_hd__buf_12_389/A sky130_fd_sc_hd__clkinv_2_30/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_221/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_232 sky130_fd_sc_hd__inv_2_124/A sky130_fd_sc_hd__inv_2_107/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_232/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_243 sky130_fd_sc_hd__clkinv_1_244/A sky130_fd_sc_hd__a22o_2_8/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_243/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_254 sky130_fd_sc_hd__inv_2_130/A sky130_fd_sc_hd__buf_2_162/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_254/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_265 sky130_fd_sc_hd__maj3_1_1/B sky130_fd_sc_hd__ha_2_149/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_265/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_276 sky130_fd_sc_hd__fa_2_80/B sky130_fd_sc_hd__fa_2_5/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_276/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o31ai_1_9 sky130_fd_sc_hd__o31ai_1_9/Y sky130_fd_sc_hd__xnor2_1_99/Y
+ sky130_fd_sc_hd__o31ai_1_9/A1 sky130_fd_sc_hd__o31ai_1_9/A3 sky130_fd_sc_hd__o31ai_1_9/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__o31ai_1
Xsky130_fd_sc_hd__clkinv_1_287 sky130_fd_sc_hd__fa_2_92/B sky130_fd_sc_hd__ha_2_99/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_287/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_298 sky130_fd_sc_hd__fa_2_258/A sky130_fd_sc_hd__ha_2_91/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_298/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_6 sky130_fd_sc_hd__nor4_1_2/A sky130_fd_sc_hd__o21ai_1_9/Y
+ sky130_fd_sc_hd__nor4_1_1/D sky130_fd_sc_hd__o21ai_1_9/A2 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__clkbuf_4_19 sky130_fd_sc_hd__clkbuf_4_19/X sky130_fd_sc_hd__clkbuf_4_19/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__a21oi_1_140 sky130_fd_sc_hd__nor2_2_10/Y sky130_fd_sc_hd__o22ai_1_140/Y
+ sky130_fd_sc_hd__a21oi_1_140/Y sky130_fd_sc_hd__fa_2_1112/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_151 sky130_fd_sc_hd__nor2_2_11/Y sky130_fd_sc_hd__o22ai_1_150/Y
+ sky130_fd_sc_hd__a21oi_1_151/Y sky130_fd_sc_hd__fa_2_1108/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_162 sky130_fd_sc_hd__nor2_2_11/Y sky130_fd_sc_hd__o22ai_1_161/Y
+ sky130_fd_sc_hd__a21oi_1_162/Y sky130_fd_sc_hd__fa_2_1119/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_173 sky130_fd_sc_hd__nand2_1_307/Y sky130_fd_sc_hd__nor2_1_99/Y
+ sky130_fd_sc_hd__xnor2_1_88/A sky130_fd_sc_hd__xnor2_1_86/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_184 sky130_fd_sc_hd__nor2_1_117/A sky130_fd_sc_hd__o21a_1_13/A1
+ sky130_fd_sc_hd__dfxtp_1_758/D sky130_fd_sc_hd__nor2_1_117/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_195 sky130_fd_sc_hd__a211o_1_9/A1 sky130_fd_sc_hd__o21ai_1_222/Y
+ sky130_fd_sc_hd__a21oi_1_195/Y sky130_fd_sc_hd__clkinv_1_698/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_103 sky130_fd_sc_hd__buf_8_103/A sky130_fd_sc_hd__buf_8_103/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_114 sky130_fd_sc_hd__buf_8_91/X sky130_fd_sc_hd__buf_6_25/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_125 sky130_fd_sc_hd__buf_8_125/A sky130_fd_sc_hd__buf_8_125/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_136 sky130_fd_sc_hd__buf_8_136/A sky130_fd_sc_hd__buf_8_136/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_147 sky130_fd_sc_hd__buf_8_147/A sky130_fd_sc_hd__buf_4_89/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_158 sky130_fd_sc_hd__buf_8_158/A sky130_fd_sc_hd__buf_8_158/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nor2_4_9 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__or2_0_5/A
+ sky130_fd_sc_hd__nor2_4_9/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_4
Xsky130_fd_sc_hd__buf_8_169 sky130_fd_sc_hd__buf_8_169/A sky130_fd_sc_hd__buf_6_47/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__a21o_2_15 sky130_fd_sc_hd__a21o_2_15/X sky130_fd_sc_hd__nor2_1_211/Y
+ sky130_fd_sc_hd__nor2_1_211/A sky130_fd_sc_hd__nor2_1_211/B VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__a21o_2_26 sky130_fd_sc_hd__a21o_2_26/X sky130_fd_sc_hd__nor2_1_295/Y
+ sky130_fd_sc_hd__fa_2_0/SUM sky130_fd_sc_hd__nor2_1_295/B VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__xor2_1_20 sky130_fd_sc_hd__xor2_1_20/B sky130_fd_sc_hd__nor4_1_3/A
+ sky130_fd_sc_hd__ha_2_151/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_31 sky130_fd_sc_hd__xor2_1_31/B sky130_fd_sc_hd__xor2_1_31/X
+ sky130_fd_sc_hd__xor2_1_31/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_42 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_985/B
+ sky130_fd_sc_hd__xor2_1_42/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_53 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_974/B
+ sky130_fd_sc_hd__xor2_1_53/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_64 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__xor2_1_64/X
+ sky130_fd_sc_hd__xor2_1_64/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_75 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__xor2_1_75/X
+ sky130_fd_sc_hd__xor2_1_75/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_86 sky130_fd_sc_hd__xor2_1_86/B sky130_fd_sc_hd__xor2_1_86/X
+ sky130_fd_sc_hd__xor2_1_87/X VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_97 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__xor2_1_97/X
+ sky130_fd_sc_hd__xor2_1_97/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2b_1_3 sky130_fd_sc_hd__nand2b_1_3/Y sky130_fd_sc_hd__xor2_1_14/A
+ sky130_fd_sc_hd__xor2_1_14/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__dfxtp_1_1308 VDD VSS sky130_fd_sc_hd__fa_2_843/B sky130_fd_sc_hd__dfxtp_1_1322/CLK
+ sky130_fd_sc_hd__a21oi_1_432/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1319 VDD VSS sky130_fd_sc_hd__fa_2_903/A sky130_fd_sc_hd__dfxtp_1_1326/CLK
+ sky130_fd_sc_hd__a21oi_1_427/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_902 VDD VSS sky130_fd_sc_hd__fa_2_937/B sky130_fd_sc_hd__dfxtp_1_902/CLK
+ sky130_fd_sc_hd__o21a_1_20/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_913 VDD VSS sky130_fd_sc_hd__fa_2_1142/A sky130_fd_sc_hd__clkinv_8_55/Y
+ sky130_fd_sc_hd__mux2_2_116/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_924 VDD VSS sky130_fd_sc_hd__fa_2_1153/A sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__mux2_2_86/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_935 VDD VSS sky130_fd_sc_hd__fa_2_1127/A sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__mux2_2_108/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_946 VDD VSS sky130_fd_sc_hd__fa_2_1138/A sky130_fd_sc_hd__clkinv_8_46/Y
+ sky130_fd_sc_hd__mux2_2_81/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_957 VDD VSS sky130_fd_sc_hd__fa_2_1166/A sky130_fd_sc_hd__clkinv_8_65/Y
+ sky130_fd_sc_hd__mux2_2_109/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a221oi_1_1 sky130_fd_sc_hd__nand4_1_83/A sky130_fd_sc_hd__o22ai_1_57/Y
+ sky130_fd_sc_hd__nor4_1_4/C sky130_fd_sc_hd__ha_2_157/B sky130_fd_sc_hd__ha_2_157/A
+ sky130_fd_sc_hd__o22ai_1_57/B2 VSS VDD VDD VSS sky130_fd_sc_hd__a221oi_1
Xsky130_fd_sc_hd__dfxtp_1_968 VDD VSS sky130_fd_sc_hd__nor2_4_15/A sky130_fd_sc_hd__clkinv_8_46/Y
+ sky130_fd_sc_hd__nor2b_1_110/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_979 VDD VSS sky130_fd_sc_hd__mux2_2_94/A0 sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__o22ai_1_216/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_500 VSS VDD sky130_fd_sc_hd__nand4_1_57/B sky130_fd_sc_hd__a22oi_1_237/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_511 VSS VDD sky130_fd_sc_hd__buf_2_165/A sky130_fd_sc_hd__nor3_2_9/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_522 VSS VDD sky130_fd_sc_hd__buf_2_148/A sky130_fd_sc_hd__clkbuf_8_3/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_533 VSS VDD sky130_fd_sc_hd__clkbuf_1_533/X sky130_fd_sc_hd__clkbuf_1_533/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_101 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_93/A sky130_fd_sc_hd__fa_2_194/B
+ sky130_fd_sc_hd__fa_2_190/A sky130_fd_sc_hd__fa_2_2/A sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_544 VSS VDD sky130_fd_sc_hd__fa_2_71/A sky130_fd_sc_hd__ha_2_99/B
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_112 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_112/A sky130_fd_sc_hd__fa_2_361/A
+ sky130_fd_sc_hd__ha_2_112/SUM sky130_fd_sc_hd__ha_2_112/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_555 VSS VDD sky130_fd_sc_hd__fa_2_31/A sky130_fd_sc_hd__ha_2_94/B
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_123 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_123/A sky130_fd_sc_hd__fa_2_531/CIN
+ sky130_fd_sc_hd__fa_2_523/A sky130_fd_sc_hd__ha_2_123/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_566 VSS VDD sky130_fd_sc_hd__buf_4_62/A sky130_fd_sc_hd__dfxtp_1_1456/Q
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_134 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_134/A sky130_fd_sc_hd__fa_2_694/A
+ sky130_fd_sc_hd__ha_2_134/SUM sky130_fd_sc_hd__ha_2_134/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_577 VSS VDD sky130_fd_sc_hd__nand3_1_13/B sky130_fd_sc_hd__a22oi_1_25/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_145 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_145/A sky130_fd_sc_hd__fa_2_834/CIN
+ sky130_fd_sc_hd__fa_2_832/B sky130_fd_sc_hd__ha_2_145/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_588 VSS VDD sky130_fd_sc_hd__nand3_1_4/B sky130_fd_sc_hd__a22oi_1_8/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_156 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_156/A sky130_fd_sc_hd__ha_2_155/B
+ sky130_fd_sc_hd__ha_2_156/SUM sky130_fd_sc_hd__ha_2_156/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_599 VSS VDD sky130_fd_sc_hd__dfxtp_1_62/D sky130_fd_sc_hd__nand4_1_32/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_807 sky130_fd_sc_hd__fa_2_808/B sky130_fd_sc_hd__fa_2_800/A
+ sky130_fd_sc_hd__fa_2_834/A sky130_fd_sc_hd__fa_2_807/B sky130_fd_sc_hd__fa_2_835/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_167 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_9/B sky130_fd_sc_hd__ha_2_166/B
+ sky130_fd_sc_hd__ha_2_167/SUM sky130_fd_sc_hd__ha_2_167/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_818 sky130_fd_sc_hd__fa_2_710/A sky130_fd_sc_hd__fa_2_711/B
+ sky130_fd_sc_hd__fa_2_818/A sky130_fd_sc_hd__fa_2_818/B sky130_fd_sc_hd__fa_2_822/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_178 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_178/A sky130_fd_sc_hd__ha_2_177/A
+ sky130_fd_sc_hd__ha_2_178/SUM sky130_fd_sc_hd__ha_2_178/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_829 sky130_fd_sc_hd__fa_2_828/CIN sky130_fd_sc_hd__fa_2_829/SUM
+ sky130_fd_sc_hd__fa_2_829/A sky130_fd_sc_hd__fa_2_832/A sky130_fd_sc_hd__ha_2_144/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_189 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_189/A sky130_fd_sc_hd__ha_2_188/A
+ sky130_fd_sc_hd__ha_2_189/SUM sky130_fd_sc_hd__ha_2_189/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__maj3_1_5 sky130_fd_sc_hd__maj3_1_6/X sky130_fd_sc_hd__maj3_1_5/X
+ sky130_fd_sc_hd__maj3_1_5/B sky130_fd_sc_hd__maj3_1_5/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__ha_2_80 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_80/A sky130_fd_sc_hd__xor2_1_8/A
+ sky130_fd_sc_hd__ha_2_80/SUM sky130_fd_sc_hd__ha_2_80/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_91 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_91/A sky130_fd_sc_hd__fa_2_49/CIN
+ sky130_fd_sc_hd__fa_2_45/B sky130_fd_sc_hd__ha_2_91/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__mux2_2_107 VSS VDD sky130_fd_sc_hd__mux2_2_107/A1 sky130_fd_sc_hd__mux2_2_107/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_107/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_118 VSS VDD sky130_fd_sc_hd__mux2_2_118/A1 sky130_fd_sc_hd__mux2_2_118/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_118/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_129 VSS VDD sky130_fd_sc_hd__mux2_2_129/A1 sky130_fd_sc_hd__mux2_2_129/A0
+ sky130_fd_sc_hd__mux2_2_135/S sky130_fd_sc_hd__mux2_2_129/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__and2_0_14 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_14/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_12/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_25 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_25/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_30/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_305 sky130_fd_sc_hd__o22ai_1_318/A2 sky130_fd_sc_hd__nor2_1_187/B
+ sky130_fd_sc_hd__o22ai_1_305/Y sky130_fd_sc_hd__nor2_1_188/B sky130_fd_sc_hd__o32ai_1_5/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_36 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_36/X sky130_fd_sc_hd__ha_2_54/A
+ sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_316 sky130_fd_sc_hd__o22ai_1_318/A2 sky130_fd_sc_hd__o22ai_1_316/B1
+ sky130_fd_sc_hd__o22ai_1_316/Y sky130_fd_sc_hd__nor2_1_192/B sky130_fd_sc_hd__o32ai_1_5/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_47 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_52/A sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__ha_2_58/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_327 sky130_fd_sc_hd__nand2_1_462/Y sky130_fd_sc_hd__nand2_1_461/Y
+ sky130_fd_sc_hd__o22ai_1_327/Y sky130_fd_sc_hd__o22ai_1_340/A1 sky130_fd_sc_hd__a21o_2_19/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_58 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_58/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_58/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_338 sky130_fd_sc_hd__nand2_1_464/Y sky130_fd_sc_hd__nand2_1_463/Y
+ sky130_fd_sc_hd__o22ai_1_338/Y sky130_fd_sc_hd__o22ai_1_338/A1 sky130_fd_sc_hd__a21o_2_18/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_69 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_76/A sky130_fd_sc_hd__nor2_4_0/Y
+ sky130_fd_sc_hd__ha_2_76/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_349 sky130_fd_sc_hd__nand2_1_464/Y sky130_fd_sc_hd__nand2_1_463/Y
+ sky130_fd_sc_hd__o22ai_1_349/Y sky130_fd_sc_hd__o22ai_1_349/A1 sky130_fd_sc_hd__o21ai_1_391/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_2_6 sky130_fd_sc_hd__nor2_2_6/B sky130_fd_sc_hd__nor2_2_6/Y
+ sky130_fd_sc_hd__nor2_2_6/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__buf_8_13 sky130_fd_sc_hd__buf_8_13/A sky130_fd_sc_hd__buf_8_13/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_24 sky130_fd_sc_hd__inv_2_25/Y sky130_fd_sc_hd__buf_8_24/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_35 sky130_fd_sc_hd__buf_8_35/A sky130_fd_sc_hd__buf_8_35/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_46 sky130_fd_sc_hd__inv_2_42/Y sky130_fd_sc_hd__buf_8_46/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_57 sky130_fd_sc_hd__inv_2_43/A sky130_fd_sc_hd__buf_8_57/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_68 sky130_fd_sc_hd__buf_8_68/A sky130_fd_sc_hd__buf_8_68/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_79 sky130_fd_sc_hd__ha_2_31/A sky130_fd_sc_hd__buf_8_79/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__dfxtp_1_209 VDD VSS sky130_fd_sc_hd__ha_2_72/A sky130_fd_sc_hd__dfxtp_1_212/CLK
+ sky130_fd_sc_hd__and2_0_79/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_2_109 VDD VSS sky130_fd_sc_hd__buf_2_109/X sky130_fd_sc_hd__buf_2_109/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__fa_2_1308 sky130_fd_sc_hd__fa_2_1309/CIN sky130_fd_sc_hd__mux2_2_226/A0
+ sky130_fd_sc_hd__fa_2_1308/A sky130_fd_sc_hd__fa_2_1308/B sky130_fd_sc_hd__fa_2_1308/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1319 sky130_fd_sc_hd__fa_2_1320/CIN sky130_fd_sc_hd__mux2_2_253/A1
+ sky130_fd_sc_hd__fa_2_1319/A sky130_fd_sc_hd__nor2_8_2/Y sky130_fd_sc_hd__fa_2_1319/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1105 VDD VSS sky130_fd_sc_hd__nor2_8_0/B sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__mux2_2_140/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1116 VDD VSS sky130_fd_sc_hd__mux2_2_153/A0 sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__o22ai_1_277/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1127 VDD VSS sky130_fd_sc_hd__mux2_2_127/A1 sky130_fd_sc_hd__clkinv_8_70/Y
+ sky130_fd_sc_hd__o31ai_1_8/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1138 VDD VSS sky130_fd_sc_hd__mux2_2_154/A0 sky130_fd_sc_hd__clkinv_8_65/Y
+ sky130_fd_sc_hd__dfxtp_1_997/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_710 VDD VSS sky130_fd_sc_hd__mux2_2_13/A1 sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__o21ai_1_50/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1149 VDD VSS sky130_fd_sc_hd__mux2_2_146/A0 sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__o22ai_1_288/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_721 VDD VSS sky130_fd_sc_hd__mux2_2_32/A0 sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__o21ai_1_58/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_732 VDD VSS sky130_fd_sc_hd__mux2_2_8/A1 sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__o21ai_1_69/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_743 VDD VSS sky130_fd_sc_hd__and2_0_170/A sky130_fd_sc_hd__dfxtp_1_744/CLK
+ sky130_fd_sc_hd__fa_2_1098/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_754 VDD VSS sky130_fd_sc_hd__fa_2_673/B sky130_fd_sc_hd__dfxtp_1_755/CLK
+ sky130_fd_sc_hd__o21a_1_15/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_765 VDD VSS sky130_fd_sc_hd__fa_2_700/A sky130_fd_sc_hd__dfxtp_1_768/CLK
+ sky130_fd_sc_hd__o21a_1_10/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_776 VDD VSS sky130_fd_sc_hd__fa_2_1075/A sky130_fd_sc_hd__clkinv_8_55/Y
+ sky130_fd_sc_hd__mux2_2_74/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__ha_2_9 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_9/A sky130_fd_sc_hd__ha_2_8/B
+ sky130_fd_sc_hd__ha_2_9/SUM sky130_fd_sc_hd__ha_2_9/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__dfxtp_1_787 VDD VSS sky130_fd_sc_hd__fa_2_1086/A sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__mux2_2_50/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_798 VDD VSS sky130_fd_sc_hd__fa_2_1050/A sky130_fd_sc_hd__clkinv_8_54/Y
+ sky130_fd_sc_hd__and2_0_313/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_330 VSS VDD sky130_fd_sc_hd__buf_8_159/A sky130_fd_sc_hd__and2_1_1/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_341 VSS VDD sky130_fd_sc_hd__buf_8_161/A sky130_fd_sc_hd__and2_1_6/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_352 VSS VDD sky130_fd_sc_hd__clkinv_1_174/A sky130_fd_sc_hd__clkinv_4_15/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_363 VSS VDD sky130_fd_sc_hd__clkbuf_1_363/X sky130_fd_sc_hd__buf_4_70/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_374 VSS VDD sky130_fd_sc_hd__clkbuf_1_374/X sky130_fd_sc_hd__nand3_1_40/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_385 VSS VDD sky130_fd_sc_hd__clkbuf_1_385/X sky130_fd_sc_hd__inv_2_135/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_396 VSS VDD sky130_fd_sc_hd__a22oi_2_14/B2 sky130_fd_sc_hd__clkbuf_1_396/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_604 sky130_fd_sc_hd__maj3_1_122/B sky130_fd_sc_hd__maj3_1_123/A
+ sky130_fd_sc_hd__fa_2_604/A sky130_fd_sc_hd__fa_2_604/B sky130_fd_sc_hd__fa_2_605/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_615 sky130_fd_sc_hd__fa_2_618/B sky130_fd_sc_hd__fa_2_615/SUM
+ sky130_fd_sc_hd__fa_2_615/A sky130_fd_sc_hd__fa_2_615/B sky130_fd_sc_hd__o22ai_1_42/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_626 sky130_fd_sc_hd__maj3_1_116/B sky130_fd_sc_hd__maj3_1_117/A
+ sky130_fd_sc_hd__fa_2_626/A sky130_fd_sc_hd__fa_2_626/B sky130_fd_sc_hd__fa_2_627/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_637 sky130_fd_sc_hd__fa_2_639/B sky130_fd_sc_hd__fa_2_633/A
+ sky130_fd_sc_hd__fa_2_698/A sky130_fd_sc_hd__ha_2_126/A sky130_fd_sc_hd__fa_2_692/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_648 sky130_fd_sc_hd__fa_2_650/B sky130_fd_sc_hd__fa_2_645/A
+ sky130_fd_sc_hd__fa_2_698/A sky130_fd_sc_hd__ha_2_126/A sky130_fd_sc_hd__ha_2_128/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_659 sky130_fd_sc_hd__fa_2_658/CIN sky130_fd_sc_hd__fa_2_659/SUM
+ sky130_fd_sc_hd__fa_2_659/A sky130_fd_sc_hd__fa_2_667/B sky130_fd_sc_hd__ha_2_135/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_350 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_350/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_350/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_190 sky130_fd_sc_hd__clkbuf_4_190/X sky130_fd_sc_hd__clkbuf_4_190/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__conb_1_3 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__conb_1_3/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__buf_12_9 sky130_fd_sc_hd__inv_2_34/Y sky130_fd_sc_hd__buf_12_9/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__o22ai_1_102 sky130_fd_sc_hd__o21a_1_8/A2 sky130_fd_sc_hd__o22ai_1_116/A1
+ sky130_fd_sc_hd__nor2_1_79/B sky130_fd_sc_hd__nor2_1_66/B sky130_fd_sc_hd__o21ai_1_92/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_113 sky130_fd_sc_hd__nand4_1_85/B sky130_fd_sc_hd__o21ai_1_92/A1
+ sky130_fd_sc_hd__o22ai_1_113/Y sky130_fd_sc_hd__o22ai_1_132/B1 sky130_fd_sc_hd__o22ai_1_121/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_124 sky130_fd_sc_hd__nor2_1_77/A sky130_fd_sc_hd__nor2_2_9/B
+ sky130_fd_sc_hd__o22ai_1_124/Y sky130_fd_sc_hd__a21oi_1_127/Y sky130_fd_sc_hd__a222oi_1_1/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_135 sky130_fd_sc_hd__nand2_1_284/Y sky130_fd_sc_hd__nand2_2_5/Y
+ sky130_fd_sc_hd__o22ai_1_135/Y sky130_fd_sc_hd__xnor2_1_62/Y sky130_fd_sc_hd__o22ai_1_149/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_146 sky130_fd_sc_hd__nand2_1_284/Y sky130_fd_sc_hd__nand2_2_5/Y
+ sky130_fd_sc_hd__o22ai_1_146/Y sky130_fd_sc_hd__xnor2_1_84/Y sky130_fd_sc_hd__o22ai_1_160/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_157 sky130_fd_sc_hd__nand2_1_338/A sky130_fd_sc_hd__nand2_1_284/Y
+ sky130_fd_sc_hd__o22ai_1_157/Y sky130_fd_sc_hd__xnor2_1_78/Y sky130_fd_sc_hd__o22ai_1_157/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_809 sky130_fd_sc_hd__o32ai_1_0/B2 sky130_fd_sc_hd__fa_2_1124/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_809/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_2_13 sky130_fd_sc_hd__nor2_2_13/B sky130_fd_sc_hd__or2_0_8/B
+ sky130_fd_sc_hd__nor2_2_13/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__o22ai_1_168 sky130_fd_sc_hd__nor2_2_13/B sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__o22ai_1_168/Y sky130_fd_sc_hd__a21oi_1_202/Y sky130_fd_sc_hd__nor2_1_133/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_179 sky130_fd_sc_hd__o22ai_1_204/B1 sky130_fd_sc_hd__nor2_1_115/B
+ sky130_fd_sc_hd__nor2_1_130/A sky130_fd_sc_hd__o22ai_1_190/A1 sky130_fd_sc_hd__o22ai_1_206/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand4_1_16 sky130_fd_sc_hd__nand4_1_16/C sky130_fd_sc_hd__nand4_1_16/B
+ sky130_fd_sc_hd__nand4_1_16/Y sky130_fd_sc_hd__nand4_1_16/D sky130_fd_sc_hd__buf_2_112/X
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__o211ai_1_3 sky130_fd_sc_hd__a31oi_1_1/Y sky130_fd_sc_hd__nand4_1_84/Y
+ sky130_fd_sc_hd__nor4_1_9/D sky130_fd_sc_hd__nor4_1_10/Y sky130_fd_sc_hd__a21oi_1_20/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__nand4_1_27 sky130_fd_sc_hd__nand4_1_27/C sky130_fd_sc_hd__nand4_1_27/B
+ sky130_fd_sc_hd__nand4_1_27/Y sky130_fd_sc_hd__nand4_1_27/D sky130_fd_sc_hd__buf_2_104/X
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_38 sky130_fd_sc_hd__nand4_1_38/C sky130_fd_sc_hd__nand4_1_38/B
+ sky130_fd_sc_hd__nand4_1_38/Y sky130_fd_sc_hd__nand4_1_38/D sky130_fd_sc_hd__nand4_1_38/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_49 sky130_fd_sc_hd__nand4_1_49/C sky130_fd_sc_hd__nand4_1_49/B
+ sky130_fd_sc_hd__nand4_1_49/Y sky130_fd_sc_hd__nand4_1_49/D sky130_fd_sc_hd__nand4_1_49/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__a31oi_1_0 VSS VDD sky130_fd_sc_hd__a31oi_1_0/Y sky130_fd_sc_hd__or2_0_0/B
+ sky130_fd_sc_hd__o21ai_1_2/Y sky130_fd_sc_hd__nor3_1_4/A sky130_fd_sc_hd__nand3_1_16/Y
+ VDD VSS sky130_fd_sc_hd__a31oi_1
Xsky130_fd_sc_hd__o21ai_1_340 VSS VDD sky130_fd_sc_hd__nor2_1_190/B sky130_fd_sc_hd__o22ai_1_322/A2
+ sky130_fd_sc_hd__a22oi_1_380/Y sky130_fd_sc_hd__o21ai_1_340/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_351 VSS VDD sky130_fd_sc_hd__o21ai_1_360/A1 sky130_fd_sc_hd__nor2_1_222/A
+ sky130_fd_sc_hd__a21oi_1_331/Y sky130_fd_sc_hd__xor2_1_222/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a211oi_1_12 sky130_fd_sc_hd__nor2b_1_105/Y sky130_fd_sc_hd__o21ai_1_303/Y
+ sky130_fd_sc_hd__nor2_1_174/Y sky130_fd_sc_hd__a211oi_1_12/Y sky130_fd_sc_hd__o21ai_1_305/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_362 VSS VDD sky130_fd_sc_hd__nor2_1_186/B sky130_fd_sc_hd__o21a_1_42/A1
+ sky130_fd_sc_hd__a21oi_1_340/Y sky130_fd_sc_hd__o21ai_1_362/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a211oi_1_23 sky130_fd_sc_hd__nor3_1_39/A sky130_fd_sc_hd__nor2_1_223/Y
+ sky130_fd_sc_hd__o22ai_1_316/Y sky130_fd_sc_hd__a211oi_1_23/Y sky130_fd_sc_hd__fa_2_1205/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_373 VSS VDD sky130_fd_sc_hd__a211oi_1_23/Y sky130_fd_sc_hd__nor2_1_214/A
+ sky130_fd_sc_hd__a21oi_1_348/Y sky130_fd_sc_hd__o21ai_1_373/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a211oi_1_34 sky130_fd_sc_hd__nor2b_2_5/Y sky130_fd_sc_hd__o22ai_1_420/Y
+ sky130_fd_sc_hd__nor2_1_302/Y sky130_fd_sc_hd__a211oi_1_34/Y sky130_fd_sc_hd__o21ai_1_469/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_384 VSS VDD sky130_fd_sc_hd__nor2_1_246/Y sky130_fd_sc_hd__or3_1_4/C
+ sky130_fd_sc_hd__xnor2_1_99/Y sky130_fd_sc_hd__o21ai_1_384/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_395 VSS VDD sky130_fd_sc_hd__xor2_1_230/X sky130_fd_sc_hd__xnor2_1_1/Y
+ sky130_fd_sc_hd__xnor2_1_99/Y sky130_fd_sc_hd__o21ai_1_395/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__mux2_2_20 VSS VDD sky130_fd_sc_hd__mux2_2_20/A1 sky130_fd_sc_hd__mux2_2_20/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_20/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_31 VSS VDD sky130_fd_sc_hd__mux2_2_31/A1 sky130_fd_sc_hd__mux2_2_31/A0
+ sky130_fd_sc_hd__mux2_2_37/S sky130_fd_sc_hd__mux2_2_31/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_42 VSS VDD sky130_fd_sc_hd__mux2_2_42/A1 sky130_fd_sc_hd__mux2_2_42/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_42/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_53 VSS VDD sky130_fd_sc_hd__mux2_2_53/A1 sky130_fd_sc_hd__mux2_2_53/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_53/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_64 VSS VDD sky130_fd_sc_hd__mux2_2_64/A1 sky130_fd_sc_hd__mux2_2_64/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_64/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_75 VSS VDD sky130_fd_sc_hd__mux2_2_75/A1 sky130_fd_sc_hd__mux2_2_75/A0
+ sky130_fd_sc_hd__mux2_2_75/S sky130_fd_sc_hd__mux2_2_75/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_86 VSS VDD sky130_fd_sc_hd__mux2_2_86/A1 sky130_fd_sc_hd__mux2_2_86/A0
+ sky130_fd_sc_hd__nor2_4_15/A sky130_fd_sc_hd__mux2_2_86/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1105 sky130_fd_sc_hd__fa_2_1106/CIN sky130_fd_sc_hd__or2_0_7/B
+ sky130_fd_sc_hd__fa_2_1105/A sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1105/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__mux2_2_97 VSS VDD sky130_fd_sc_hd__mux2_2_97/A1 sky130_fd_sc_hd__mux2_2_97/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_97/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1116 sky130_fd_sc_hd__fa_2_1117/CIN sky130_fd_sc_hd__fa_2_1116/SUM
+ sky130_fd_sc_hd__fa_2_1116/A sky130_fd_sc_hd__fa_2_1116/B sky130_fd_sc_hd__fa_2_1116/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1127 sky130_fd_sc_hd__fa_2_1128/CIN sky130_fd_sc_hd__mux2_2_108/A1
+ sky130_fd_sc_hd__fa_2_1127/A sky130_fd_sc_hd__fa_2_1127/B sky130_fd_sc_hd__fa_2_1127/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1138 sky130_fd_sc_hd__fa_2_1139/CIN sky130_fd_sc_hd__mux2_2_81/A0
+ sky130_fd_sc_hd__fa_2_1138/A sky130_fd_sc_hd__fa_2_1138/B sky130_fd_sc_hd__fa_2_1138/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1149 sky130_fd_sc_hd__fa_2_1150/CIN sky130_fd_sc_hd__mux2_2_95/A1
+ sky130_fd_sc_hd__fa_2_1149/A sky130_fd_sc_hd__fa_2_1149/B sky130_fd_sc_hd__fa_2_1149/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_540 VDD VSS sky130_fd_sc_hd__fa_2_951/A sky130_fd_sc_hd__dfxtp_1_544/CLK
+ sky130_fd_sc_hd__a22o_1_45/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_551 VDD VSS sky130_fd_sc_hd__and2_0_183/A sky130_fd_sc_hd__dfxtp_1_571/CLK
+ sky130_fd_sc_hd__dfxtp_1_552/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_562 VDD VSS sky130_fd_sc_hd__dfxtp_1_562/Q sky130_fd_sc_hd__dfxtp_1_576/CLK
+ sky130_fd_sc_hd__dfxtp_1_562/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_573 VDD VSS sky130_fd_sc_hd__and2_0_202/A sky130_fd_sc_hd__dfxtp_1_577/CLK
+ sky130_fd_sc_hd__a22o_1_36/B1 VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_584 VDD VSS sky130_fd_sc_hd__nor4_1_6/B sky130_fd_sc_hd__dfxtp_1_594/CLK
+ sky130_fd_sc_hd__and2_0_251/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_595 VDD VSS sky130_fd_sc_hd__or4_1_2/C sky130_fd_sc_hd__dfxtp_1_595/CLK
+ sky130_fd_sc_hd__nor2_1_29/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_160 VSS VDD sky130_fd_sc_hd__clkbuf_1_160/X sky130_fd_sc_hd__clkbuf_1_160/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_171 VSS VDD sky130_fd_sc_hd__a22oi_1_90/A2 sky130_fd_sc_hd__clkbuf_1_171/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_182 VSS VDD sky130_fd_sc_hd__nand4_1_24/B sky130_fd_sc_hd__a22oi_1_118/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_193 VSS VDD sky130_fd_sc_hd__buf_12_127/A sky130_fd_sc_hd__clkbuf_1_193/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_401 sky130_fd_sc_hd__fa_2_403/CIN sky130_fd_sc_hd__fa_2_396/A
+ sky130_fd_sc_hd__fa_2_401/A sky130_fd_sc_hd__fa_2_401/B sky130_fd_sc_hd__fa_2_401/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_412 sky130_fd_sc_hd__fa_2_413/CIN sky130_fd_sc_hd__fa_2_407/A
+ sky130_fd_sc_hd__fa_2_412/A sky130_fd_sc_hd__fa_2_425/A sky130_fd_sc_hd__fa_2_401/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_423 sky130_fd_sc_hd__fa_2_321/B sky130_fd_sc_hd__fa_2_423/SUM
+ sky130_fd_sc_hd__fa_2_423/A sky130_fd_sc_hd__fa_2_423/B sky130_fd_sc_hd__fa_2_423/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_434 sky130_fd_sc_hd__fa_2_431/CIN sky130_fd_sc_hd__fa_2_434/SUM
+ sky130_fd_sc_hd__fa_2_434/A sky130_fd_sc_hd__fa_2_434/B sky130_fd_sc_hd__fa_2_434/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_445 sky130_fd_sc_hd__fa_2_442/CIN sky130_fd_sc_hd__nor2_1_170/A
+ sky130_fd_sc_hd__fa_2_445/A sky130_fd_sc_hd__fa_2_445/B sky130_fd_sc_hd__fa_2_445/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_456 sky130_fd_sc_hd__fa_2_452/CIN sky130_fd_sc_hd__or3_1_2/A
+ sky130_fd_sc_hd__fa_2_456/A sky130_fd_sc_hd__fa_2_456/B sky130_fd_sc_hd__fa_2_456/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_467 sky130_fd_sc_hd__fa_2_468/CIN sky130_fd_sc_hd__maj3_1_106/A
+ sky130_fd_sc_hd__ha_2_123/A sky130_fd_sc_hd__ha_2_121/B sky130_fd_sc_hd__ha_2_122/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_478 sky130_fd_sc_hd__fa_2_480/CIN sky130_fd_sc_hd__fa_2_476/A
+ sky130_fd_sc_hd__ha_2_125/B sky130_fd_sc_hd__ha_2_123/B sky130_fd_sc_hd__fa_2_567/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_489 sky130_fd_sc_hd__maj3_1_96/B sky130_fd_sc_hd__maj3_1_97/A
+ sky130_fd_sc_hd__fa_2_489/A sky130_fd_sc_hd__fa_2_489/B sky130_fd_sc_hd__fa_2_490/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_180 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_180/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_180/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_191 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_191/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__ha_2_161/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_406 sky130_fd_sc_hd__buf_8_186/X sky130_fd_sc_hd__buf_12_461/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_417 sky130_fd_sc_hd__buf_8_180/X sky130_fd_sc_hd__buf_12_514/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_428 sky130_fd_sc_hd__buf_8_184/X sky130_fd_sc_hd__buf_12_428/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_439 sky130_fd_sc_hd__buf_2_246/X sky130_fd_sc_hd__buf_12_439/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_309 sky130_fd_sc_hd__clkbuf_4_165/X sky130_fd_sc_hd__clkinv_2_23/Y
+ sky130_fd_sc_hd__clkbuf_1_400/X sky130_fd_sc_hd__a22oi_1_309/A2 sky130_fd_sc_hd__a22oi_1_309/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__fa_2_990 sky130_fd_sc_hd__fa_2_991/CIN sky130_fd_sc_hd__mux2_2_7/A0
+ sky130_fd_sc_hd__fa_2_990/A sky130_fd_sc_hd__fa_2_990/B sky130_fd_sc_hd__fa_2_990/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_1_606 sky130_fd_sc_hd__ha_2_182/B sky130_fd_sc_hd__fa_2_1033/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_606/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_617 sky130_fd_sc_hd__nor2_2_6/B sky130_fd_sc_hd__nor2_1_41/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_617/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_628 sky130_fd_sc_hd__nand2_1_338/A sky130_fd_sc_hd__nor2_2_10/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_628/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_639 sky130_fd_sc_hd__o22ai_1_157/B2 sky130_fd_sc_hd__ha_2_192/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_639/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_170 VSS VDD sky130_fd_sc_hd__o21ai_1_171/A2 sky130_fd_sc_hd__xnor2_1_87/Y
+ sky130_fd_sc_hd__a21oi_1_147/Y sky130_fd_sc_hd__o21ai_1_170/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_181 VSS VDD sky130_fd_sc_hd__nand2_2_5/Y sky130_fd_sc_hd__xnor2_1_75/Y
+ sky130_fd_sc_hd__a21oi_1_156/Y sky130_fd_sc_hd__o21ai_1_181/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_192 VSS VDD sky130_fd_sc_hd__xnor2_1_89/A sky130_fd_sc_hd__o21ai_1_192/A1
+ sky130_fd_sc_hd__nand2_1_293/B sky130_fd_sc_hd__a22o_1_72/B2 VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_15 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1174/A sky130_fd_sc_hd__nor2_2_16/Y
+ sky130_fd_sc_hd__nor3_1_39/A sky130_fd_sc_hd__fa_2_1176/A sky130_fd_sc_hd__nor3_1_39/B
+ sky130_fd_sc_hd__a222oi_1_15/Y sky130_fd_sc_hd__fa_2_1173/B sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_26 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1241/A sky130_fd_sc_hd__nor2_2_17/Y
+ sky130_fd_sc_hd__nor3_1_40/A sky130_fd_sc_hd__nor2_4_18/B sky130_fd_sc_hd__xor2_1_254/A
+ sky130_fd_sc_hd__a222oi_1_26/Y sky130_fd_sc_hd__fa_2_1240/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_37 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1279/A sky130_fd_sc_hd__nor2_2_18/Y
+ sky130_fd_sc_hd__nor3_1_41/A sky130_fd_sc_hd__fa_2_1281/A sky130_fd_sc_hd__nor3_1_41/B
+ sky130_fd_sc_hd__a222oi_1_37/Y sky130_fd_sc_hd__fa_2_1278/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2_1_530 sky130_fd_sc_hd__nand2_1_530/Y sky130_fd_sc_hd__nand2_1_543/B
+ sky130_fd_sc_hd__o21ai_1_463/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_17 VSS VDD sky130_fd_sc_hd__maj3_1_2/A sky130_fd_sc_hd__xnor2_1_17/Y
+ sky130_fd_sc_hd__ha_2_154/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_541 sky130_fd_sc_hd__nand2_1_541/Y sky130_fd_sc_hd__nand2_1_543/B
+ sky130_fd_sc_hd__o21ai_1_488/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_28 VSS VDD sky130_fd_sc_hd__xnor2_1_28/B sky130_fd_sc_hd__xnor2_1_28/Y
+ sky130_fd_sc_hd__nor4_1_7/B VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_552 sky130_fd_sc_hd__nor4_1_13/A sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__dfxtp_1_82/Q VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_39 VSS VDD sky130_fd_sc_hd__xnor2_1_40/B sky130_fd_sc_hd__xnor2_1_39/Y
+ sky130_fd_sc_hd__xnor2_1_39/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_563 sky130_fd_sc_hd__nand2_1_563/Y sky130_fd_sc_hd__buf_4_122/A
+ sky130_fd_sc_hd__nand2_1_563/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_1110 sky130_fd_sc_hd__o31ai_1_0/A3 sky130_fd_sc_hd__nor4_1_4/C
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1110/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1121 sky130_fd_sc_hd__nor2_1_322/A sky130_fd_sc_hd__nor2_1_318/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1121/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1132 sky130_fd_sc_hd__clkinv_4_41/A sky130_fd_sc_hd__nand2_1_567/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1132/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_370 VDD VSS sky130_fd_sc_hd__fa_2_1114/A sky130_fd_sc_hd__clkinv_4_32/Y
+ sky130_fd_sc_hd__and2_0_139/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a211oi_1_8 sky130_fd_sc_hd__nor2_2_12/Y sky130_fd_sc_hd__nor2_1_136/Y
+ sky130_fd_sc_hd__o22ai_1_202/Y sky130_fd_sc_hd__a211oi_1_8/Y sky130_fd_sc_hd__fa_2_1089/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__dfxtp_1_381 VDD VSS sky130_fd_sc_hd__fa_2_1109/B sky130_fd_sc_hd__dfxtp_1_393/CLK
+ sky130_fd_sc_hd__and2_0_188/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_1 sky130_fd_sc_hd__nand3_1_1/C sky130_fd_sc_hd__nand2_1_1/B
+ sky130_fd_sc_hd__nand2_1_9/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_392 VDD VSS sky130_fd_sc_hd__fa_2_1120/B sky130_fd_sc_hd__dfxtp_1_393/CLK
+ sky130_fd_sc_hd__and2_0_103/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_220 sky130_fd_sc_hd__maj3_1_39/B sky130_fd_sc_hd__maj3_1_40/A
+ sky130_fd_sc_hd__fa_2_220/A sky130_fd_sc_hd__fa_2_220/B sky130_fd_sc_hd__fa_2_221/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_16_9 sky130_fd_sc_hd__buf_12_368/A sky130_fd_sc_hd__bufbuf_8_0/X
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__fa_2_231 sky130_fd_sc_hd__maj3_1_37/B sky130_fd_sc_hd__maj3_1_38/A
+ sky130_fd_sc_hd__fa_2_231/A sky130_fd_sc_hd__fa_2_231/B sky130_fd_sc_hd__fa_2_232/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_242 sky130_fd_sc_hd__fa_2_239/B sky130_fd_sc_hd__fa_2_235/B
+ sky130_fd_sc_hd__fa_2_242/A sky130_fd_sc_hd__fa_2_242/B sky130_fd_sc_hd__fa_2_273/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_253 sky130_fd_sc_hd__fa_2_252/A sky130_fd_sc_hd__fa_2_246/B
+ sky130_fd_sc_hd__fa_2_5/B sky130_fd_sc_hd__fa_2_281/A sky130_fd_sc_hd__fa_2_265/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_264 sky130_fd_sc_hd__fa_2_267/B sky130_fd_sc_hd__fa_2_264/SUM
+ sky130_fd_sc_hd__fa_2_264/A sky130_fd_sc_hd__fa_2_264/B sky130_fd_sc_hd__fa_2_264/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_275 sky130_fd_sc_hd__fa_2_168/A sky130_fd_sc_hd__fa_2_169/B
+ sky130_fd_sc_hd__fa_2_275/A sky130_fd_sc_hd__fa_2_275/B sky130_fd_sc_hd__fa_2_279/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_286 sky130_fd_sc_hd__xnor2_1_2/A sky130_fd_sc_hd__fa_2_286/SUM
+ sky130_fd_sc_hd__ha_2_115/A sky130_fd_sc_hd__fa_2_286/B sky130_fd_sc_hd__fa_2_286/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_2 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_2/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__and2_0_2/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__fa_2_297 sky130_fd_sc_hd__fa_2_296/B sky130_fd_sc_hd__fa_2_297/SUM
+ sky130_fd_sc_hd__ha_2_116/A sky130_fd_sc_hd__ha_2_114/B sky130_fd_sc_hd__fa_2_425/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor4_1_9 sky130_fd_sc_hd__nor4_1_9/D sky130_fd_sc_hd__nor4_1_9/C
+ sky130_fd_sc_hd__nor4_1_9/Y sky130_fd_sc_hd__nor4_1_9/A sky130_fd_sc_hd__nor4_1_9/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__nor4_1
Xsky130_fd_sc_hd__a22oi_1_8 sky130_fd_sc_hd__nor2_2_0/Y sky130_fd_sc_hd__clkinv_1_4/Y
+ sky130_fd_sc_hd__nand4_1_27/Y sky130_fd_sc_hd__nand4_1_11/Y sky130_fd_sc_hd__a22oi_1_8/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__diode_2_103 sky130_fd_sc_hd__inv_2_135/Y VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_114 sky130_fd_sc_hd__buf_2_225/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_125 sky130_fd_sc_hd__buf_2_250/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_136 sky130_fd_sc_hd__clkbuf_1_526/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_147 sky130_fd_sc_hd__buf_2_247/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_158 sky130_fd_sc_hd__clkbuf_4_173/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_169 sky130_fd_sc_hd__clkbuf_4_178/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__buf_2_270 VDD VSS sky130_fd_sc_hd__buf_2_270/X sky130_fd_sc_hd__buf_2_270/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_281 VDD VSS sky130_fd_sc_hd__buf_2_281/X sig_frequency[0]
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_12_203 sky130_fd_sc_hd__buf_6_23/X sky130_fd_sc_hd__buf_12_203/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_50 sky130_fd_sc_hd__nor2_2_6/Y sky130_fd_sc_hd__o22ai_1_82/Y
+ sky130_fd_sc_hd__a21oi_1_50/Y sky130_fd_sc_hd__fa_2_1038/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_214 sky130_fd_sc_hd__buf_12_214/A sky130_fd_sc_hd__buf_12_214/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_61 sky130_fd_sc_hd__a21oi_1_61/A1 sky130_fd_sc_hd__nor2_1_46/B
+ sky130_fd_sc_hd__xnor2_1_52/A sky130_fd_sc_hd__xnor2_1_50/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_225 sky130_fd_sc_hd__buf_12_225/A sky130_fd_sc_hd__buf_12_261/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_72 sky130_fd_sc_hd__xnor2_1_33/B sky130_fd_sc_hd__nor2_1_55/Y
+ sky130_fd_sc_hd__xnor2_1_35/A sky130_fd_sc_hd__nand2_1_244/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_236 sky130_fd_sc_hd__buf_12_236/A sky130_fd_sc_hd__buf_12_236/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_83 sky130_fd_sc_hd__a21o_2_3/A2 sky130_fd_sc_hd__o21ai_1_92/Y
+ sky130_fd_sc_hd__a21oi_1_83/Y sky130_fd_sc_hd__fa_2_1001/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_247 sky130_fd_sc_hd__buf_12_247/A sky130_fd_sc_hd__buf_12_247/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_94 sky130_fd_sc_hd__a21oi_1_94/A1 sky130_fd_sc_hd__o22ai_1_98/Y
+ sky130_fd_sc_hd__a21oi_1_94/Y sky130_fd_sc_hd__a211o_1_6/A1 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_1_106 sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__a22oi_2_12/A1
+ sky130_fd_sc_hd__buf_2_76/X sky130_fd_sc_hd__clkbuf_1_167/X sky130_fd_sc_hd__a22oi_1_106/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_258 sky130_fd_sc_hd__buf_12_258/A sky130_fd_sc_hd__buf_12_258/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_117 sky130_fd_sc_hd__a22oi_1_97/B1 sky130_fd_sc_hd__a22oi_1_97/A1
+ sky130_fd_sc_hd__buf_2_57/X sky130_fd_sc_hd__clkbuf_4_81/X sky130_fd_sc_hd__nand4_1_24/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_269 sky130_fd_sc_hd__buf_12_269/A sky130_fd_sc_hd__buf_12_269/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_128 sky130_fd_sc_hd__a22oi_1_96/B1 sky130_fd_sc_hd__a22oi_1_96/A1
+ sky130_fd_sc_hd__clkbuf_1_143/X sky130_fd_sc_hd__a22oi_1_128/A2 sky130_fd_sc_hd__nand4_1_27/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_139 sky130_fd_sc_hd__a22oi_1_96/B1 sky130_fd_sc_hd__a22oi_1_96/A1
+ sky130_fd_sc_hd__clkbuf_1_140/X sky130_fd_sc_hd__a22oi_1_139/A2 sky130_fd_sc_hd__nand4_1_30/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_403 sky130_fd_sc_hd__nor3_1_32/C sky130_fd_sc_hd__nor4_1_9/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_403/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_414 sky130_fd_sc_hd__o21ai_1_35/A2 sky130_fd_sc_hd__fa_2_944/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_414/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_425 sky130_fd_sc_hd__o22ai_1_60/B2 sky130_fd_sc_hd__dfxtp_1_483/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_425/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_436 sky130_fd_sc_hd__fa_2_961/B sky130_fd_sc_hd__nor2_1_37/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_436/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_447 sky130_fd_sc_hd__fa_2_954/B sky130_fd_sc_hd__dfxtp_1_494/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_447/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_458 sky130_fd_sc_hd__nor2_1_66/B sky130_fd_sc_hd__fa_2_983/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_458/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_469 sky130_fd_sc_hd__a21oi_1_42/A1 sky130_fd_sc_hd__o22ai_1_88/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_469/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_300 sky130_fd_sc_hd__or2_0_9/B sky130_fd_sc_hd__nor3_1_38/C
+ sky130_fd_sc_hd__o21bai_1_2/A2 sky130_fd_sc_hd__nor3_1_38/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_311 sky130_fd_sc_hd__o21a_1_39/B1 sky130_fd_sc_hd__o21a_1_38/A1
+ sky130_fd_sc_hd__a21oi_1_311/Y sky130_fd_sc_hd__o21a_1_42/A2 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_322 sky130_fd_sc_hd__xor2_1_185/X sky130_fd_sc_hd__o21ai_1_341/Y
+ sky130_fd_sc_hd__a21oi_1_322/Y sky130_fd_sc_hd__nand2_1_418/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_333 sky130_fd_sc_hd__nor2_2_16/Y sky130_fd_sc_hd__o21ai_1_354/Y
+ sky130_fd_sc_hd__nor2_1_214/B sky130_fd_sc_hd__fa_2_1189/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_344 sky130_fd_sc_hd__clkinv_1_921/Y sky130_fd_sc_hd__nor2_1_219/Y
+ sky130_fd_sc_hd__a21oi_1_344/Y sky130_fd_sc_hd__nor2b_2_3/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_70 sky130_fd_sc_hd__clkbuf_4_81/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_355 sky130_fd_sc_hd__nor3_1_39/A sky130_fd_sc_hd__o22ai_1_317/Y
+ sky130_fd_sc_hd__a21oi_1_355/Y sky130_fd_sc_hd__fa_2_1201/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_81 sky130_fd_sc_hd__buf_2_134/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_366 sky130_fd_sc_hd__o21a_1_48/B1 sky130_fd_sc_hd__nor2_1_232/Y
+ sky130_fd_sc_hd__a21oi_1_366/Y sky130_fd_sc_hd__nor2_1_232/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_92 sky130_fd_sc_hd__clkbuf_4_208/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_377 sky130_fd_sc_hd__nor3_1_40/B sky130_fd_sc_hd__nor2b_1_119/Y
+ sky130_fd_sc_hd__a21oi_1_377/Y sky130_fd_sc_hd__nor2b_2_4/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_388 sky130_fd_sc_hd__fa_2_1238/A sky130_fd_sc_hd__o22ai_1_357/Y
+ sky130_fd_sc_hd__a21oi_1_388/Y sky130_fd_sc_hd__clkinv_1_946/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_399 sky130_fd_sc_hd__nor3_1_40/A sky130_fd_sc_hd__o22ai_1_365/Y
+ sky130_fd_sc_hd__a21oi_1_399/Y sky130_fd_sc_hd__fa_2_1229/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_3 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1091/A sky130_fd_sc_hd__nor2_4_13/Y
+ sky130_fd_sc_hd__nor2_4_12/Y sky130_fd_sc_hd__xor2_1_88/A sky130_fd_sc_hd__nor2_4_13/A
+ sky130_fd_sc_hd__a222oi_1_3/Y sky130_fd_sc_hd__fa_2_1090/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2_1_360 sky130_fd_sc_hd__nand2_1_360/Y sky130_fd_sc_hd__nor2_1_163/B
+ sky130_fd_sc_hd__o31ai_1_6/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_371 sky130_fd_sc_hd__a21o_2_9/A2 sky130_fd_sc_hd__nand2_1_371/B
+ sky130_fd_sc_hd__nor2_1_170/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_970 sky130_fd_sc_hd__o22ai_1_348/A1 sky130_fd_sc_hd__nor2_1_256/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_970/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_382 sky130_fd_sc_hd__nand2_1_382/Y sky130_fd_sc_hd__xor2_1_163/A
+ sky130_fd_sc_hd__nor2_1_182/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_981 sky130_fd_sc_hd__nand2_1_472/B sky130_fd_sc_hd__fa_2_146/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_981/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_393 sky130_fd_sc_hd__nor2_1_224/A sky130_fd_sc_hd__nand2_1_393/B
+ sky130_fd_sc_hd__o32ai_1_5/B2 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_992 sky130_fd_sc_hd__o22ai_1_361/A1 sky130_fd_sc_hd__fa_2_1234/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_992/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_2_15 VDD VSS sky130_fd_sc_hd__buf_2_15/X sky130_fd_sc_hd__ha_2_17/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_26 VDD VSS sky130_fd_sc_hd__buf_8_1/A sky130_fd_sc_hd__inv_2_3/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_37 VDD VSS sky130_fd_sc_hd__buf_2_37/X sky130_fd_sc_hd__buf_4_36/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_48 VDD VSS sky130_fd_sc_hd__buf_2_48/X sky130_fd_sc_hd__buf_2_48/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_59 VDD VSS sky130_fd_sc_hd__buf_2_59/X sky130_fd_sc_hd__buf_2_59/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o211ai_1_20 sky130_fd_sc_hd__nor2_1_135/Y sky130_fd_sc_hd__nor2_1_127/A
+ sky130_fd_sc_hd__xor2_1_137/A sky130_fd_sc_hd__a22oi_1_357/Y sky130_fd_sc_hd__nand2_1_329/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_31 sky130_fd_sc_hd__o21ai_1_311/A2 sky130_fd_sc_hd__nor2_1_180/A
+ sky130_fd_sc_hd__xor2_1_150/A sky130_fd_sc_hd__nand2_1_384/Y sky130_fd_sc_hd__nand2_1_386/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_42 sky130_fd_sc_hd__nor2_1_222/A sky130_fd_sc_hd__a21oi_1_350/Y
+ sky130_fd_sc_hd__xor2_1_193/A sky130_fd_sc_hd__nand2_1_435/Y sky130_fd_sc_hd__nand2_1_438/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_53 sky130_fd_sc_hd__a21oi_1_395/Y sky130_fd_sc_hd__nor2_1_265/A
+ sky130_fd_sc_hd__xor2_1_269/A sky130_fd_sc_hd__a21oi_1_392/Y sky130_fd_sc_hd__nand2_1_485/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_64 sky130_fd_sc_hd__a21oi_1_455/Y sky130_fd_sc_hd__nor2_1_309/A
+ sky130_fd_sc_hd__xor2_1_310/A sky130_fd_sc_hd__a211oi_1_32/Y sky130_fd_sc_hd__nand2_1_535/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__nor4_1_12 sky130_fd_sc_hd__nor4_1_12/D sky130_fd_sc_hd__nor4_1_12/C
+ sky130_fd_sc_hd__nor4_1_12/Y sky130_fd_sc_hd__nor4_1_12/A sky130_fd_sc_hd__nor4_1_12/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__nor4_1
Xsky130_fd_sc_hd__clkinv_1_200 sky130_fd_sc_hd__inv_2_107/A sky130_fd_sc_hd__a22o_2_8/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_200/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_211 sky130_fd_sc_hd__clkinv_2_25/A sky130_fd_sc_hd__a22oi_1_297/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_211/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_222 sky130_fd_sc_hd__inv_2_113/A sky130_fd_sc_hd__a22o_1_25/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_222/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_233 sky130_fd_sc_hd__inv_2_125/A sky130_fd_sc_hd__inv_2_106/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_233/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_244 sky130_fd_sc_hd__buf_8_210/A sky130_fd_sc_hd__clkinv_1_244/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_244/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_255 sky130_fd_sc_hd__inv_2_133/A sky130_fd_sc_hd__inv_2_128/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_255/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_266 sky130_fd_sc_hd__o21ai_1_29/B1 sky130_fd_sc_hd__ha_2_154/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_266/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_277 sky130_fd_sc_hd__fa_2_91/A sky130_fd_sc_hd__fa_2_82/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_277/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_288 sky130_fd_sc_hd__fa_2_87/B sky130_fd_sc_hd__ha_2_99/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_288/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_299 sky130_fd_sc_hd__fa_2_281/B sky130_fd_sc_hd__ha_2_104/B
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_2_0 sky130_fd_sc_hd__nor2_1_7/Y sky130_fd_sc_hd__o21ai_2_0/Y
+ sky130_fd_sc_hd__or2_1_2/B sky130_fd_sc_hd__or2_1_2/A VSS VDD VDD VSS sky130_fd_sc_hd__o21ai_2
Xsky130_fd_sc_hd__a21oi_1_7 sky130_fd_sc_hd__or4_1_1/C sky130_fd_sc_hd__o21ai_1_10/Y
+ sky130_fd_sc_hd__nor4_1_1/C sky130_fd_sc_hd__nor2b_1_52/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_130 sky130_fd_sc_hd__clkinv_1_585/Y sky130_fd_sc_hd__o22ai_1_134/Y
+ sky130_fd_sc_hd__a21oi_1_130/Y sky130_fd_sc_hd__a211o_1_6/A1 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_141 sky130_fd_sc_hd__nor2_2_10/Y sky130_fd_sc_hd__o22ai_1_141/Y
+ sky130_fd_sc_hd__a21oi_1_141/Y sky130_fd_sc_hd__fa_2_1113/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_152 sky130_fd_sc_hd__nor2_2_11/Y sky130_fd_sc_hd__o22ai_1_151/Y
+ sky130_fd_sc_hd__a21oi_1_152/Y sky130_fd_sc_hd__fa_2_1109/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_163 sky130_fd_sc_hd__nor2_2_11/Y sky130_fd_sc_hd__o22ai_1_162/Y
+ sky130_fd_sc_hd__a21oi_1_163/Y sky130_fd_sc_hd__fa_2_1120/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_174 sky130_fd_sc_hd__nand2_1_306/Y sky130_fd_sc_hd__nor2_1_97/A
+ sky130_fd_sc_hd__xnor2_1_84/A sky130_fd_sc_hd__xnor2_1_82/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_185 sky130_fd_sc_hd__o21a_1_14/B1 sky130_fd_sc_hd__nor2_1_118/Y
+ sky130_fd_sc_hd__dfxtp_1_757/D sky130_fd_sc_hd__nor2_1_118/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_196 sky130_fd_sc_hd__clkinv_1_705/Y sky130_fd_sc_hd__o21ai_1_224/Y
+ sky130_fd_sc_hd__a21oi_1_196/Y sky130_fd_sc_hd__nand2_1_331/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_104 sky130_fd_sc_hd__buf_8_104/A sky130_fd_sc_hd__buf_4_55/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_115 sky130_fd_sc_hd__buf_8_74/X sky130_fd_sc_hd__buf_6_26/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_126 sky130_fd_sc_hd__buf_6_31/X sky130_fd_sc_hd__buf_4_81/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_137 sky130_fd_sc_hd__buf_8_137/A sky130_fd_sc_hd__buf_8_137/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_148 sky130_fd_sc_hd__buf_8_148/A sky130_fd_sc_hd__buf_4_85/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_159 sky130_fd_sc_hd__buf_8_159/A sky130_fd_sc_hd__buf_8_159/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nand2_1_190 sky130_fd_sc_hd__fa_2_664/B sky130_fd_sc_hd__fa_2_700/B
+ sky130_fd_sc_hd__ha_2_130/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__a21o_2_16 sky130_fd_sc_hd__a21o_2_16/X sky130_fd_sc_hd__nor2_1_212/Y
+ sky130_fd_sc_hd__nor2_1_212/A sky130_fd_sc_hd__nor2_1_212/B VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__a21o_2_27 sky130_fd_sc_hd__a21o_2_27/X sky130_fd_sc_hd__nor2_1_296/Y
+ sky130_fd_sc_hd__fa_2_8/SUM sky130_fd_sc_hd__nor2_1_296/B VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__xor2_1_10 sky130_fd_sc_hd__nor4_1_2/B sky130_fd_sc_hd__xor2_1_10/X
+ sky130_fd_sc_hd__nor4_1_4/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_21 sky130_fd_sc_hd__xor2_1_21/B sky130_fd_sc_hd__xor2_1_21/X
+ sky130_fd_sc_hd__nor4_1_4/B VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_32 sky130_fd_sc_hd__xor2_1_32/B sky130_fd_sc_hd__xor2_1_32/X
+ sky130_fd_sc_hd__xor2_1_33/X VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_43 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_984/B
+ sky130_fd_sc_hd__xor2_1_43/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_54 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_973/B
+ sky130_fd_sc_hd__xor2_1_54/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_65 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__xor2_1_65/X
+ sky130_fd_sc_hd__xor2_1_65/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_76 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__xor2_1_76/X
+ sky130_fd_sc_hd__xor2_1_76/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_87 sky130_fd_sc_hd__xor2_1_88/X sky130_fd_sc_hd__xor2_1_87/X
+ sky130_fd_sc_hd__xor2_1_87/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_98 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__xor2_1_98/X
+ sky130_fd_sc_hd__xor2_1_98/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2b_1_4 sky130_fd_sc_hd__nand2b_1_4/Y sky130_fd_sc_hd__nor4_1_5/D
+ sky130_fd_sc_hd__nor3_1_32/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a21o_2_0 sky130_fd_sc_hd__a21o_2_0/X sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__a21o_2_0/A1 sky130_fd_sc_hd__a21o_2_2/A2 VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__dfxtp_1_1309 VDD VSS sky130_fd_sc_hd__fa_2_842/B sky130_fd_sc_hd__dfxtp_1_1322/CLK
+ sky130_fd_sc_hd__o21a_1_65/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_903 VDD VSS sky130_fd_sc_hd__fa_2_938/B sky130_fd_sc_hd__dfxtp_1_904/CLK
+ sky130_fd_sc_hd__dfxtp_1_903/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_914 VDD VSS sky130_fd_sc_hd__fa_2_1143/A sky130_fd_sc_hd__clkinv_8_55/Y
+ sky130_fd_sc_hd__mux2_2_113/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_925 VDD VSS sky130_fd_sc_hd__fa_2_1154/A sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__mux2_2_84/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_936 VDD VSS sky130_fd_sc_hd__fa_2_1128/A sky130_fd_sc_hd__clkinv_8_55/Y
+ sky130_fd_sc_hd__mux2_2_105/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_947 VDD VSS sky130_fd_sc_hd__fa_2_1139/A sky130_fd_sc_hd__clkinv_8_46/Y
+ sky130_fd_sc_hd__mux2_2_79/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_958 VDD VSS sky130_fd_sc_hd__fa_2_1167/A sky130_fd_sc_hd__clkinv_8_65/Y
+ sky130_fd_sc_hd__mux2_2_106/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a221oi_1_2 sky130_fd_sc_hd__a221oi_1_2/Y sky130_fd_sc_hd__xnor2_1_93/Y
+ sky130_fd_sc_hd__xor2_1_185/B sky130_fd_sc_hd__nand2_1_366/Y sky130_fd_sc_hd__o31ai_1_6/A3
+ sky130_fd_sc_hd__nor2_1_163/B VSS VDD VDD VSS sky130_fd_sc_hd__a221oi_1
Xsky130_fd_sc_hd__dfxtp_1_969 VDD VSS sky130_fd_sc_hd__nor3_1_38/C sky130_fd_sc_hd__clkinv_8_46/Y
+ sky130_fd_sc_hd__o21bai_1_2/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_501 VSS VDD sky130_fd_sc_hd__buf_8_208/A sky130_fd_sc_hd__clkbuf_4_203/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_512 VSS VDD sky130_fd_sc_hd__buf_12_398/A sky130_fd_sc_hd__clkbuf_1_516/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_523 VSS VDD sky130_fd_sc_hd__clkbuf_1_523/X sky130_fd_sc_hd__clkbuf_1_523/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_534 VSS VDD sky130_fd_sc_hd__clkbuf_4_207/A sky130_fd_sc_hd__clkbuf_1_534/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_102 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_93/A sky130_fd_sc_hd__fa_2_210/A
+ sky130_fd_sc_hd__ha_2_102/SUM sky130_fd_sc_hd__ha_2_99/A sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_545 VSS VDD sky130_fd_sc_hd__fa_2_242/B sky130_fd_sc_hd__ha_2_96/B
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_113 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_114/B sky130_fd_sc_hd__fa_2_384/CIN
+ sky130_fd_sc_hd__fa_2_376/A sky130_fd_sc_hd__ha_2_113/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_556 VSS VDD sky130_fd_sc_hd__nand2_1_83/B sky130_fd_sc_hd__nand4_1_63/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_124 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_124/A sky130_fd_sc_hd__fa_2_547/B
+ sky130_fd_sc_hd__fa_2_543/B sky130_fd_sc_hd__ha_2_124/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_567 VSS VDD sky130_fd_sc_hd__a22oi_1_13/A2 sig_amplitude[1]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_135 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_135/A sky130_fd_sc_hd__fa_2_700/CIN
+ sky130_fd_sc_hd__fa_2_698/B sky130_fd_sc_hd__ha_2_135/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_578 VSS VDD sky130_fd_sc_hd__nand3_1_12/B sky130_fd_sc_hd__a22oi_1_23/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_146 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_146/A sky130_fd_sc_hd__fa_2_849/CIN
+ sky130_fd_sc_hd__ha_2_146/SUM sky130_fd_sc_hd__ha_2_146/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_589 VSS VDD sky130_fd_sc_hd__nand3_1_3/B sky130_fd_sc_hd__a22oi_1_6/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_157 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_157/A sky130_fd_sc_hd__ha_2_156/B
+ sky130_fd_sc_hd__ha_2_157/SUM sky130_fd_sc_hd__ha_2_157/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_808 sky130_fd_sc_hd__fa_2_810/CIN sky130_fd_sc_hd__fa_2_799/A
+ sky130_fd_sc_hd__ha_2_138/A sky130_fd_sc_hd__fa_2_808/B sky130_fd_sc_hd__fa_2_808/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_168 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_168/A sky130_fd_sc_hd__fa_2_900/A
+ sky130_fd_sc_hd__fa_2_901/B sky130_fd_sc_hd__ha_2_168/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_819 sky130_fd_sc_hd__fa_2_818/B sky130_fd_sc_hd__fa_2_819/SUM
+ sky130_fd_sc_hd__fa_2_819/A sky130_fd_sc_hd__fa_2_819/B sky130_fd_sc_hd__fa_2_823/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_179 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_179/A sky130_fd_sc_hd__ha_2_178/A
+ sky130_fd_sc_hd__ha_2_179/SUM sky130_fd_sc_hd__ha_2_179/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__maj3_1_6 sky130_fd_sc_hd__maj3_1_7/X sky130_fd_sc_hd__maj3_1_6/X
+ sky130_fd_sc_hd__maj3_1_6/B sky130_fd_sc_hd__maj3_1_6/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__ha_2_70 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_70/A sky130_fd_sc_hd__xor2_1_7/A
+ sky130_fd_sc_hd__ha_2_70/SUM sky130_fd_sc_hd__ha_2_70/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_81 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_81/A sky130_fd_sc_hd__ha_2_80/B
+ sky130_fd_sc_hd__ha_2_81/SUM sky130_fd_sc_hd__ha_2_81/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_92 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_93/A sky130_fd_sc_hd__fa_2_52/B
+ sky130_fd_sc_hd__fa_2_48/A sky130_fd_sc_hd__fa_2_2/A sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_0 VSS VDD sky130_fd_sc_hd__clkbuf_1_0/X sky130_fd_sc_hd__nor3_1_4/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__mux2_2_108 VSS VDD sky130_fd_sc_hd__mux2_2_108/A1 sky130_fd_sc_hd__mux2_2_108/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_108/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_119 VSS VDD sky130_fd_sc_hd__mux2_2_119/A1 sky130_fd_sc_hd__mux2_2_119/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_119/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__clkinv_1_0 sky130_fd_sc_hd__nor3_1_1/B sky130_fd_sc_hd__nand2_1_19/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_0/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_190 sky130_fd_sc_hd__nor2_1_190/B sky130_fd_sc_hd__o21a_1_35/A1
+ sky130_fd_sc_hd__nor2_1_190/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__and2_0_15 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_15/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_16/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_26 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_26/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_35/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_306 sky130_fd_sc_hd__nor2_1_191/B sky130_fd_sc_hd__nor2_1_224/A
+ sky130_fd_sc_hd__o22ai_1_306/Y sky130_fd_sc_hd__o22ai_1_319/A1 sky130_fd_sc_hd__a222oi_1_19/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_37 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_37/X sky130_fd_sc_hd__ha_2_50/A
+ sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_317 sky130_fd_sc_hd__o32ai_1_5/A3 sky130_fd_sc_hd__o22ai_1_322/B1
+ sky130_fd_sc_hd__o22ai_1_317/Y sky130_fd_sc_hd__nor2_1_193/B sky130_fd_sc_hd__o21a_1_42/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_48 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_51/A sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__ha_2_52/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_328 sky130_fd_sc_hd__nand2_1_462/Y sky130_fd_sc_hd__nand2_1_461/Y
+ sky130_fd_sc_hd__o22ai_1_328/Y sky130_fd_sc_hd__nand2_1_473/B sky130_fd_sc_hd__o21ai_1_387/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_59 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_59/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_59/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_339 sky130_fd_sc_hd__nand2_1_464/Y sky130_fd_sc_hd__nand2_1_463/Y
+ sky130_fd_sc_hd__o22ai_1_339/Y sky130_fd_sc_hd__nand2_1_472/B sky130_fd_sc_hd__o21ai_1_386/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_2_7 sky130_fd_sc_hd__nor2_2_8/B sky130_fd_sc_hd__nor2_2_7/Y
+ sky130_fd_sc_hd__nor2_2_7/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__buf_8_14 sky130_fd_sc_hd__inv_2_5/Y sky130_fd_sc_hd__buf_8_14/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_25 sky130_fd_sc_hd__ha_2_21/A sky130_fd_sc_hd__buf_8_25/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_36 sky130_fd_sc_hd__buf_8_36/A sky130_fd_sc_hd__buf_8_36/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_47 sky130_fd_sc_hd__inv_2_14/Y sky130_fd_sc_hd__buf_8_47/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_58 sky130_fd_sc_hd__buf_8_58/A sky130_fd_sc_hd__buf_8_58/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_69 sky130_fd_sc_hd__buf_8_69/A sky130_fd_sc_hd__buf_8_69/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__o21ai_1_500 VSS VDD sky130_fd_sc_hd__nand2_1_561/A sky130_fd_sc_hd__o21ai_1_507/A1
+ sky130_fd_sc_hd__nand2_1_561/Y sky130_fd_sc_hd__and2_0_350/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__fa_2_1309 sky130_fd_sc_hd__fa_2_1310/CIN sky130_fd_sc_hd__mux2_2_224/A0
+ sky130_fd_sc_hd__fa_2_1309/A sky130_fd_sc_hd__fa_2_1309/B sky130_fd_sc_hd__fa_2_1309/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1106 VDD VSS sky130_fd_sc_hd__nor2b_2_3/A sky130_fd_sc_hd__clkinv_4_23/Y
+ sky130_fd_sc_hd__nor2b_1_118/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1117 VDD VSS sky130_fd_sc_hd__mux2_2_150/A0 sky130_fd_sc_hd__clkinv_8_49/Y
+ sky130_fd_sc_hd__o22ai_1_276/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1128 VDD VSS sky130_fd_sc_hd__mux2_2_125/A1 sky130_fd_sc_hd__clkinv_8_70/Y
+ sky130_fd_sc_hd__a21oi_1_322/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_700 VDD VSS sky130_fd_sc_hd__mux2_2_35/A0 sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__o21ai_1_40/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1139 VDD VSS sky130_fd_sc_hd__mux2_2_151/A0 sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__dfxtp_1_998/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_711 VDD VSS sky130_fd_sc_hd__mux2_2_11/A1 sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__o21ai_1_51/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_722 VDD VSS sky130_fd_sc_hd__mux2_2_29/A0 sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__o21ai_1_59/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_733 VDD VSS sky130_fd_sc_hd__mux2_2_6/A1 sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__o21ai_1_70/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_744 VDD VSS sky130_fd_sc_hd__and2_0_167/A sky130_fd_sc_hd__dfxtp_1_744/CLK
+ sky130_fd_sc_hd__fa_2_1099/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_755 VDD VSS sky130_fd_sc_hd__fa_2_678/B sky130_fd_sc_hd__dfxtp_1_755/CLK
+ sky130_fd_sc_hd__dfxtp_1_755/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_766 VDD VSS sky130_fd_sc_hd__ha_2_135/A sky130_fd_sc_hd__dfxtp_1_768/CLK
+ sky130_fd_sc_hd__dfxtp_1_766/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_777 VDD VSS sky130_fd_sc_hd__fa_2_1076/A sky130_fd_sc_hd__clkinv_8_55/Y
+ sky130_fd_sc_hd__mux2_2_72/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_788 VDD VSS sky130_fd_sc_hd__fa_2_1087/A sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__mux2_2_48/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_799 VDD VSS sky130_fd_sc_hd__fa_2_1051/A sky130_fd_sc_hd__clkinv_8_54/Y
+ sky130_fd_sc_hd__and2_0_314/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_320 VSS VDD sky130_fd_sc_hd__clkinv_1_156/A sky130_fd_sc_hd__and2_1_5/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_331 VSS VDD sky130_fd_sc_hd__buf_4_58/A sky130_fd_sc_hd__buf_2_274/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_342 VSS VDD sky130_fd_sc_hd__buf_8_137/A sky130_fd_sc_hd__and2_4_0/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_353 VSS VDD sky130_fd_sc_hd__clkbuf_1_353/X sky130_fd_sc_hd__nor3_1_15/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_364 VSS VDD sky130_fd_sc_hd__buf_8_147/A sky130_fd_sc_hd__buf_8_156/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_375 VSS VDD sky130_fd_sc_hd__clkbuf_1_375/X sky130_fd_sc_hd__nand3_1_38/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_386 VSS VDD sky130_fd_sc_hd__clkbuf_1_386/X sky130_fd_sc_hd__clkbuf_1_386/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_397 VSS VDD sky130_fd_sc_hd__a22oi_2_13/B2 sky130_fd_sc_hd__clkbuf_1_397/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_605 sky130_fd_sc_hd__fa_2_607/B sky130_fd_sc_hd__fa_2_605/SUM
+ sky130_fd_sc_hd__fa_2_605/A sky130_fd_sc_hd__fa_2_605/B sky130_fd_sc_hd__fa_2_609/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_616 sky130_fd_sc_hd__fa_2_619/B sky130_fd_sc_hd__fa_2_614/B
+ sky130_fd_sc_hd__fa_2_695/A sky130_fd_sc_hd__fa_2_689/B sky130_fd_sc_hd__fa_2_616/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_627 sky130_fd_sc_hd__fa_2_630/CIN sky130_fd_sc_hd__fa_2_627/SUM
+ sky130_fd_sc_hd__fa_2_627/A sky130_fd_sc_hd__fa_2_627/B sky130_fd_sc_hd__fa_2_627/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_638 sky130_fd_sc_hd__maj3_1_113/B sky130_fd_sc_hd__maj3_1_114/A
+ sky130_fd_sc_hd__fa_2_638/A sky130_fd_sc_hd__fa_2_638/B sky130_fd_sc_hd__fa_2_639/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_649 sky130_fd_sc_hd__maj3_1_110/B sky130_fd_sc_hd__maj3_1_111/A
+ sky130_fd_sc_hd__fa_2_649/A sky130_fd_sc_hd__fa_2_649/B sky130_fd_sc_hd__fa_2_650/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_90 VDD VSS sky130_fd_sc_hd__a22o_1_6/B2 sky130_fd_sc_hd__dfxtp_1_93/CLK
+ sky130_fd_sc_hd__buf_6_52/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_340 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_340/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_340/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_180 sky130_fd_sc_hd__clkbuf_4_180/X sky130_fd_sc_hd__clkbuf_4_180/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_351 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_351/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_351/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_191 sky130_fd_sc_hd__clkbuf_4_191/X sky130_fd_sc_hd__clkbuf_4_191/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__conb_1_4 sky130_fd_sc_hd__conb_1_4/LO sky130_fd_sc_hd__conb_1_4/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__inv_2_140 sky130_fd_sc_hd__nor2_8_2/A sky130_fd_sc_hd__inv_2_140/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__o22ai_1_103 sky130_fd_sc_hd__o22ai_1_130/B1 sky130_fd_sc_hd__o22ai_1_117/A1
+ sky130_fd_sc_hd__nor2_1_79/A sky130_fd_sc_hd__nor2_1_67/B sky130_fd_sc_hd__o22ai_1_132/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_114 sky130_fd_sc_hd__o21a_1_8/A2 sky130_fd_sc_hd__nor2_1_69/B
+ sky130_fd_sc_hd__nor2_1_83/B sky130_fd_sc_hd__o22ai_1_120/B1 sky130_fd_sc_hd__o21ai_1_92/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_125 sky130_fd_sc_hd__nor2_2_9/B sky130_fd_sc_hd__nor2_1_77/A
+ sky130_fd_sc_hd__o22ai_1_125/Y sky130_fd_sc_hd__o21a_1_8/X sky130_fd_sc_hd__a21oi_1_132/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_136 sky130_fd_sc_hd__nand2_1_284/Y sky130_fd_sc_hd__nand2_2_5/Y
+ sky130_fd_sc_hd__o22ai_1_136/Y sky130_fd_sc_hd__xnor2_1_64/Y sky130_fd_sc_hd__o22ai_1_150/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_147 sky130_fd_sc_hd__nand2_1_284/Y sky130_fd_sc_hd__nand2_2_5/Y
+ sky130_fd_sc_hd__o22ai_1_147/Y sky130_fd_sc_hd__xnor2_1_86/Y sky130_fd_sc_hd__o22ai_1_161/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_158 sky130_fd_sc_hd__nand2_1_338/A sky130_fd_sc_hd__nand2_1_284/Y
+ sky130_fd_sc_hd__o22ai_1_158/Y sky130_fd_sc_hd__xnor2_1_80/Y sky130_fd_sc_hd__o22ai_1_158/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_2_14 sky130_fd_sc_hd__nor2_2_15/A sky130_fd_sc_hd__nor3_1_38/A
+ sky130_fd_sc_hd__nor2_2_14/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__o22ai_1_169 sky130_fd_sc_hd__nor2_2_13/B sky130_fd_sc_hd__nor2_1_127/A
+ sky130_fd_sc_hd__o22ai_1_169/Y sky130_fd_sc_hd__a21oi_1_199/Y sky130_fd_sc_hd__nor2_1_131/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand4_1_17 sky130_fd_sc_hd__nand4_1_17/C sky130_fd_sc_hd__nand4_1_17/B
+ sky130_fd_sc_hd__nand4_1_17/Y sky130_fd_sc_hd__nand4_1_17/D sky130_fd_sc_hd__buf_2_111/X
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__o211ai_1_4 sky130_fd_sc_hd__a21oi_1_93/Y sky130_fd_sc_hd__nor2_1_77/A
+ sky130_fd_sc_hd__xor2_1_65/A sky130_fd_sc_hd__o211ai_1_4/C1 sky130_fd_sc_hd__o211ai_1_5/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__nand4_1_28 sky130_fd_sc_hd__nand4_1_28/C sky130_fd_sc_hd__nand4_1_28/B
+ sky130_fd_sc_hd__nand4_1_28/Y sky130_fd_sc_hd__nand4_1_28/D sky130_fd_sc_hd__buf_2_103/X
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand4_1_39 sky130_fd_sc_hd__nand4_1_39/C sky130_fd_sc_hd__nand4_1_39/B
+ sky130_fd_sc_hd__nand4_1_39/Y sky130_fd_sc_hd__nand4_1_39/D sky130_fd_sc_hd__nand4_1_39/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__a31oi_1_1 VSS VDD sky130_fd_sc_hd__a31oi_1_1/Y sky130_fd_sc_hd__a211o_1_2/X
+ sky130_fd_sc_hd__o31ai_1_4/Y sky130_fd_sc_hd__a31oi_1_1/A1 sky130_fd_sc_hd__a31oi_1_1/A3
+ VDD VSS sky130_fd_sc_hd__a31oi_1
Xsky130_fd_sc_hd__o21ai_1_330 VSS VDD sky130_fd_sc_hd__nor2_1_203/Y sky130_fd_sc_hd__or3_1_3/C
+ sky130_fd_sc_hd__o31ai_1_7/A2 sky130_fd_sc_hd__o21ai_1_330/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_341 VSS VDD sky130_fd_sc_hd__xor2_1_185/X sky130_fd_sc_hd__xnor2_1_2/Y
+ sky130_fd_sc_hd__o31ai_1_7/A2 sky130_fd_sc_hd__o21ai_1_341/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_352 VSS VDD sky130_fd_sc_hd__nor3_1_39/A sky130_fd_sc_hd__nor2_1_215/A
+ sky130_fd_sc_hd__nand2_1_432/Y sky130_fd_sc_hd__o21ai_1_352/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a211oi_1_13 sky130_fd_sc_hd__nor2b_1_104/Y sky130_fd_sc_hd__o22ai_1_249/Y
+ sky130_fd_sc_hd__nor2_1_175/Y sky130_fd_sc_hd__a211oi_1_13/Y sky130_fd_sc_hd__o21ai_1_307/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__a211oi_1_24 sky130_fd_sc_hd__nor2b_2_3/Y sky130_fd_sc_hd__o22ai_1_319/Y
+ sky130_fd_sc_hd__nor2_1_225/Y sky130_fd_sc_hd__a211oi_1_24/Y sky130_fd_sc_hd__o21ai_1_383/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_363 VSS VDD sky130_fd_sc_hd__a21oi_1_350/Y sky130_fd_sc_hd__nor2_1_224/A
+ sky130_fd_sc_hd__nand2_1_434/Y sky130_fd_sc_hd__xor2_1_189/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_374 VSS VDD sky130_fd_sc_hd__o21a_1_42/X sky130_fd_sc_hd__nor2_1_222/A
+ sky130_fd_sc_hd__a21oi_1_349/Y sky130_fd_sc_hd__xor2_1_201/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a211oi_1_35 sky130_fd_sc_hd__nor2_2_18/Y sky130_fd_sc_hd__nor2_1_303/Y
+ sky130_fd_sc_hd__o22ai_1_421/Y sky130_fd_sc_hd__nor2_1_302/B sky130_fd_sc_hd__fa_2_1289/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_385 VSS VDD sky130_fd_sc_hd__nand2_1_471/B sky130_fd_sc_hd__nor2_1_251/Y
+ sky130_fd_sc_hd__o31ai_1_9/A1 sky130_fd_sc_hd__o21ai_1_385/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_396 VSS VDD sky130_fd_sc_hd__o22ai_1_358/A1 sky130_fd_sc_hd__nor2_1_267/A
+ sky130_fd_sc_hd__nand2_1_477/Y sky130_fd_sc_hd__xor2_1_255/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__mux2_2_10 VSS VDD sky130_fd_sc_hd__mux2_2_10/A1 sky130_fd_sc_hd__mux2_2_10/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_10/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_21 VSS VDD sky130_fd_sc_hd__mux2_2_21/A1 sky130_fd_sc_hd__mux2_2_21/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_21/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_32 VSS VDD sky130_fd_sc_hd__mux2_2_32/A1 sky130_fd_sc_hd__mux2_2_32/A0
+ sky130_fd_sc_hd__mux2_2_37/S sky130_fd_sc_hd__mux2_2_32/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_43 VSS VDD sky130_fd_sc_hd__mux2_2_43/A1 sky130_fd_sc_hd__mux2_2_43/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_43/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_54 VSS VDD sky130_fd_sc_hd__mux2_2_54/A1 sky130_fd_sc_hd__mux2_2_54/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_54/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_65 VSS VDD sky130_fd_sc_hd__mux2_2_65/A1 sky130_fd_sc_hd__mux2_2_65/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_65/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_76 VSS VDD sky130_fd_sc_hd__mux2_2_76/A1 sky130_fd_sc_hd__xor2_1_162/X
+ sky130_fd_sc_hd__nor2_4_15/A sky130_fd_sc_hd__mux2_2_76/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_87 VSS VDD sky130_fd_sc_hd__mux2_2_87/A1 sky130_fd_sc_hd__mux2_2_87/A0
+ sky130_fd_sc_hd__nor2_4_15/A sky130_fd_sc_hd__mux2_2_87/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1106 sky130_fd_sc_hd__xor2_1_138/B sky130_fd_sc_hd__mux2_2_68/A0
+ sky130_fd_sc_hd__fa_2_1106/A sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1106/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__mux2_2_98 VSS VDD sky130_fd_sc_hd__mux2_2_98/A1 sky130_fd_sc_hd__mux2_2_98/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_98/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1117 sky130_fd_sc_hd__fa_2_1118/CIN sky130_fd_sc_hd__fa_2_1117/SUM
+ sky130_fd_sc_hd__fa_2_1117/A sky130_fd_sc_hd__fa_2_1117/B sky130_fd_sc_hd__fa_2_1117/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1128 sky130_fd_sc_hd__fa_2_1129/CIN sky130_fd_sc_hd__mux2_2_105/A1
+ sky130_fd_sc_hd__fa_2_1128/A sky130_fd_sc_hd__fa_2_1128/B sky130_fd_sc_hd__fa_2_1128/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1139 sky130_fd_sc_hd__xor2_1_141/B sky130_fd_sc_hd__mux2_2_79/A0
+ sky130_fd_sc_hd__fa_2_1139/A sky130_fd_sc_hd__fa_2_1139/B sky130_fd_sc_hd__fa_2_1139/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__xor2_1_190 sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__fa_2_1189/B
+ sky130_fd_sc_hd__xor2_1_190/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_530 VDD VSS sky130_fd_sc_hd__fa_2_961/A sky130_fd_sc_hd__dfxtp_1_533/CLK
+ sky130_fd_sc_hd__and2_0_260/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_541 VDD VSS sky130_fd_sc_hd__or3_1_0/B sky130_fd_sc_hd__dfxtp_1_544/CLK
+ sky130_fd_sc_hd__a22o_1_44/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_552 VDD VSS sky130_fd_sc_hd__dfxtp_1_552/Q sky130_fd_sc_hd__dfxtp_1_594/CLK
+ sky130_fd_sc_hd__dfxtp_1_552/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_563 VDD VSS sky130_fd_sc_hd__and2_0_218/A sky130_fd_sc_hd__dfxtp_1_571/CLK
+ sky130_fd_sc_hd__dfxtp_1_564/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_574 VDD VSS sky130_fd_sc_hd__a22o_1_36/B1 sky130_fd_sc_hd__dfxtp_1_576/CLK
+ sky130_fd_sc_hd__a22o_1_36/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_585 VDD VSS sky130_fd_sc_hd__nor4_1_8/A sky130_fd_sc_hd__dfxtp_1_591/CLK
+ sky130_fd_sc_hd__and2_0_252/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_596 VDD VSS sky130_fd_sc_hd__and2_0_206/A sky130_fd_sc_hd__dfxtp_1_601/CLK
+ sky130_fd_sc_hd__fa_2_1016/B VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_150 VSS VDD sky130_fd_sc_hd__clkbuf_1_150/X sky130_fd_sc_hd__clkbuf_1_250/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_161 VSS VDD sky130_fd_sc_hd__a22oi_2_12/A2 sky130_fd_sc_hd__clkbuf_1_161/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_172 VSS VDD sky130_fd_sc_hd__a22oi_1_86/A2 sky130_fd_sc_hd__clkbuf_1_172/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_183 VSS VDD sky130_fd_sc_hd__nand4_1_23/B sky130_fd_sc_hd__a22oi_1_114/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_194 VSS VDD sky130_fd_sc_hd__buf_12_135/A sky130_fd_sc_hd__clkbuf_1_228/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_402 sky130_fd_sc_hd__maj3_1_59/B sky130_fd_sc_hd__maj3_1_60/A
+ sky130_fd_sc_hd__fa_2_402/A sky130_fd_sc_hd__fa_2_402/B sky130_fd_sc_hd__fa_2_403/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_413 sky130_fd_sc_hd__fa_2_415/CIN sky130_fd_sc_hd__fa_2_410/A
+ sky130_fd_sc_hd__fa_2_413/A sky130_fd_sc_hd__fa_2_413/B sky130_fd_sc_hd__fa_2_413/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_424 sky130_fd_sc_hd__fa_2_423/B sky130_fd_sc_hd__fa_2_420/B
+ sky130_fd_sc_hd__fa_2_424/A sky130_fd_sc_hd__fa_2_424/B sky130_fd_sc_hd__fa_2_412/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_435 sky130_fd_sc_hd__fa_2_426/CIN sky130_fd_sc_hd__a21o_2_9/A1
+ sky130_fd_sc_hd__fa_2_435/A sky130_fd_sc_hd__fa_2_435/B sky130_fd_sc_hd__fa_2_435/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_446 sky130_fd_sc_hd__fa_2_442/B sky130_fd_sc_hd__fa_2_445/B
+ sky130_fd_sc_hd__fa_2_446/A sky130_fd_sc_hd__fa_2_446/B sky130_fd_sc_hd__fa_2_446/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_457 sky130_fd_sc_hd__fa_2_454/CIN sky130_fd_sc_hd__fa_2_459/A
+ sky130_fd_sc_hd__fa_2_546/B sky130_fd_sc_hd__fa_2_555/A sky130_fd_sc_hd__fa_2_531/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_468 sky130_fd_sc_hd__maj3_1_104/B sky130_fd_sc_hd__maj3_1_105/A
+ sky130_fd_sc_hd__fa_2_502/B sky130_fd_sc_hd__fa_2_558/B sky130_fd_sc_hd__fa_2_468/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_479 sky130_fd_sc_hd__maj3_1_99/B sky130_fd_sc_hd__maj3_1_100/A
+ sky130_fd_sc_hd__fa_2_479/A sky130_fd_sc_hd__fa_2_479/B sky130_fd_sc_hd__fa_2_480/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nand3_1_50 sky130_fd_sc_hd__nand3_1_50/Y sky130_fd_sc_hd__nand3_1_50/A
+ sky130_fd_sc_hd__nand3_1_50/C sky130_fd_sc_hd__nand3_1_50/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__and2_0_170 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_170/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_170/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_181 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_181/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_181/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_192 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_192/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_899/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_407 sky130_fd_sc_hd__buf_8_204/X sky130_fd_sc_hd__buf_12_407/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_418 sky130_fd_sc_hd__buf_8_223/X sky130_fd_sc_hd__buf_12_504/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_429 sky130_fd_sc_hd__buf_8_215/X sky130_fd_sc_hd__buf_12_496/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__fa_2_980 sky130_fd_sc_hd__fa_2_981/CIN sky130_fd_sc_hd__mux2_2_27/A0
+ sky130_fd_sc_hd__fa_2_980/A sky130_fd_sc_hd__fa_2_980/B sky130_fd_sc_hd__fa_2_980/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_991 sky130_fd_sc_hd__fa_2_992/CIN sky130_fd_sc_hd__mux2_2_5/A0
+ sky130_fd_sc_hd__fa_2_991/A sky130_fd_sc_hd__fa_2_991/B sky130_fd_sc_hd__fa_2_991/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_1_607 sky130_fd_sc_hd__ha_2_183/B sky130_fd_sc_hd__fa_2_1032/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_607/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_618 sky130_fd_sc_hd__nand2_2_6/A sky130_fd_sc_hd__nand2_1_339/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_618/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_629 sky130_fd_sc_hd__a211o_1_9/A1 sky130_fd_sc_hd__nor2_1_126/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_629/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_160 VSS VDD sky130_fd_sc_hd__o21ai_1_171/A2 sky130_fd_sc_hd__xnor2_1_67/Y
+ sky130_fd_sc_hd__a21oi_1_137/Y sky130_fd_sc_hd__o21ai_1_160/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_171 VSS VDD sky130_fd_sc_hd__o21ai_1_171/A2 sky130_fd_sc_hd__xnor2_1_89/Y
+ sky130_fd_sc_hd__a21oi_1_148/Y sky130_fd_sc_hd__o21ai_1_171/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_182 VSS VDD sky130_fd_sc_hd__nand2_2_5/Y sky130_fd_sc_hd__xnor2_1_77/Y
+ sky130_fd_sc_hd__a21oi_1_157/Y sky130_fd_sc_hd__o21ai_1_182/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_193 VSS VDD sky130_fd_sc_hd__xnor2_1_85/A sky130_fd_sc_hd__o21ai_1_193/A1
+ sky130_fd_sc_hd__nand2_1_292/B sky130_fd_sc_hd__xnor2_1_87/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__edfxtp_1_0 VDD VSS sky130_fd_sc_hd__edfxtp_1_0/CLK sky130_fd_sc_hd__nor2_1_29/A
+ sky130_fd_sc_hd__xor2_1_27/X sky130_fd_sc_hd__edfxtp_1_0/Q VDD VSS sky130_fd_sc_hd__edfxtp_1
Xsky130_fd_sc_hd__a222oi_1_16 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1190/A sky130_fd_sc_hd__nor2_2_16/Y
+ sky130_fd_sc_hd__nor3_1_39/A sky130_fd_sc_hd__nor2_4_16/B sky130_fd_sc_hd__xor2_1_209/A
+ sky130_fd_sc_hd__a222oi_1_16/Y sky130_fd_sc_hd__fa_2_1189/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_27 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1228/A sky130_fd_sc_hd__nor2_2_17/Y
+ sky130_fd_sc_hd__nor3_1_40/A sky130_fd_sc_hd__fa_2_1230/A sky130_fd_sc_hd__nor3_1_40/B
+ sky130_fd_sc_hd__a222oi_1_27/Y sky130_fd_sc_hd__fa_2_1227/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_38 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1278/A sky130_fd_sc_hd__nor2_2_18/Y
+ sky130_fd_sc_hd__nor3_1_41/A sky130_fd_sc_hd__fa_2_1280/A sky130_fd_sc_hd__nor3_1_41/B
+ sky130_fd_sc_hd__a222oi_1_38/Y sky130_fd_sc_hd__fa_2_1277/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2_1_520 sky130_fd_sc_hd__nand2_1_520/Y sky130_fd_sc_hd__nand2_1_520/B
+ sky130_fd_sc_hd__nor2_8_2/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_531 sky130_fd_sc_hd__nand2_1_531/Y sky130_fd_sc_hd__nand2_1_543/B
+ sky130_fd_sc_hd__o21ai_1_467/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_18 VSS VDD sky130_fd_sc_hd__nor2_1_20/B sky130_fd_sc_hd__maj3_1_0/A
+ sky130_fd_sc_hd__nor2_1_9/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_542 sky130_fd_sc_hd__nand2_1_542/Y sky130_fd_sc_hd__nor2b_2_5/A
+ sky130_fd_sc_hd__xor2_1_298/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_29 VSS VDD sky130_fd_sc_hd__or4_1_2/X sky130_fd_sc_hd__a21o_2_0/A1
+ sky130_fd_sc_hd__nor4_1_6/C VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_553 sky130_fd_sc_hd__nand2_1_553/Y sky130_fd_sc_hd__buf_6_49/A
+ sky130_fd_sc_hd__nor2_1_316/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_564 sky130_fd_sc_hd__nand2_1_564/Y sky130_fd_sc_hd__buf_4_121/X
+ sky130_fd_sc_hd__nand2_1_564/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_0 sky130_fd_sc_hd__nor3_1_1/Y sky130_fd_sc_hd__nor2b_1_0/Y
+ sky130_fd_sc_hd__nor2_1_2/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1100 sky130_fd_sc_hd__o32ai_1_11/B2 sky130_fd_sc_hd__o32ai_1_11/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1100/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1111 sky130_fd_sc_hd__nor4_1_13/B sky130_fd_sc_hd__o22ai_1_437/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1111/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1122 sky130_fd_sc_hd__inv_8_0/A sky130_fd_sc_hd__buf_2_143/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1122/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1133 sky130_fd_sc_hd__clkinv_1_1134/A sky130_fd_sc_hd__nand2_1_568/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1133/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_360 VDD VSS sky130_fd_sc_hd__a22o_2_5/B2 sky130_fd_sc_hd__dfxtp_1_360/CLK
+ sky130_fd_sc_hd__xor2_1_17/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_371 VDD VSS sky130_fd_sc_hd__fa_2_1115/A sky130_fd_sc_hd__dfxtp_1_391/CLK
+ sky130_fd_sc_hd__and2_0_133/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a211oi_1_9 sky130_fd_sc_hd__nor2_2_12/Y sky130_fd_sc_hd__nor2_1_137/Y
+ sky130_fd_sc_hd__o22ai_1_204/Y sky130_fd_sc_hd__a211oi_1_9/Y sky130_fd_sc_hd__fa_2_1088/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__dfxtp_1_382 VDD VSS sky130_fd_sc_hd__fa_2_1110/B sky130_fd_sc_hd__clkinv_4_32/Y
+ sky130_fd_sc_hd__and2_0_155/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_2 sky130_fd_sc_hd__nand3_1_2/C sky130_fd_sc_hd__nand2_1_2/B
+ sky130_fd_sc_hd__nand2_1_9/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_393 VDD VSS sky130_fd_sc_hd__nor2_2_11/A sky130_fd_sc_hd__dfxtp_1_393/CLK
+ sky130_fd_sc_hd__and2_0_101/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_210 sky130_fd_sc_hd__fa_2_212/CIN sky130_fd_sc_hd__fa_2_205/A
+ sky130_fd_sc_hd__fa_2_210/A sky130_fd_sc_hd__fa_2_210/B sky130_fd_sc_hd__fa_2_217/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_221 sky130_fd_sc_hd__fa_2_226/B sky130_fd_sc_hd__fa_2_221/SUM
+ sky130_fd_sc_hd__fa_2_221/A sky130_fd_sc_hd__fa_2_221/B sky130_fd_sc_hd__fa_2_221/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_232 sky130_fd_sc_hd__fa_2_236/B sky130_fd_sc_hd__fa_2_232/SUM
+ sky130_fd_sc_hd__fa_2_232/A sky130_fd_sc_hd__fa_2_232/B sky130_fd_sc_hd__fa_2_232/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_243 sky130_fd_sc_hd__fa_2_244/CIN sky130_fd_sc_hd__fa_2_237/A
+ sky130_fd_sc_hd__ha_2_104/B sky130_fd_sc_hd__fa_2_281/A sky130_fd_sc_hd__fa_2_277/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_254 sky130_fd_sc_hd__fa_2_256/B sky130_fd_sc_hd__fa_2_251/A
+ sky130_fd_sc_hd__fa_2_281/B sky130_fd_sc_hd__fa_2_254/B sky130_fd_sc_hd__ha_2_106/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_265 sky130_fd_sc_hd__fa_2_264/A sky130_fd_sc_hd__fa_2_260/A
+ sky130_fd_sc_hd__fa_2_274/A sky130_fd_sc_hd__fa_2_265/B sky130_fd_sc_hd__fa_2_277/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_276 sky130_fd_sc_hd__fa_2_275/B sky130_fd_sc_hd__fa_2_276/SUM
+ sky130_fd_sc_hd__fa_2_276/A sky130_fd_sc_hd__fa_2_276/B sky130_fd_sc_hd__fa_2_280/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_287 sky130_fd_sc_hd__fa_2_286/CIN sky130_fd_sc_hd__nor2_1_208/A
+ sky130_fd_sc_hd__fa_2_389/B sky130_fd_sc_hd__fa_2_287/B sky130_fd_sc_hd__fa_2_287/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_3 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_3/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_8/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__fa_2_298 sky130_fd_sc_hd__fa_2_294/B sky130_fd_sc_hd__fa_2_298/SUM
+ sky130_fd_sc_hd__ha_2_115/A sky130_fd_sc_hd__fa_2_393/A sky130_fd_sc_hd__fa_2_424/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22oi_1_9 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__a22oi_1_9/A1
+ sky130_fd_sc_hd__buf_2_287/X sky130_fd_sc_hd__a22oi_1_9/A2 sky130_fd_sc_hd__nand3_1_4/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__diode_2_104 sky130_fd_sc_hd__inv_2_135/Y VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_115 sky130_fd_sc_hd__buf_2_225/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_126 sky130_fd_sc_hd__buf_2_250/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_137 sky130_fd_sc_hd__clkbuf_1_526/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_148 sky130_fd_sc_hd__clkbuf_1_541/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__fa_2_90 sky130_fd_sc_hd__fa_2_94/B sky130_fd_sc_hd__fa_2_90/SUM
+ sky130_fd_sc_hd__fa_2_90/A sky130_fd_sc_hd__fa_2_90/B sky130_fd_sc_hd__fa_2_90/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__diode_2_159 sky130_fd_sc_hd__clkbuf_4_173/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__buf_2_260 VDD VSS sky130_fd_sc_hd__fa_2_5/B sky130_fd_sc_hd__fa_2_82/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_271 VDD VSS sky130_fd_sc_hd__buf_2_271/X sky130_fd_sc_hd__buf_2_271/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_282 VDD VSS sky130_fd_sc_hd__buf_2_282/X sig_amplitude[0]
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__a21oi_1_40 sky130_fd_sc_hd__nor2_1_41/Y sky130_fd_sc_hd__o22ai_1_73/Y
+ sky130_fd_sc_hd__a21oi_1_40/Y sky130_fd_sc_hd__fa_2_1043/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_204 sky130_fd_sc_hd__buf_4_45/X sky130_fd_sc_hd__buf_12_262/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_51 sky130_fd_sc_hd__nor2_2_6/Y sky130_fd_sc_hd__o22ai_1_83/Y
+ sky130_fd_sc_hd__a21oi_1_51/Y sky130_fd_sc_hd__fa_2_1039/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_215 sky130_fd_sc_hd__buf_4_52/X sky130_fd_sc_hd__buf_12_215/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_62 sky130_fd_sc_hd__a21oi_1_62/A1 sky130_fd_sc_hd__nor2_1_45/B
+ sky130_fd_sc_hd__xnor2_1_48/A sky130_fd_sc_hd__xnor2_1_46/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_226 sky130_fd_sc_hd__buf_12_226/A sky130_fd_sc_hd__buf_12_265/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_73 sky130_fd_sc_hd__o21a_1_2/B1 sky130_fd_sc_hd__o21a_1_1/A1
+ sky130_fd_sc_hd__a21oi_1_73/Y sky130_fd_sc_hd__nor2_1_63/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_237 sky130_fd_sc_hd__buf_12_237/A sky130_fd_sc_hd__buf_12_237/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_84 sky130_fd_sc_hd__a21oi_1_88/A2 sky130_fd_sc_hd__a21oi_1_85/B1
+ sky130_fd_sc_hd__a21oi_1_84/Y sky130_fd_sc_hd__a211o_1_6/A1 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_248 sky130_fd_sc_hd__buf_12_248/A sky130_fd_sc_hd__buf_12_248/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_95 sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__o21ai_1_110/Y
+ sky130_fd_sc_hd__a21oi_1_95/Y sky130_fd_sc_hd__fa_2_987/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_1_107 sky130_fd_sc_hd__clkbuf_4_72/X sky130_fd_sc_hd__clkbuf_4_73/X
+ sky130_fd_sc_hd__a22oi_1_107/B2 sky130_fd_sc_hd__buf_2_92/X sky130_fd_sc_hd__buf_2_107/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_259 sky130_fd_sc_hd__buf_12_259/A sky130_fd_sc_hd__buf_12_259/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_118 sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__a22oi_2_12/A1
+ sky130_fd_sc_hd__buf_2_73/X sky130_fd_sc_hd__clkbuf_1_164/X sky130_fd_sc_hd__a22oi_1_118/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_129 sky130_fd_sc_hd__a22oi_1_97/B1 sky130_fd_sc_hd__a22oi_1_97/A1
+ sky130_fd_sc_hd__buf_2_54/X sky130_fd_sc_hd__clkbuf_4_78/X sky130_fd_sc_hd__nand4_1_27/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkinv_1_404 sky130_fd_sc_hd__nor3_1_31/B sky130_fd_sc_hd__or4_1_2/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_404/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_415 sky130_fd_sc_hd__nor2_1_36/A sky130_fd_sc_hd__fa_2_945/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_415/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_426 sky130_fd_sc_hd__o21ai_1_38/A2 sky130_fd_sc_hd__fa_2_969/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_426/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_437 sky130_fd_sc_hd__fa_2_955/B sky130_fd_sc_hd__dfxtp_1_493/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_437/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_448 sky130_fd_sc_hd__fa_2_953/B sky130_fd_sc_hd__nor2b_1_85/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_448/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_459 sky130_fd_sc_hd__nor2_1_67/B sky130_fd_sc_hd__fa_2_981/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_459/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_6_80 VDD VSS sky130_fd_sc_hd__buf_6_80/X sky130_fd_sc_hd__buf_6_80/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__a21oi_1_301 sky130_fd_sc_hd__o21a_1_31/B1 sky130_fd_sc_hd__o21a_1_30/A1
+ sky130_fd_sc_hd__a21oi_1_301/Y sky130_fd_sc_hd__nor2_1_218/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_312 sky130_fd_sc_hd__o21a_1_40/B1 sky130_fd_sc_hd__o21a_1_39/A1
+ sky130_fd_sc_hd__a21oi_1_312/Y sky130_fd_sc_hd__nor2_1_195/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_323 sky130_fd_sc_hd__o21ai_1_352/Y sky130_fd_sc_hd__clkinv_1_901/Y
+ sky130_fd_sc_hd__a21oi_1_323/Y sky130_fd_sc_hd__nor2b_2_3/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_334 sky130_fd_sc_hd__fa_2_1187/A sky130_fd_sc_hd__o22ai_1_302/Y
+ sky130_fd_sc_hd__a21oi_1_334/Y sky130_fd_sc_hd__nor3_1_39/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_60 sky130_fd_sc_hd__buf_2_102/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_345 sky130_fd_sc_hd__fa_2_1205/A sky130_fd_sc_hd__o22ai_1_311/Y
+ sky130_fd_sc_hd__a21oi_1_345/Y sky130_fd_sc_hd__clkinv_1_861/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_71 sky130_fd_sc_hd__clkbuf_4_81/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_356 sky130_fd_sc_hd__fa_2_1197/A sky130_fd_sc_hd__o22ai_1_318/Y
+ sky130_fd_sc_hd__a21oi_1_356/Y sky130_fd_sc_hd__nor3_1_39/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_82 sky130_fd_sc_hd__nand4_1_42/B VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_367 sky130_fd_sc_hd__nor2_1_233/A sky130_fd_sc_hd__o21a_1_48/A1
+ sky130_fd_sc_hd__a21oi_1_367/Y sky130_fd_sc_hd__nor2_1_233/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_93 sky130_fd_sc_hd__clkbuf_4_208/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_378 sky130_fd_sc_hd__or3_1_4/C sky130_fd_sc_hd__o21ai_1_384/Y
+ sky130_fd_sc_hd__a21oi_1_378/Y sky130_fd_sc_hd__nor2_1_246/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_389 sky130_fd_sc_hd__nor2b_2_4/Y sky130_fd_sc_hd__o21ai_1_404/Y
+ sky130_fd_sc_hd__a21oi_1_389/Y sky130_fd_sc_hd__o21ai_1_413/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_4 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1141/A sky130_fd_sc_hd__nor2_2_15/Y
+ sky130_fd_sc_hd__nor3_1_38/A sky130_fd_sc_hd__fa_2_1143/A sky130_fd_sc_hd__nor3_1_38/B
+ sky130_fd_sc_hd__a222oi_1_4/Y sky130_fd_sc_hd__fa_2_1140/B sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2_1_350 sky130_fd_sc_hd__o21a_1_24/B1 sky130_fd_sc_hd__fa_2_1154/A
+ sky130_fd_sc_hd__o21a_1_24/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_361 sky130_fd_sc_hd__nand2_1_361/Y sky130_fd_sc_hd__nand2_1_364/Y
+ sky130_fd_sc_hd__nand2_1_362/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_960 sky130_fd_sc_hd__nor2_1_239/A sky130_fd_sc_hd__nor2_1_240/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_960/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_372 sky130_fd_sc_hd__nor2_1_170/B sky130_fd_sc_hd__nand2_1_372/B
+ sky130_fd_sc_hd__nor2_1_171/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_971 sky130_fd_sc_hd__o22ai_1_349/A1 sky130_fd_sc_hd__or3_1_4/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_971/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_383 sky130_fd_sc_hd__nand2_1_383/Y sky130_fd_sc_hd__nand2_1_387/B
+ sky130_fd_sc_hd__o21ai_1_328/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_982 sky130_fd_sc_hd__nand2_1_473/B sky130_fd_sc_hd__fa_2_148/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_982/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_394 sky130_fd_sc_hd__xnor2_1_94/B sky130_fd_sc_hd__fa_2_1189/A
+ sky130_fd_sc_hd__o21a_1_30/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_993 sky130_fd_sc_hd__nor2_1_234/B sky130_fd_sc_hd__fa_2_1227/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_993/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand3_4_0 sky130_fd_sc_hd__nand3_4_0/Y sky130_fd_sc_hd__nand3_4_1/A
+ sky130_fd_sc_hd__nand3_4_0/B sky130_fd_sc_hd__nand3_4_1/B VSS VDD VSS VDD sky130_fd_sc_hd__nand3_4
Xsky130_fd_sc_hd__dfxtp_1_190 VDD VSS sky130_fd_sc_hd__ha_2_66/A sky130_fd_sc_hd__dfxtp_1_197/CLK
+ sky130_fd_sc_hd__nor2b_1_27/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_2_16 VDD VSS sky130_fd_sc_hd__buf_2_16/X sky130_fd_sc_hd__ha_2_18/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_27 VDD VSS sky130_fd_sc_hd__buf_8_54/A sky130_fd_sc_hd__ha_2_29/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_38 VDD VSS sky130_fd_sc_hd__buf_4_39/A sky130_fd_sc_hd__buf_2_38/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_49 VDD VSS sky130_fd_sc_hd__buf_8_91/A sky130_fd_sc_hd__ha_2_44/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__a21boi_1_0 sky130_fd_sc_hd__a21boi_1_0/Y sky130_fd_sc_hd__fa_2_995/A
+ sky130_fd_sc_hd__a21oi_1_131/Y sky130_fd_sc_hd__a21o_2_3/A2 VDD VSS VDD VSS sky130_fd_sc_hd__a21boi_1
Xsky130_fd_sc_hd__o211ai_1_10 sky130_fd_sc_hd__nor2_1_85/Y sky130_fd_sc_hd__nor2_1_77/A
+ sky130_fd_sc_hd__xor2_1_83/A sky130_fd_sc_hd__a22oi_1_333/Y sky130_fd_sc_hd__nand2_1_272/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_21 sky130_fd_sc_hd__nand2_2_6/Y sky130_fd_sc_hd__a21oi_1_220/Y
+ sky130_fd_sc_hd__xor2_1_93/A sky130_fd_sc_hd__nand2_1_331/Y sky130_fd_sc_hd__nand2_1_334/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_32 sky130_fd_sc_hd__nor2_1_180/A sky130_fd_sc_hd__a211oi_1_16/Y
+ sky130_fd_sc_hd__xor2_1_151/A sky130_fd_sc_hd__nand2_1_385/Y sky130_fd_sc_hd__nand2_1_386/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_43 sky130_fd_sc_hd__o21ai_1_365/A2 sky130_fd_sc_hd__nor2_1_222/A
+ sky130_fd_sc_hd__xor2_1_195/A sky130_fd_sc_hd__nand2_1_436/Y sky130_fd_sc_hd__nand2_1_438/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_54 sky130_fd_sc_hd__nor2_1_265/A sky130_fd_sc_hd__a21oi_1_410/Y
+ sky130_fd_sc_hd__xor2_1_238/A sky130_fd_sc_hd__nand2_1_487/Y sky130_fd_sc_hd__nand2_1_490/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_65 sky130_fd_sc_hd__a21oi_1_455/Y sky130_fd_sc_hd__nor2_1_307/A
+ sky130_fd_sc_hd__xor2_1_314/A sky130_fd_sc_hd__a21oi_1_452/Y sky130_fd_sc_hd__nand2_1_537/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__clkinv_1_201 sky130_fd_sc_hd__buf_8_209/A sky130_fd_sc_hd__clkinv_1_201/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_201/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor4_1_13 sky130_fd_sc_hd__nor4_1_13/D sky130_fd_sc_hd__nor4_1_13/C
+ sky130_fd_sc_hd__nor4_1_13/Y sky130_fd_sc_hd__nor4_1_13/A sky130_fd_sc_hd__nor4_1_13/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__nor4_1
Xsky130_fd_sc_hd__clkinv_1_212 sky130_fd_sc_hd__clkinv_2_26/A sky130_fd_sc_hd__a22oi_1_293/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_212/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_223 sky130_fd_sc_hd__buf_8_199/A sky130_fd_sc_hd__inv_4_0/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_223/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_234 sky130_fd_sc_hd__inv_2_126/A sky130_fd_sc_hd__inv_2_106/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_234/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_245 sky130_fd_sc_hd__clkinv_1_246/A sky130_fd_sc_hd__buf_8_214/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_245/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_256 sky130_fd_sc_hd__buf_8_219/A sky130_fd_sc_hd__inv_2_134/Y
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_267 sky130_fd_sc_hd__o22ai_1_0/B2 sky130_fd_sc_hd__ha_2_150/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_267/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_278 sky130_fd_sc_hd__fa_2_2/B sky130_fd_sc_hd__ha_2_97/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_278/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_289 sky130_fd_sc_hd__fa_2_91/B sky130_fd_sc_hd__ha_2_93/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_289/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_8 sky130_fd_sc_hd__or4_1_1/D sky130_fd_sc_hd__o21ai_1_11/Y
+ sky130_fd_sc_hd__a21oi_1_8/Y sky130_fd_sc_hd__o31ai_1_1/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_120 sky130_fd_sc_hd__clkinv_1_461/Y sky130_fd_sc_hd__o22ai_1_127/Y
+ sky130_fd_sc_hd__a21oi_1_120/Y sky130_fd_sc_hd__a211o_1_8/A2 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_131 sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__a22o_1_70/X
+ sky130_fd_sc_hd__a21oi_1_131/Y sky130_fd_sc_hd__fa_2_993/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_142 sky130_fd_sc_hd__nor2_2_10/Y sky130_fd_sc_hd__o22ai_1_142/Y
+ sky130_fd_sc_hd__a21oi_1_142/Y sky130_fd_sc_hd__fa_2_1114/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_153 sky130_fd_sc_hd__nor2_2_11/Y sky130_fd_sc_hd__o22ai_1_152/Y
+ sky130_fd_sc_hd__a21oi_1_153/Y sky130_fd_sc_hd__fa_2_1110/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_164 sky130_fd_sc_hd__nor2_2_11/Y sky130_fd_sc_hd__o22ai_1_163/Y
+ sky130_fd_sc_hd__a21oi_1_164/Y sky130_fd_sc_hd__a22o_1_72/A2 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_175 sky130_fd_sc_hd__nand2_1_305/Y sky130_fd_sc_hd__nor2_1_96/A
+ sky130_fd_sc_hd__xnor2_1_80/A sky130_fd_sc_hd__xnor2_1_78/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_186 sky130_fd_sc_hd__o21a_1_15/B1 sky130_fd_sc_hd__o21a_1_14/A1
+ sky130_fd_sc_hd__dfxtp_1_755/D sky130_fd_sc_hd__nor2_1_119/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_197 sky130_fd_sc_hd__a21o_2_5/A2 sky130_fd_sc_hd__o21ai_1_225/Y
+ sky130_fd_sc_hd__a21oi_1_197/Y sky130_fd_sc_hd__fa_2_1067/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_105 sky130_fd_sc_hd__buf_8_105/A sky130_fd_sc_hd__buf_8_105/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_116 sky130_fd_sc_hd__buf_8_124/A sky130_fd_sc_hd__buf_4_76/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_127 sky130_fd_sc_hd__buf_8_127/A sky130_fd_sc_hd__buf_4_75/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_138 sky130_fd_sc_hd__and2_4_0/X sky130_fd_sc_hd__buf_4_70/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_149 sky130_fd_sc_hd__buf_8_149/A sky130_fd_sc_hd__buf_8_149/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nand2_1_180 sky130_fd_sc_hd__fa_2_512/A sky130_fd_sc_hd__fa_2_546/B
+ sky130_fd_sc_hd__fa_2_564/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_191 sky130_fd_sc_hd__fa_2_683/CIN sky130_fd_sc_hd__ha_2_131/A
+ sky130_fd_sc_hd__ha_2_132/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_790 sky130_fd_sc_hd__nor2_1_148/A sky130_fd_sc_hd__nor2_1_149/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_790/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21o_2_17 sky130_fd_sc_hd__a21o_2_17/X sky130_fd_sc_hd__nor2_1_213/Y
+ sky130_fd_sc_hd__nor2_1_213/A sky130_fd_sc_hd__or3_1_3/X VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__a21o_2_28 sky130_fd_sc_hd__a21o_2_28/X sky130_fd_sc_hd__nor2_1_297/Y
+ sky130_fd_sc_hd__fa_2_19/SUM sky130_fd_sc_hd__nor2_1_297/B VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__xor2_1_11 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__xor2_1_11/X
+ sky130_fd_sc_hd__xor2_1_11/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_22 sky130_fd_sc_hd__xor2_1_22/B sky130_fd_sc_hd__maj3_1_3/B
+ sky130_fd_sc_hd__nor4_1_4/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_33 sky130_fd_sc_hd__xor2_1_34/X sky130_fd_sc_hd__xor2_1_33/X
+ sky130_fd_sc_hd__xor2_1_60/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_44 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_983/B
+ sky130_fd_sc_hd__xor2_1_44/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_55 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_972/B
+ sky130_fd_sc_hd__xor2_1_55/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_66 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__xor2_1_66/X
+ sky130_fd_sc_hd__xor2_1_66/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_77 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__fa_2_999/B
+ sky130_fd_sc_hd__xor2_1_77/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_88 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__xor2_1_88/X
+ sky130_fd_sc_hd__xor2_1_88/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_99 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__xor2_1_99/X
+ sky130_fd_sc_hd__xor2_1_99/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2b_1_5 sky130_fd_sc_hd__nand2b_1_5/Y sky130_fd_sc_hd__buf_2_263/X
+ sky130_fd_sc_hd__nor2_1_29/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a21o_2_1 sky130_fd_sc_hd__a21o_2_1/X sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__xor2_1_29/X sky130_fd_sc_hd__a21o_2_2/A2 VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__dfxtp_1_904 VDD VSS sky130_fd_sc_hd__fa_2_939/B sky130_fd_sc_hd__dfxtp_1_904/CLK
+ sky130_fd_sc_hd__o21a_1_19/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_915 VDD VSS sky130_fd_sc_hd__fa_2_1144/A sky130_fd_sc_hd__clkinv_8_55/Y
+ sky130_fd_sc_hd__mux2_2_110/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_926 VDD VSS sky130_fd_sc_hd__fa_2_1155/A sky130_fd_sc_hd__clkinv_8_46/Y
+ sky130_fd_sc_hd__mux2_2_82/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_937 VDD VSS sky130_fd_sc_hd__fa_2_1129/A sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__mux2_2_102/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_948 VDD VSS sky130_fd_sc_hd__xor2_1_164/A sky130_fd_sc_hd__clkinv_8_46/Y
+ sky130_fd_sc_hd__mux2_2_77/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_959 VDD VSS sky130_fd_sc_hd__fa_2_1168/A sky130_fd_sc_hd__clkinv_8_65/Y
+ sky130_fd_sc_hd__mux2_2_103/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a221oi_1_3 sky130_fd_sc_hd__a221oi_1_3/Y sky130_fd_sc_hd__o31ai_1_7/A2
+ sky130_fd_sc_hd__xor2_1_185/B sky130_fd_sc_hd__nand2_1_418/Y sky130_fd_sc_hd__o31ai_1_8/A3
+ sky130_fd_sc_hd__nor2_1_205/B VSS VDD VDD VSS sky130_fd_sc_hd__a221oi_1
Xsky130_fd_sc_hd__clkbuf_1_502 VSS VDD sky130_fd_sc_hd__buf_12_386/A sky130_fd_sc_hd__clkbuf_1_513/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_513 VSS VDD sky130_fd_sc_hd__clkbuf_1_513/X sky130_fd_sc_hd__buf_8_187/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_524 VSS VDD sky130_fd_sc_hd__clkbuf_1_524/X sky130_fd_sc_hd__clkbuf_1_524/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_535 VSS VDD sky130_fd_sc_hd__clkbuf_1_535/X sky130_fd_sc_hd__clkbuf_4_208/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_103 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_104/B sky130_fd_sc_hd__fa_2_233/CIN
+ sky130_fd_sc_hd__fa_2_225/A sky130_fd_sc_hd__fa_2_31/A sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_546 VSS VDD sky130_fd_sc_hd__fa_2_242/A sky130_fd_sc_hd__fa_2_87/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_114 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_114/A sky130_fd_sc_hd__fa_2_389/CIN
+ sky130_fd_sc_hd__fa_2_381/A sky130_fd_sc_hd__ha_2_114/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_557 VSS VDD sky130_fd_sc_hd__nand2_1_87/B sky130_fd_sc_hd__nand4_1_61/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_125 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_125/A sky130_fd_sc_hd__fa_2_551/B
+ sky130_fd_sc_hd__ha_2_125/SUM sky130_fd_sc_hd__ha_2_125/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_568 VSS VDD sky130_fd_sc_hd__a22oi_1_9/A1 sky130_fd_sc_hd__nor3_2_0/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_136 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_136/A sky130_fd_sc_hd__maj3_1_160/B
+ sky130_fd_sc_hd__maj3_1_161/A sky130_fd_sc_hd__ha_2_140/A sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_579 VSS VDD sky130_fd_sc_hd__nand3_1_11/B sky130_fd_sc_hd__a22oi_1_22/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_147 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_147/A sky130_fd_sc_hd__fa_2_863/CIN
+ sky130_fd_sc_hd__ha_2_147/SUM sky130_fd_sc_hd__ha_2_147/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_158 VSS VDD VSS VDD sky130_fd_sc_hd__or4_1_0/A sky130_fd_sc_hd__xor2_1_13/A
+ sky130_fd_sc_hd__ha_2_158/SUM sky130_fd_sc_hd__ha_2_158/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__fa_2_809 sky130_fd_sc_hd__fa_2_712/A sky130_fd_sc_hd__fa_2_713/B
+ sky130_fd_sc_hd__fa_2_809/A sky130_fd_sc_hd__fa_2_809/B sky130_fd_sc_hd__fa_2_815/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__ha_2_169 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_169/A sky130_fd_sc_hd__fa_2_928/A
+ sky130_fd_sc_hd__fa_2_929/B sky130_fd_sc_hd__ha_2_169/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__maj3_1_7 sky130_fd_sc_hd__maj3_1_8/X sky130_fd_sc_hd__maj3_1_7/X
+ sky130_fd_sc_hd__maj3_1_7/B sky130_fd_sc_hd__maj3_1_7/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__ha_2_60 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_60/A sky130_fd_sc_hd__xor2_1_6/A
+ sky130_fd_sc_hd__ha_2_60/SUM sky130_fd_sc_hd__ha_2_60/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_71 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_71/A sky130_fd_sc_hd__ha_2_70/B
+ sky130_fd_sc_hd__ha_2_71/SUM sky130_fd_sc_hd__ha_2_71/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_82 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_82/A sky130_fd_sc_hd__ha_2_81/B
+ sky130_fd_sc_hd__ha_2_82/SUM sky130_fd_sc_hd__ha_2_82/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__o22a_1_0 sky130_fd_sc_hd__o22a_1_0/A2 sky130_fd_sc_hd__o22a_1_0/X
+ sky130_fd_sc_hd__xor2_1_31/A sky130_fd_sc_hd__fa_2_944/A sky130_fd_sc_hd__o22a_1_0/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22a_1
Xsky130_fd_sc_hd__ha_2_93 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_93/A sky130_fd_sc_hd__fa_2_68/A
+ sky130_fd_sc_hd__ha_2_93/SUM sky130_fd_sc_hd__ha_2_99/A sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_1 VSS VDD sky130_fd_sc_hd__clkbuf_1_1/X sky130_fd_sc_hd__nand2b_1_0/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__mux2_2_109 VSS VDD sky130_fd_sc_hd__mux2_2_109/A1 sky130_fd_sc_hd__mux2_2_109/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_109/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__clkinv_1_1 sky130_fd_sc_hd__nor3_1_4/B sky130_fd_sc_hd__nor3_1_3/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_180 sky130_fd_sc_hd__o21a_1_29/A1 sky130_fd_sc_hd__nor2_1_180/Y
+ sky130_fd_sc_hd__nor2_1_180/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_191 sky130_fd_sc_hd__nor2_1_191/B sky130_fd_sc_hd__nor2_1_191/Y
+ sky130_fd_sc_hd__nor2_1_191/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__and2_0_16 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_16/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_13/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_27 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_27/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_34/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_307 sky130_fd_sc_hd__o22ai_1_322/A2 sky130_fd_sc_hd__o22ai_1_307/B1
+ sky130_fd_sc_hd__o22ai_1_307/Y sky130_fd_sc_hd__nor2_1_185/B sky130_fd_sc_hd__o32ai_1_5/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_38 VSS VDD VDD VSS sky130_fd_sc_hd__nand3_2_3/B sky130_fd_sc_hd__xor2_1_5/B
+ sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_318 sky130_fd_sc_hd__o22ai_1_318/A2 sky130_fd_sc_hd__nor2_1_195/B
+ sky130_fd_sc_hd__o22ai_1_318/Y sky130_fd_sc_hd__nor2_1_196/B sky130_fd_sc_hd__o32ai_1_5/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_49 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_50/A sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__ha_2_57/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_329 sky130_fd_sc_hd__nand2_1_462/Y sky130_fd_sc_hd__nand2_1_461/Y
+ sky130_fd_sc_hd__o22ai_1_329/Y sky130_fd_sc_hd__o22ai_1_342/A1 sky130_fd_sc_hd__a21o_2_20/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_2_8 sky130_fd_sc_hd__nor2_2_8/B sky130_fd_sc_hd__nor2_2_8/Y
+ sky130_fd_sc_hd__nor2_2_9/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__a22oi_1_290 sky130_fd_sc_hd__clkbuf_1_378/X sky130_fd_sc_hd__clkbuf_1_379/X
+ sky130_fd_sc_hd__clkbuf_4_170/X sky130_fd_sc_hd__buf_2_194/X sky130_fd_sc_hd__nand4_1_72/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_8_15 sky130_fd_sc_hd__buf_8_15/A sky130_fd_sc_hd__buf_8_15/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_26 sky130_fd_sc_hd__inv_2_3/A sky130_fd_sc_hd__buf_8_26/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_37 sky130_fd_sc_hd__inv_2_9/Y sky130_fd_sc_hd__buf_8_37/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_48 sky130_fd_sc_hd__buf_8_48/A sky130_fd_sc_hd__buf_8_48/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_59 sky130_fd_sc_hd__buf_8_59/A sky130_fd_sc_hd__buf_8_59/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__o21ai_1_501 VSS VDD sky130_fd_sc_hd__nand2_1_562/A sky130_fd_sc_hd__o21ai_1_507/A1
+ sky130_fd_sc_hd__nand2_1_562/Y sky130_fd_sc_hd__and2_0_349/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1107 VDD VSS sky130_fd_sc_hd__o32ai_1_5/A1 sky130_fd_sc_hd__clkinv_4_23/Y
+ sky130_fd_sc_hd__nor2b_1_116/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1118 VDD VSS sky130_fd_sc_hd__mux2_2_147/A0 sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__o22ai_1_275/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1129 VDD VSS sky130_fd_sc_hd__mux2_2_171/A0 sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__dfxtp_1_988/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_701 VDD VSS sky130_fd_sc_hd__mux2_2_33/A0 sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__o21ai_1_41/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_712 VDD VSS sky130_fd_sc_hd__mux2_2_9/A1 sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__o21ai_1_52/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_723 VDD VSS sky130_fd_sc_hd__mux2_2_26/A1 sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__o21ai_1_60/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_734 VDD VSS sky130_fd_sc_hd__mux2_2_4/A1 sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__o21ai_1_71/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_745 VDD VSS sky130_fd_sc_hd__and2_0_181/A sky130_fd_sc_hd__dfxtp_1_747/CLK
+ sky130_fd_sc_hd__fa_2_1100/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_756 VDD VSS sky130_fd_sc_hd__fa_2_672/A sky130_fd_sc_hd__dfxtp_1_764/CLK
+ sky130_fd_sc_hd__o21a_1_14/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_767 VDD VSS sky130_fd_sc_hd__fa_2_701/B sky130_fd_sc_hd__dfxtp_1_768/CLK
+ sky130_fd_sc_hd__o21a_1_9/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_778 VDD VSS sky130_fd_sc_hd__fa_2_1077/A sky130_fd_sc_hd__clkinv_8_55/Y
+ sky130_fd_sc_hd__mux2_2_70/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_789 VDD VSS sky130_fd_sc_hd__fa_2_1088/A sky130_fd_sc_hd__clkinv_8_45/Y
+ sky130_fd_sc_hd__mux2_2_46/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_310 VSS VDD sky130_fd_sc_hd__nand4_1_35/D sky130_fd_sc_hd__a22oi_1_159/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_321 VSS VDD sky130_fd_sc_hd__clkbuf_1_321/X sky130_fd_sc_hd__nand3_2_4/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_332 VSS VDD sky130_fd_sc_hd__buf_4_63/A sky130_fd_sc_hd__buf_4_122/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_343 VSS VDD sky130_fd_sc_hd__buf_8_136/A sky130_fd_sc_hd__and2_4_0/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_354 VSS VDD sky130_fd_sc_hd__buf_8_165/A sky130_fd_sc_hd__buf_4_84/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_365 VSS VDD sky130_fd_sc_hd__clkbuf_4_155/A sky130_fd_sc_hd__inv_8_0/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_376 VSS VDD sky130_fd_sc_hd__clkbuf_1_376/X sky130_fd_sc_hd__nor3_1_25/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_387 VSS VDD sky130_fd_sc_hd__a22oi_2_25/B2 sky130_fd_sc_hd__clkbuf_1_387/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_398 VSS VDD sky130_fd_sc_hd__clkbuf_1_398/X sky130_fd_sc_hd__clkbuf_1_398/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_606 sky130_fd_sc_hd__fa_2_608/B sky130_fd_sc_hd__fa_2_604/A
+ sky130_fd_sc_hd__fa_2_698/A sky130_fd_sc_hd__fa_2_689/B sky130_fd_sc_hd__fa_2_692/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_617 sky130_fd_sc_hd__fa_2_616/CIN sky130_fd_sc_hd__fa_2_617/SUM
+ sky130_fd_sc_hd__fa_2_701/B sky130_fd_sc_hd__fa_2_667/B sky130_fd_sc_hd__fa_2_678/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_628 sky130_fd_sc_hd__fa_2_627/A sky130_fd_sc_hd__fa_2_623/A
+ sky130_fd_sc_hd__fa_2_698/A sky130_fd_sc_hd__ha_2_130/A sky130_fd_sc_hd__fa_2_683/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_639 sky130_fd_sc_hd__fa_2_641/B sky130_fd_sc_hd__fa_2_639/SUM
+ sky130_fd_sc_hd__fa_2_639/A sky130_fd_sc_hd__fa_2_639/B sky130_fd_sc_hd__fa_2_643/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_80 VDD VSS sky130_fd_sc_hd__nand2_1_19/A sky130_fd_sc_hd__dfxtp_1_83/CLK
+ sky130_fd_sc_hd__o21a_1_0/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_91 VDD VSS sky130_fd_sc_hd__a22o_1_7/B2 sky130_fd_sc_hd__dfxtp_1_93/CLK
+ sky130_fd_sc_hd__dfxtp_1_91/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_330 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_330/X sky130_fd_sc_hd__inv_2_139/Y
+ sky130_fd_sc_hd__and2_0_330/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_170 sky130_fd_sc_hd__clkbuf_4_170/X sky130_fd_sc_hd__clkbuf_4_170/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_341 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_341/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_341/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_181 sky130_fd_sc_hd__clkbuf_4_181/X sky130_fd_sc_hd__clkbuf_4_181/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_352 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_352/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_352/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_192 sky130_fd_sc_hd__clkbuf_4_192/X sky130_fd_sc_hd__clkbuf_4_192/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__conb_1_5 sky130_fd_sc_hd__conb_1_5/LO sky130_fd_sc_hd__conb_1_5/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__inv_2_130 sky130_fd_sc_hd__inv_2_130/A sky130_fd_sc_hd__inv_2_130/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_141 sky130_fd_sc_hd__nor4_1_13/A sky130_fd_sc_hd__inv_2_141/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__o22ai_1_104 sky130_fd_sc_hd__o21a_1_8/A2 sky130_fd_sc_hd__nor2_1_64/B
+ sky130_fd_sc_hd__nor2_1_80/B sky130_fd_sc_hd__o22ai_1_110/B1 sky130_fd_sc_hd__o21ai_1_92/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_115 sky130_fd_sc_hd__o22ai_1_130/B1 sky130_fd_sc_hd__nor2_1_70/B
+ sky130_fd_sc_hd__nor2_1_83/A sky130_fd_sc_hd__nor2_1_70/A sky130_fd_sc_hd__o22ai_1_132/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_126 sky130_fd_sc_hd__a21oi_1_119/Y sky130_fd_sc_hd__nor2_1_76/A
+ sky130_fd_sc_hd__o22ai_1_126/Y sky130_fd_sc_hd__nor2_2_9/B sky130_fd_sc_hd__a211oi_1_7/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_137 sky130_fd_sc_hd__nand2_1_284/Y sky130_fd_sc_hd__nand2_2_5/Y
+ sky130_fd_sc_hd__o22ai_1_137/Y sky130_fd_sc_hd__xnor2_1_66/Y sky130_fd_sc_hd__o22ai_1_151/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_148 sky130_fd_sc_hd__nand2_1_284/Y sky130_fd_sc_hd__nand2_2_5/Y
+ sky130_fd_sc_hd__o22ai_1_148/Y sky130_fd_sc_hd__xnor2_1_88/Y sky130_fd_sc_hd__o22ai_1_162/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_159 sky130_fd_sc_hd__nand2_1_338/A sky130_fd_sc_hd__nand2_1_284/Y
+ sky130_fd_sc_hd__o22ai_1_159/Y sky130_fd_sc_hd__xnor2_1_82/Y sky130_fd_sc_hd__o22ai_1_159/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_2_15 sky130_fd_sc_hd__nor2_2_15/B sky130_fd_sc_hd__nor2_2_15/Y
+ sky130_fd_sc_hd__nor2_2_15/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__nand4_1_18 sky130_fd_sc_hd__nand4_1_18/C sky130_fd_sc_hd__nand4_1_18/B
+ sky130_fd_sc_hd__nand4_1_18/Y sky130_fd_sc_hd__nand4_1_18/D sky130_fd_sc_hd__buf_2_110/X
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__o211ai_1_5 sky130_fd_sc_hd__a21oi_1_95/Y sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__xor2_1_66/A sky130_fd_sc_hd__o211ai_1_5/C1 sky130_fd_sc_hd__o211ai_1_5/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__nand4_1_29 sky130_fd_sc_hd__nand4_1_29/C sky130_fd_sc_hd__nand4_1_29/B
+ sky130_fd_sc_hd__nand4_1_29/Y sky130_fd_sc_hd__nand4_1_29/D sky130_fd_sc_hd__buf_2_102/X
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__nand3b_2_0 sky130_fd_sc_hd__nor2_4_2/A sky130_fd_sc_hd__nor3_1_0/A
+ sky130_fd_sc_hd__nor4_1_0/A sky130_fd_sc_hd__nor4_1_0/B VSS VDD VSS VDD sky130_fd_sc_hd__nand3b_2
Xsky130_fd_sc_hd__a31oi_1_2 VSS VDD sky130_fd_sc_hd__a31oi_1_2/Y sky130_fd_sc_hd__o22ai_1_60/Y
+ sky130_fd_sc_hd__a31oi_1_2/A2 sky130_fd_sc_hd__a221o_1_0/X sky130_fd_sc_hd__nand2b_1_9/Y
+ VDD VSS sky130_fd_sc_hd__a31oi_1
Xsky130_fd_sc_hd__o21ai_1_320 VSS VDD sky130_fd_sc_hd__o21a_1_29/X sky130_fd_sc_hd__nor2_1_180/A
+ sky130_fd_sc_hd__a21oi_1_289/Y sky130_fd_sc_hd__xor2_1_156/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_331 VSS VDD sky130_fd_sc_hd__nand2_1_419/B sky130_fd_sc_hd__nor2_1_208/Y
+ sky130_fd_sc_hd__o31ai_1_8/A2 sky130_fd_sc_hd__o21ai_1_331/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_342 VSS VDD sky130_fd_sc_hd__o22ai_1_301/A1 sky130_fd_sc_hd__nor2_1_224/A
+ sky130_fd_sc_hd__nand2_1_425/Y sky130_fd_sc_hd__xor2_1_210/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_353 VSS VDD sky130_fd_sc_hd__a222oi_1_17/Y sky130_fd_sc_hd__nor2_1_224/A
+ sky130_fd_sc_hd__a22oi_1_381/Y sky130_fd_sc_hd__o21ai_1_353/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a211oi_1_14 sky130_fd_sc_hd__nor2_2_15/Y sky130_fd_sc_hd__nor2_1_176/Y
+ sky130_fd_sc_hd__o22ai_1_250/Y sky130_fd_sc_hd__nor2_1_175/B sky130_fd_sc_hd__fa_2_1136/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_364 VSS VDD sky130_fd_sc_hd__a222oi_1_20/Y sky130_fd_sc_hd__nor2_1_224/A
+ sky130_fd_sc_hd__nand2_1_434/Y sky130_fd_sc_hd__xor2_1_190/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a211oi_1_25 sky130_fd_sc_hd__nor2_1_267/Y sky130_fd_sc_hd__nor2_1_257/Y
+ sky130_fd_sc_hd__nor2_1_258/Y sky130_fd_sc_hd__a211oi_1_25/Y sky130_fd_sc_hd__fa_2_1233/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_375 VSS VDD sky130_fd_sc_hd__a222oi_1_21/Y sky130_fd_sc_hd__nor2_1_224/A
+ sky130_fd_sc_hd__a22oi_1_385/Y sky130_fd_sc_hd__o21ai_1_375/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a211oi_1_36 sky130_fd_sc_hd__nor2b_1_126/Y sky130_fd_sc_hd__nor2_1_306/Y
+ sky130_fd_sc_hd__o21ai_1_487/Y sky130_fd_sc_hd__a211oi_1_36/Y sky130_fd_sc_hd__o21ai_1_488/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_386 VSS VDD sky130_fd_sc_hd__nand2_1_472/B sky130_fd_sc_hd__nor2_1_252/Y
+ sky130_fd_sc_hd__nor2_1_251/B sky130_fd_sc_hd__o21ai_1_386/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_397 VSS VDD sky130_fd_sc_hd__a222oi_1_26/Y sky130_fd_sc_hd__nor2_1_267/A
+ sky130_fd_sc_hd__nand2_1_477/Y sky130_fd_sc_hd__xor2_1_256/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__mux2_2_11 VSS VDD sky130_fd_sc_hd__mux2_2_11/A1 sky130_fd_sc_hd__mux2_2_11/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_11/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_22 VSS VDD sky130_fd_sc_hd__mux2_2_22/A1 sky130_fd_sc_hd__mux2_2_22/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_22/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_33 VSS VDD sky130_fd_sc_hd__mux2_2_33/A1 sky130_fd_sc_hd__mux2_2_33/A0
+ sky130_fd_sc_hd__mux2_2_37/S sky130_fd_sc_hd__mux2_2_33/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_44 VSS VDD sky130_fd_sc_hd__mux2_2_44/A1 sky130_fd_sc_hd__mux2_2_44/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_44/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_55 VSS VDD sky130_fd_sc_hd__mux2_2_55/A1 sky130_fd_sc_hd__mux2_2_55/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_55/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_66 VSS VDD sky130_fd_sc_hd__mux2_2_66/A1 sky130_fd_sc_hd__xor2_1_138/X
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_66/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_77 VSS VDD sky130_fd_sc_hd__mux2_2_77/A1 sky130_fd_sc_hd__xor2_1_141/X
+ sky130_fd_sc_hd__nor2_4_15/A sky130_fd_sc_hd__mux2_2_77/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_88 VSS VDD sky130_fd_sc_hd__mux2_2_88/A1 sky130_fd_sc_hd__mux2_2_88/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_88/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1107 sky130_fd_sc_hd__fa_2_1108/CIN sky130_fd_sc_hd__fa_2_1107/SUM
+ sky130_fd_sc_hd__fa_2_1107/A sky130_fd_sc_hd__fa_2_1107/B sky130_fd_sc_hd__ha_2_201/COUT
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__mux2_2_99 VSS VDD sky130_fd_sc_hd__mux2_2_99/A1 sky130_fd_sc_hd__mux2_2_99/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_99/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1118 sky130_fd_sc_hd__fa_2_1119/CIN sky130_fd_sc_hd__fa_2_1118/SUM
+ sky130_fd_sc_hd__fa_2_1118/A sky130_fd_sc_hd__fa_2_1118/B sky130_fd_sc_hd__fa_2_1118/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1129 sky130_fd_sc_hd__fa_2_1130/CIN sky130_fd_sc_hd__mux2_2_102/A1
+ sky130_fd_sc_hd__fa_2_1129/A sky130_fd_sc_hd__fa_2_1129/B sky130_fd_sc_hd__fa_2_1129/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_520 VDD VSS sky130_fd_sc_hd__nor4_1_10/D sky130_fd_sc_hd__dfxtp_1_520/CLK
+ sky130_fd_sc_hd__and2_0_256/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_180 sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__fa_2_1142/B
+ sky130_fd_sc_hd__xor2_1_180/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_191 sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__fa_2_1188/B
+ sky130_fd_sc_hd__xor2_1_191/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_531 VDD VSS sky130_fd_sc_hd__fa_2_960/A sky130_fd_sc_hd__dfxtp_1_533/CLK
+ sky130_fd_sc_hd__and2_0_259/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_542 VDD VSS sky130_fd_sc_hd__fa_2_949/A sky130_fd_sc_hd__dfxtp_1_544/CLK
+ sky130_fd_sc_hd__a22o_1_43/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_553 VDD VSS sky130_fd_sc_hd__and2_0_223/A sky130_fd_sc_hd__dfxtp_1_571/CLK
+ sky130_fd_sc_hd__dfxtp_1_554/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_564 VDD VSS sky130_fd_sc_hd__dfxtp_1_564/Q sky130_fd_sc_hd__dfxtp_1_594/CLK
+ sky130_fd_sc_hd__dfxtp_1_564/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_575 VDD VSS sky130_fd_sc_hd__and2_0_201/A sky130_fd_sc_hd__dfxtp_1_577/CLK
+ sky130_fd_sc_hd__dfxtp_1_576/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_586 VDD VSS sky130_fd_sc_hd__nor4_1_8/D sky130_fd_sc_hd__dfxtp_1_591/CLK
+ sky130_fd_sc_hd__and2_0_244/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_597 VDD VSS sky130_fd_sc_hd__and2_0_207/A sky130_fd_sc_hd__dfxtp_1_601/CLK
+ sky130_fd_sc_hd__fa_2_1017/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_140 VSS VDD sky130_fd_sc_hd__clkbuf_1_140/X sky130_fd_sc_hd__clkbuf_1_140/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_151 VSS VDD sky130_fd_sc_hd__a22oi_1_96/B2 sky130_fd_sc_hd__clkbuf_1_151/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_162 VSS VDD sky130_fd_sc_hd__clkbuf_1_162/X sky130_fd_sc_hd__clkbuf_1_162/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_173 VSS VDD sky130_fd_sc_hd__clkbuf_1_173/X sky130_fd_sc_hd__nand3_1_28/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_184 VSS VDD sky130_fd_sc_hd__nand4_1_22/B sky130_fd_sc_hd__a22oi_1_110/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_195 VSS VDD sky130_fd_sc_hd__clkbuf_1_196/A sky130_fd_sc_hd__clkbuf_4_95/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_403 sky130_fd_sc_hd__fa_2_406/B sky130_fd_sc_hd__fa_2_403/SUM
+ sky130_fd_sc_hd__fa_2_403/A sky130_fd_sc_hd__fa_2_403/B sky130_fd_sc_hd__fa_2_403/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_414 sky130_fd_sc_hd__maj3_1_56/B sky130_fd_sc_hd__maj3_1_57/A
+ sky130_fd_sc_hd__fa_2_414/A sky130_fd_sc_hd__fa_2_414/B sky130_fd_sc_hd__fa_2_415/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_425 sky130_fd_sc_hd__fa_2_423/A sky130_fd_sc_hd__fa_2_425/SUM
+ sky130_fd_sc_hd__fa_2_425/A sky130_fd_sc_hd__fa_2_425/B sky130_fd_sc_hd__fa_2_404/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_436 sky130_fd_sc_hd__fa_2_433/A sky130_fd_sc_hd__fa_2_426/B
+ sky130_fd_sc_hd__fa_2_531/B sky130_fd_sc_hd__fa_2_436/B sky130_fd_sc_hd__fa_2_439/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_447 sky130_fd_sc_hd__fa_2_444/B sky130_fd_sc_hd__fa_2_446/B
+ sky130_fd_sc_hd__ha_2_125/B sky130_fd_sc_hd__ha_2_122/B sky130_fd_sc_hd__fa_2_555/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_458 sky130_fd_sc_hd__fa_2_455/B sky130_fd_sc_hd__fa_2_459/CIN
+ sky130_fd_sc_hd__fa_2_458/A sky130_fd_sc_hd__fa_2_458/B sky130_fd_sc_hd__fa_2_458/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_469 sky130_fd_sc_hd__maj3_1_103/B sky130_fd_sc_hd__maj3_1_104/A
+ sky130_fd_sc_hd__fa_2_535/A sky130_fd_sc_hd__fa_2_469/B sky130_fd_sc_hd__fa_2_470/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nand3_1_40 sky130_fd_sc_hd__nand3_1_40/Y sky130_fd_sc_hd__a22o_1_28/X
+ sky130_fd_sc_hd__nand3_2_8/C sky130_fd_sc_hd__or2_1_1/X VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_51 sky130_fd_sc_hd__nand3_1_51/Y sky130_fd_sc_hd__nand3_1_51/A
+ sky130_fd_sc_hd__nand3_1_51/C sky130_fd_sc_hd__nand3_1_52/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__dfxtp_1_1460 VDD VSS sky130_fd_sc_hd__buf_2_143/A sky130_fd_sc_hd__dfxtp_1_1461/CLK
+ sky130_fd_sc_hd__and2_0_341/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_160 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_160/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__ha_2_159/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_171 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_171/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__fa_2_862/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_182 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_182/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_182/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_90 sky130_fd_sc_hd__buf_8_66/A sky130_fd_sc_hd__inv_2_56/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_90/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_193 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_193/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_900/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_408 sky130_fd_sc_hd__buf_8_203/X sky130_fd_sc_hd__buf_6_82/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_419 sky130_fd_sc_hd__buf_12_419/A sky130_fd_sc_hd__buf_12_481/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__fa_2_970 sky130_fd_sc_hd__fa_2_971/CIN sky130_fd_sc_hd__fa_2_970/SUM
+ sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_970/B sky130_fd_sc_hd__xor2_1_57/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_981 sky130_fd_sc_hd__fa_2_982/CIN sky130_fd_sc_hd__mux2_2_25/A0
+ sky130_fd_sc_hd__fa_2_981/A sky130_fd_sc_hd__fa_2_981/B sky130_fd_sc_hd__fa_2_981/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_992 sky130_fd_sc_hd__xor2_1_32/B sky130_fd_sc_hd__mux2_2_3/A0
+ sky130_fd_sc_hd__fa_2_992/A sky130_fd_sc_hd__fa_2_992/B sky130_fd_sc_hd__fa_2_992/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_1_608 sky130_fd_sc_hd__ha_2_184/B sky130_fd_sc_hd__fa_2_1031/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_608/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_619 sky130_fd_sc_hd__o21ai_1_274/A2 sky130_fd_sc_hd__fa_2_1076/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_619/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o21ai_1_150 VSS VDD sky130_fd_sc_hd__nor2_1_76/A sky130_fd_sc_hd__a21oi_1_129/Y
+ sky130_fd_sc_hd__a21oi_1_125/Y sky130_fd_sc_hd__xor2_1_56/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_161 VSS VDD sky130_fd_sc_hd__o21ai_1_171/A2 sky130_fd_sc_hd__xnor2_1_69/Y
+ sky130_fd_sc_hd__a21oi_1_138/Y sky130_fd_sc_hd__o21ai_1_161/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_172 VSS VDD sky130_fd_sc_hd__o21ai_1_189/A2 sky130_fd_sc_hd__nand2_2_5/Y
+ sky130_fd_sc_hd__a21oi_1_149/Y sky130_fd_sc_hd__o21ai_1_172/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_183 VSS VDD sky130_fd_sc_hd__nand2_2_5/Y sky130_fd_sc_hd__xnor2_1_79/Y
+ sky130_fd_sc_hd__a21oi_1_158/Y sky130_fd_sc_hd__o21ai_1_183/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_194 VSS VDD sky130_fd_sc_hd__xnor2_1_81/A sky130_fd_sc_hd__o21ai_1_194/A1
+ sky130_fd_sc_hd__nand2_1_291/B sky130_fd_sc_hd__xnor2_1_83/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_17 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1177/A sky130_fd_sc_hd__nor2_2_16/Y
+ sky130_fd_sc_hd__nor3_1_39/A sky130_fd_sc_hd__fa_2_1179/A sky130_fd_sc_hd__nor3_1_39/B
+ sky130_fd_sc_hd__a222oi_1_17/Y sky130_fd_sc_hd__fa_2_1176/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_28 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1227/A sky130_fd_sc_hd__nor2_2_17/Y
+ sky130_fd_sc_hd__nor3_1_40/A sky130_fd_sc_hd__fa_2_1229/A sky130_fd_sc_hd__nor3_1_40/B
+ sky130_fd_sc_hd__a222oi_1_28/Y sky130_fd_sc_hd__fa_2_1226/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_39 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1277/A sky130_fd_sc_hd__nor2_2_18/Y
+ sky130_fd_sc_hd__nor3_1_41/A sky130_fd_sc_hd__fa_2_1279/A sky130_fd_sc_hd__nor3_1_41/B
+ sky130_fd_sc_hd__a222oi_1_39/Y sky130_fd_sc_hd__fa_2_1276/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2_1_510 sky130_fd_sc_hd__o21a_1_67/B1 sky130_fd_sc_hd__fa_2_1298/A
+ sky130_fd_sc_hd__o21a_1_67/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_521 sky130_fd_sc_hd__nand2_1_521/Y sky130_fd_sc_hd__inv_2_140/Y
+ sky130_fd_sc_hd__nand2_1_521/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_532 sky130_fd_sc_hd__nand2_1_532/Y sky130_fd_sc_hd__nor2b_2_5/A
+ sky130_fd_sc_hd__xor2_1_299/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__xnor2_1_19 VSS VDD sky130_fd_sc_hd__nor2_1_21/B sky130_fd_sc_hd__xnor2_1_19/Y
+ sky130_fd_sc_hd__nor2_1_21/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__nand2_1_543 sky130_fd_sc_hd__nand2_1_543/Y sky130_fd_sc_hd__nand2_1_543/B
+ sky130_fd_sc_hd__o21ai_1_478/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_554 sky130_fd_sc_hd__nand2_1_554/Y sky130_fd_sc_hd__buf_6_50/A
+ sky130_fd_sc_hd__nand2_1_554/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_565 sky130_fd_sc_hd__nand2_1_565/Y sky130_fd_sc_hd__buf_6_85/X
+ sky130_fd_sc_hd__nand2_1_565/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_1 sky130_fd_sc_hd__nor2_2_0/Y sky130_fd_sc_hd__nor2b_1_1/Y
+ sky130_fd_sc_hd__inv_2_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1101 sky130_fd_sc_hd__nor2_1_310/B sky130_fd_sc_hd__o21ai_1_490/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1101/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1112 sky130_fd_sc_hd__nor2_1_311/A sky130_fd_sc_hd__nor2_1_312/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1112/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1123 sky130_fd_sc_hd__inv_8_1/A sky130_fd_sc_hd__buf_6_86/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1123/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1134 sky130_fd_sc_hd__dfxtp_1_84/D sky130_fd_sc_hd__clkinv_1_1134/A
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_350 VDD VSS sky130_fd_sc_hd__a22o_1_23/B2 sky130_fd_sc_hd__dfxtp_1_354/CLK
+ sky130_fd_sc_hd__ha_2_152/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_361 VDD VSS sky130_fd_sc_hd__xor2_1_17/A sky130_fd_sc_hd__dfxtp_1_361/CLK
+ sky130_fd_sc_hd__dfxtp_1_361/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_372 VDD VSS sky130_fd_sc_hd__fa_2_1116/A sky130_fd_sc_hd__dfxtp_1_391/CLK
+ sky130_fd_sc_hd__and2_0_129/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_383 VDD VSS sky130_fd_sc_hd__fa_2_1111/B sky130_fd_sc_hd__clkinv_4_32/Y
+ sky130_fd_sc_hd__and2_0_150/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_3 sky130_fd_sc_hd__nand3_1_3/C sky130_fd_sc_hd__nand2_1_3/B
+ sky130_fd_sc_hd__nand2_1_9/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_394 VDD VSS sky130_fd_sc_hd__ha_2_185/A sky130_fd_sc_hd__dfxtp_1_411/CLK
+ sky130_fd_sc_hd__and2_0_233/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_200 sky130_fd_sc_hd__fa_2_198/B sky130_fd_sc_hd__fa_2_193/A
+ sky130_fd_sc_hd__fa_2_2/A sky130_fd_sc_hd__ha_2_93/A sky130_fd_sc_hd__fa_2_281/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_211 sky130_fd_sc_hd__maj3_1_41/B sky130_fd_sc_hd__maj3_1_42/A
+ sky130_fd_sc_hd__fa_2_211/A sky130_fd_sc_hd__fa_2_211/B sky130_fd_sc_hd__fa_2_212/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_222 sky130_fd_sc_hd__fa_2_219/B sky130_fd_sc_hd__fa_2_222/SUM
+ sky130_fd_sc_hd__fa_2_32/A sky130_fd_sc_hd__fa_2_261/A sky130_fd_sc_hd__fa_2_274/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_233 sky130_fd_sc_hd__fa_2_235/CIN sky130_fd_sc_hd__fa_2_227/B
+ sky130_fd_sc_hd__fa_2_280/A sky130_fd_sc_hd__fa_2_266/B sky130_fd_sc_hd__fa_2_233/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_244 sky130_fd_sc_hd__fa_2_246/CIN sky130_fd_sc_hd__fa_2_240/A
+ sky130_fd_sc_hd__fa_2_283/A sky130_fd_sc_hd__fa_2_244/B sky130_fd_sc_hd__fa_2_244/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_255 sky130_fd_sc_hd__maj3_1_32/B sky130_fd_sc_hd__maj3_1_33/A
+ sky130_fd_sc_hd__fa_2_255/A sky130_fd_sc_hd__fa_2_255/B sky130_fd_sc_hd__fa_2_256/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_266 sky130_fd_sc_hd__fa_2_267/A sky130_fd_sc_hd__fa_2_263/A
+ sky130_fd_sc_hd__fa_2_280/B sky130_fd_sc_hd__fa_2_266/B sky130_fd_sc_hd__fa_2_266/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_277 sky130_fd_sc_hd__fa_2_276/B sky130_fd_sc_hd__fa_2_277/SUM
+ sky130_fd_sc_hd__fa_2_277/A sky130_fd_sc_hd__fa_2_277/B sky130_fd_sc_hd__fa_2_283/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_288 sky130_fd_sc_hd__fa_2_287/CIN sky130_fd_sc_hd__fa_2_288/SUM
+ sky130_fd_sc_hd__fa_2_288/A sky130_fd_sc_hd__fa_2_288/B sky130_fd_sc_hd__fa_2_288/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_4 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_4/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__fa_2_299 sky130_fd_sc_hd__fa_2_290/B sky130_fd_sc_hd__fa_2_292/B
+ sky130_fd_sc_hd__ha_2_115/A sky130_fd_sc_hd__ha_2_115/B sky130_fd_sc_hd__fa_2_401/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__diode_2_105 sky130_fd_sc_hd__inv_2_135/Y VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_116 sky130_fd_sc_hd__buf_2_225/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_127 sky130_fd_sc_hd__buf_2_250/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_138 sky130_fd_sc_hd__clkbuf_1_526/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__fa_2_80 sky130_fd_sc_hd__fa_2_77/B sky130_fd_sc_hd__fa_2_80/SUM
+ sky130_fd_sc_hd__ha_2_95/A sky130_fd_sc_hd__fa_2_80/B sky130_fd_sc_hd__fa_2_81/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__diode_2_149 sky130_fd_sc_hd__buf_2_192/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__fa_2_91 sky130_fd_sc_hd__fa_2_93/CIN sky130_fd_sc_hd__fa_2_85/B
+ sky130_fd_sc_hd__fa_2_91/A sky130_fd_sc_hd__fa_2_91/B sky130_fd_sc_hd__fa_2_91/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_250 VDD VSS sky130_fd_sc_hd__buf_2_250/X sky130_fd_sc_hd__buf_2_250/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_261 VDD VSS sky130_fd_sc_hd__fa_2_15/B sky130_fd_sc_hd__ha_2_97/B
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_272 VDD VSS sky130_fd_sc_hd__buf_2_272/X sky130_fd_sc_hd__nor2_2_19/Y
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_283 VDD VSS serial_out sky130_fd_sc_hd__buf_2_283/A VDD VSS
+ sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1290 VDD VSS sky130_fd_sc_hd__mux2_2_194/A0 sky130_fd_sc_hd__clkinv_8_75/Y
+ sky130_fd_sc_hd__o22ai_1_345/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a21oi_1_30 sky130_fd_sc_hd__nor2_1_41/Y sky130_fd_sc_hd__o22ai_1_63/Y
+ sky130_fd_sc_hd__a21oi_1_30/Y sky130_fd_sc_hd__fa_2_1033/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_41 sky130_fd_sc_hd__nor2_1_41/Y sky130_fd_sc_hd__o22ai_1_74/Y
+ sky130_fd_sc_hd__a21oi_1_41/Y sky130_fd_sc_hd__fa_2_1044/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_205 sky130_fd_sc_hd__buf_4_50/X sky130_fd_sc_hd__buf_12_205/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_52 sky130_fd_sc_hd__nor2_2_6/Y sky130_fd_sc_hd__o22ai_1_84/Y
+ sky130_fd_sc_hd__a21oi_1_52/Y sky130_fd_sc_hd__fa_2_1040/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_216 sky130_fd_sc_hd__buf_6_25/X sky130_fd_sc_hd__buf_12_216/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_63 sky130_fd_sc_hd__a21oi_1_63/A1 sky130_fd_sc_hd__nor2_1_44/B
+ sky130_fd_sc_hd__xnor2_1_44/A sky130_fd_sc_hd__xnor2_1_42/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_227 sky130_fd_sc_hd__buf_12_227/A sky130_fd_sc_hd__buf_12_258/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_74 sky130_fd_sc_hd__o21a_1_3/B1 sky130_fd_sc_hd__o21a_1_2/A1
+ sky130_fd_sc_hd__a21oi_1_74/Y sky130_fd_sc_hd__nor2_1_64/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_238 sky130_fd_sc_hd__buf_12_238/A sky130_fd_sc_hd__buf_12_238/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_85 sky130_fd_sc_hd__a21oi_1_85/A1 sky130_fd_sc_hd__a21oi_1_85/B1
+ sky130_fd_sc_hd__a21oi_1_85/Y sky130_fd_sc_hd__a211o_1_6/A1 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_249 sky130_fd_sc_hd__buf_12_249/A sky130_fd_sc_hd__buf_12_249/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_96 sky130_fd_sc_hd__a21oi_1_96/A1 sky130_fd_sc_hd__o22ai_1_99/Y
+ sky130_fd_sc_hd__a21oi_1_96/Y sky130_fd_sc_hd__a211o_1_6/A1 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_1_108 sky130_fd_sc_hd__a22oi_1_96/B1 sky130_fd_sc_hd__a22oi_1_96/A1
+ sky130_fd_sc_hd__clkbuf_1_148/X sky130_fd_sc_hd__a22oi_1_108/A2 sky130_fd_sc_hd__nand4_1_22/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_119 sky130_fd_sc_hd__clkbuf_4_72/X sky130_fd_sc_hd__clkbuf_4_73/X
+ sky130_fd_sc_hd__a22oi_1_119/B2 sky130_fd_sc_hd__buf_2_89/X sky130_fd_sc_hd__clkbuf_4_91/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor3_1_0 sky130_fd_sc_hd__inv_2_1/Y sky130_fd_sc_hd__nor3_1_0/Y
+ sky130_fd_sc_hd__nor3_1_0/A sky130_fd_sc_hd__or2_0_0/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__clkinv_1_405 sky130_fd_sc_hd__nand2_1_212/B sky130_fd_sc_hd__nor4_1_6/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_405/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_416 sky130_fd_sc_hd__nor3_1_34/A sky130_fd_sc_hd__dfxtp_1_502/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_416/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_427 sky130_fd_sc_hd__nor3_1_37/A sky130_fd_sc_hd__dfxtp_1_480/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_427/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_438 sky130_fd_sc_hd__fa_2_969/B sky130_fd_sc_hd__o21ai_1_38/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_438/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_449 sky130_fd_sc_hd__fa_2_952/B sky130_fd_sc_hd__nand2b_1_7/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_449/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_6_70 VDD VSS sky130_fd_sc_hd__buf_6_70/X sky130_fd_sc_hd__buf_6_70/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_81 VDD VSS sky130_fd_sc_hd__buf_6_81/X sky130_fd_sc_hd__buf_6_81/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__a21oi_1_302 sky130_fd_sc_hd__o21a_1_32/B1 sky130_fd_sc_hd__o21a_1_31/A1
+ sky130_fd_sc_hd__a21oi_1_302/Y sky130_fd_sc_hd__nor2_1_185/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_313 sky130_fd_sc_hd__nor2_1_196/A sky130_fd_sc_hd__o21a_1_40/A1
+ sky130_fd_sc_hd__a21oi_1_313/Y sky130_fd_sc_hd__nor2_1_196/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_324 sky130_fd_sc_hd__clkinv_1_902/Y sky130_fd_sc_hd__clkinv_1_901/Y
+ sky130_fd_sc_hd__a21oi_1_324/Y sky130_fd_sc_hd__nand2_1_439/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_50 sky130_fd_sc_hd__buf_2_75/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_335 sky130_fd_sc_hd__fa_2_1181/A sky130_fd_sc_hd__o22ai_1_303/Y
+ sky130_fd_sc_hd__a21oi_1_335/Y sky130_fd_sc_hd__nor2_2_16/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_61 sky130_fd_sc_hd__buf_2_102/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_346 sky130_fd_sc_hd__o21ai_1_376/Y sky130_fd_sc_hd__o21ai_1_371/Y
+ sky130_fd_sc_hd__a21oi_1_346/Y sky130_fd_sc_hd__nor2b_1_112/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_72 sky130_fd_sc_hd__clkbuf_4_86/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_357 sky130_fd_sc_hd__clkinv_1_861/Y sky130_fd_sc_hd__o22ai_1_320/Y
+ sky130_fd_sc_hd__a21oi_1_357/Y sky130_fd_sc_hd__fa_2_1206/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_83 sky130_fd_sc_hd__nand4_1_45/B VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_368 sky130_fd_sc_hd__nor2_1_234/A sky130_fd_sc_hd__nor2_1_234/Y
+ sky130_fd_sc_hd__a21oi_1_368/Y sky130_fd_sc_hd__nor2_1_234/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_94 sky130_fd_sc_hd__clkbuf_1_535/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_379 sky130_fd_sc_hd__or3_1_4/C sky130_fd_sc_hd__o21ai_1_392/Y
+ sky130_fd_sc_hd__a21oi_1_379/Y sky130_fd_sc_hd__nor2_1_248/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a222oi_1_5 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1123/A sky130_fd_sc_hd__nor2_2_15/Y
+ sky130_fd_sc_hd__nor3_1_38/A sky130_fd_sc_hd__fa_2_1125/A sky130_fd_sc_hd__nor3_1_38/B
+ sky130_fd_sc_hd__a222oi_1_5/Y sky130_fd_sc_hd__fa_2_1122/B sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2_1_340 sky130_fd_sc_hd__o32ai_1_2/A3 sky130_fd_sc_hd__nor2_2_15/A
+ sky130_fd_sc_hd__nor2_2_14/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_351 sky130_fd_sc_hd__o21a_1_25/B1 sky130_fd_sc_hd__fa_2_1152/A
+ sky130_fd_sc_hd__o21a_1_25/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_950 sky130_fd_sc_hd__o22ai_1_379/A2 sky130_fd_sc_hd__nor3_1_40/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_950/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_362 sky130_fd_sc_hd__nand2_1_362/Y sky130_fd_sc_hd__mux2_2_99/S
+ sky130_fd_sc_hd__nand2_1_362/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_961 sky130_fd_sc_hd__nor2_1_241/A sky130_fd_sc_hd__nor2_1_242/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_961/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_373 sky130_fd_sc_hd__nand2_1_373/Y sky130_fd_sc_hd__xor2_1_164/A
+ sky130_fd_sc_hd__nor2_1_182/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_972 sky130_fd_sc_hd__nor2_1_245/A sky130_fd_sc_hd__xnor2_1_99/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_972/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_384 sky130_fd_sc_hd__nand2_1_384/Y sky130_fd_sc_hd__nand2_1_387/B
+ sky130_fd_sc_hd__o21ai_1_323/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_983 sky130_fd_sc_hd__nand2_1_474/B sky130_fd_sc_hd__fa_2_143/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_983/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_395 sky130_fd_sc_hd__o21a_1_31/B1 sky130_fd_sc_hd__fa_2_1187/A
+ sky130_fd_sc_hd__o21a_1_31/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_994 sky130_fd_sc_hd__nor2_1_261/A sky130_fd_sc_hd__fa_2_1239/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_994/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand3_4_1 sky130_fd_sc_hd__nand3_4_1/Y sky130_fd_sc_hd__nand3_4_1/A
+ sky130_fd_sc_hd__nand3_4_1/B sky130_fd_sc_hd__nand3_4_1/C VSS VDD VSS VDD sky130_fd_sc_hd__nand3_4
Xsky130_fd_sc_hd__dfxtp_1_180 VDD VSS sky130_fd_sc_hd__ha_2_54/A sky130_fd_sc_hd__dfxtp_1_182/CLK
+ sky130_fd_sc_hd__and2_0_60/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_191 VDD VSS sky130_fd_sc_hd__ha_2_65/A sky130_fd_sc_hd__dfxtp_1_195/CLK
+ sky130_fd_sc_hd__nor2b_1_31/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_2_17 VDD VSS sky130_fd_sc_hd__buf_8_43/A sky130_fd_sc_hd__buf_2_33/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_28 VDD VSS sky130_fd_sc_hd__buf_8_49/A sky130_fd_sc_hd__ha_2_15/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_39 VDD VSS sky130_fd_sc_hd__buf_2_39/X sky130_fd_sc_hd__buf_2_39/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__a21boi_1_1 sky130_fd_sc_hd__a21boi_1_1/Y sky130_fd_sc_hd__nor2_2_15/Y
+ sky130_fd_sc_hd__a21oi_1_268/Y sky130_fd_sc_hd__fa_2_1135/A VDD VSS VDD VSS sky130_fd_sc_hd__a21boi_1
Xsky130_fd_sc_hd__o211ai_1_11 sky130_fd_sc_hd__nor2_1_74/A sky130_fd_sc_hd__o22ai_1_92/A1
+ sky130_fd_sc_hd__xor2_1_39/A sky130_fd_sc_hd__nand2_1_274/Y sky130_fd_sc_hd__nand2_1_277/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_22 sky130_fd_sc_hd__nor2_1_127/A sky130_fd_sc_hd__a222oi_1_3/Y
+ sky130_fd_sc_hd__xor2_1_94/A sky130_fd_sc_hd__nand2_1_334/Y sky130_fd_sc_hd__nand2_1_332/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_33 sky130_fd_sc_hd__nor2_1_172/A sky130_fd_sc_hd__a222oi_1_10/Y
+ sky130_fd_sc_hd__xor2_1_153/A sky130_fd_sc_hd__nand2_1_387/Y sky130_fd_sc_hd__a21oi_1_284/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_44 sky130_fd_sc_hd__nor2_1_222/A sky130_fd_sc_hd__a211oi_1_23/Y
+ sky130_fd_sc_hd__xor2_1_196/A sky130_fd_sc_hd__nand2_1_437/Y sky130_fd_sc_hd__nand2_1_438/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_55 sky130_fd_sc_hd__o21ai_1_419/A2 sky130_fd_sc_hd__nor2_1_265/A
+ sky130_fd_sc_hd__xor2_1_240/A sky130_fd_sc_hd__nand2_1_488/Y sky130_fd_sc_hd__nand2_1_490/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_66 sky130_fd_sc_hd__nor2_1_307/A sky130_fd_sc_hd__a21oi_1_470/Y
+ sky130_fd_sc_hd__xor2_1_283/A sky130_fd_sc_hd__nand2_1_539/Y sky130_fd_sc_hd__nand2_1_542/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__fa_2_1290 sky130_fd_sc_hd__fa_2_1291/CIN sky130_fd_sc_hd__mux2_2_227/A0
+ sky130_fd_sc_hd__fa_2_1290/A sky130_fd_sc_hd__fa_2_1290/B sky130_fd_sc_hd__fa_2_1290/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_1_202 sky130_fd_sc_hd__clkinv_2_21/A sky130_fd_sc_hd__a22o_1_31/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_202/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_213 sky130_fd_sc_hd__clkinv_2_27/A sky130_fd_sc_hd__a22oi_1_281/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_213/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_224 sky130_fd_sc_hd__clkinv_1_225/A sky130_fd_sc_hd__o21ai_2_0/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_224/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_235 sky130_fd_sc_hd__clkinv_1_236/A sky130_fd_sc_hd__buf_8_185/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_235/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_246 sky130_fd_sc_hd__buf_12_395/A sky130_fd_sc_hd__clkinv_1_246/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_246/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_257 sky130_fd_sc_hd__o21ai_1_8/A1 sky130_fd_sc_hd__o21ai_1_9/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_257/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_268 sky130_fd_sc_hd__maj3_1_2/B sky130_fd_sc_hd__ha_2_155/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_268/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_279 sky130_fd_sc_hd__fa_2_9/A sky130_fd_sc_hd__fa_2_2/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_279/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_9 sky130_fd_sc_hd__or4_1_1/B sky130_fd_sc_hd__a21oi_1_9/B1
+ sky130_fd_sc_hd__a21oi_1_9/Y sky130_fd_sc_hd__o21ai_1_13/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_110 sky130_fd_sc_hd__clkinv_1_565/Y sky130_fd_sc_hd__o21ai_1_132/Y
+ sky130_fd_sc_hd__a21oi_1_110/Y sky130_fd_sc_hd__a211o_1_8/A2 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_121 sky130_fd_sc_hd__clkinv_1_585/Y sky130_fd_sc_hd__o22ai_1_129/Y
+ sky130_fd_sc_hd__a21oi_1_121/Y sky130_fd_sc_hd__a211o_1_8/A2 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_132 sky130_fd_sc_hd__fa_2_1005/A sky130_fd_sc_hd__o21ai_1_155/Y
+ sky130_fd_sc_hd__a21oi_1_132/Y sky130_fd_sc_hd__nor2_4_10/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_143 sky130_fd_sc_hd__nor2_2_10/Y sky130_fd_sc_hd__o22ai_1_143/Y
+ sky130_fd_sc_hd__a21oi_1_143/Y sky130_fd_sc_hd__fa_2_1115/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_154 sky130_fd_sc_hd__nor2_2_11/Y sky130_fd_sc_hd__o22ai_1_153/Y
+ sky130_fd_sc_hd__a21oi_1_154/Y sky130_fd_sc_hd__fa_2_1111/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_165 sky130_fd_sc_hd__nor2_2_11/Y sky130_fd_sc_hd__o22ai_1_163/Y
+ sky130_fd_sc_hd__a21oi_1_165/Y sky130_fd_sc_hd__nor2_1_141/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_176 sky130_fd_sc_hd__nand2_1_304/Y sky130_fd_sc_hd__nor2_1_95/A
+ sky130_fd_sc_hd__xnor2_1_76/A sky130_fd_sc_hd__xnor2_1_74/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_187 sky130_fd_sc_hd__nor2_1_120/B sky130_fd_sc_hd__o21a_1_15/A1
+ sky130_fd_sc_hd__dfxtp_1_753/D sky130_fd_sc_hd__o21ai_1_206/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_198 sky130_fd_sc_hd__clkinv_1_700/Y sky130_fd_sc_hd__o22ai_1_171/Y
+ sky130_fd_sc_hd__a21oi_1_198/Y sky130_fd_sc_hd__nand2_1_333/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_106 sky130_fd_sc_hd__buf_8_106/A sky130_fd_sc_hd__buf_8_106/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_117 sky130_fd_sc_hd__buf_8_117/A sky130_fd_sc_hd__buf_8_117/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_128 sky130_fd_sc_hd__buf_8_128/A sky130_fd_sc_hd__buf_8_128/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_139 sky130_fd_sc_hd__buf_8_139/A sky130_fd_sc_hd__buf_4_86/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nand2_1_170 sky130_fd_sc_hd__fa_2_355/A sky130_fd_sc_hd__fa_2_422/B
+ sky130_fd_sc_hd__fa_2_425/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_181 sky130_fd_sc_hd__fa_2_532/A sky130_fd_sc_hd__fa_2_551/A
+ sky130_fd_sc_hd__fa_2_554/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_780 sky130_fd_sc_hd__o22ai_1_261/A2 sky130_fd_sc_hd__nor2_2_15/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_780/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_192 sky130_fd_sc_hd__fa_2_568/B sky130_fd_sc_hd__fa_2_698/A
+ sky130_fd_sc_hd__fa_2_700/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_791 sky130_fd_sc_hd__o32ai_1_1/A3 sky130_fd_sc_hd__fa_2_1141/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_791/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21o_2_18 sky130_fd_sc_hd__a21o_2_18/X sky130_fd_sc_hd__nor2_1_251/Y
+ sky130_fd_sc_hd__nor2_1_251/A sky130_fd_sc_hd__nor2_1_251/B VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__a21o_2_29 sky130_fd_sc_hd__a21o_2_29/X sky130_fd_sc_hd__nor2_1_298/Y
+ sky130_fd_sc_hd__fa_2_26/SUM sky130_fd_sc_hd__or3_1_5/X VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__xor2_1_12 sky130_fd_sc_hd__xor2_1_17/A sky130_fd_sc_hd__xor2_1_12/X
+ sky130_fd_sc_hd__xor2_1_12/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_23 sky130_fd_sc_hd__xor2_1_23/B sky130_fd_sc_hd__xor2_1_23/X
+ sky130_fd_sc_hd__xor2_1_23/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_34 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__xor2_1_34/X
+ sky130_fd_sc_hd__nor2_4_9/B VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_45 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_982/B
+ sky130_fd_sc_hd__xor2_1_45/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_56 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_971/B
+ sky130_fd_sc_hd__xor2_1_56/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_67 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__xor2_1_67/X
+ sky130_fd_sc_hd__xor2_1_67/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_78 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__fa_2_998/B
+ sky130_fd_sc_hd__xor2_1_78/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_89 sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__xor2_1_89/X
+ sky130_fd_sc_hd__xor2_1_89/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2b_1_6 sky130_fd_sc_hd__nand2b_1_6/Y sky130_fd_sc_hd__fa_2_949/A
+ sky130_fd_sc_hd__nor2b_1_87/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a21o_2_2 sky130_fd_sc_hd__a21o_2_2/X sky130_fd_sc_hd__a21o_2_2/B1
+ sky130_fd_sc_hd__xor2_1_28/X sky130_fd_sc_hd__a21o_2_2/A2 VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__dfxtp_1_905 VDD VSS sky130_fd_sc_hd__fa_2_940/B sky130_fd_sc_hd__clkinv_4_22/Y
+ sky130_fd_sc_hd__dfxtp_1_905/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_916 VDD VSS sky130_fd_sc_hd__fa_2_1145/A sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__mux2_2_107/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_927 VDD VSS sky130_fd_sc_hd__fa_2_1156/A sky130_fd_sc_hd__clkinv_8_46/Y
+ sky130_fd_sc_hd__mux2_2_80/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_938 VDD VSS sky130_fd_sc_hd__fa_2_1130/A sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__mux2_2_99/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_949 VDD VSS sky130_fd_sc_hd__fa_2_1158/B sky130_fd_sc_hd__clkinv_8_64/Y
+ sky130_fd_sc_hd__mux2_2_123/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a221oi_1_4 sky130_fd_sc_hd__a221oi_1_4/Y sky130_fd_sc_hd__xnor2_1_99/Y
+ sky130_fd_sc_hd__xor2_1_275/B sky130_fd_sc_hd__nand2_1_470/Y sky130_fd_sc_hd__o31ai_1_9/A3
+ sky130_fd_sc_hd__nor2_1_248/B VSS VDD VDD VSS sky130_fd_sc_hd__a221oi_1
Xsky130_fd_sc_hd__clkbuf_1_503 VSS VDD sky130_fd_sc_hd__buf_12_392/A sky130_fd_sc_hd__inv_2_121/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_514 VSS VDD sky130_fd_sc_hd__buf_4_110/A sky130_fd_sc_hd__buf_8_202/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_525 VSS VDD sky130_fd_sc_hd__clkbuf_1_525/X sky130_fd_sc_hd__clkbuf_1_525/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_536 VSS VDD sky130_fd_sc_hd__clkbuf_4_208/A sky130_fd_sc_hd__clkbuf_1_536/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_104 VSS VDD VSS VDD sky130_fd_sc_hd__fa_2_32/A sky130_fd_sc_hd__fa_2_238/CIN
+ sky130_fd_sc_hd__fa_2_230/A sky130_fd_sc_hd__ha_2_104/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_547 VSS VDD sky130_fd_sc_hd__fa_2_209/B sky130_fd_sc_hd__fa_2_67/B
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_115 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_115/A sky130_fd_sc_hd__fa_2_405/B
+ sky130_fd_sc_hd__fa_2_401/B sky130_fd_sc_hd__ha_2_115/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_558 VSS VDD sky130_fd_sc_hd__nand2_1_89/B sky130_fd_sc_hd__nand4_1_60/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_126 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_126/A sky130_fd_sc_hd__maj3_1_133/B
+ sky130_fd_sc_hd__maj3_1_134/A sky130_fd_sc_hd__ha_2_130/A sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_569 VSS VDD sky130_fd_sc_hd__and2_0_1/A sky130_fd_sc_hd__nor4_1_0/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_137 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_140/A sky130_fd_sc_hd__fa_2_719/B
+ sky130_fd_sc_hd__ha_2_137/SUM sky130_fd_sc_hd__ha_2_141/A sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_148 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_148/A sky130_fd_sc_hd__xor2_1_12/A
+ sky130_fd_sc_hd__ha_2_148/SUM sky130_fd_sc_hd__ha_2_148/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_159 VSS VDD VSS VDD sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__ha_2_158/B
+ sky130_fd_sc_hd__ha_2_159/SUM sky130_fd_sc_hd__ha_2_159/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__maj3_1_8 sky130_fd_sc_hd__maj3_1_9/X sky130_fd_sc_hd__maj3_1_8/X
+ sky130_fd_sc_hd__maj3_1_8/B sky130_fd_sc_hd__maj3_1_8/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__ha_2_50 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_50/A sky130_fd_sc_hd__xor2_1_5/A
+ sky130_fd_sc_hd__ha_2_50/SUM sky130_fd_sc_hd__ha_2_50/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_61 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_61/A sky130_fd_sc_hd__ha_2_60/B
+ sky130_fd_sc_hd__ha_2_61/SUM sky130_fd_sc_hd__ha_2_61/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_72 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_72/A sky130_fd_sc_hd__ha_2_71/B
+ sky130_fd_sc_hd__ha_2_72/SUM sky130_fd_sc_hd__ha_2_72/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_83 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_83/A sky130_fd_sc_hd__ha_2_82/B
+ sky130_fd_sc_hd__ha_2_83/SUM sky130_fd_sc_hd__ha_2_83/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_94 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_95/B sky130_fd_sc_hd__fa_2_91/CIN
+ sky130_fd_sc_hd__fa_2_83/A sky130_fd_sc_hd__ha_2_94/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_2 VSS VDD sky130_fd_sc_hd__buf_4_0/A sky130_fd_sc_hd__clkbuf_1_2/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__a221o_1_0 sky130_fd_sc_hd__a221o_1_0/X sky130_fd_sc_hd__a221o_1_0/B1
+ sky130_fd_sc_hd__nor2_1_40/B sky130_fd_sc_hd__a221o_1_0/B2 sky130_fd_sc_hd__nor2_1_40/A
+ VSS VDD sky130_fd_sc_hd__nor3_1_37/Y VDD VSS sky130_fd_sc_hd__a221o_1
Xsky130_fd_sc_hd__sdlclkp_4_90 sky130_fd_sc_hd__conb_1_28/LO sky130_fd_sc_hd__clkinv_8_47/A
+ sky130_fd_sc_hd__dfxtp_1_1322/CLK sky130_fd_sc_hd__or2_0_12/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__clkinv_1_2 sky130_fd_sc_hd__nor2_1_1/B sky130_fd_sc_hd__nand3_1_17/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_2/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_170 sky130_fd_sc_hd__nor2_1_170/B sky130_fd_sc_hd__nor2_1_170/Y
+ sky130_fd_sc_hd__nor2_1_170/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_181 sky130_fd_sc_hd__o21a_1_29/A1 sky130_fd_sc_hd__nor2_1_181/Y
+ sky130_fd_sc_hd__nor2_1_181/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_192 sky130_fd_sc_hd__nor2_1_192/B sky130_fd_sc_hd__o21a_1_36/A1
+ sky130_fd_sc_hd__o21a_1_37/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_90 sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__a22oi_2_12/A1
+ sky130_fd_sc_hd__buf_2_80/X sky130_fd_sc_hd__a22oi_1_90/A2 sky130_fd_sc_hd__a22oi_1_90/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__and2_0_17 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_17/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__and2_0_17/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_28 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_28/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_36/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_308 sky130_fd_sc_hd__o32ai_1_5/A3 sky130_fd_sc_hd__nor2_1_188/B
+ sky130_fd_sc_hd__o22ai_1_308/Y sky130_fd_sc_hd__o22ai_1_308/A1 sky130_fd_sc_hd__o21a_1_42/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__and2_0_39 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_60/A sky130_fd_sc_hd__nor2_4_1/Y
+ sky130_fd_sc_hd__ha_2_54/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_319 sky130_fd_sc_hd__nor2_1_199/B sky130_fd_sc_hd__nor2_1_224/A
+ sky130_fd_sc_hd__o22ai_1_319/Y sky130_fd_sc_hd__o22ai_1_319/A1 sky130_fd_sc_hd__a222oi_1_23/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_2_9 sky130_fd_sc_hd__nor2_2_9/B sky130_fd_sc_hd__or2_0_6/B
+ sky130_fd_sc_hd__nor2_2_9/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__a22oi_1_280 sky130_fd_sc_hd__clkbuf_1_376/X sky130_fd_sc_hd__nor2_2_5/Y
+ sky130_fd_sc_hd__buf_2_212/X sky130_fd_sc_hd__clkbuf_1_468/X sky130_fd_sc_hd__nand4_1_69/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_291 sky130_fd_sc_hd__nor2_2_4/Y sky130_fd_sc_hd__clkbuf_1_377/X
+ sky130_fd_sc_hd__a22oi_1_291/B2 sky130_fd_sc_hd__clkbuf_4_184/X sky130_fd_sc_hd__nand4_1_72/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_4_120 VDD VSS sky130_fd_sc_hd__buf_4_120/X sky130_fd_sc_hd__buf_4_120/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_8_16 sky130_fd_sc_hd__inv_2_28/Y sky130_fd_sc_hd__buf_8_16/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_27 sky130_fd_sc_hd__inv_2_23/Y sky130_fd_sc_hd__buf_8_27/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_38 sky130_fd_sc_hd__inv_2_6/A sky130_fd_sc_hd__buf_8_38/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_49 sky130_fd_sc_hd__buf_8_49/A sky130_fd_sc_hd__buf_8_49/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__o21ai_1_502 VSS VDD sky130_fd_sc_hd__nand2_1_563/A sky130_fd_sc_hd__o21ai_1_507/A1
+ sky130_fd_sc_hd__nand2_1_563/Y sky130_fd_sc_hd__and2_0_355/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1108 VDD VSS sky130_fd_sc_hd__nor2_4_16/B sky130_fd_sc_hd__clkinv_4_23/Y
+ sky130_fd_sc_hd__nor2b_1_114/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1119 VDD VSS sky130_fd_sc_hd__mux2_2_144/A0 sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__o22ai_1_274/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_702 VDD VSS sky130_fd_sc_hd__mux2_2_31/A0 sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__o21ai_1_42/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_713 VDD VSS sky130_fd_sc_hd__mux2_2_7/A1 sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__o21ai_1_53/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_724 VDD VSS sky130_fd_sc_hd__mux2_2_24/A1 sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__o21ai_1_61/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_735 VDD VSS sky130_fd_sc_hd__mux2_2_1/A1 sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__o21ai_1_72/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_746 VDD VSS sky130_fd_sc_hd__and2_0_182/A sky130_fd_sc_hd__dfxtp_1_747/CLK
+ sky130_fd_sc_hd__fa_2_1101/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_757 VDD VSS sky130_fd_sc_hd__fa_2_677/A sky130_fd_sc_hd__dfxtp_1_764/CLK
+ sky130_fd_sc_hd__dfxtp_1_757/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_768 VDD VSS sky130_fd_sc_hd__fa_2_699/A sky130_fd_sc_hd__dfxtp_1_768/CLK
+ sky130_fd_sc_hd__xnor2_1_90/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_779 VDD VSS sky130_fd_sc_hd__fa_2_1078/A sky130_fd_sc_hd__clkinv_8_55/Y
+ sky130_fd_sc_hd__mux2_2_67/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_300 VSS VDD sky130_fd_sc_hd__nand4_1_45/D sky130_fd_sc_hd__a22oi_1_199/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_311 VSS VDD sky130_fd_sc_hd__nand4_1_34/D sky130_fd_sc_hd__a22oi_1_155/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_322 VSS VDD sky130_fd_sc_hd__clkbuf_1_322/X sky130_fd_sc_hd__nand3_1_32/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_333 VSS VDD sky130_fd_sc_hd__buf_12_286/A sky130_fd_sc_hd__buf_4_69/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_344 VSS VDD sky130_fd_sc_hd__buf_12_276/A sky130_fd_sc_hd__and2_4_0/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_355 VSS VDD sky130_fd_sc_hd__buf_8_167/A sky130_fd_sc_hd__clkinv_4_15/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_366 VSS VDD sky130_fd_sc_hd__clkbuf_1_366/X sky130_fd_sc_hd__a22o_2_3/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_377 VSS VDD sky130_fd_sc_hd__clkbuf_1_377/X sky130_fd_sc_hd__nor3_1_24/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_388 VSS VDD sky130_fd_sc_hd__a22oi_2_24/B2 sky130_fd_sc_hd__clkbuf_1_388/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_607 sky130_fd_sc_hd__maj3_1_121/B sky130_fd_sc_hd__maj3_1_122/A
+ sky130_fd_sc_hd__fa_2_607/A sky130_fd_sc_hd__fa_2_607/B sky130_fd_sc_hd__fa_2_608/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_399 VSS VDD sky130_fd_sc_hd__clkbuf_1_399/X sky130_fd_sc_hd__clkbuf_1_399/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_618 sky130_fd_sc_hd__maj3_1_118/B sky130_fd_sc_hd__maj3_1_119/A
+ sky130_fd_sc_hd__fa_2_618/A sky130_fd_sc_hd__fa_2_618/B sky130_fd_sc_hd__fa_2_619/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_629 sky130_fd_sc_hd__fa_2_630/A sky130_fd_sc_hd__fa_2_626/A
+ sky130_fd_sc_hd__fa_2_695/A sky130_fd_sc_hd__fa_2_689/B sky130_fd_sc_hd__fa_2_683/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_70 VDD VSS sky130_fd_sc_hd__ha_2_104/B sky130_fd_sc_hd__dfxtp_1_73/CLK
+ sky130_fd_sc_hd__buf_2_290/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_81 VDD VSS sky130_fd_sc_hd__dfxtp_1_81/Q sky130_fd_sc_hd__dfxtp_1_8/CLK
+ sky130_fd_sc_hd__nand3_1_17/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_92 VDD VSS sky130_fd_sc_hd__a22o_1_8/B2 sky130_fd_sc_hd__dfxtp_1_93/CLK
+ sky130_fd_sc_hd__dfxtp_1_92/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_320 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_320/X sky130_fd_sc_hd__mux2_2_99/S
+ sky130_fd_sc_hd__and2_0_320/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_160 sky130_fd_sc_hd__clkbuf_4_160/X sky130_fd_sc_hd__buf_2_138/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_331 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_331/X sky130_fd_sc_hd__inv_2_139/Y
+ sky130_fd_sc_hd__and2_0_331/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_171 sky130_fd_sc_hd__clkbuf_4_171/X sky130_fd_sc_hd__clkbuf_4_171/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_342 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_342/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_342/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_182 sky130_fd_sc_hd__clkbuf_4_182/X sky130_fd_sc_hd__clkbuf_4_182/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_353 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_353/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_353/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_193 sky130_fd_sc_hd__nand4_1_79/D sky130_fd_sc_hd__a22oi_1_317/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__conb_1_6 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__conb_1_6/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__or2_0_0 sky130_fd_sc_hd__or2_0_0/A sky130_fd_sc_hd__or2_0_0/X sky130_fd_sc_hd__or2_0_0/B
+ VSS VDD VSS VDD sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__inv_2_120 sky130_fd_sc_hd__inv_2_120/A sky130_fd_sc_hd__inv_2_120/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_131 sky130_fd_sc_hd__inv_2_131/A sky130_fd_sc_hd__inv_2_132/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__o22ai_1_105 sky130_fd_sc_hd__o22ai_1_130/B1 sky130_fd_sc_hd__nor2_1_65/B
+ sky130_fd_sc_hd__nor2_1_80/A sky130_fd_sc_hd__o22ai_1_116/A1 sky130_fd_sc_hd__o22ai_1_132/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_116 sky130_fd_sc_hd__o21a_1_8/A2 sky130_fd_sc_hd__nor2_1_65/B
+ sky130_fd_sc_hd__nor2_1_84/B sky130_fd_sc_hd__o22ai_1_116/A1 sky130_fd_sc_hd__o21ai_1_92/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_127 sky130_fd_sc_hd__nor2_1_76/A sky130_fd_sc_hd__nor2_2_9/B
+ sky130_fd_sc_hd__o22ai_1_127/Y sky130_fd_sc_hd__a21oi_1_127/Y sky130_fd_sc_hd__a211oi_1_5/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_138 sky130_fd_sc_hd__nand2_1_284/Y sky130_fd_sc_hd__nand2_2_5/Y
+ sky130_fd_sc_hd__o22ai_1_138/Y sky130_fd_sc_hd__xnor2_1_68/Y sky130_fd_sc_hd__o22ai_1_152/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_149 sky130_fd_sc_hd__nand2_1_338/A sky130_fd_sc_hd__nand2_1_284/Y
+ sky130_fd_sc_hd__o22ai_1_149/Y sky130_fd_sc_hd__xnor2_1_62/Y sky130_fd_sc_hd__o22ai_1_149/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_2_16 sky130_fd_sc_hd__nor2_2_16/B sky130_fd_sc_hd__nor2_2_16/Y
+ sky130_fd_sc_hd__nor2_4_16/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__nand4_1_19 sky130_fd_sc_hd__nand4_1_19/C sky130_fd_sc_hd__nand4_1_19/B
+ sky130_fd_sc_hd__nand4_1_19/Y sky130_fd_sc_hd__nand4_1_19/D sky130_fd_sc_hd__buf_2_109/X
+ VDD VSS VDD VSS sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__o211ai_1_6 sky130_fd_sc_hd__o211ai_1_6/A1 sky130_fd_sc_hd__o21a_1_8/A2
+ sky130_fd_sc_hd__o211ai_1_6/Y sky130_fd_sc_hd__o211ai_1_6/C1 sky130_fd_sc_hd__o211ai_1_6/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__a31oi_1_3 VSS VDD sky130_fd_sc_hd__a31oi_1_3/Y sky130_fd_sc_hd__a31oi_1_3/B1
+ sky130_fd_sc_hd__a31oi_1_3/A2 sky130_fd_sc_hd__a31oi_1_3/A1 sky130_fd_sc_hd__a31oi_1_3/A3
+ VDD VSS sky130_fd_sc_hd__a31oi_1
Xsky130_fd_sc_hd__o21ai_1_310 VSS VDD sky130_fd_sc_hd__a222oi_1_10/Y sky130_fd_sc_hd__nor2_1_182/A
+ sky130_fd_sc_hd__nand2_1_382/Y sky130_fd_sc_hd__xor2_1_145/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_321 VSS VDD sky130_fd_sc_hd__a222oi_1_11/Y sky130_fd_sc_hd__nor2_1_182/A
+ sky130_fd_sc_hd__a22oi_1_377/Y sky130_fd_sc_hd__o21ai_1_321/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_332 VSS VDD sky130_fd_sc_hd__nand2_1_420/B sky130_fd_sc_hd__nor2_1_209/Y
+ sky130_fd_sc_hd__nor2_1_208/B sky130_fd_sc_hd__o21ai_1_332/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_343 VSS VDD sky130_fd_sc_hd__a222oi_1_16/Y sky130_fd_sc_hd__nor2_1_224/A
+ sky130_fd_sc_hd__nand2_1_425/Y sky130_fd_sc_hd__xor2_1_211/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_354 VSS VDD sky130_fd_sc_hd__o22ai_1_322/A2 sky130_fd_sc_hd__nor2_1_218/A
+ sky130_fd_sc_hd__a22oi_1_382/Y sky130_fd_sc_hd__o21ai_1_354/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a211oi_1_15 sky130_fd_sc_hd__nor2b_1_105/Y sky130_fd_sc_hd__nor2_1_179/Y
+ sky130_fd_sc_hd__o21ai_1_325/Y sky130_fd_sc_hd__a211oi_1_15/Y sky130_fd_sc_hd__o21ai_1_326/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_365 VSS VDD sky130_fd_sc_hd__o21ai_1_365/A2 sky130_fd_sc_hd__nor2_1_224/A
+ sky130_fd_sc_hd__nand2_1_434/Y sky130_fd_sc_hd__xor2_1_191/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a211oi_1_26 sky130_fd_sc_hd__nor2b_1_119/Y sky130_fd_sc_hd__o21ai_1_411/Y
+ sky130_fd_sc_hd__nor2_1_259/Y sky130_fd_sc_hd__a211oi_1_26/Y sky130_fd_sc_hd__o21ai_1_413/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_376 VSS VDD sky130_fd_sc_hd__o22ai_1_318/A2 sky130_fd_sc_hd__nor2_1_223/A
+ sky130_fd_sc_hd__a21oi_1_352/Y sky130_fd_sc_hd__o21ai_1_376/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a211oi_1_37 sky130_fd_sc_hd__nor3_1_41/A sky130_fd_sc_hd__nor2_1_308/Y
+ sky130_fd_sc_hd__o22ai_1_430/Y sky130_fd_sc_hd__a211oi_1_37/Y sky130_fd_sc_hd__fa_2_1307/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_387 VSS VDD sky130_fd_sc_hd__nand2_1_473/B sky130_fd_sc_hd__nor2_1_253/Y
+ sky130_fd_sc_hd__nor2_1_252/B sky130_fd_sc_hd__o21ai_1_387/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_398 VSS VDD sky130_fd_sc_hd__nor2_1_257/B sky130_fd_sc_hd__nor2_1_267/A
+ sky130_fd_sc_hd__nand2_1_477/Y sky130_fd_sc_hd__xor2_1_257/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__mux2_2_12 VSS VDD sky130_fd_sc_hd__mux2_2_12/A1 sky130_fd_sc_hd__mux2_2_12/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_12/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_23 VSS VDD sky130_fd_sc_hd__mux2_2_23/A1 sky130_fd_sc_hd__mux2_2_23/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_23/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_34 VSS VDD sky130_fd_sc_hd__mux2_2_34/A1 sky130_fd_sc_hd__mux2_2_34/A0
+ sky130_fd_sc_hd__mux2_2_37/S sky130_fd_sc_hd__mux2_2_34/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_45 VSS VDD sky130_fd_sc_hd__mux2_2_45/A1 sky130_fd_sc_hd__mux2_2_45/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_45/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_56 VSS VDD sky130_fd_sc_hd__mux2_2_56/A1 sky130_fd_sc_hd__mux2_2_56/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_56/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_67 VSS VDD sky130_fd_sc_hd__mux2_2_67/A1 sky130_fd_sc_hd__mux2_2_67/A0
+ sky130_fd_sc_hd__mux2_2_75/S sky130_fd_sc_hd__mux2_2_67/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_78 VSS VDD sky130_fd_sc_hd__mux2_2_78/A1 sky130_fd_sc_hd__mux2_2_78/A0
+ sky130_fd_sc_hd__nor2_4_15/A sky130_fd_sc_hd__mux2_2_78/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_89 VSS VDD sky130_fd_sc_hd__mux2_2_89/A1 sky130_fd_sc_hd__mux2_2_89/A0
+ sky130_fd_sc_hd__mux2_2_99/S sky130_fd_sc_hd__mux2_2_89/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1108 sky130_fd_sc_hd__fa_2_1109/CIN sky130_fd_sc_hd__fa_2_1108/SUM
+ sky130_fd_sc_hd__fa_2_1108/A sky130_fd_sc_hd__fa_2_1108/B sky130_fd_sc_hd__fa_2_1108/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1119 sky130_fd_sc_hd__fa_2_1120/CIN sky130_fd_sc_hd__fa_2_1119/SUM
+ sky130_fd_sc_hd__fa_2_1119/A sky130_fd_sc_hd__nor2_1_99/A sky130_fd_sc_hd__fa_2_1119/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_510 VDD VSS sky130_fd_sc_hd__nor4_1_11/D sky130_fd_sc_hd__edfxtp_1_0/CLK
+ sky130_fd_sc_hd__a22o_1_61/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_170 sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__fa_2_1152/B
+ sky130_fd_sc_hd__xor2_1_170/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_521 VDD VSS sky130_fd_sc_hd__xor2_1_30/A sky130_fd_sc_hd__dfxtp_1_526/CLK
+ sky130_fd_sc_hd__and2_0_255/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_181 sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__fa_2_1141/B
+ sky130_fd_sc_hd__xor2_1_181/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_192 sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__fa_2_1187/B
+ sky130_fd_sc_hd__xor2_1_192/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_532 VDD VSS sky130_fd_sc_hd__fa_2_959/A sky130_fd_sc_hd__dfxtp_1_533/CLK
+ sky130_fd_sc_hd__and2_0_258/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_543 VDD VSS sky130_fd_sc_hd__fa_2_948/A sky130_fd_sc_hd__dfxtp_1_544/CLK
+ sky130_fd_sc_hd__a22o_1_42/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_554 VDD VSS sky130_fd_sc_hd__dfxtp_1_554/Q sky130_fd_sc_hd__dfxtp_1_576/CLK
+ sky130_fd_sc_hd__dfxtp_1_554/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_565 VDD VSS sky130_fd_sc_hd__and2_0_235/A sky130_fd_sc_hd__dfxtp_1_577/CLK
+ sky130_fd_sc_hd__a22o_1_34/B1 VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_576 VDD VSS sky130_fd_sc_hd__dfxtp_1_576/Q sky130_fd_sc_hd__dfxtp_1_576/CLK
+ sky130_fd_sc_hd__nor2_1_27/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_587 VDD VSS sky130_fd_sc_hd__nor4_1_8/B sky130_fd_sc_hd__dfxtp_1_594/CLK
+ sky130_fd_sc_hd__and2_0_243/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_598 VDD VSS sky130_fd_sc_hd__and2_0_208/A sky130_fd_sc_hd__dfxtp_1_601/CLK
+ sky130_fd_sc_hd__fa_2_1018/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_130 VSS VDD sky130_fd_sc_hd__ha_2_10/A sky130_fd_sc_hd__dfxtp_1_130/Q
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_141 VSS VDD sky130_fd_sc_hd__clkbuf_1_141/X sky130_fd_sc_hd__clkbuf_1_141/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_152 VSS VDD sky130_fd_sc_hd__a22oi_1_92/B2 sky130_fd_sc_hd__clkbuf_1_152/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_163 VSS VDD sky130_fd_sc_hd__clkbuf_1_163/X sky130_fd_sc_hd__clkbuf_1_163/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_174 VSS VDD sky130_fd_sc_hd__clkbuf_1_174/X sky130_fd_sc_hd__nand3_2_2/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_185 VSS VDD sky130_fd_sc_hd__nand4_1_20/B sky130_fd_sc_hd__clkbuf_1_244/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_196 VSS VDD sky130_fd_sc_hd__buf_4_40/A sky130_fd_sc_hd__clkbuf_1_196/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_404 sky130_fd_sc_hd__fa_2_403/A sky130_fd_sc_hd__fa_2_397/B
+ sky130_fd_sc_hd__fa_2_404/A sky130_fd_sc_hd__fa_2_404/B sky130_fd_sc_hd__fa_2_416/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_415 sky130_fd_sc_hd__fa_2_418/B sky130_fd_sc_hd__fa_2_415/SUM
+ sky130_fd_sc_hd__fa_2_415/A sky130_fd_sc_hd__fa_2_415/B sky130_fd_sc_hd__fa_2_415/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_426 sky130_fd_sc_hd__fa_2_433/CIN sky130_fd_sc_hd__fa_2_426/SUM
+ sky130_fd_sc_hd__fa_2_426/A sky130_fd_sc_hd__fa_2_426/B sky130_fd_sc_hd__fa_2_426/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_437 sky130_fd_sc_hd__fa_2_426/A sky130_fd_sc_hd__fa_2_435/B
+ sky130_fd_sc_hd__fa_2_566/B sky130_fd_sc_hd__fa_2_437/B sky130_fd_sc_hd__fa_2_440/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_448 sky130_fd_sc_hd__fa_2_445/CIN sky130_fd_sc_hd__fa_2_448/SUM
+ sky130_fd_sc_hd__fa_2_448/A sky130_fd_sc_hd__fa_2_448/B sky130_fd_sc_hd__fa_2_448/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_459 sky130_fd_sc_hd__fa_2_452/A sky130_fd_sc_hd__fa_2_456/B
+ sky130_fd_sc_hd__fa_2_459/A sky130_fd_sc_hd__fa_2_459/B sky130_fd_sc_hd__fa_2_459/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nand3_1_30 sky130_fd_sc_hd__buf_2_120/A sky130_fd_sc_hd__nand3_2_2/A
+ sky130_fd_sc_hd__nand3_1_30/C sky130_fd_sc_hd__nand3_2_2/C VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_41 sky130_fd_sc_hd__inv_4_1/A sky130_fd_sc_hd__nor3_1_26/A
+ sky130_fd_sc_hd__nor3_1_26/C sky130_fd_sc_hd__nor3_1_27/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_52 sky130_fd_sc_hd__nand3_1_52/Y sky130_fd_sc_hd__nand3_1_52/A
+ sky130_fd_sc_hd__nand3_1_52/C sky130_fd_sc_hd__nand3_1_52/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__dfxtp_1_1450 VDD VSS sky130_fd_sc_hd__dfxtp_1_1450/Q sky130_fd_sc_hd__sdlclkp_1_6/GCLK
+ sky130_fd_sc_hd__and2_0_347/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1461 VDD VSS sky130_fd_sc_hd__buf_2_275/A sky130_fd_sc_hd__dfxtp_1_1461/CLK
+ sky130_fd_sc_hd__and2_0_345/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_150 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_150/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_925/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_161 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_161/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__fa_2_860/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_172 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_172/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_172/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_80 sky130_fd_sc_hd__clkinv_1_81/A sky130_fd_sc_hd__buf_2_44/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_80/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_183 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_183/X sky130_fd_sc_hd__and2_0_235/B
+ sky130_fd_sc_hd__and2_0_183/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_91 sky130_fd_sc_hd__clkinv_1_92/A sky130_fd_sc_hd__nand3_1_26/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_91/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_194 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_194/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_901/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_409 sky130_fd_sc_hd__bufbuf_8_5/X sky130_fd_sc_hd__buf_12_409/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__fa_2_960 sky130_fd_sc_hd__fa_2_959/CIN sky130_fd_sc_hd__fa_2_960/SUM
+ sky130_fd_sc_hd__fa_2_960/A sky130_fd_sc_hd__fa_2_960/B sky130_fd_sc_hd__fa_2_960/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_971 sky130_fd_sc_hd__fa_2_972/CIN sky130_fd_sc_hd__fa_2_971/SUM
+ sky130_fd_sc_hd__fa_2_971/A sky130_fd_sc_hd__fa_2_971/B sky130_fd_sc_hd__fa_2_971/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_982 sky130_fd_sc_hd__fa_2_983/CIN sky130_fd_sc_hd__mux2_2_23/A0
+ sky130_fd_sc_hd__fa_2_982/A sky130_fd_sc_hd__fa_2_982/B sky130_fd_sc_hd__fa_2_982/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_993 sky130_fd_sc_hd__fa_2_994/CIN sky130_fd_sc_hd__fa_2_993/SUM
+ sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__fa_2_993/B sky130_fd_sc_hd__xor2_1_83/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_1_0 sky130_fd_sc_hd__conb_1_8/LO sky130_fd_sc_hd__clkinv_4_1/Y
+ sky130_fd_sc_hd__dfxtp_1_126/CLK sky130_fd_sc_hd__clkbuf_1_1/X VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_1
Xsky130_fd_sc_hd__clkinv_1_609 sky130_fd_sc_hd__ha_2_184/A sky130_fd_sc_hd__ha_2_185/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_609/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__mux2_2_260 VSS VDD sky130_fd_sc_hd__mux2_2_260/A1 sky130_fd_sc_hd__mux2_2_260/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_260/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__o21ai_1_140 VSS VDD sky130_fd_sc_hd__a21oi_1_129/Y sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__a21oi_1_116/Y sky130_fd_sc_hd__xor2_1_48/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_151 VSS VDD sky130_fd_sc_hd__o22ai_1_132/B2 sky130_fd_sc_hd__o21ai_1_92/A1
+ sky130_fd_sc_hd__a22oi_1_341/Y sky130_fd_sc_hd__o21ai_1_151/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_162 VSS VDD sky130_fd_sc_hd__o21ai_1_171/A2 sky130_fd_sc_hd__xnor2_1_71/Y
+ sky130_fd_sc_hd__a21oi_1_139/Y sky130_fd_sc_hd__o21ai_1_162/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_173 VSS VDD sky130_fd_sc_hd__nand2_2_5/Y sky130_fd_sc_hd__o21ai_1_190/A2
+ sky130_fd_sc_hd__nand2_1_285/Y sky130_fd_sc_hd__o21ai_1_173/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_184 VSS VDD sky130_fd_sc_hd__nand2_2_5/Y sky130_fd_sc_hd__xnor2_1_81/Y
+ sky130_fd_sc_hd__a21oi_1_159/Y sky130_fd_sc_hd__o21ai_1_184/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_195 VSS VDD sky130_fd_sc_hd__xnor2_1_77/A sky130_fd_sc_hd__o21ai_1_195/A1
+ sky130_fd_sc_hd__nand2_1_290/B sky130_fd_sc_hd__xnor2_1_79/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_18 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1176/A sky130_fd_sc_hd__nor2_2_16/Y
+ sky130_fd_sc_hd__nor3_1_39/A sky130_fd_sc_hd__fa_2_1178/A sky130_fd_sc_hd__nor3_1_39/B
+ sky130_fd_sc_hd__a222oi_1_18/Y sky130_fd_sc_hd__fa_2_1175/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__a222oi_1_29 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1226/A sky130_fd_sc_hd__nor2_2_17/Y
+ sky130_fd_sc_hd__nor3_1_40/A sky130_fd_sc_hd__fa_2_1228/A sky130_fd_sc_hd__nor3_1_40/B
+ sky130_fd_sc_hd__a222oi_1_29/Y sky130_fd_sc_hd__fa_2_1225/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2_1_500 sky130_fd_sc_hd__o21a_1_58/B1 sky130_fd_sc_hd__fa_2_1287/A
+ sky130_fd_sc_hd__o21a_1_58/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_511 sky130_fd_sc_hd__nor2_1_284/A sky130_fd_sc_hd__fa_2_1295/A
+ sky130_fd_sc_hd__fa_2_1294/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_522 sky130_fd_sc_hd__nand2_1_522/Y sky130_fd_sc_hd__o31ai_1_12/A3
+ sky130_fd_sc_hd__o31ai_1_12/A2 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_90 sky130_fd_sc_hd__maj3_1_91/X sky130_fd_sc_hd__maj3_1_90/X
+ sky130_fd_sc_hd__maj3_1_90/B sky130_fd_sc_hd__maj3_1_90/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_533 sky130_fd_sc_hd__nand2_1_533/Y sky130_fd_sc_hd__nand2_1_543/B
+ sky130_fd_sc_hd__o21ai_1_470/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_544 sky130_fd_sc_hd__nand2_1_544/Y sky130_fd_sc_hd__nor2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_485/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_555 sky130_fd_sc_hd__nand2_1_555/Y sky130_fd_sc_hd__buf_2_274/X
+ sky130_fd_sc_hd__nand2_1_555/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_566 sky130_fd_sc_hd__nand2_1_566/Y sky130_fd_sc_hd__nand2_1_566/B
+ sky130_fd_sc_hd__nand2_1_566/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_2 sky130_fd_sc_hd__xor2_1_2/X sky130_fd_sc_hd__nor2b_1_2/Y
+ sky130_fd_sc_hd__or2_0_1/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1102 sky130_fd_sc_hd__o21ai_1_490/A1 sky130_fd_sc_hd__fa_2_1307/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1102/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1113 sky130_fd_sc_hd__nor2_1_314/B sky130_fd_sc_hd__nor2_1_315/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1113/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1124 sky130_fd_sc_hd__clkinv_2_42/A sky130_fd_sc_hd__buf_2_285/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1124/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_340 VDD VSS sky130_fd_sc_hd__a22o_1_21/B2 sky130_fd_sc_hd__dfxtp_1_354/CLK
+ sky130_fd_sc_hd__ha_2_157/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_351 VDD VSS sky130_fd_sc_hd__ha_2_152/A sky130_fd_sc_hd__dfxtp_1_361/CLK
+ sky130_fd_sc_hd__o2bb2ai_1_7/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_362 VDD VSS sky130_fd_sc_hd__ha_2_201/A sky130_fd_sc_hd__dfxtp_1_380/CLK
+ sky130_fd_sc_hd__and2_0_178/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_373 VDD VSS sky130_fd_sc_hd__fa_2_1117/A sky130_fd_sc_hd__clkinv_4_32/Y
+ sky130_fd_sc_hd__and2_0_124/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_384 VDD VSS sky130_fd_sc_hd__fa_2_1112/B sky130_fd_sc_hd__clkinv_4_32/Y
+ sky130_fd_sc_hd__and2_0_145/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_4 sky130_fd_sc_hd__nand3_1_4/C sky130_fd_sc_hd__nand2_1_4/B
+ sky130_fd_sc_hd__nand2_1_9/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_395 VDD VSS sky130_fd_sc_hd__fa_2_1031/A sky130_fd_sc_hd__dfxtp_1_411/CLK
+ sky130_fd_sc_hd__and2_0_232/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_201 sky130_fd_sc_hd__maj3_1_43/B sky130_fd_sc_hd__maj3_1_44/A
+ sky130_fd_sc_hd__fa_2_201/A sky130_fd_sc_hd__fa_2_201/B sky130_fd_sc_hd__fa_2_202/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_212 sky130_fd_sc_hd__fa_2_215/B sky130_fd_sc_hd__fa_2_212/SUM
+ sky130_fd_sc_hd__fa_2_212/A sky130_fd_sc_hd__fa_2_212/B sky130_fd_sc_hd__fa_2_212/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_223 sky130_fd_sc_hd__fa_2_225/CIN sky130_fd_sc_hd__fa_2_216/B
+ sky130_fd_sc_hd__fa_2_242/A sky130_fd_sc_hd__fa_2_274/A sky130_fd_sc_hd__fa_2_266/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_234 sky130_fd_sc_hd__fa_2_235/A sky130_fd_sc_hd__fa_2_227/A
+ sky130_fd_sc_hd__ha_2_91/B sky130_fd_sc_hd__fa_2_277/B sky130_fd_sc_hd__fa_2_144/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_245 sky130_fd_sc_hd__maj3_1_34/B sky130_fd_sc_hd__maj3_1_35/A
+ sky130_fd_sc_hd__fa_2_245/A sky130_fd_sc_hd__fa_2_245/B sky130_fd_sc_hd__fa_2_246/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_256 sky130_fd_sc_hd__fa_2_259/B sky130_fd_sc_hd__fa_2_256/SUM
+ sky130_fd_sc_hd__fa_2_256/A sky130_fd_sc_hd__fa_2_256/B sky130_fd_sc_hd__o22ai_1_17/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_267 sky130_fd_sc_hd__fa_2_170/A sky130_fd_sc_hd__maj3_1_30/A
+ sky130_fd_sc_hd__fa_2_267/A sky130_fd_sc_hd__fa_2_267/B sky130_fd_sc_hd__fa_2_269/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_278 sky130_fd_sc_hd__fa_2_164/A sky130_fd_sc_hd__fa_2_168/B
+ sky130_fd_sc_hd__fa_2_278/A sky130_fd_sc_hd__fa_2_278/B sky130_fd_sc_hd__fa_2_283/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_289 sky130_fd_sc_hd__fa_2_287/B sky130_fd_sc_hd__fa_2_288/B
+ sky130_fd_sc_hd__ha_2_108/B sky130_fd_sc_hd__fa_2_404/A sky130_fd_sc_hd__fa_2_286/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_5 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_5/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_0/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__diode_2_106 sky130_fd_sc_hd__inv_2_135/Y VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_117 sky130_fd_sc_hd__buf_2_225/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_128 sky130_fd_sc_hd__buf_2_250/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__fa_2_70 sky130_fd_sc_hd__fa_2_73/B sky130_fd_sc_hd__fa_2_70/SUM
+ sky130_fd_sc_hd__fa_2_70/A sky130_fd_sc_hd__fa_2_70/B sky130_fd_sc_hd__fa_2_70/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__diode_2_139 sky130_fd_sc_hd__clkbuf_1_526/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__fa_2_81 sky130_fd_sc_hd__fa_2_83/CIN sky130_fd_sc_hd__fa_2_74/B
+ sky130_fd_sc_hd__fa_2_87/A sky130_fd_sc_hd__fa_2_81/B sky130_fd_sc_hd__fa_2_91/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_92 sky130_fd_sc_hd__fa_2_93/A sky130_fd_sc_hd__fa_2_85/A sky130_fd_sc_hd__ha_2_91/B
+ sky130_fd_sc_hd__fa_2_92/B sky130_fd_sc_hd__fa_2_2/B VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_240 VDD VSS sky130_fd_sc_hd__buf_2_240/X sky130_fd_sc_hd__buf_6_60/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_251 VDD VSS sky130_fd_sc_hd__buf_2_251/X sky130_fd_sc_hd__buf_2_251/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_262 VDD VSS sky130_fd_sc_hd__buf_2_262/X sky130_fd_sc_hd__buf_2_262/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_273 VDD VSS sky130_fd_sc_hd__buf_6_49/A sky130_fd_sc_hd__buf_4_56/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_284 VDD VSS sky130_fd_sc_hd__nand3_2_2/A sky130_fd_sc_hd__buf_2_284/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1280 VDD VSS sky130_fd_sc_hd__mux2_2_199/A0 sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__dfxtp_1_436/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1291 VDD VSS sky130_fd_sc_hd__mux2_2_191/A0 sky130_fd_sc_hd__clkinv_8_75/Y
+ sky130_fd_sc_hd__o22ai_1_344/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a21oi_1_20 sky130_fd_sc_hd__nand4_1_84/B sky130_fd_sc_hd__o2111ai_1_1/Y
+ sky130_fd_sc_hd__a21oi_1_20/Y sky130_fd_sc_hd__a211o_1_1/X VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_31 sky130_fd_sc_hd__nor2_1_41/Y sky130_fd_sc_hd__o22ai_1_64/Y
+ sky130_fd_sc_hd__a21oi_1_31/Y sky130_fd_sc_hd__fa_2_1034/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_42 sky130_fd_sc_hd__a21oi_1_42/A1 sky130_fd_sc_hd__a22o_1_67/X
+ sky130_fd_sc_hd__a21oi_1_42/Y sky130_fd_sc_hd__o21ai_1_81/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_206 sky130_fd_sc_hd__buf_4_48/X sky130_fd_sc_hd__buf_12_224/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_53 sky130_fd_sc_hd__nor2_2_6/Y sky130_fd_sc_hd__o22ai_1_85/Y
+ sky130_fd_sc_hd__a21oi_1_53/Y sky130_fd_sc_hd__fa_2_1041/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_217 sky130_fd_sc_hd__buf_6_24/X sky130_fd_sc_hd__buf_12_217/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_64 sky130_fd_sc_hd__a21oi_1_64/A1 sky130_fd_sc_hd__nor2_1_43/B
+ sky130_fd_sc_hd__xnor2_1_40/A sky130_fd_sc_hd__xnor2_1_38/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_228 sky130_fd_sc_hd__buf_12_228/A sky130_fd_sc_hd__buf_12_228/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_75 sky130_fd_sc_hd__o21a_1_4/B1 sky130_fd_sc_hd__o21a_1_3/A1
+ sky130_fd_sc_hd__a21oi_1_75/Y sky130_fd_sc_hd__nor2_1_65/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_239 sky130_fd_sc_hd__buf_12_239/A sky130_fd_sc_hd__buf_12_239/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_86 sky130_fd_sc_hd__a211o_1_6/A1 sky130_fd_sc_hd__o21ai_1_100/Y
+ sky130_fd_sc_hd__a21oi_1_86/Y sky130_fd_sc_hd__nand2_1_261/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_97 sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__o21ai_1_112/Y
+ sky130_fd_sc_hd__a21oi_1_97/Y sky130_fd_sc_hd__fa_2_990/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_1_109 sky130_fd_sc_hd__a22oi_1_97/B1 sky130_fd_sc_hd__a22oi_1_97/A1
+ sky130_fd_sc_hd__buf_2_59/X sky130_fd_sc_hd__clkbuf_4_83/X sky130_fd_sc_hd__nand4_1_22/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__fa_2_790 sky130_fd_sc_hd__maj3_1_135/B sky130_fd_sc_hd__maj3_1_136/A
+ sky130_fd_sc_hd__fa_2_790/A sky130_fd_sc_hd__fa_2_790/B sky130_fd_sc_hd__fa_2_791/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor3_1_1 sky130_fd_sc_hd__nor3_1_4/B sky130_fd_sc_hd__nor3_1_1/Y
+ sky130_fd_sc_hd__nor3_2_1/A sky130_fd_sc_hd__nor3_1_1/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__clkinv_1_406 sky130_fd_sc_hd__nand2_1_213/B sky130_fd_sc_hd__nor4_1_7/D
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_406/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_417 sky130_fd_sc_hd__o22ai_1_58/A2 sky130_fd_sc_hd__dfxtp_1_501/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_417/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_428 sky130_fd_sc_hd__nor2_1_40/A sky130_fd_sc_hd__fa_2_967/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_428/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_439 sky130_fd_sc_hd__fa_2_965/B sky130_fd_sc_hd__dfxtp_1_483/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_439/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_6_60 VDD VSS sky130_fd_sc_hd__buf_6_66/A sky130_fd_sc_hd__buf_6_60/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_71 VDD VSS sky130_fd_sc_hd__buf_6_71/X sky130_fd_sc_hd__buf_6_71/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_82 VDD VSS sky130_fd_sc_hd__buf_6_82/X sky130_fd_sc_hd__buf_6_82/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__a21oi_1_303 sky130_fd_sc_hd__o21a_1_33/B1 sky130_fd_sc_hd__o21a_1_32/A1
+ sky130_fd_sc_hd__a21oi_1_303/Y sky130_fd_sc_hd__nor2_1_186/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_314 sky130_fd_sc_hd__o21a_1_41/B1 sky130_fd_sc_hd__nor2_1_197/Y
+ sky130_fd_sc_hd__a21oi_1_314/Y sky130_fd_sc_hd__nor2_1_197/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_40 sky130_fd_sc_hd__buf_2_104/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_325 sky130_fd_sc_hd__o21ai_1_352/Y sky130_fd_sc_hd__nor2_1_215/Y
+ sky130_fd_sc_hd__a21oi_1_325/Y sky130_fd_sc_hd__nor2b_1_112/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_51 sky130_fd_sc_hd__buf_2_75/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_336 sky130_fd_sc_hd__nor2_2_16/Y sky130_fd_sc_hd__o21ai_1_358/Y
+ sky130_fd_sc_hd__nor2_1_216/B sky130_fd_sc_hd__fa_2_1188/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_62 sky130_fd_sc_hd__buf_2_110/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_347 sky130_fd_sc_hd__nor2b_2_3/Y sky130_fd_sc_hd__o21ai_1_373/Y
+ sky130_fd_sc_hd__a21oi_1_347/Y sky130_fd_sc_hd__o21ai_1_380/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_73 sky130_fd_sc_hd__clkbuf_4_86/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_358 sky130_fd_sc_hd__nor3_1_39/A sky130_fd_sc_hd__o22ai_1_321/Y
+ sky130_fd_sc_hd__a21oi_1_358/Y sky130_fd_sc_hd__fa_2_1196/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_84 sky130_fd_sc_hd__nand4_1_45/B VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_369 sky130_fd_sc_hd__o21a_1_50/B1 sky130_fd_sc_hd__o21a_1_49/A1
+ sky130_fd_sc_hd__a21oi_1_369/Y sky130_fd_sc_hd__nor2_1_235/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_95 sky130_fd_sc_hd__clkbuf_1_535/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a222oi_1_6 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1139/A sky130_fd_sc_hd__nor2_2_15/Y
+ sky130_fd_sc_hd__nor3_1_38/A sky130_fd_sc_hd__nor2_2_15/A sky130_fd_sc_hd__xor2_1_164/A
+ sky130_fd_sc_hd__a222oi_1_6/Y sky130_fd_sc_hd__fa_2_1138/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__o221ai_1_0 sky130_fd_sc_hd__nand2b_1_7/Y sky130_fd_sc_hd__o221ai_1_0/Y
+ sky130_fd_sc_hd__fa_2_951/A sky130_fd_sc_hd__o21ai_1_34/Y sky130_fd_sc_hd__fa_2_952/A
+ sky130_fd_sc_hd__o221ai_1_0/B2 VDD VSS VSS VDD sky130_fd_sc_hd__o221ai_1
Xsky130_fd_sc_hd__nand2_1_330 sky130_fd_sc_hd__nand2_1_330/Y sky130_fd_sc_hd__xor2_1_88/A
+ sky130_fd_sc_hd__nand2_2_6/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_341 sky130_fd_sc_hd__nor2_1_182/A sky130_fd_sc_hd__nand2_1_341/B
+ sky130_fd_sc_hd__o32ai_1_2/B2 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_940 sky130_fd_sc_hd__o21a_1_42/A2 sky130_fd_sc_hd__fa_2_1202/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_940/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_352 sky130_fd_sc_hd__o21a_1_26/B1 sky130_fd_sc_hd__fa_2_1150/A
+ sky130_fd_sc_hd__o21a_1_26/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_951 sky130_fd_sc_hd__nor3_1_40/B sky130_fd_sc_hd__o32ai_1_8/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_951/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_363 sky130_fd_sc_hd__nand2_1_363/Y sky130_fd_sc_hd__nand2_1_364/Y
+ sky130_fd_sc_hd__nand2_1_365/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_962 sky130_fd_sc_hd__o31ai_1_9/B1 sky130_fd_sc_hd__a221oi_1_4/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_962/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_374 sky130_fd_sc_hd__nand2_1_374/Y sky130_fd_sc_hd__nand2_1_387/B
+ sky130_fd_sc_hd__o21ai_1_301/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_973 sky130_fd_sc_hd__nor2_1_248/A sky130_fd_sc_hd__or3_1_4/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_973/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_385 sky130_fd_sc_hd__nand2_1_385/Y sky130_fd_sc_hd__nand2_1_387/B
+ sky130_fd_sc_hd__o21ai_1_326/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_984 sky130_fd_sc_hd__nand2_1_475/B sky130_fd_sc_hd__fa_2_158/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_984/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_396 sky130_fd_sc_hd__o21a_1_32/B1 sky130_fd_sc_hd__fa_2_1185/A
+ sky130_fd_sc_hd__o21a_1_32/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_995 sky130_fd_sc_hd__o22ai_1_364/B1 sky130_fd_sc_hd__fa_2_1240/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_995/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_170 VDD VSS sky130_fd_sc_hd__xor2_1_4/B sky130_fd_sc_hd__dfxtp_1_170/CLK
+ sky130_fd_sc_hd__nor2b_1_15/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_181 VDD VSS sky130_fd_sc_hd__ha_2_53/A sky130_fd_sc_hd__dfxtp_1_182/CLK
+ sky130_fd_sc_hd__and2_0_55/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_192 VDD VSS sky130_fd_sc_hd__ha_2_64/A sky130_fd_sc_hd__dfxtp_1_195/CLK
+ sky130_fd_sc_hd__nor2b_1_33/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_2_18 VDD VSS sky130_fd_sc_hd__buf_8_19/A sky130_fd_sc_hd__ha_2_22/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_29 VDD VSS sky130_fd_sc_hd__buf_8_2/A sky130_fd_sc_hd__ha_2_28/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__a21boi_1_2 sky130_fd_sc_hd__a21boi_1_2/Y sky130_fd_sc_hd__nor2_2_15/Y
+ sky130_fd_sc_hd__a21oi_1_285/Y sky130_fd_sc_hd__fa_2_1153/A VDD VSS VDD VSS sky130_fd_sc_hd__a21boi_1
Xsky130_fd_sc_hd__o211ai_1_12 sky130_fd_sc_hd__nor2_1_77/A sky130_fd_sc_hd__a222oi_1_1/Y
+ sky130_fd_sc_hd__xor2_1_40/A sky130_fd_sc_hd__nand2_1_277/Y sky130_fd_sc_hd__nand2_1_275/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_23 sky130_fd_sc_hd__o21a_1_16/X sky130_fd_sc_hd__nor2_1_127/A
+ sky130_fd_sc_hd__xor2_1_95/A sky130_fd_sc_hd__nand2_1_333/Y sky130_fd_sc_hd__nand2_1_334/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_34 sky130_fd_sc_hd__nor2_1_182/A sky130_fd_sc_hd__a21oi_1_294/Y
+ sky130_fd_sc_hd__xor2_1_154/A sky130_fd_sc_hd__nand2_1_388/Y sky130_fd_sc_hd__a21oi_1_286/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_45 sky130_fd_sc_hd__nor2_1_214/A sky130_fd_sc_hd__a222oi_1_20/Y
+ sky130_fd_sc_hd__xor2_1_198/A sky130_fd_sc_hd__nand2_1_439/Y sky130_fd_sc_hd__a21oi_1_344/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_56 sky130_fd_sc_hd__nor2_1_265/A sky130_fd_sc_hd__a211oi_1_30/Y
+ sky130_fd_sc_hd__xor2_1_241/A sky130_fd_sc_hd__nand2_1_489/Y sky130_fd_sc_hd__nand2_1_490/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__fa_2_1280 sky130_fd_sc_hd__fa_2_1281/CIN sky130_fd_sc_hd__mux2_2_252/A1
+ sky130_fd_sc_hd__fa_2_1280/A sky130_fd_sc_hd__fa_2_1280/B sky130_fd_sc_hd__fa_2_1280/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o211ai_1_67 sky130_fd_sc_hd__o21ai_1_473/A2 sky130_fd_sc_hd__nor2_1_307/A
+ sky130_fd_sc_hd__xor2_1_285/A sky130_fd_sc_hd__nand2_1_540/Y sky130_fd_sc_hd__nand2_1_542/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__fa_2_1291 sky130_fd_sc_hd__fa_2_1292/CIN sky130_fd_sc_hd__mux2_2_225/A0
+ sky130_fd_sc_hd__fa_2_1291/A sky130_fd_sc_hd__fa_2_1291/B sky130_fd_sc_hd__fa_2_1291/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_1_203 sky130_fd_sc_hd__clkinv_1_204/A sky130_fd_sc_hd__a22o_4_0/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_203/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_214 sky130_fd_sc_hd__clkinv_2_28/A sky130_fd_sc_hd__a22oi_1_269/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_214/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_225 sky130_fd_sc_hd__clkinv_1_225/Y sky130_fd_sc_hd__clkinv_1_225/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_225/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_236 sky130_fd_sc_hd__buf_12_380/A sky130_fd_sc_hd__clkinv_1_236/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_236/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_247 sky130_fd_sc_hd__clkinv_1_248/A sky130_fd_sc_hd__buf_8_214/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_247/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_258 sky130_fd_sc_hd__nor2_1_8/A sky130_fd_sc_hd__nor2b_1_52/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_258/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_269 sky130_fd_sc_hd__nor2_1_11/B sky130_fd_sc_hd__ha_2_152/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_269/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_100 sky130_fd_sc_hd__a21o_2_3/A2 sky130_fd_sc_hd__o22ai_1_101/Y
+ sky130_fd_sc_hd__a21oi_1_100/Y sky130_fd_sc_hd__fa_2_975/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_111 sky130_fd_sc_hd__clkinv_1_566/Y sky130_fd_sc_hd__o21ai_1_134/Y
+ sky130_fd_sc_hd__a21oi_1_111/Y sky130_fd_sc_hd__a211o_1_6/A1 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_122 sky130_fd_sc_hd__a21o_2_3/X sky130_fd_sc_hd__o22ai_1_131/Y
+ sky130_fd_sc_hd__a21oi_1_122/Y sky130_fd_sc_hd__a211o_1_3/A1 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_133 sky130_fd_sc_hd__a21o_2_3/A2 sky130_fd_sc_hd__o21ai_1_156/Y
+ sky130_fd_sc_hd__a21oi_1_133/Y sky130_fd_sc_hd__fa_2_999/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_144 sky130_fd_sc_hd__nor2_2_10/Y sky130_fd_sc_hd__o22ai_1_144/Y
+ sky130_fd_sc_hd__a21oi_1_144/Y sky130_fd_sc_hd__fa_2_1116/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_155 sky130_fd_sc_hd__nor2_2_11/Y sky130_fd_sc_hd__o22ai_1_154/Y
+ sky130_fd_sc_hd__a21oi_1_155/Y sky130_fd_sc_hd__fa_2_1112/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_166 sky130_fd_sc_hd__clkinv_1_673/Y sky130_fd_sc_hd__nor2_1_98/B
+ sky130_fd_sc_hd__xnor2_1_89/A sky130_fd_sc_hd__xnor2_1_87/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_177 sky130_fd_sc_hd__nand2_1_303/Y sky130_fd_sc_hd__nor2_1_94/A
+ sky130_fd_sc_hd__xnor2_1_72/A sky130_fd_sc_hd__xnor2_1_70/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_188 sky130_fd_sc_hd__nor2_2_13/A sky130_fd_sc_hd__a32o_1_1/B2
+ sky130_fd_sc_hd__a21oi_1_188/Y sky130_fd_sc_hd__a32o_1_1/A3 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_199 sky130_fd_sc_hd__nor2_2_12/Y sky130_fd_sc_hd__o211ai_1_16/Y
+ sky130_fd_sc_hd__a21oi_1_199/Y sky130_fd_sc_hd__fa_2_1067/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_107 sky130_fd_sc_hd__buf_8_107/A sky130_fd_sc_hd__buf_8_107/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_118 sky130_fd_sc_hd__buf_4_69/A sky130_fd_sc_hd__buf_4_73/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_129 sky130_fd_sc_hd__inv_2_89/Y sky130_fd_sc_hd__buf_8_129/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nand2_1_160 sky130_fd_sc_hd__fa_2_204/A sky130_fd_sc_hd__fa_2_277/B
+ sky130_fd_sc_hd__fa_2_273/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_171 sky130_fd_sc_hd__fa_2_370/A sky130_fd_sc_hd__fa_2_404/B
+ sky130_fd_sc_hd__fa_2_422/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_770 sky130_fd_sc_hd__fa_2_1121/B sky130_fd_sc_hd__nor2_2_11/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_770/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_182 sky130_fd_sc_hd__fa_2_555/B sky130_fd_sc_hd__fa_2_566/B
+ sky130_fd_sc_hd__fa_2_427/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_781 sky130_fd_sc_hd__nand2_1_387/B sky130_fd_sc_hd__nor2_1_182/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_781/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_193 sky130_fd_sc_hd__fa_2_745/A sky130_fd_sc_hd__ha_2_140/A
+ sky130_fd_sc_hd__ha_2_145/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_792 sky130_fd_sc_hd__o32ai_1_1/A2 sky130_fd_sc_hd__fa_2_1140/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_792/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21o_2_19 sky130_fd_sc_hd__a21o_2_19/X sky130_fd_sc_hd__nor2_1_252/Y
+ sky130_fd_sc_hd__nor2_1_252/A sky130_fd_sc_hd__nor2_1_252/B VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__xor2_1_13 sky130_fd_sc_hd__or4_1_1/A sky130_fd_sc_hd__xor2_1_13/X
+ sky130_fd_sc_hd__xor2_1_13/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_24 sky130_fd_sc_hd__xor2_1_24/B sky130_fd_sc_hd__xor2_1_24/X
+ sky130_fd_sc_hd__xor2_1_24/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_35 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_992/B
+ sky130_fd_sc_hd__xor2_1_35/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_46 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_981/B
+ sky130_fd_sc_hd__xor2_1_46/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_57 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__xor2_1_57/X
+ sky130_fd_sc_hd__xor2_1_57/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_68 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__xor2_1_68/X
+ sky130_fd_sc_hd__xor2_1_68/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_79 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__fa_2_997/B
+ sky130_fd_sc_hd__xor2_1_79/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2b_1_7 sky130_fd_sc_hd__nand2b_1_7/Y sky130_fd_sc_hd__nor2b_1_86/Y
+ sky130_fd_sc_hd__nand2b_1_7/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a21o_2_3 sky130_fd_sc_hd__a21o_2_3/X sky130_fd_sc_hd__a21o_2_3/B1
+ sky130_fd_sc_hd__fa_2_1006/A sky130_fd_sc_hd__a21o_2_3/A2 VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__dfxtp_1_906 VDD VSS sky130_fd_sc_hd__fa_2_941/B sky130_fd_sc_hd__clkinv_4_22/Y
+ sky130_fd_sc_hd__o21a_1_18/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_917 VDD VSS sky130_fd_sc_hd__fa_2_1146/A sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__mux2_2_104/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_928 VDD VSS sky130_fd_sc_hd__fa_2_1157/A sky130_fd_sc_hd__clkinv_8_46/Y
+ sky130_fd_sc_hd__mux2_2_78/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_939 VDD VSS sky130_fd_sc_hd__fa_2_1131/A sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__mux2_2_96/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a221oi_1_5 sky130_fd_sc_hd__a221oi_1_5/Y sky130_fd_sc_hd__nor2_1_286/A
+ sky130_fd_sc_hd__xor2_1_275/B sky130_fd_sc_hd__nand2_1_522/Y sky130_fd_sc_hd__o31ai_1_12/A3
+ sky130_fd_sc_hd__nor2_1_290/B VSS VDD VDD VSS sky130_fd_sc_hd__a221oi_1
Xsky130_fd_sc_hd__clkbuf_1_504 VSS VDD sky130_fd_sc_hd__buf_8_213/A sky130_fd_sc_hd__a22o_4_0/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_515 VSS VDD sky130_fd_sc_hd__clkbuf_1_515/X sky130_fd_sc_hd__buf_8_197/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_526 VSS VDD sky130_fd_sc_hd__clkbuf_1_526/X sky130_fd_sc_hd__clkbuf_1_527/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_537 VSS VDD sky130_fd_sc_hd__clkbuf_4_170/A sky130_fd_sc_hd__clkbuf_1_538/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_105 VSS VDD VSS VDD sky130_fd_sc_hd__fa_2_2/A sky130_fd_sc_hd__fa_2_254/B
+ sky130_fd_sc_hd__fa_2_250/B sky130_fd_sc_hd__ha_2_96/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_548 VSS VDD sky130_fd_sc_hd__ha_2_107/A sky130_fd_sc_hd__ha_2_99/B
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_116 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_116/A sky130_fd_sc_hd__fa_2_409/B
+ sky130_fd_sc_hd__ha_2_116/SUM sky130_fd_sc_hd__ha_2_116/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_559 VSS VDD sky130_fd_sc_hd__nand2_1_91/B sky130_fd_sc_hd__nand4_1_59/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_127 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_130/A sky130_fd_sc_hd__fa_2_585/B
+ sky130_fd_sc_hd__ha_2_127/SUM sky130_fd_sc_hd__ha_2_131/A sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_138 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_138/A sky130_fd_sc_hd__fa_2_720/B
+ sky130_fd_sc_hd__ha_2_138/SUM sky130_fd_sc_hd__ha_2_141/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_149 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_149/A sky130_fd_sc_hd__ha_2_148/B
+ sky130_fd_sc_hd__ha_2_149/SUM sky130_fd_sc_hd__ha_2_149/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_40 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_40/A sky130_fd_sc_hd__xor2_1_4/A
+ sky130_fd_sc_hd__ha_2_40/SUM sky130_fd_sc_hd__ha_2_40/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__maj3_1_9 sky130_fd_sc_hd__maj3_1_9/C sky130_fd_sc_hd__maj3_1_9/X
+ sky130_fd_sc_hd__maj3_1_9/B sky130_fd_sc_hd__maj3_1_9/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__ha_2_51 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_51/A sky130_fd_sc_hd__ha_2_50/B
+ sky130_fd_sc_hd__ha_2_51/SUM sky130_fd_sc_hd__ha_2_51/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_62 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_62/A sky130_fd_sc_hd__ha_2_61/B
+ sky130_fd_sc_hd__ha_2_62/SUM sky130_fd_sc_hd__ha_2_62/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_73 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_73/A sky130_fd_sc_hd__ha_2_72/B
+ sky130_fd_sc_hd__ha_2_73/SUM sky130_fd_sc_hd__ha_2_73/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_84 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_84/A sky130_fd_sc_hd__ha_2_83/B
+ sky130_fd_sc_hd__ha_2_84/SUM sky130_fd_sc_hd__ha_2_84/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_95 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_95/A sky130_fd_sc_hd__fa_2_96/CIN
+ sky130_fd_sc_hd__fa_2_88/A sky130_fd_sc_hd__ha_2_95/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_3 VSS VDD sky130_fd_sc_hd__buf_4_1/A sky130_fd_sc_hd__clkbuf_1_3/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__sdlclkp_4_80 sky130_fd_sc_hd__conb_1_25/LO sky130_fd_sc_hd__clkinv_8_72/A
+ sky130_fd_sc_hd__dfxtp_1_899/CLK sky130_fd_sc_hd__or2_0_9/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_91 sky130_fd_sc_hd__conb_1_28/LO sky130_fd_sc_hd__clkinv_8_47/A
+ sky130_fd_sc_hd__dfxtp_1_1326/CLK sky130_fd_sc_hd__or2_0_12/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__clkinv_1_3 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__nor2_4_2/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_3/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_160 sky130_fd_sc_hd__nor2_1_163/A sky130_fd_sc_hd__nor2_1_160/Y
+ sky130_fd_sc_hd__o31ai_1_6/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_171 sky130_fd_sc_hd__or3_1_2/X sky130_fd_sc_hd__nor2_1_171/Y
+ sky130_fd_sc_hd__nor2_1_171/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_182 sky130_fd_sc_hd__o21a_1_29/A1 sky130_fd_sc_hd__nor2_1_182/Y
+ sky130_fd_sc_hd__nor2_1_182/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_193 sky130_fd_sc_hd__nor2_1_193/B sky130_fd_sc_hd__o21a_1_37/A1
+ sky130_fd_sc_hd__o21a_1_38/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_80 sky130_fd_sc_hd__clkbuf_4_8/X sky130_fd_sc_hd__clkbuf_4_9/X
+ sky130_fd_sc_hd__clkbuf_1_19/X sky130_fd_sc_hd__a22oi_1_80/A2 sky130_fd_sc_hd__a22oi_1_80/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_91 sky130_fd_sc_hd__clkbuf_4_72/X sky130_fd_sc_hd__clkbuf_4_73/X
+ sky130_fd_sc_hd__a22oi_1_91/B2 sky130_fd_sc_hd__buf_2_96/X sky130_fd_sc_hd__buf_2_111/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__and2_0_18 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_18/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_15/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_29 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_29/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__xor2_1_3/X sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__o22ai_1_309 sky130_fd_sc_hd__o22ai_1_322/A2 sky130_fd_sc_hd__o22ai_1_309/B1
+ sky130_fd_sc_hd__o22ai_1_309/Y sky130_fd_sc_hd__nor2_1_187/B sky130_fd_sc_hd__o32ai_1_5/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__a22oi_1_270 sky130_fd_sc_hd__clkbuf_1_378/X sky130_fd_sc_hd__clkbuf_1_379/X
+ sky130_fd_sc_hd__clkbuf_4_173/X sky130_fd_sc_hd__buf_2_199/X sky130_fd_sc_hd__nand4_1_67/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_281 sky130_fd_sc_hd__clkbuf_4_165/X sky130_fd_sc_hd__clkinv_2_23/Y
+ sky130_fd_sc_hd__clkbuf_1_407/X sky130_fd_sc_hd__a22oi_1_281/A2 sky130_fd_sc_hd__a22oi_1_281/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_292 sky130_fd_sc_hd__clkbuf_1_376/X sky130_fd_sc_hd__nor2_2_5/Y
+ sky130_fd_sc_hd__buf_2_209/X sky130_fd_sc_hd__clkbuf_1_465/X sky130_fd_sc_hd__nand4_1_72/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_4_110 VDD VSS sky130_fd_sc_hd__buf_4_119/A sky130_fd_sc_hd__buf_4_110/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_121 VDD VSS sky130_fd_sc_hd__buf_4_121/X sky130_fd_sc_hd__buf_4_64/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_8_17 sky130_fd_sc_hd__inv_2_10/Y sky130_fd_sc_hd__buf_8_17/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_28 sky130_fd_sc_hd__ha_2_27/A sky130_fd_sc_hd__buf_8_28/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_39 sky130_fd_sc_hd__inv_2_37/Y sky130_fd_sc_hd__buf_8_39/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__clkinv_4_80 sky130_fd_sc_hd__clkinv_4_80/A sky130_fd_sc_hd__clkinv_4_80/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_80/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__o21ai_1_503 VSS VDD sky130_fd_sc_hd__nand2_1_564/A sky130_fd_sc_hd__o21ai_1_507/A1
+ sky130_fd_sc_hd__nand2_1_564/Y sky130_fd_sc_hd__and2_0_348/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1109 VDD VSS sky130_fd_sc_hd__mux2_2_135/S sky130_fd_sc_hd__clkinv_4_23/Y
+ sky130_fd_sc_hd__nor2b_1_117/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_703 VDD VSS sky130_fd_sc_hd__mux2_2_27/A1 sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__o21ai_1_43/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_714 VDD VSS sky130_fd_sc_hd__mux2_2_5/A1 sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__o21ai_1_54/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_725 VDD VSS sky130_fd_sc_hd__mux2_2_22/A1 sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__o21ai_1_62/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_736 VDD VSS sky130_fd_sc_hd__mux2_2_0/A1 sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__o21ai_1_73/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_747 VDD VSS sky130_fd_sc_hd__and2_0_168/A sky130_fd_sc_hd__dfxtp_1_747/CLK
+ sky130_fd_sc_hd__fa_2_1102/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_758 VDD VSS sky130_fd_sc_hd__ha_2_133/A sky130_fd_sc_hd__dfxtp_1_764/CLK
+ sky130_fd_sc_hd__dfxtp_1_758/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_769 VDD VSS sky130_fd_sc_hd__or2_0_8/A sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__nor2b_1_98/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_301 VSS VDD sky130_fd_sc_hd__nand4_1_44/D sky130_fd_sc_hd__a22oi_1_195/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_312 VSS VDD sky130_fd_sc_hd__nand4_1_33/D sky130_fd_sc_hd__a22oi_1_151/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_323 VSS VDD sky130_fd_sc_hd__buf_8_125/A sky130_fd_sc_hd__and2_1_5/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_334 VSS VDD sky130_fd_sc_hd__buf_8_130/A sky130_fd_sc_hd__buf_8_155/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_345 VSS VDD sky130_fd_sc_hd__buf_8_150/A sky130_fd_sc_hd__buf_2_126/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_356 VSS VDD sky130_fd_sc_hd__buf_8_141/A sky130_fd_sc_hd__buf_6_37/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_367 VSS VDD sky130_fd_sc_hd__clkinv_4_16/A sky130_fd_sc_hd__buf_8_149/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_378 VSS VDD sky130_fd_sc_hd__clkbuf_1_378/X sky130_fd_sc_hd__nor3_1_22/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_389 VSS VDD sky130_fd_sc_hd__a22oi_2_22/B2 sky130_fd_sc_hd__clkbuf_1_389/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_608 sky130_fd_sc_hd__fa_2_610/B sky130_fd_sc_hd__fa_2_608/SUM
+ sky130_fd_sc_hd__fa_2_608/A sky130_fd_sc_hd__fa_2_608/B sky130_fd_sc_hd__fa_2_612/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_619 sky130_fd_sc_hd__fa_2_622/B sky130_fd_sc_hd__fa_2_619/SUM
+ sky130_fd_sc_hd__fa_2_619/A sky130_fd_sc_hd__fa_2_619/B sky130_fd_sc_hd__o22ai_1_43/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_60 VDD VSS sky130_fd_sc_hd__ha_2_125/A sky130_fd_sc_hd__dfxtp_1_60/CLK
+ sky130_fd_sc_hd__dfxtp_1_60/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_71 VDD VSS sky130_fd_sc_hd__ha_2_91/B sky130_fd_sc_hd__dfxtp_1_73/CLK
+ sky130_fd_sc_hd__buf_2_289/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_82 VDD VSS sky130_fd_sc_hd__dfxtp_1_82/Q sky130_fd_sc_hd__dfxtp_1_83/CLK
+ sky130_fd_sc_hd__dfxtp_1_83/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_93 VDD VSS sky130_fd_sc_hd__a22o_1_9/B2 sky130_fd_sc_hd__dfxtp_1_93/CLK
+ sky130_fd_sc_hd__dfxtp_1_93/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_310 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_310/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_310/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_150 sky130_fd_sc_hd__nand4_1_35/B sky130_fd_sc_hd__a22oi_1_161/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_321 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_321/X sky130_fd_sc_hd__mux2_2_99/S
+ sky130_fd_sc_hd__and2_0_321/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_161 sky130_fd_sc_hd__clkbuf_4_161/X sky130_fd_sc_hd__buf_2_139/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_332 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_332/X sky130_fd_sc_hd__inv_2_139/Y
+ sky130_fd_sc_hd__and2_0_332/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_172 sky130_fd_sc_hd__clkbuf_4_172/X sky130_fd_sc_hd__clkbuf_4_172/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_343 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_343/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_343/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_183 sky130_fd_sc_hd__clkbuf_4_183/X sky130_fd_sc_hd__clkbuf_4_183/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_354 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_354/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_354/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_194 sky130_fd_sc_hd__nand4_1_78/D sky130_fd_sc_hd__a22oi_1_313/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__conb_1_7 sky130_fd_sc_hd__conb_1_7/LO sky130_fd_sc_hd__conb_1_7/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__inv_2_110 sky130_fd_sc_hd__inv_2_110/A sky130_fd_sc_hd__inv_2_131/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__or2_0_1 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__or2_0_1/X sky130_fd_sc_hd__or2_0_1/B
+ VSS VDD VSS VDD sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__inv_2_121 sky130_fd_sc_hd__inv_2_121/A sky130_fd_sc_hd__inv_2_121/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_132 sky130_fd_sc_hd__inv_2_132/A sky130_fd_sc_hd__inv_2_132/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__o22ai_1_106 sky130_fd_sc_hd__o22ai_1_132/B1 sky130_fd_sc_hd__o22ai_1_119/A1
+ sky130_fd_sc_hd__o22ai_1_106/Y sky130_fd_sc_hd__o22ai_1_120/B1 sky130_fd_sc_hd__o21ai_1_92/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_117 sky130_fd_sc_hd__o22ai_1_130/B1 sky130_fd_sc_hd__nor2_1_66/B
+ sky130_fd_sc_hd__nor2_1_84/A sky130_fd_sc_hd__o22ai_1_117/A1 sky130_fd_sc_hd__o22ai_1_132/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_128 sky130_fd_sc_hd__nor2_1_87/A sky130_fd_sc_hd__o22ai_1_130/B1
+ sky130_fd_sc_hd__o22ai_1_128/Y sky130_fd_sc_hd__o22ai_1_132/B1 sky130_fd_sc_hd__nor2_1_88/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_139 sky130_fd_sc_hd__nand2_1_284/Y sky130_fd_sc_hd__nand2_2_5/Y
+ sky130_fd_sc_hd__o22ai_1_139/Y sky130_fd_sc_hd__xnor2_1_70/Y sky130_fd_sc_hd__o22ai_1_153/B2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_2_17 sky130_fd_sc_hd__nor2_2_17/B sky130_fd_sc_hd__nor2_2_17/Y
+ sky130_fd_sc_hd__nor2_4_18/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__o211ai_1_7 sky130_fd_sc_hd__nor2_1_76/A sky130_fd_sc_hd__nor2_1_79/Y
+ sky130_fd_sc_hd__xor2_1_80/A sky130_fd_sc_hd__o211ai_1_7/C1 sky130_fd_sc_hd__o211ai_1_7/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__a31oi_1_4 VSS VDD sky130_fd_sc_hd__a31oi_1_4/Y sky130_fd_sc_hd__a31oi_1_4/B1
+ sky130_fd_sc_hd__a31oi_1_4/A2 sky130_fd_sc_hd__a31oi_1_4/A1 sky130_fd_sc_hd__a31oi_1_4/A3
+ VDD VSS sky130_fd_sc_hd__a31oi_1
Xsky130_fd_sc_hd__a211o_1_0 VSS VDD VSS VDD sky130_fd_sc_hd__a211o_1_0/X sky130_fd_sc_hd__nor3_1_27/A
+ sky130_fd_sc_hd__nor2_1_16/Y sky130_fd_sc_hd__nor3_1_27/C sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o21ai_1_300 VSS VDD sky130_fd_sc_hd__o22ai_1_265/A2 sky130_fd_sc_hd__nor2_1_176/A
+ sky130_fd_sc_hd__a22oi_1_374/Y sky130_fd_sc_hd__o21ai_1_300/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_311 VSS VDD sky130_fd_sc_hd__o21ai_1_311/A2 sky130_fd_sc_hd__nor2_1_182/A
+ sky130_fd_sc_hd__nand2_1_382/Y sky130_fd_sc_hd__xor2_1_146/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_322 VSS VDD sky130_fd_sc_hd__o22ai_1_261/A2 sky130_fd_sc_hd__nor2_1_181/A
+ sky130_fd_sc_hd__a21oi_1_292/Y sky130_fd_sc_hd__o21ai_1_322/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_333 VSS VDD sky130_fd_sc_hd__nand2_1_421/B sky130_fd_sc_hd__nor2_1_210/Y
+ sky130_fd_sc_hd__nor2_1_209/B sky130_fd_sc_hd__o21ai_1_333/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_344 VSS VDD sky130_fd_sc_hd__nor2_1_214/B sky130_fd_sc_hd__nor2_1_224/A
+ sky130_fd_sc_hd__nand2_1_425/Y sky130_fd_sc_hd__xor2_1_212/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_355 VSS VDD sky130_fd_sc_hd__nor2_1_185/B sky130_fd_sc_hd__o21a_1_42/A1
+ sky130_fd_sc_hd__a21oi_1_334/Y sky130_fd_sc_hd__o21ai_1_355/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_60 sky130_fd_sc_hd__o21a_1_60/X sky130_fd_sc_hd__o21a_1_60/A1
+ sky130_fd_sc_hd__o21a_1_60/B1 sky130_fd_sc_hd__fa_2_1283/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__a211oi_1_16 sky130_fd_sc_hd__nor3_1_38/A sky130_fd_sc_hd__nor2_1_181/Y
+ sky130_fd_sc_hd__o22ai_1_259/Y sky130_fd_sc_hd__a211oi_1_16/Y sky130_fd_sc_hd__fa_2_1154/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_366 VSS VDD sky130_fd_sc_hd__a211oi_1_23/Y sky130_fd_sc_hd__nor2_1_224/A
+ sky130_fd_sc_hd__nand2_1_434/Y sky130_fd_sc_hd__xor2_1_192/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a211oi_1_27 sky130_fd_sc_hd__nor2b_2_4/Y sky130_fd_sc_hd__o22ai_1_363/Y
+ sky130_fd_sc_hd__nor2_1_260/Y sky130_fd_sc_hd__a211oi_1_27/Y sky130_fd_sc_hd__o21ai_1_415/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_377 VSS VDD sky130_fd_sc_hd__nor2_1_193/B sky130_fd_sc_hd__o21a_1_42/A1
+ sky130_fd_sc_hd__a21oi_1_353/Y sky130_fd_sc_hd__o21ai_1_377/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a211oi_1_38 sky130_fd_sc_hd__nor2b_2_5/Y sky130_fd_sc_hd__o22ai_1_433/Y
+ sky130_fd_sc_hd__nor2_1_310/Y sky130_fd_sc_hd__a211oi_1_38/Y sky130_fd_sc_hd__o21ai_1_491/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_388 VSS VDD sky130_fd_sc_hd__nand2_1_474/B sky130_fd_sc_hd__nor2_1_254/Y
+ sky130_fd_sc_hd__nor2_1_253/B sky130_fd_sc_hd__o21ai_1_388/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_399 VSS VDD sky130_fd_sc_hd__nor2_1_259/B sky130_fd_sc_hd__nor2_1_267/A
+ sky130_fd_sc_hd__nand2_1_477/Y sky130_fd_sc_hd__xor2_1_258/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__mux2_2_13 VSS VDD sky130_fd_sc_hd__mux2_2_13/A1 sky130_fd_sc_hd__mux2_2_13/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_13/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_24 VSS VDD sky130_fd_sc_hd__mux2_2_24/A1 sky130_fd_sc_hd__mux2_2_24/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_24/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_35 VSS VDD sky130_fd_sc_hd__mux2_2_35/A1 sky130_fd_sc_hd__mux2_2_35/A0
+ sky130_fd_sc_hd__mux2_2_37/S sky130_fd_sc_hd__mux2_2_35/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_46 VSS VDD sky130_fd_sc_hd__mux2_2_46/A1 sky130_fd_sc_hd__mux2_2_46/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_46/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_57 VSS VDD sky130_fd_sc_hd__mux2_2_57/A1 sky130_fd_sc_hd__mux2_2_57/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_57/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_68 VSS VDD sky130_fd_sc_hd__mux2_2_68/A1 sky130_fd_sc_hd__mux2_2_68/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_68/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_79 VSS VDD sky130_fd_sc_hd__mux2_2_79/A1 sky130_fd_sc_hd__mux2_2_79/A0
+ sky130_fd_sc_hd__nor2_4_15/A sky130_fd_sc_hd__mux2_2_79/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__fa_2_1109 sky130_fd_sc_hd__fa_2_1110/CIN sky130_fd_sc_hd__fa_2_1109/SUM
+ sky130_fd_sc_hd__fa_2_1109/A sky130_fd_sc_hd__fa_2_1109/B sky130_fd_sc_hd__fa_2_1109/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_500 VDD VSS sky130_fd_sc_hd__o21ai_1_36/A1 sky130_fd_sc_hd__dfxtp_1_502/CLK
+ sky130_fd_sc_hd__nor2b_1_77/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_160 sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__fa_2_1123/B
+ sky130_fd_sc_hd__xor2_1_160/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_511 VDD VSS sky130_fd_sc_hd__nor4_1_11/A sky130_fd_sc_hd__dfxtp_1_520/CLK
+ sky130_fd_sc_hd__a22o_1_60/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_171 sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__fa_2_1151/B
+ sky130_fd_sc_hd__xor2_1_171/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_522 VDD VSS sky130_fd_sc_hd__fa_2_969/A sky130_fd_sc_hd__dfxtp_1_538/CLK
+ sky130_fd_sc_hd__and2_0_266/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_182 sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__xor2_1_182/X
+ sky130_fd_sc_hd__xor2_1_182/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_193 sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__fa_2_1186/B
+ sky130_fd_sc_hd__xor2_1_193/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_533 VDD VSS sky130_fd_sc_hd__or3_1_1/B sky130_fd_sc_hd__dfxtp_1_533/CLK
+ sky130_fd_sc_hd__and2_0_257/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_544 VDD VSS sky130_fd_sc_hd__fa_2_947/A sky130_fd_sc_hd__dfxtp_1_544/CLK
+ sky130_fd_sc_hd__a22o_1_41/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_555 VDD VSS sky130_fd_sc_hd__and2_0_222/A sky130_fd_sc_hd__dfxtp_1_571/CLK
+ sky130_fd_sc_hd__dfxtp_1_556/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_566 VDD VSS sky130_fd_sc_hd__a22o_1_34/B1 sky130_fd_sc_hd__dfxtp_1_576/CLK
+ sky130_fd_sc_hd__a22o_1_34/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_577 VDD VSS sky130_fd_sc_hd__and2_0_200/A sky130_fd_sc_hd__dfxtp_1_577/CLK
+ sky130_fd_sc_hd__nand2_1_206/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_588 VDD VSS sky130_fd_sc_hd__nor4_1_8/C sky130_fd_sc_hd__dfxtp_1_594/CLK
+ sky130_fd_sc_hd__and2_0_253/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_599 VDD VSS sky130_fd_sc_hd__and2_0_209/A sky130_fd_sc_hd__dfxtp_1_601/CLK
+ sky130_fd_sc_hd__fa_2_1019/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_120 VSS VDD sky130_fd_sc_hd__buf_4_3/A sky130_fd_sc_hd__buf_6_2/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_131 VSS VDD sky130_fd_sc_hd__buf_6_19/A sky130_fd_sc_hd__buf_4_32/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_142 VSS VDD sky130_fd_sc_hd__clkbuf_1_142/X sky130_fd_sc_hd__clkbuf_1_142/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_0 VDD VSS sky130_fd_sc_hd__dfxtp_1_0/Q sky130_fd_sc_hd__dfxtp_1_8/CLK
+ sky130_fd_sc_hd__nor2b_1_0/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_153 VSS VDD sky130_fd_sc_hd__a22oi_1_88/B2 sky130_fd_sc_hd__clkbuf_1_153/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_164 VSS VDD sky130_fd_sc_hd__clkbuf_1_164/X sky130_fd_sc_hd__clkbuf_1_248/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_175 VSS VDD sky130_fd_sc_hd__nand4_1_31/B sky130_fd_sc_hd__a22oi_1_145/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_186 VSS VDD sky130_fd_sc_hd__nand4_1_19/B sky130_fd_sc_hd__a22oi_1_98/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_197 VSS VDD sky130_fd_sc_hd__buf_8_105/A sky130_fd_sc_hd__buf_8_86/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_405 sky130_fd_sc_hd__fa_2_407/B sky130_fd_sc_hd__fa_2_402/A
+ sky130_fd_sc_hd__fa_2_413/A sky130_fd_sc_hd__fa_2_405/B sky130_fd_sc_hd__ha_2_116/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_416 sky130_fd_sc_hd__fa_2_415/A sky130_fd_sc_hd__fa_2_411/A
+ sky130_fd_sc_hd__fa_2_424/A sky130_fd_sc_hd__fa_2_416/B sky130_fd_sc_hd__fa_2_422/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_427 sky130_fd_sc_hd__xnor2_1_3/A sky130_fd_sc_hd__fa_2_427/SUM
+ sky130_fd_sc_hd__ha_2_124/A sky130_fd_sc_hd__fa_2_427/B sky130_fd_sc_hd__fa_2_427/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_438 sky130_fd_sc_hd__fa_2_434/A sky130_fd_sc_hd__fa_2_433/B
+ sky130_fd_sc_hd__fa_2_566/B sky130_fd_sc_hd__fa_2_438/B sky130_fd_sc_hd__fa_2_534/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_449 sky130_fd_sc_hd__fa_2_446/CIN sky130_fd_sc_hd__fa_2_451/CIN
+ sky130_fd_sc_hd__fa_2_566/A sky130_fd_sc_hd__fa_2_543/A sky130_fd_sc_hd__fa_2_449/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nand3_1_20 sky130_fd_sc_hd__nand3_1_20/Y sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__ha_2_20/A VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_31 sky130_fd_sc_hd__nand3_1_31/Y sky130_fd_sc_hd__nand2_2_0/B
+ sky130_fd_sc_hd__nand3_1_31/C sky130_fd_sc_hd__nand3_1_31/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_42 sky130_fd_sc_hd__o31ai_1_0/B1 sky130_fd_sc_hd__ha_2_167/B
+ sky130_fd_sc_hd__o31ai_1_0/A3 sky130_fd_sc_hd__xor2_1_9/X VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__dfxtp_1_1440 VDD VSS sky130_fd_sc_hd__mux2_2_222/A1 sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__o31ai_1_11/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1451 VDD VSS sky130_fd_sc_hd__buf_4_66/A sky130_fd_sc_hd__sdlclkp_1_6/GCLK
+ sky130_fd_sc_hd__and2_0_354/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1462 VDD VSS sky130_fd_sc_hd__buf_2_274/A sky130_fd_sc_hd__dfxtp_1_1464/CLK
+ sky130_fd_sc_hd__and2_0_343/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_140 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_140/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_923/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_151 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_151/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__fa_2_872/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_162 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_162/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_846/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_70 sky130_fd_sc_hd__clkinv_1_71/A sky130_fd_sc_hd__dfxtp_1_255/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_70/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_173 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_173/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_173/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_81 sky130_fd_sc_hd__buf_8_81/A sky130_fd_sc_hd__clkinv_1_81/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_81/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_184 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_184/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_184/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_92 sky130_fd_sc_hd__clkinv_1_92/Y sky130_fd_sc_hd__clkinv_1_92/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_92/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_195 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_195/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_902/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__fa_2_950 sky130_fd_sc_hd__fa_2_949/CIN sky130_fd_sc_hd__fa_2_950/SUM
+ sky130_fd_sc_hd__or3_1_0/B sky130_fd_sc_hd__fa_2_950/B sky130_fd_sc_hd__fa_2_950/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_961 sky130_fd_sc_hd__fa_2_960/CIN sky130_fd_sc_hd__fa_2_961/SUM
+ sky130_fd_sc_hd__fa_2_961/A sky130_fd_sc_hd__fa_2_961/B sky130_fd_sc_hd__fa_2_961/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_972 sky130_fd_sc_hd__fa_2_973/CIN sky130_fd_sc_hd__fa_2_972/SUM
+ sky130_fd_sc_hd__fa_2_972/A sky130_fd_sc_hd__fa_2_972/B sky130_fd_sc_hd__fa_2_972/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_983 sky130_fd_sc_hd__fa_2_984/CIN sky130_fd_sc_hd__mux2_2_21/A0
+ sky130_fd_sc_hd__fa_2_983/A sky130_fd_sc_hd__fa_2_983/B sky130_fd_sc_hd__fa_2_983/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_994 sky130_fd_sc_hd__fa_2_995/CIN sky130_fd_sc_hd__fa_2_994/SUM
+ sky130_fd_sc_hd__fa_2_994/A sky130_fd_sc_hd__fa_2_994/B sky130_fd_sc_hd__fa_2_994/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_1_1 sky130_fd_sc_hd__conb_1_11/LO sky130_fd_sc_hd__clkinv_4_74/A
+ sky130_fd_sc_hd__dfxtp_1_166/CLK sky130_fd_sc_hd__or2_1_0/X VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_1
Xsky130_fd_sc_hd__mux2_2_250 VSS VDD sky130_fd_sc_hd__mux2_2_250/A1 sky130_fd_sc_hd__mux2_2_250/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_250/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_261 VSS VDD sky130_fd_sc_hd__mux2_2_261/A1 sky130_fd_sc_hd__mux2_2_261/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_261/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__o21ai_1_130 VSS VDD sky130_fd_sc_hd__a21oi_1_127/Y sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__nand2b_1_13/Y sky130_fd_sc_hd__o21ai_1_130/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_141 VSS VDD sky130_fd_sc_hd__a21oi_1_134/Y sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__a21oi_1_117/Y sky130_fd_sc_hd__xor2_1_49/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_152 VSS VDD sky130_fd_sc_hd__o21ai_1_152/A2 sky130_fd_sc_hd__o21ai_1_92/A1
+ sky130_fd_sc_hd__a22oi_1_342/Y sky130_fd_sc_hd__o21ai_1_152/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_163 VSS VDD sky130_fd_sc_hd__o21ai_1_171/A2 sky130_fd_sc_hd__xnor2_1_73/Y
+ sky130_fd_sc_hd__a21oi_1_140/Y sky130_fd_sc_hd__o21ai_1_163/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_174 VSS VDD sky130_fd_sc_hd__nand2_2_5/Y sky130_fd_sc_hd__o21ai_1_191/A2
+ sky130_fd_sc_hd__nand2_1_285/Y sky130_fd_sc_hd__o21ai_1_174/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_185 VSS VDD sky130_fd_sc_hd__nand2_2_5/Y sky130_fd_sc_hd__xnor2_1_83/Y
+ sky130_fd_sc_hd__a21oi_1_160/Y sky130_fd_sc_hd__o21ai_1_185/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_196 VSS VDD sky130_fd_sc_hd__xnor2_1_73/A sky130_fd_sc_hd__o21ai_1_196/A1
+ sky130_fd_sc_hd__nand2_1_289/B sky130_fd_sc_hd__xnor2_1_75/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a222oi_1_19 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1175/A sky130_fd_sc_hd__nor2_2_16/Y
+ sky130_fd_sc_hd__nor3_1_39/A sky130_fd_sc_hd__fa_2_1177/A sky130_fd_sc_hd__nor3_1_39/B
+ sky130_fd_sc_hd__a222oi_1_19/Y sky130_fd_sc_hd__fa_2_1174/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2_1_501 sky130_fd_sc_hd__o21a_1_59/B1 sky130_fd_sc_hd__fa_2_1285/A
+ sky130_fd_sc_hd__o21a_1_59/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_512 sky130_fd_sc_hd__o32ai_1_11/B1 sky130_fd_sc_hd__o32ai_1_11/A3
+ sky130_fd_sc_hd__o21bai_1_5/A2 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_80 sky130_fd_sc_hd__maj3_1_81/X sky130_fd_sc_hd__maj3_1_80/X
+ sky130_fd_sc_hd__maj3_1_80/B sky130_fd_sc_hd__maj3_1_80/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_523 sky130_fd_sc_hd__o31ai_1_12/A2 sky130_fd_sc_hd__nand2_1_523/B
+ sky130_fd_sc_hd__nor2_1_293/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_91 sky130_fd_sc_hd__maj3_1_92/X sky130_fd_sc_hd__maj3_1_91/X
+ sky130_fd_sc_hd__maj3_1_91/B sky130_fd_sc_hd__maj3_1_91/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_534 sky130_fd_sc_hd__nand2_1_534/Y sky130_fd_sc_hd__nand2_1_543/B
+ sky130_fd_sc_hd__o21ai_1_456/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_545 sky130_fd_sc_hd__nand2_1_545/Y sky130_fd_sc_hd__nor2b_1_126/Y
+ sky130_fd_sc_hd__o21ai_1_485/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_556 sky130_fd_sc_hd__nand2_1_556/Y sky130_fd_sc_hd__buf_2_275/X
+ sky130_fd_sc_hd__nand2_1_556/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_567 sky130_fd_sc_hd__nand2_1_567/Y sky130_fd_sc_hd__nand2_1_567/B
+ sky130_fd_sc_hd__nand2_1_567/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_3 sky130_fd_sc_hd__nor2b_1_3/B_N sky130_fd_sc_hd__nor2b_1_3/Y
+ sky130_fd_sc_hd__or2_0_1/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1103 sky130_fd_sc_hd__nor2_1_281/B sky130_fd_sc_hd__fa_2_1300/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1103/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1114 sky130_fd_sc_hd__nor4_1_13/D sky130_fd_sc_hd__nand3_1_52/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1114/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1125 sky130_fd_sc_hd__clkinv_4_35/A sky130_fd_sc_hd__buf_6_89/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1125/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_330 VDD VSS sky130_fd_sc_hd__a22o_1_30/B2 sky130_fd_sc_hd__clkinv_4_27/Y
+ sky130_fd_sc_hd__o21ai_1_22/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_341 VDD VSS sky130_fd_sc_hd__ha_2_157/A sky130_fd_sc_hd__dfxtp_1_347/CLK
+ sky130_fd_sc_hd__o21ai_1_31/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_352 VDD VSS sky130_fd_sc_hd__a22o_1_19/B2 sky130_fd_sc_hd__dfxtp_1_354/CLK
+ sky130_fd_sc_hd__ha_2_151/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_363 VDD VSS sky130_fd_sc_hd__fa_2_1107/A sky130_fd_sc_hd__dfxtp_1_380/CLK
+ sky130_fd_sc_hd__and2_0_176/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_374 VDD VSS sky130_fd_sc_hd__fa_2_1118/A sky130_fd_sc_hd__clkinv_4_32/Y
+ sky130_fd_sc_hd__and2_0_119/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_385 VDD VSS sky130_fd_sc_hd__fa_2_1113/B sky130_fd_sc_hd__clkinv_4_32/Y
+ sky130_fd_sc_hd__and2_0_140/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_5 sky130_fd_sc_hd__nand3_1_5/C sky130_fd_sc_hd__nand2_1_5/B
+ sky130_fd_sc_hd__nand2_1_9/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_396 VDD VSS sky130_fd_sc_hd__nor2_1_56/A sky130_fd_sc_hd__dfxtp_1_411/CLK
+ sky130_fd_sc_hd__and2_0_231/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_202 sky130_fd_sc_hd__fa_2_205/B sky130_fd_sc_hd__fa_2_202/SUM
+ sky130_fd_sc_hd__fa_2_202/A sky130_fd_sc_hd__fa_2_202/B sky130_fd_sc_hd__fa_2_202/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_213 sky130_fd_sc_hd__fa_2_214/B sky130_fd_sc_hd__fa_2_206/A
+ sky130_fd_sc_hd__ha_2_107/A sky130_fd_sc_hd__fa_2_31/A sky130_fd_sc_hd__fa_2_281/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_224 sky130_fd_sc_hd__fa_2_225/B sky130_fd_sc_hd__fa_2_216/A
+ sky130_fd_sc_hd__fa_2_5/B sky130_fd_sc_hd__fa_2_32/A sky130_fd_sc_hd__fa_2_209/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_235 sky130_fd_sc_hd__fa_2_237/CIN sky130_fd_sc_hd__fa_2_231/A
+ sky130_fd_sc_hd__fa_2_235/A sky130_fd_sc_hd__fa_2_235/B sky130_fd_sc_hd__fa_2_235/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_246 sky130_fd_sc_hd__fa_2_251/B sky130_fd_sc_hd__fa_2_246/SUM
+ sky130_fd_sc_hd__fa_2_246/A sky130_fd_sc_hd__fa_2_246/B sky130_fd_sc_hd__fa_2_246/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_257 sky130_fd_sc_hd__fa_2_258/CIN sky130_fd_sc_hd__fa_2_252/B
+ sky130_fd_sc_hd__fa_2_2/A sky130_fd_sc_hd__fa_2_266/B sky130_fd_sc_hd__fa_2_283/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_268 sky130_fd_sc_hd__fa_2_171/A sky130_fd_sc_hd__fa_2_170/B
+ sky130_fd_sc_hd__fa_2_268/A sky130_fd_sc_hd__fa_2_268/B sky130_fd_sc_hd__fa_2_272/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_279 sky130_fd_sc_hd__fa_2_278/B sky130_fd_sc_hd__fa_2_279/SUM
+ sky130_fd_sc_hd__fa_2_279/A sky130_fd_sc_hd__fa_2_279/B sky130_fd_sc_hd__fa_2_279/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_6 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_6/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_1/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__diode_2_107 sky130_fd_sc_hd__inv_2_135/Y VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_118 sky130_fd_sc_hd__buf_2_225/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__fa_2_60 sky130_fd_sc_hd__fa_2_63/B sky130_fd_sc_hd__fa_2_60/SUM
+ sky130_fd_sc_hd__fa_2_60/A sky130_fd_sc_hd__fa_2_60/B sky130_fd_sc_hd__fa_2_60/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_71 sky130_fd_sc_hd__fa_2_72/B sky130_fd_sc_hd__fa_2_64/A sky130_fd_sc_hd__fa_2_71/A
+ sky130_fd_sc_hd__ha_2_94/B sky130_fd_sc_hd__fa_2_139/B VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__diode_2_129 sky130_fd_sc_hd__buf_2_250/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__fa_2_82 sky130_fd_sc_hd__fa_2_83/B sky130_fd_sc_hd__fa_2_74/A sky130_fd_sc_hd__fa_2_82/A
+ sky130_fd_sc_hd__ha_2_95/A sky130_fd_sc_hd__fa_2_67/B VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_93 sky130_fd_sc_hd__fa_2_95/CIN sky130_fd_sc_hd__fa_2_89/A
+ sky130_fd_sc_hd__fa_2_93/A sky130_fd_sc_hd__fa_2_93/B sky130_fd_sc_hd__fa_2_93/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_230 VDD VSS sky130_fd_sc_hd__buf_2_230/X sky130_fd_sc_hd__buf_2_230/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_241 VDD VSS sky130_fd_sc_hd__buf_8_214/A sky130_fd_sc_hd__buf_6_59/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_252 VDD VSS sky130_fd_sc_hd__nor2_1_29/A sky130_fd_sc_hd__buf_2_252/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_263 VDD VSS sky130_fd_sc_hd__buf_2_263/X sky130_fd_sc_hd__buf_2_263/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_274 VDD VSS sky130_fd_sc_hd__buf_2_274/X sky130_fd_sc_hd__buf_2_274/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_285 VDD VSS sky130_fd_sc_hd__buf_2_285/X sky130_fd_sc_hd__buf_2_285/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1270 VDD VSS sky130_fd_sc_hd__mux2_2_219/A0 sky130_fd_sc_hd__clkinv_8_63/Y
+ sky130_fd_sc_hd__dfxtp_1_426/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1281 VDD VSS sky130_fd_sc_hd__mux2_2_196/A0 sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__dfxtp_1_437/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1292 VDD VSS sky130_fd_sc_hd__mux2_2_189/A0 sky130_fd_sc_hd__clkinv_8_75/Y
+ sky130_fd_sc_hd__o22ai_1_343/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a21oi_1_10 sky130_fd_sc_hd__a21oi_1_11/Y sky130_fd_sc_hd__nor2_1_11/Y
+ sky130_fd_sc_hd__nor2_1_10/B sky130_fd_sc_hd__nand2_1_48/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_21 sky130_fd_sc_hd__nor2_1_36/B sky130_fd_sc_hd__nor3_1_34/Y
+ sky130_fd_sc_hd__a21oi_1_21/Y sky130_fd_sc_hd__nor2_1_36/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_32 sky130_fd_sc_hd__nor2_1_41/Y sky130_fd_sc_hd__o22ai_1_65/Y
+ sky130_fd_sc_hd__a21oi_1_32/Y sky130_fd_sc_hd__fa_2_1035/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_43 sky130_fd_sc_hd__nor2_2_6/Y sky130_fd_sc_hd__o22ai_1_75/Y
+ sky130_fd_sc_hd__a21oi_1_43/Y sky130_fd_sc_hd__fa_2_1031/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_207 sky130_fd_sc_hd__buf_12_207/A sky130_fd_sc_hd__buf_12_230/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_54 sky130_fd_sc_hd__nor2_2_6/Y sky130_fd_sc_hd__o22ai_1_86/Y
+ sky130_fd_sc_hd__a21oi_1_54/Y sky130_fd_sc_hd__fa_2_1042/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_218 sky130_fd_sc_hd__buf_6_26/X sky130_fd_sc_hd__buf_12_245/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_65 sky130_fd_sc_hd__a21oi_1_65/A1 sky130_fd_sc_hd__nor2_1_42/B
+ sky130_fd_sc_hd__xnor2_1_36/A sky130_fd_sc_hd__xnor2_1_34/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_229 sky130_fd_sc_hd__buf_12_229/A sky130_fd_sc_hd__buf_12_229/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_76 sky130_fd_sc_hd__o21a_1_5/B1 sky130_fd_sc_hd__o21a_1_4/A1
+ sky130_fd_sc_hd__a21oi_1_76/Y sky130_fd_sc_hd__nor2_1_66/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_87 sky130_fd_sc_hd__nand2_1_262/A sky130_fd_sc_hd__o21ai_1_102/Y
+ sky130_fd_sc_hd__a21oi_1_87/Y sky130_fd_sc_hd__a211o_1_3/A1 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_98 sky130_fd_sc_hd__fa_2_978/A sky130_fd_sc_hd__o22ai_1_100/Y
+ sky130_fd_sc_hd__a21oi_1_98/Y sky130_fd_sc_hd__nor2_2_7/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__fa_2_780 sky130_fd_sc_hd__fa_2_783/B sky130_fd_sc_hd__fa_2_780/SUM
+ sky130_fd_sc_hd__fa_2_780/A sky130_fd_sc_hd__fa_2_780/B sky130_fd_sc_hd__fa_2_785/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_791 sky130_fd_sc_hd__fa_2_794/B sky130_fd_sc_hd__fa_2_791/SUM
+ sky130_fd_sc_hd__fa_2_791/A sky130_fd_sc_hd__fa_2_791/B sky130_fd_sc_hd__o22ai_1_54/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor3_1_2 sky130_fd_sc_hd__nor3_1_2/C sky130_fd_sc_hd__nor3_1_2/Y
+ sky130_fd_sc_hd__nor3_2_1/A sky130_fd_sc_hd__or2_0_0/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__clkinv_1_407 sky130_fd_sc_hd__nand2_1_215/B sky130_fd_sc_hd__nor4_1_8/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_407/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_418 sky130_fd_sc_hd__o21ai_1_36/A2 sky130_fd_sc_hd__fa_2_948/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_418/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_429 sky130_fd_sc_hd__o22ai_1_59/A2 sky130_fd_sc_hd__dfxtp_1_493/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_429/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_6_50 VDD VSS sky130_fd_sc_hd__buf_6_50/X sky130_fd_sc_hd__buf_6_50/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_61 VDD VSS sky130_fd_sc_hd__buf_6_61/X sky130_fd_sc_hd__buf_6_61/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_72 VDD VSS sky130_fd_sc_hd__buf_6_72/X sky130_fd_sc_hd__buf_6_72/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_83 VDD VSS sky130_fd_sc_hd__buf_6_83/X sky130_fd_sc_hd__buf_6_83/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__a21oi_1_304 sky130_fd_sc_hd__o21a_1_34/B1 sky130_fd_sc_hd__o21a_1_33/A1
+ sky130_fd_sc_hd__a21oi_1_304/Y sky130_fd_sc_hd__nor2_1_187/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_30 sky130_fd_sc_hd__buf_2_77/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_315 sky130_fd_sc_hd__nor2_1_198/A sky130_fd_sc_hd__o21a_1_41/A1
+ sky130_fd_sc_hd__a21oi_1_315/Y sky130_fd_sc_hd__nor2_1_198/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_41 sky130_fd_sc_hd__buf_2_104/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_326 sky130_fd_sc_hd__fa_2_1181/A sky130_fd_sc_hd__o22ai_1_299/Y
+ sky130_fd_sc_hd__a21oi_1_326/Y sky130_fd_sc_hd__nor3_1_39/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_52 sky130_fd_sc_hd__buf_2_109/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_337 sky130_fd_sc_hd__fa_2_1184/A sky130_fd_sc_hd__o22ai_1_304/Y
+ sky130_fd_sc_hd__a21oi_1_337/Y sky130_fd_sc_hd__nor2_2_16/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_63 sky130_fd_sc_hd__buf_2_110/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_348 sky130_fd_sc_hd__nor2_1_224/Y sky130_fd_sc_hd__nor2_1_219/Y
+ sky130_fd_sc_hd__a21oi_1_348/Y sky130_fd_sc_hd__fa_2_1199/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_74 sky130_fd_sc_hd__clkbuf_4_83/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_359 sky130_fd_sc_hd__fa_2_1201/A sky130_fd_sc_hd__o22ai_1_322/Y
+ sky130_fd_sc_hd__o21a_1_42/B1 sky130_fd_sc_hd__nor2_2_16/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_85 sky130_fd_sc_hd__nand4_1_45/B VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_96 sky130_fd_sc_hd__clkbuf_4_208/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a222oi_1_7 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1126/A sky130_fd_sc_hd__nor2_2_15/Y
+ sky130_fd_sc_hd__nor3_1_38/A sky130_fd_sc_hd__fa_2_1128/A sky130_fd_sc_hd__nor3_1_38/B
+ sky130_fd_sc_hd__a222oi_1_7/Y sky130_fd_sc_hd__fa_2_1125/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__o221ai_1_1 sky130_fd_sc_hd__o221ai_1_1/A2 sky130_fd_sc_hd__o221ai_1_1/Y
+ sky130_fd_sc_hd__a21oi_1_26/Y sky130_fd_sc_hd__nand3_1_48/Y sky130_fd_sc_hd__fa_2_959/A
+ sky130_fd_sc_hd__o21ai_1_37/Y VDD VSS VSS VDD sky130_fd_sc_hd__o221ai_1
Xsky130_fd_sc_hd__nand2_1_320 sky130_fd_sc_hd__nand2_1_320/Y sky130_fd_sc_hd__nand2_1_339/B
+ sky130_fd_sc_hd__xor2_1_87/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_331 sky130_fd_sc_hd__nand2_1_331/Y sky130_fd_sc_hd__nand2_1_331/B
+ sky130_fd_sc_hd__o21ai_1_254/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_930 sky130_fd_sc_hd__o32ai_1_5/B2 sky130_fd_sc_hd__o32ai_1_5/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_930/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_342 sky130_fd_sc_hd__xnor2_1_91/B sky130_fd_sc_hd__fa_2_1138/A
+ sky130_fd_sc_hd__o21a_1_17/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_941 sky130_fd_sc_hd__nor2_2_16/B sky130_fd_sc_hd__nor2_4_16/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_941/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_353 sky130_fd_sc_hd__o21a_1_27/B1 sky130_fd_sc_hd__fa_2_1148/A
+ sky130_fd_sc_hd__o21a_1_27/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_952 sky130_fd_sc_hd__nor2_1_257/A sky130_fd_sc_hd__nor2b_1_119/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_952/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_364 sky130_fd_sc_hd__nand2_1_364/Y sky130_fd_sc_hd__mux2_2_92/A0
+ sky130_fd_sc_hd__nor2_4_15/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_963 sky130_fd_sc_hd__o31ai_1_10/B1 sky130_fd_sc_hd__a21oi_1_382/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_963/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_375 sky130_fd_sc_hd__nand2_1_375/Y sky130_fd_sc_hd__nand2_1_387/B
+ sky130_fd_sc_hd__o21ai_1_305/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_974 sky130_fd_sc_hd__o32ai_1_7/B2 sky130_fd_sc_hd__fa_2_1244/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_974/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_386 sky130_fd_sc_hd__nand2_1_386/Y sky130_fd_sc_hd__nor2b_1_104/A
+ sky130_fd_sc_hd__xor2_1_163/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_985 sky130_fd_sc_hd__nand2_1_476/B sky130_fd_sc_hd__fa_2_164/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_985/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_397 sky130_fd_sc_hd__o21a_1_33/B1 sky130_fd_sc_hd__fa_2_1183/A
+ sky130_fd_sc_hd__o21a_1_33/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_996 sky130_fd_sc_hd__nor2_1_228/B sky130_fd_sc_hd__fa_2_1237/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_996/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_160 VDD VSS sky130_fd_sc_hd__ha_2_49/A sky130_fd_sc_hd__dfxtp_1_170/CLK
+ sky130_fd_sc_hd__nor2b_1_19/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_171 VDD VSS sky130_fd_sc_hd__nor3_2_4/A sky130_fd_sc_hd__clkinv_4_9/Y
+ sky130_fd_sc_hd__ha_2_49/B VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_182 VDD VSS sky130_fd_sc_hd__ha_2_52/A sky130_fd_sc_hd__dfxtp_1_182/CLK
+ sky130_fd_sc_hd__and2_0_51/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_193 VDD VSS sky130_fd_sc_hd__ha_2_63/A sky130_fd_sc_hd__dfxtp_1_195/CLK
+ sky130_fd_sc_hd__nor2b_1_28/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__buf_2_19 VDD VSS sky130_fd_sc_hd__buf_8_23/A sky130_fd_sc_hd__ha_2_22/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__a21boi_1_3 sky130_fd_sc_hd__a21boi_1_3/Y sky130_fd_sc_hd__nor2_2_16/Y
+ sky130_fd_sc_hd__a21oi_1_328/Y sky130_fd_sc_hd__fa_2_1186/A VDD VSS VDD VSS sky130_fd_sc_hd__a21boi_1
Xsky130_fd_sc_hd__o211ai_1_13 sky130_fd_sc_hd__o21a_1_8/X sky130_fd_sc_hd__nor2_1_77/A
+ sky130_fd_sc_hd__xor2_1_41/A sky130_fd_sc_hd__nand2_1_276/Y sky130_fd_sc_hd__nand2_1_277/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_24 sky130_fd_sc_hd__nor2_1_180/A sky130_fd_sc_hd__nor2_1_172/B
+ sky130_fd_sc_hd__xor2_1_171/A sky130_fd_sc_hd__nand2_1_374/Y sky130_fd_sc_hd__nand2_1_376/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_35 sky130_fd_sc_hd__a21oi_1_294/Y sky130_fd_sc_hd__nor2_1_180/A
+ sky130_fd_sc_hd__xor2_1_158/A sky130_fd_sc_hd__a21oi_1_291/Y sky130_fd_sc_hd__nand2_1_389/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_46 sky130_fd_sc_hd__nor2_1_224/A sky130_fd_sc_hd__a21oi_1_354/Y
+ sky130_fd_sc_hd__xor2_1_199/A sky130_fd_sc_hd__nand2_1_440/Y sky130_fd_sc_hd__a21oi_1_346/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_57 sky130_fd_sc_hd__nor2_1_257/A sky130_fd_sc_hd__a222oi_1_30/Y
+ sky130_fd_sc_hd__xor2_1_243/A sky130_fd_sc_hd__nand2_1_491/Y sky130_fd_sc_hd__a21oi_1_404/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__fa_2_1270 sky130_fd_sc_hd__fa_2_1271/CIN sky130_fd_sc_hd__mux2_2_199/A1
+ sky130_fd_sc_hd__fa_2_1270/A sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1270/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o211ai_1_68 sky130_fd_sc_hd__nor2_1_307/A sky130_fd_sc_hd__a211oi_1_37/Y
+ sky130_fd_sc_hd__xor2_1_286/A sky130_fd_sc_hd__nand2_1_541/Y sky130_fd_sc_hd__nand2_1_542/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__fa_2_1281 sky130_fd_sc_hd__fa_2_1282/CIN sky130_fd_sc_hd__mux2_2_249/A1
+ sky130_fd_sc_hd__fa_2_1281/A sky130_fd_sc_hd__fa_2_1281/B sky130_fd_sc_hd__fa_2_1281/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1292 sky130_fd_sc_hd__xor2_1_276/B sky130_fd_sc_hd__mux2_2_223/A0
+ sky130_fd_sc_hd__fa_2_1292/A sky130_fd_sc_hd__fa_2_1292/B sky130_fd_sc_hd__fa_2_1292/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_1_204 sky130_fd_sc_hd__buf_8_200/A sky130_fd_sc_hd__clkinv_1_204/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_204/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_215 sky130_fd_sc_hd__clkinv_2_29/A sky130_fd_sc_hd__a22oi_1_265/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_215/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_226 sky130_fd_sc_hd__inv_2_118/A sky130_fd_sc_hd__buf_8_199/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_226/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_237 sky130_fd_sc_hd__clkinv_1_238/A sky130_fd_sc_hd__buf_8_214/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_237/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_248 sky130_fd_sc_hd__clkinv_1_248/Y sky130_fd_sc_hd__clkinv_1_248/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_248/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_259 sky130_fd_sc_hd__nor2_1_9/B sky130_fd_sc_hd__nand2_1_33/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_259/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_101 sky130_fd_sc_hd__fa_2_976/A sky130_fd_sc_hd__o22ai_1_106/Y
+ sky130_fd_sc_hd__a21oi_1_101/Y sky130_fd_sc_hd__nor2_4_10/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_112 sky130_fd_sc_hd__clkinv_1_569/Y sky130_fd_sc_hd__o22ai_1_122/Y
+ sky130_fd_sc_hd__a21oi_1_112/Y sky130_fd_sc_hd__a211o_1_6/A1 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_123 sky130_fd_sc_hd__a21o_2_3/A2 sky130_fd_sc_hd__o21ai_1_147/Y
+ sky130_fd_sc_hd__a21oi_1_123/Y sky130_fd_sc_hd__fa_2_998/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_134 sky130_fd_sc_hd__a21o_2_3/A2 sky130_fd_sc_hd__o21ai_1_157/Y
+ sky130_fd_sc_hd__a21oi_1_134/Y sky130_fd_sc_hd__fa_2_1003/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_145 sky130_fd_sc_hd__nor2_2_10/Y sky130_fd_sc_hd__o22ai_1_145/Y
+ sky130_fd_sc_hd__a21oi_1_145/Y sky130_fd_sc_hd__fa_2_1117/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_156 sky130_fd_sc_hd__nor2_2_11/Y sky130_fd_sc_hd__o22ai_1_155/Y
+ sky130_fd_sc_hd__a21oi_1_156/Y sky130_fd_sc_hd__fa_2_1113/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nor2_1_320 sky130_fd_sc_hd__nor2_1_322/A sky130_fd_sc_hd__nor2_1_320/Y
+ sky130_fd_sc_hd__nor2_1_320/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a21oi_1_167 sky130_fd_sc_hd__clkinv_1_671/Y sky130_fd_sc_hd__nor2_1_97/B
+ sky130_fd_sc_hd__xnor2_1_85/A sky130_fd_sc_hd__xnor2_1_83/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_178 sky130_fd_sc_hd__nand2_1_302/Y sky130_fd_sc_hd__nor2_1_93/A
+ sky130_fd_sc_hd__xnor2_1_68/A sky130_fd_sc_hd__xnor2_1_66/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_189 sky130_fd_sc_hd__a21o_2_5/A2 sky130_fd_sc_hd__o21ai_1_209/Y
+ sky130_fd_sc_hd__a21oi_1_189/Y sky130_fd_sc_hd__fa_2_1073/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_108 sky130_fd_sc_hd__buf_8_91/A sky130_fd_sc_hd__buf_8_113/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_119 sky130_fd_sc_hd__buf_8_119/A sky130_fd_sc_hd__buf_6_39/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nand2_1_150 sky130_fd_sc_hd__fa_2_39/CIN sky130_fd_sc_hd__fa_2_139/B
+ sky130_fd_sc_hd__fa_2_76/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_161 sky130_fd_sc_hd__fa_2_219/A sky130_fd_sc_hd__fa_2_281/A
+ sky130_fd_sc_hd__fa_2_277/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_760 sky130_fd_sc_hd__ha_2_192/B sky130_fd_sc_hd__fa_2_1115/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_760/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_172 sky130_fd_sc_hd__fa_2_390/A sky130_fd_sc_hd__fa_2_409/A
+ sky130_fd_sc_hd__fa_2_412/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_771 sky130_fd_sc_hd__o22ai_1_206/A1 sky130_fd_sc_hd__nor2_2_12/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_771/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_183 sky130_fd_sc_hd__fa_2_559/CIN sky130_fd_sc_hd__fa_2_531/B
+ sky130_fd_sc_hd__ha_2_117/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_782 sky130_fd_sc_hd__or2_0_9/B sky130_fd_sc_hd__nor2_1_183/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_782/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_194 sky130_fd_sc_hd__fa_2_755/B sky130_fd_sc_hd__ha_2_140/A
+ sky130_fd_sc_hd__ha_2_142/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_793 sky130_fd_sc_hd__nor2_1_154/A sky130_fd_sc_hd__nor2_1_155/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_793/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand3_2_0 sky130_fd_sc_hd__nor2_4_3/Y sky130_fd_sc_hd__nand3_2_0/Y
+ sky130_fd_sc_hd__nand3_2_0/B sky130_fd_sc_hd__nand3_2_0/C VSS VDD VSS VDD sky130_fd_sc_hd__nand3_2
Xsky130_fd_sc_hd__xor2_1_14 sky130_fd_sc_hd__xor2_1_14/B sky130_fd_sc_hd__xor2_1_14/X
+ sky130_fd_sc_hd__xor2_1_14/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_25 sky130_fd_sc_hd__xor2_1_25/B sky130_fd_sc_hd__xor2_1_25/X
+ sky130_fd_sc_hd__xor2_1_25/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_36 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_991/B
+ sky130_fd_sc_hd__xor2_1_36/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_47 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_980/B
+ sky130_fd_sc_hd__xor2_1_47/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_58 sky130_fd_sc_hd__xor2_1_58/B sky130_fd_sc_hd__xor2_1_58/X
+ sky130_fd_sc_hd__xor2_1_59/X VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_69 sky130_fd_sc_hd__nor2_4_9/Y sky130_fd_sc_hd__xor2_1_69/X
+ sky130_fd_sc_hd__xor2_1_69/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2b_1_8 sky130_fd_sc_hd__nand2b_1_8/Y sky130_fd_sc_hd__fa_2_957/A
+ sky130_fd_sc_hd__nor2b_1_89/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a21o_2_4 sky130_fd_sc_hd__a21o_2_4/X sky130_fd_sc_hd__a21o_2_4/B1
+ sky130_fd_sc_hd__a21o_2_5/A2 sky130_fd_sc_hd__fa_2_1076/A VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__dfxtp_1_907 VDD VSS sky130_fd_sc_hd__fa_2_942/B sky130_fd_sc_hd__clkinv_4_22/Y
+ sky130_fd_sc_hd__dfxtp_1_907/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_918 VDD VSS sky130_fd_sc_hd__fa_2_1147/A sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__mux2_2_101/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_929 VDD VSS sky130_fd_sc_hd__xor2_1_163/A sky130_fd_sc_hd__clkinv_8_46/Y
+ sky130_fd_sc_hd__mux2_2_76/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_505 VSS VDD sky130_fd_sc_hd__nand4_1_55/D sky130_fd_sc_hd__a22oi_1_231/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_516 VSS VDD sky130_fd_sc_hd__clkbuf_1_516/X sky130_fd_sc_hd__buf_8_209/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_527 VSS VDD sky130_fd_sc_hd__clkbuf_1_527/X sky130_fd_sc_hd__clkbuf_1_527/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_538 VSS VDD sky130_fd_sc_hd__clkbuf_1_538/X sky130_fd_sc_hd__clkbuf_1_538/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_106 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_97/A sky130_fd_sc_hd__fa_2_258/B
+ sky130_fd_sc_hd__ha_2_106/SUM sky130_fd_sc_hd__fa_2_15/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_549 VSS VDD sky130_fd_sc_hd__fa_2_1173/A sky130_fd_sc_hd__nor2_8_0/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_117 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_118/B sky130_fd_sc_hd__fa_2_454/B
+ sky130_fd_sc_hd__fa_2_458/A sky130_fd_sc_hd__ha_2_117/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_128 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_128/A sky130_fd_sc_hd__fa_2_586/B
+ sky130_fd_sc_hd__ha_2_128/SUM sky130_fd_sc_hd__ha_2_131/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_139 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_140/A sky130_fd_sc_hd__fa_2_725/CIN
+ sky130_fd_sc_hd__fa_2_722/A sky130_fd_sc_hd__ha_2_139/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_30 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_30/A sky130_fd_sc_hd__xor2_1_3/A
+ sky130_fd_sc_hd__ha_2_30/SUM sky130_fd_sc_hd__ha_2_30/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_41 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_41/A sky130_fd_sc_hd__ha_2_40/B
+ sky130_fd_sc_hd__ha_2_41/SUM sky130_fd_sc_hd__ha_2_41/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_52 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_52/A sky130_fd_sc_hd__ha_2_51/B
+ sky130_fd_sc_hd__ha_2_52/SUM sky130_fd_sc_hd__ha_2_52/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_63 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_63/A sky130_fd_sc_hd__ha_2_62/B
+ sky130_fd_sc_hd__ha_2_63/SUM sky130_fd_sc_hd__ha_2_63/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_74 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_74/A sky130_fd_sc_hd__ha_2_73/B
+ sky130_fd_sc_hd__ha_2_74/SUM sky130_fd_sc_hd__ha_2_74/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_85 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_85/A sky130_fd_sc_hd__ha_2_84/B
+ sky130_fd_sc_hd__ha_2_85/SUM sky130_fd_sc_hd__ha_2_85/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_96 VSS VDD VSS VDD sky130_fd_sc_hd__fa_2_2/A sky130_fd_sc_hd__fa_2_112/B
+ sky130_fd_sc_hd__fa_2_108/B sky130_fd_sc_hd__ha_2_96/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_4 VSS VDD sky130_fd_sc_hd__buf_4_2/A sky130_fd_sc_hd__buf_4_1/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__sdlclkp_4_70 sky130_fd_sc_hd__conb_1_23/LO sky130_fd_sc_hd__clkinv_8_40/A
+ sky130_fd_sc_hd__dfxtp_1_626/CLK sky130_fd_sc_hd__or2_0_6/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_81 sky130_fd_sc_hd__conb_1_26/LO sky130_fd_sc_hd__clkinv_8_68/Y
+ sky130_fd_sc_hd__dfxtp_1_1047/CLK sky130_fd_sc_hd__or2_0_10/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_92 sky130_fd_sc_hd__conb_1_29/LO sky130_fd_sc_hd__clkinv_4_33/Y
+ sky130_fd_sc_hd__dfxtp_1_1464/CLK sky130_fd_sc_hd__nand2b_1_18/Y VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_150 sky130_fd_sc_hd__nor2_1_150/B sky130_fd_sc_hd__o21a_1_23/A1
+ sky130_fd_sc_hd__o21a_1_24/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_1_4 sky130_fd_sc_hd__clkinv_1_4/Y sky130_fd_sc_hd__nor2_4_3/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_4/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_161 sky130_fd_sc_hd__nor2_1_161/B sky130_fd_sc_hd__nor2_1_161/Y
+ sky130_fd_sc_hd__nor2_1_163/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_172 sky130_fd_sc_hd__nor2_1_172/B sky130_fd_sc_hd__nor2_1_172/Y
+ sky130_fd_sc_hd__nor2_1_172/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_183 sky130_fd_sc_hd__nor2_1_183/B sky130_fd_sc_hd__nor2_1_183/Y
+ sky130_fd_sc_hd__nor2_1_183/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_194 sky130_fd_sc_hd__o21a_1_42/A2 sky130_fd_sc_hd__o21a_1_38/A1
+ sky130_fd_sc_hd__o21a_1_39/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_70 sky130_fd_sc_hd__nor2_2_2/Y sky130_fd_sc_hd__a22oi_1_82/A1
+ sky130_fd_sc_hd__clkbuf_1_58/X sky130_fd_sc_hd__clkbuf_1_54/X sky130_fd_sc_hd__nand4_1_12/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_81 sky130_fd_sc_hd__a22oi_1_81/B1 sky130_fd_sc_hd__clkbuf_1_99/X
+ sky130_fd_sc_hd__clkbuf_1_35/X sky130_fd_sc_hd__clkbuf_4_10/X sky130_fd_sc_hd__nand4_1_15/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_92 sky130_fd_sc_hd__a22oi_1_96/B1 sky130_fd_sc_hd__a22oi_1_96/A1
+ sky130_fd_sc_hd__a22oi_1_92/B2 sky130_fd_sc_hd__a22oi_1_92/A2 sky130_fd_sc_hd__nand4_1_18/D
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__and2_0_19 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_19/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_19/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__buf_12_390 sky130_fd_sc_hd__buf_8_188/X sky130_fd_sc_hd__buf_12_390/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_260 sky130_fd_sc_hd__clkbuf_1_376/X sky130_fd_sc_hd__nor2_2_5/Y
+ sky130_fd_sc_hd__buf_2_217/X sky130_fd_sc_hd__clkbuf_1_473/X sky130_fd_sc_hd__nand4_1_64/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_271 sky130_fd_sc_hd__nor2_2_4/Y sky130_fd_sc_hd__clkbuf_1_377/X
+ sky130_fd_sc_hd__a22oi_1_271/B2 sky130_fd_sc_hd__clkbuf_4_189/X sky130_fd_sc_hd__nand4_1_67/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_282 sky130_fd_sc_hd__clkbuf_1_378/X sky130_fd_sc_hd__clkbuf_1_379/X
+ sky130_fd_sc_hd__buf_2_222/X sky130_fd_sc_hd__buf_2_196/X sky130_fd_sc_hd__nand4_1_70/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_4_100 VDD VSS sky130_fd_sc_hd__buf_4_100/X sky130_fd_sc_hd__buf_4_100/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__a22oi_1_293 sky130_fd_sc_hd__clkbuf_4_165/X sky130_fd_sc_hd__clkinv_2_23/Y
+ sky130_fd_sc_hd__clkbuf_1_404/X sky130_fd_sc_hd__a22oi_1_293/A2 sky130_fd_sc_hd__a22oi_1_293/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_4_111 VDD VSS sky130_fd_sc_hd__buf_4_111/X sky130_fd_sc_hd__buf_8_209/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_122 VDD VSS sky130_fd_sc_hd__buf_4_122/X sky130_fd_sc_hd__buf_4_122/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_8_18 sky130_fd_sc_hd__inv_2_26/Y sky130_fd_sc_hd__buf_8_18/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_29 sky130_fd_sc_hd__buf_8_29/A sky130_fd_sc_hd__buf_8_29/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__clkinv_1_590 sky130_fd_sc_hd__a22o_1_68/A1 sky130_fd_sc_hd__a22o_1_68/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_590/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_4_70 sky130_fd_sc_hd__clkinv_4_70/A sky130_fd_sc_hd__clkinv_4_71/A
+ VSS VDD VDD VSS VSS sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__inv_16_0/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__o21ai_1_504 VSS VDD sky130_fd_sc_hd__nand2_1_565/A sky130_fd_sc_hd__o21ai_1_507/A1
+ sky130_fd_sc_hd__nand2_1_565/Y sky130_fd_sc_hd__and2_0_353/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_704 VDD VSS sky130_fd_sc_hd__mux2_2_25/A1 sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__o21ai_1_44/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_715 VDD VSS sky130_fd_sc_hd__mux2_2_3/A1 sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__o21ai_1_55/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_726 VDD VSS sky130_fd_sc_hd__mux2_2_20/A1 sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__o21ai_1_63/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_737 VDD VSS sky130_fd_sc_hd__and2_0_163/A sky130_fd_sc_hd__dfxtp_1_747/CLK
+ sky130_fd_sc_hd__fa_2_1092/B VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_748 VDD VSS sky130_fd_sc_hd__and2_0_172/A sky130_fd_sc_hd__dfxtp_1_755/CLK
+ sky130_fd_sc_hd__fa_2_1103/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_759 VDD VSS sky130_fd_sc_hd__fa_2_686/B sky130_fd_sc_hd__dfxtp_1_764/CLK
+ sky130_fd_sc_hd__o21a_1_13/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_302 VSS VDD sky130_fd_sc_hd__nand4_1_43/D sky130_fd_sc_hd__a22oi_1_191/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_313 VSS VDD sky130_fd_sc_hd__nand4_1_32/D sky130_fd_sc_hd__a22oi_1_147/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_324 VSS VDD sky130_fd_sc_hd__buf_8_128/A sky130_fd_sc_hd__and2_1_1/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_335 VSS VDD sky130_fd_sc_hd__buf_8_123/A sky130_fd_sc_hd__and2_1_7/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_346 VSS VDD sky130_fd_sc_hd__buf_8_160/A sky130_fd_sc_hd__inv_2_93/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_357 VSS VDD sky130_fd_sc_hd__inv_16_5/A sky130_fd_sc_hd__inv_2_104/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_368 VSS VDD sky130_fd_sc_hd__buf_4_82/A sky130_fd_sc_hd__buf_4_81/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_379 VSS VDD sky130_fd_sc_hd__clkbuf_1_379/X sky130_fd_sc_hd__nor3_1_23/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_609 sky130_fd_sc_hd__fa_2_608/A sky130_fd_sc_hd__fa_2_609/SUM
+ sky130_fd_sc_hd__fa_2_667/B sky130_fd_sc_hd__ha_2_128/A sky130_fd_sc_hd__ha_2_126/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_50 VDD VSS sky130_fd_sc_hd__fa_2_502/B sky130_fd_sc_hd__dfxtp_1_60/CLK
+ sky130_fd_sc_hd__dfxtp_1_66/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_61 VDD VSS sky130_fd_sc_hd__ha_2_117/B sky130_fd_sc_hd__dfxtp_1_61/CLK
+ sky130_fd_sc_hd__dfxtp_1_77/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_72 VDD VSS sky130_fd_sc_hd__ha_2_96/B sky130_fd_sc_hd__dfxtp_1_77/CLK
+ sky130_fd_sc_hd__buf_2_288/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_83 VDD VSS sky130_fd_sc_hd__dfxtp_1_83/Q sky130_fd_sc_hd__dfxtp_1_83/CLK
+ sky130_fd_sc_hd__inv_2_2/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_94 VDD VSS sky130_fd_sc_hd__ha_2_9/B sky130_fd_sc_hd__dfxtp_1_95/CLK
+ sky130_fd_sc_hd__and2_0_2/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_300 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_300/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_300/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_140 sky130_fd_sc_hd__nand4_1_45/B sky130_fd_sc_hd__a22oi_1_201/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_311 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_311/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_311/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_151 sky130_fd_sc_hd__nand4_1_34/B sky130_fd_sc_hd__a22oi_1_157/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_322 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_322/X sky130_fd_sc_hd__mux2_2_99/S
+ sky130_fd_sc_hd__and2_0_322/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_162 sky130_fd_sc_hd__clkbuf_4_162/X sky130_fd_sc_hd__buf_2_142/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_333 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_333/X sky130_fd_sc_hd__buf_2_263/X
+ sky130_fd_sc_hd__nor3_1_40/C sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_173 sky130_fd_sc_hd__clkbuf_4_173/X sky130_fd_sc_hd__clkbuf_4_173/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_344 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_344/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_344/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_184 sky130_fd_sc_hd__clkbuf_4_184/X sky130_fd_sc_hd__clkbuf_4_184/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_355 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_355/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_355/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_195 sky130_fd_sc_hd__nand4_1_77/D sky130_fd_sc_hd__a22oi_1_309/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__conb_1_8 sky130_fd_sc_hd__conb_1_8/LO sky130_fd_sc_hd__conb_1_8/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__inv_2_100 sky130_fd_sc_hd__inv_2_100/A sky130_fd_sc_hd__inv_2_100/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_111 sky130_fd_sc_hd__inv_2_111/A sky130_fd_sc_hd__inv_2_111/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__or2_0_2 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__or2_0_2/X sky130_fd_sc_hd__or2_0_2/B
+ VSS VDD VSS VDD sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__inv_2_122 sky130_fd_sc_hd__inv_2_122/A sky130_fd_sc_hd__inv_2_122/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_133 sky130_fd_sc_hd__inv_2_133/A sky130_fd_sc_hd__inv_2_133/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__o22ai_1_107 sky130_fd_sc_hd__nand4_1_85/A sky130_fd_sc_hd__o21ai_1_92/A1
+ sky130_fd_sc_hd__o22ai_1_107/Y sky130_fd_sc_hd__o22ai_1_132/B1 sky130_fd_sc_hd__nor2_1_70/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_118 sky130_fd_sc_hd__nand4_1_85/A sky130_fd_sc_hd__o22ai_1_132/B1
+ sky130_fd_sc_hd__o22ai_1_118/Y sky130_fd_sc_hd__o21ai_1_92/A1 sky130_fd_sc_hd__nand4_1_85/C
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_129 sky130_fd_sc_hd__nor2_1_76/A sky130_fd_sc_hd__nor2_2_9/B
+ sky130_fd_sc_hd__o22ai_1_129/Y sky130_fd_sc_hd__a21oi_1_132/Y sky130_fd_sc_hd__a211oi_1_6/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_2_18 sky130_fd_sc_hd__nor2_2_18/B sky130_fd_sc_hd__nor2_2_18/Y
+ sky130_fd_sc_hd__nor2_4_19/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__o211ai_1_8 sky130_fd_sc_hd__nor2_1_81/Y sky130_fd_sc_hd__nor2_1_76/A
+ sky130_fd_sc_hd__xor2_1_81/A sky130_fd_sc_hd__o211ai_1_8/C1 sky130_fd_sc_hd__o211ai_1_8/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__a211o_1_1 VSS VDD VSS VDD sky130_fd_sc_hd__a211o_1_1/X sky130_fd_sc_hd__nand4_1_84/A
+ sky130_fd_sc_hd__o22ai_1_58/Y sky130_fd_sc_hd__o221ai_1_0/Y sky130_fd_sc_hd__a21oi_1_22/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o21ai_1_301 VSS VDD sky130_fd_sc_hd__nor2_1_143/B sky130_fd_sc_hd__o21a_1_29/A1
+ sky130_fd_sc_hd__a21oi_1_274/Y sky130_fd_sc_hd__o21ai_1_301/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_312 VSS VDD sky130_fd_sc_hd__a211oi_1_16/Y sky130_fd_sc_hd__nor2_1_182/A
+ sky130_fd_sc_hd__nand2_1_382/Y sky130_fd_sc_hd__xor2_1_147/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_323 VSS VDD sky130_fd_sc_hd__nor2_1_151/B sky130_fd_sc_hd__o21a_1_29/A1
+ sky130_fd_sc_hd__a21oi_1_293/Y sky130_fd_sc_hd__o21ai_1_323/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_334 VSS VDD sky130_fd_sc_hd__nand2_1_422/B sky130_fd_sc_hd__nor2_1_211/Y
+ sky130_fd_sc_hd__nor2_1_210/B sky130_fd_sc_hd__o21ai_1_334/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_345 VSS VDD sky130_fd_sc_hd__nor2_1_216/B sky130_fd_sc_hd__nor2_1_224/A
+ sky130_fd_sc_hd__nand2_1_425/Y sky130_fd_sc_hd__xor2_1_213/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_50 sky130_fd_sc_hd__o21a_1_50/X sky130_fd_sc_hd__o21a_1_50/A1
+ sky130_fd_sc_hd__o21a_1_50/B1 sky130_fd_sc_hd__fa_2_1256/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_61 sky130_fd_sc_hd__o21a_1_61/X sky130_fd_sc_hd__o21a_1_61/A1
+ sky130_fd_sc_hd__o21a_1_61/B1 sky130_fd_sc_hd__fa_2_1280/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21ai_1_356 VSS VDD sky130_fd_sc_hd__nor2_1_222/A sky130_fd_sc_hd__a21oi_1_338/Y
+ sky130_fd_sc_hd__a211oi_1_19/Y sky130_fd_sc_hd__xor2_1_225/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a211oi_1_17 sky130_fd_sc_hd__nor2b_1_104/Y sky130_fd_sc_hd__o22ai_1_262/Y
+ sky130_fd_sc_hd__nor2_1_183/Y sky130_fd_sc_hd__a211oi_1_17/Y sky130_fd_sc_hd__o21ai_1_329/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_367 VSS VDD sky130_fd_sc_hd__a222oi_1_20/Y sky130_fd_sc_hd__nor2_1_222/A
+ sky130_fd_sc_hd__a21oi_1_341/Y sky130_fd_sc_hd__xor2_1_194/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a211oi_1_28 sky130_fd_sc_hd__nor2_2_17/Y sky130_fd_sc_hd__nor2_1_261/Y
+ sky130_fd_sc_hd__o22ai_1_364/Y sky130_fd_sc_hd__nor2_1_260/B sky130_fd_sc_hd__fa_2_1238/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_378 VSS VDD sky130_fd_sc_hd__nor2_1_222/A sky130_fd_sc_hd__a21oi_1_356/Y
+ sky130_fd_sc_hd__a211oi_1_22/Y sky130_fd_sc_hd__xor2_1_204/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_389 VSS VDD sky130_fd_sc_hd__nand2_1_475/B sky130_fd_sc_hd__nor2_1_255/Y
+ sky130_fd_sc_hd__nor2_1_254/B sky130_fd_sc_hd__o21ai_1_389/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__mux2_2_14 VSS VDD sky130_fd_sc_hd__mux2_2_14/A1 sky130_fd_sc_hd__mux2_2_14/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_14/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_25 VSS VDD sky130_fd_sc_hd__mux2_2_25/A1 sky130_fd_sc_hd__mux2_2_25/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_25/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_36 VSS VDD sky130_fd_sc_hd__mux2_2_36/A1 sky130_fd_sc_hd__mux2_2_36/A0
+ sky130_fd_sc_hd__mux2_2_37/S sky130_fd_sc_hd__mux2_2_36/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_47 VSS VDD sky130_fd_sc_hd__mux2_2_47/A1 sky130_fd_sc_hd__mux2_2_47/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_47/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_58 VSS VDD sky130_fd_sc_hd__mux2_2_58/A1 sky130_fd_sc_hd__mux2_2_58/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_58/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_69 VSS VDD sky130_fd_sc_hd__mux2_2_69/A1 sky130_fd_sc_hd__mux2_2_69/A0
+ sky130_fd_sc_hd__mux2_2_75/S sky130_fd_sc_hd__mux2_2_69/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__xor2_1_150 sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__fa_2_1133/B
+ sky130_fd_sc_hd__xor2_1_150/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_501 VDD VSS sky130_fd_sc_hd__dfxtp_1_501/Q sky130_fd_sc_hd__dfxtp_1_502/CLK
+ sky130_fd_sc_hd__nor2b_1_61/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_161 sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__xor2_1_161/X
+ sky130_fd_sc_hd__xor2_1_161/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_512 VDD VSS sky130_fd_sc_hd__nor4_1_11/C sky130_fd_sc_hd__dfxtp_1_520/CLK
+ sky130_fd_sc_hd__a22o_1_59/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_172 sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__fa_2_1150/B
+ sky130_fd_sc_hd__xor2_1_172/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_523 VDD VSS sky130_fd_sc_hd__fa_2_968/A sky130_fd_sc_hd__dfxtp_1_526/CLK
+ sky130_fd_sc_hd__and2_0_267/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_183 sky130_fd_sc_hd__xor2_1_183/B sky130_fd_sc_hd__xor2_1_183/X
+ sky130_fd_sc_hd__xor2_1_184/X VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_194 sky130_fd_sc_hd__nor2_8_0/Y sky130_fd_sc_hd__fa_2_1185/B
+ sky130_fd_sc_hd__xor2_1_194/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_534 VDD VSS sky130_fd_sc_hd__fa_2_957/A sky130_fd_sc_hd__dfxtp_1_538/CLK
+ sky130_fd_sc_hd__a22o_1_51/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_545 VDD VSS sky130_fd_sc_hd__fa_2_946/A sky130_fd_sc_hd__dfxtp_1_548/CLK
+ sky130_fd_sc_hd__a22o_1_40/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_556 VDD VSS sky130_fd_sc_hd__dfxtp_1_556/Q sky130_fd_sc_hd__dfxtp_1_576/CLK
+ sky130_fd_sc_hd__dfxtp_1_556/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_567 VDD VSS sky130_fd_sc_hd__and2_0_217/A sky130_fd_sc_hd__dfxtp_1_577/CLK
+ sky130_fd_sc_hd__dfxtp_1_568/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_578 VDD VSS sky130_fd_sc_hd__nand2_1_206/A sky130_fd_sc_hd__dfxtp_1_595/CLK
+ sky130_fd_sc_hd__o31ai_1_2/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_589 VDD VSS sky130_fd_sc_hd__nor4_1_6/D sky130_fd_sc_hd__dfxtp_1_594/CLK
+ sky130_fd_sc_hd__and2_0_246/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_110 VSS VDD sky130_fd_sc_hd__buf_8_36/A sky130_fd_sc_hd__buf_8_2/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_121 VSS VDD sky130_fd_sc_hd__buf_8_42/A sky130_fd_sc_hd__buf_12_92/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_132 VSS VDD sky130_fd_sc_hd__buf_12_128/A sky130_fd_sc_hd__buf_2_48/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_143 VSS VDD sky130_fd_sc_hd__clkbuf_1_143/X sky130_fd_sc_hd__clkbuf_1_143/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_154 VSS VDD sky130_fd_sc_hd__a22oi_1_84/B2 sky130_fd_sc_hd__clkbuf_1_154/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_1 VDD VSS sky130_fd_sc_hd__dfxtp_1_1/Q sky130_fd_sc_hd__dfxtp_1_8/CLK
+ sky130_fd_sc_hd__o21ai_1_0/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_165 VSS VDD sky130_fd_sc_hd__clkbuf_1_165/X sky130_fd_sc_hd__clkbuf_1_165/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_176 VSS VDD sky130_fd_sc_hd__nand4_1_30/B sky130_fd_sc_hd__a22oi_1_141/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_187 VSS VDD sky130_fd_sc_hd__nand4_1_18/B sky130_fd_sc_hd__a22oi_1_94/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_198 VSS VDD sky130_fd_sc_hd__clkbuf_1_198/X sky130_fd_sc_hd__buf_2_116/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_406 sky130_fd_sc_hd__maj3_1_58/B sky130_fd_sc_hd__maj3_1_59/A
+ sky130_fd_sc_hd__fa_2_406/A sky130_fd_sc_hd__fa_2_406/B sky130_fd_sc_hd__fa_2_407/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_417 sky130_fd_sc_hd__fa_2_418/A sky130_fd_sc_hd__fa_2_414/A
+ sky130_fd_sc_hd__fa_2_417/A sky130_fd_sc_hd__fa_2_417/B sky130_fd_sc_hd__fa_2_417/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_428 sky130_fd_sc_hd__fa_2_427/CIN sky130_fd_sc_hd__a21o_2_6/A1
+ sky130_fd_sc_hd__fa_2_531/B sky130_fd_sc_hd__fa_2_428/B sky130_fd_sc_hd__fa_2_428/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_439 sky130_fd_sc_hd__fa_2_438/B sky130_fd_sc_hd__fa_2_439/SUM
+ sky130_fd_sc_hd__ha_2_125/A sky130_fd_sc_hd__ha_2_123/B sky130_fd_sc_hd__fa_2_567/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nand3_1_10 sky130_fd_sc_hd__nand3_1_10/Y sky130_fd_sc_hd__nand3_1_10/A
+ sky130_fd_sc_hd__nand3_1_10/C sky130_fd_sc_hd__nand3_1_10/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_21 sky130_fd_sc_hd__buf_2_23/A sky130_fd_sc_hd__nand3_2_2/A
+ sky130_fd_sc_hd__nand3_1_25/B sky130_fd_sc_hd__xor2_1_1/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_32 sky130_fd_sc_hd__nand3_1_32/Y sky130_fd_sc_hd__nor2_4_2/Y
+ sky130_fd_sc_hd__nand3_2_3/B sky130_fd_sc_hd__and2_0_37/X VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_43 sky130_fd_sc_hd__nand3_1_43/Y sky130_fd_sc_hd__nor3_1_27/A
+ sky130_fd_sc_hd__inv_8_1/Y sky130_fd_sc_hd__nor3_1_26/A VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__dfxtp_1_1430 VDD VSS sky130_fd_sc_hd__mux2_2_245/A0 sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__o22ai_1_403/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1441 VDD VSS sky130_fd_sc_hd__mux2_2_220/A1 sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__a221oi_1_5/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1452 VDD VSS sky130_fd_sc_hd__buf_6_85/A sky130_fd_sc_hd__dfxtp_1_1464/CLK
+ sky130_fd_sc_hd__and2_0_353/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1463 VDD VSS sky130_fd_sc_hd__dfxtp_1_1463/Q sky130_fd_sc_hd__dfxtp_1_1464/CLK
+ sky130_fd_sc_hd__and2_0_344/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_130 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_130/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_921/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_141 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_141/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__fa_2_870/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_152 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_152/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_897/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_60 sky130_fd_sc_hd__and2_0_34/A sky130_fd_sc_hd__ha_2_39/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_60/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_163 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_163/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_163/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_71 sky130_fd_sc_hd__buf_2_116/A sky130_fd_sc_hd__clkinv_1_71/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_71/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_174 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_174/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_174/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_82 sky130_fd_sc_hd__inv_2_68/A sky130_fd_sc_hd__inv_2_54/Y
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_185 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_185/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__fa_2_930/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_93 sky130_fd_sc_hd__inv_2_57/A sky130_fd_sc_hd__buf_2_48/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_93/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_196 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_196/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__ha_2_162/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__fa_2_940 sky130_fd_sc_hd__fa_2_918/A sky130_fd_sc_hd__fa_2_919/B
+ sky130_fd_sc_hd__fa_2_940/A sky130_fd_sc_hd__fa_2_940/B sky130_fd_sc_hd__ha_2_125/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_951 sky130_fd_sc_hd__fa_2_950/CIN sky130_fd_sc_hd__fa_2_951/SUM
+ sky130_fd_sc_hd__fa_2_951/A sky130_fd_sc_hd__fa_2_951/B sky130_fd_sc_hd__fa_2_951/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_962 sky130_fd_sc_hd__fa_2_961/CIN sky130_fd_sc_hd__fa_2_962/SUM
+ sky130_fd_sc_hd__fa_2_962/A sky130_fd_sc_hd__fa_2_962/B sky130_fd_sc_hd__fa_2_962/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_973 sky130_fd_sc_hd__fa_2_974/CIN sky130_fd_sc_hd__fa_2_973/SUM
+ sky130_fd_sc_hd__fa_2_973/A sky130_fd_sc_hd__fa_2_973/B sky130_fd_sc_hd__fa_2_973/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_984 sky130_fd_sc_hd__fa_2_985/CIN sky130_fd_sc_hd__mux2_2_19/A0
+ sky130_fd_sc_hd__fa_2_984/A sky130_fd_sc_hd__fa_2_984/B sky130_fd_sc_hd__fa_2_984/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_995 sky130_fd_sc_hd__fa_2_996/CIN sky130_fd_sc_hd__fa_2_995/SUM
+ sky130_fd_sc_hd__fa_2_995/A sky130_fd_sc_hd__fa_2_995/B sky130_fd_sc_hd__fa_2_995/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_1_2 sky130_fd_sc_hd__conb_1_17/LO sky130_fd_sc_hd__clkinv_4_48/A
+ sky130_fd_sc_hd__clkinv_2_38/A sky130_fd_sc_hd__nor2_1_14/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_1
Xsky130_fd_sc_hd__mux2_2_240 VSS VDD sky130_fd_sc_hd__mux2_2_240/A1 sky130_fd_sc_hd__mux2_2_240/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_240/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_251 VSS VDD sky130_fd_sc_hd__mux2_2_251/A1 sky130_fd_sc_hd__mux2_2_251/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_251/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_262 VSS VDD sky130_fd_sc_hd__mux2_2_262/A1 sky130_fd_sc_hd__mux2_2_262/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_262/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__o21ai_1_120 VSS VDD sky130_fd_sc_hd__o22ai_1_130/B1 sky130_fd_sc_hd__nand4_1_85/D
+ sky130_fd_sc_hd__a21oi_1_105/Y sky130_fd_sc_hd__o21ai_1_120/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_131 VSS VDD sky130_fd_sc_hd__a211oi_1_6/Y sky130_fd_sc_hd__nor2_1_77/A
+ sky130_fd_sc_hd__a21oi_1_110/Y sky130_fd_sc_hd__xor2_1_45/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_142 VSS VDD sky130_fd_sc_hd__a21oi_1_124/Y sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__a21oi_1_118/Y sky130_fd_sc_hd__xor2_1_50/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_153 VSS VDD sky130_fd_sc_hd__o21ai_1_153/A2 sky130_fd_sc_hd__o21ai_1_92/A1
+ sky130_fd_sc_hd__a22oi_1_343/Y sky130_fd_sc_hd__o21ai_1_153/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_164 VSS VDD sky130_fd_sc_hd__o21ai_1_171/A2 sky130_fd_sc_hd__xnor2_1_75/Y
+ sky130_fd_sc_hd__a21oi_1_141/Y sky130_fd_sc_hd__o21ai_1_164/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_175 VSS VDD sky130_fd_sc_hd__nand2_2_5/Y sky130_fd_sc_hd__xnor2_1_63/Y
+ sky130_fd_sc_hd__a21oi_1_150/Y sky130_fd_sc_hd__o21ai_1_175/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_186 VSS VDD sky130_fd_sc_hd__nand2_2_5/Y sky130_fd_sc_hd__xnor2_1_85/Y
+ sky130_fd_sc_hd__a21oi_1_161/Y sky130_fd_sc_hd__o21ai_1_186/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_197 VSS VDD sky130_fd_sc_hd__xnor2_1_69/A sky130_fd_sc_hd__o21ai_1_197/A1
+ sky130_fd_sc_hd__nand2_1_288/B sky130_fd_sc_hd__xnor2_1_71/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__maj3_1_70 sky130_fd_sc_hd__maj3_1_71/X sky130_fd_sc_hd__maj3_1_70/X
+ sky130_fd_sc_hd__maj3_1_70/B sky130_fd_sc_hd__maj3_1_70/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_502 sky130_fd_sc_hd__o21a_1_60/B1 sky130_fd_sc_hd__fa_2_1283/A
+ sky130_fd_sc_hd__o21a_1_60/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_513 sky130_fd_sc_hd__nand2_1_513/Y sky130_fd_sc_hd__nor2_1_286/A
+ sky130_fd_sc_hd__xor2_1_275/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_81 sky130_fd_sc_hd__maj3_1_81/C sky130_fd_sc_hd__maj3_1_81/X
+ sky130_fd_sc_hd__maj3_1_81/B sky130_fd_sc_hd__maj3_1_81/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_524 sky130_fd_sc_hd__nor2_1_293/B sky130_fd_sc_hd__nand2_1_524/B
+ sky130_fd_sc_hd__nor2_1_294/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_92 sky130_fd_sc_hd__maj3_1_93/X sky130_fd_sc_hd__maj3_1_92/X
+ sky130_fd_sc_hd__maj3_1_92/B sky130_fd_sc_hd__maj3_1_92/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_535 sky130_fd_sc_hd__nand2_1_535/Y sky130_fd_sc_hd__nor2b_2_5/Y
+ sky130_fd_sc_hd__o21ai_1_463/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_546 sky130_fd_sc_hd__o21a_1_68/A1 sky130_fd_sc_hd__nor2_2_18/B
+ sky130_fd_sc_hd__nor2_4_19/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_557 sky130_fd_sc_hd__nand2_1_557/Y sky130_fd_sc_hd__inv_8_0/Y
+ sky130_fd_sc_hd__nand2_1_557/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_568 sky130_fd_sc_hd__nand2_1_568/Y sky130_fd_sc_hd__nand2_1_568/B
+ sky130_fd_sc_hd__nand2_1_568/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_4 sky130_fd_sc_hd__ha_2_25/SUM sky130_fd_sc_hd__nor2b_1_4/Y
+ sky130_fd_sc_hd__or2_0_1/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1104 sky130_fd_sc_hd__o22ai_1_435/A1 sky130_fd_sc_hd__fa_2_1301/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1104/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1115 sky130_fd_sc_hd__nor4_1_13/C sky130_fd_sc_hd__nor2_1_315/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1115/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1126 sky130_fd_sc_hd__clkinv_4_36/A sky130_fd_sc_hd__clkbuf_4_227/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1126/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_320 VDD VSS sky130_fd_sc_hd__or4_1_0/D sky130_fd_sc_hd__dfxtp_1_325/CLK
+ sky130_fd_sc_hd__and2_0_196/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_331 VDD VSS sky130_fd_sc_hd__a22o_2_8/B2 sky130_fd_sc_hd__clkinv_4_27/Y
+ sky130_fd_sc_hd__o21ai_1_23/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_342 VDD VSS sky130_fd_sc_hd__a22o_1_26/B2 sky130_fd_sc_hd__dfxtp_1_354/CLK
+ sky130_fd_sc_hd__ha_2_156/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_353 VDD VSS sky130_fd_sc_hd__ha_2_151/A sky130_fd_sc_hd__dfxtp_1_361/CLK
+ sky130_fd_sc_hd__o2bb2ai_1_8/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_364 VDD VSS sky130_fd_sc_hd__fa_2_1108/A sky130_fd_sc_hd__dfxtp_1_380/CLK
+ sky130_fd_sc_hd__and2_0_171/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_375 VDD VSS sky130_fd_sc_hd__fa_2_1119/A sky130_fd_sc_hd__clkinv_4_32/Y
+ sky130_fd_sc_hd__and2_0_113/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_386 VDD VSS sky130_fd_sc_hd__fa_2_1114/B sky130_fd_sc_hd__dfxtp_1_391/CLK
+ sky130_fd_sc_hd__and2_0_135/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_6 sky130_fd_sc_hd__nand3_1_6/C sky130_fd_sc_hd__nand2_1_6/B
+ sky130_fd_sc_hd__nand2_1_9/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_397 VDD VSS sky130_fd_sc_hd__fa_2_1033/A sky130_fd_sc_hd__dfxtp_1_411/CLK
+ sky130_fd_sc_hd__and2_0_230/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_203 sky130_fd_sc_hd__fa_2_204/CIN sky130_fd_sc_hd__fa_2_197/A
+ sky130_fd_sc_hd__ha_2_91/A sky130_fd_sc_hd__fa_2_261/A sky130_fd_sc_hd__fa_2_281/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_214 sky130_fd_sc_hd__fa_2_216/CIN sky130_fd_sc_hd__fa_2_211/A
+ sky130_fd_sc_hd__fa_2_214/A sky130_fd_sc_hd__fa_2_214/B sky130_fd_sc_hd__fa_2_222/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_225 sky130_fd_sc_hd__fa_2_227/CIN sky130_fd_sc_hd__fa_2_220/A
+ sky130_fd_sc_hd__fa_2_225/A sky130_fd_sc_hd__fa_2_225/B sky130_fd_sc_hd__fa_2_225/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_236 sky130_fd_sc_hd__maj3_1_36/B sky130_fd_sc_hd__maj3_1_37/A
+ sky130_fd_sc_hd__fa_2_236/A sky130_fd_sc_hd__fa_2_236/B sky130_fd_sc_hd__fa_2_237/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_247 sky130_fd_sc_hd__fa_2_244/B sky130_fd_sc_hd__fa_2_247/SUM
+ sky130_fd_sc_hd__fa_2_247/A sky130_fd_sc_hd__fa_2_15/B sky130_fd_sc_hd__fa_2_242/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_258 sky130_fd_sc_hd__fa_2_260/CIN sky130_fd_sc_hd__fa_2_255/A
+ sky130_fd_sc_hd__fa_2_258/A sky130_fd_sc_hd__fa_2_258/B sky130_fd_sc_hd__fa_2_258/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_269 sky130_fd_sc_hd__fa_2_268/B sky130_fd_sc_hd__fa_2_269/SUM
+ sky130_fd_sc_hd__fa_2_269/A sky130_fd_sc_hd__fa_2_269/B sky130_fd_sc_hd__fa_2_273/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_7 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_7/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_2/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__diode_2_108 sky130_fd_sc_hd__inv_2_135/Y VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__fa_2_50 sky130_fd_sc_hd__maj3_1_19/B sky130_fd_sc_hd__maj3_1_20/A
+ sky130_fd_sc_hd__fa_2_50/A sky130_fd_sc_hd__fa_2_50/B sky130_fd_sc_hd__fa_2_51/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__diode_2_119 sky130_fd_sc_hd__buf_2_225/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__fa_2_61 sky130_fd_sc_hd__fa_2_62/CIN sky130_fd_sc_hd__fa_2_55/A
+ sky130_fd_sc_hd__ha_2_91/A sky130_fd_sc_hd__fa_2_80/B sky130_fd_sc_hd__fa_2_139/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_72 sky130_fd_sc_hd__fa_2_74/CIN sky130_fd_sc_hd__fa_2_69/A
+ sky130_fd_sc_hd__fa_2_72/A sky130_fd_sc_hd__fa_2_72/B sky130_fd_sc_hd__fa_2_80/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_83 sky130_fd_sc_hd__fa_2_85/CIN sky130_fd_sc_hd__fa_2_78/A
+ sky130_fd_sc_hd__fa_2_83/A sky130_fd_sc_hd__fa_2_83/B sky130_fd_sc_hd__fa_2_83/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_94 sky130_fd_sc_hd__maj3_1_10/B sky130_fd_sc_hd__maj3_1_11/A
+ sky130_fd_sc_hd__fa_2_94/A sky130_fd_sc_hd__fa_2_94/B sky130_fd_sc_hd__fa_2_95/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_220 VDD VSS sky130_fd_sc_hd__buf_2_220/X sky130_fd_sc_hd__buf_2_220/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_231 VDD VSS sky130_fd_sc_hd__buf_2_231/X sky130_fd_sc_hd__buf_2_231/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_242 VDD VSS sky130_fd_sc_hd__buf_2_242/X sky130_fd_sc_hd__buf_2_242/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_253 VDD VSS sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__buf_2_253/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_264 VDD VSS sky130_fd_sc_hd__buf_2_264/X sky130_fd_sc_hd__nand2_2_2/Y
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_275 VDD VSS sky130_fd_sc_hd__buf_2_275/X sky130_fd_sc_hd__buf_2_275/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_286 VDD VSS sky130_fd_sc_hd__buf_2_286/X sky130_fd_sc_hd__buf_2_286/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1260 VDD VSS sky130_fd_sc_hd__mux2_2_192/A0 sky130_fd_sc_hd__clkinv_8_75/Y
+ sky130_fd_sc_hd__o22ai_1_331/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1271 VDD VSS sky130_fd_sc_hd__mux2_2_218/A0 sky130_fd_sc_hd__clkinv_8_63/Y
+ sky130_fd_sc_hd__dfxtp_1_427/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1282 VDD VSS sky130_fd_sc_hd__mux2_2_193/A0 sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__dfxtp_1_438/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1293 VDD VSS sky130_fd_sc_hd__mux2_2_186/A0 sky130_fd_sc_hd__clkinv_8_75/Y
+ sky130_fd_sc_hd__o22ai_1_342/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a21oi_1_11 sky130_fd_sc_hd__xor2_1_20/B sky130_fd_sc_hd__a21oi_1_12/Y
+ sky130_fd_sc_hd__a21oi_1_11/Y sky130_fd_sc_hd__nor2_1_11/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_22 sky130_fd_sc_hd__nand2b_1_6/Y sky130_fd_sc_hd__o21ai_1_36/Y
+ sky130_fd_sc_hd__a21oi_1_22/Y sky130_fd_sc_hd__or3_1_0/X VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_33 sky130_fd_sc_hd__nor2_1_41/Y sky130_fd_sc_hd__o22ai_1_66/Y
+ sky130_fd_sc_hd__a21oi_1_33/Y sky130_fd_sc_hd__fa_2_1036/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_44 sky130_fd_sc_hd__nor2_2_6/Y sky130_fd_sc_hd__o22ai_1_76/Y
+ sky130_fd_sc_hd__a21oi_1_44/Y sky130_fd_sc_hd__fa_2_1032/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_208 sky130_fd_sc_hd__buf_6_27/X sky130_fd_sc_hd__buf_12_208/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_55 sky130_fd_sc_hd__nor2_2_6/Y sky130_fd_sc_hd__o22ai_1_87/Y
+ sky130_fd_sc_hd__a21oi_1_55/Y sky130_fd_sc_hd__fa_2_1043/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_219 sky130_fd_sc_hd__buf_12_219/A sky130_fd_sc_hd__buf_12_249/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_66 sky130_fd_sc_hd__nand2_1_250/Y sky130_fd_sc_hd__nor2_1_49/Y
+ sky130_fd_sc_hd__xnor2_1_59/A sky130_fd_sc_hd__xnor2_1_57/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_77 sky130_fd_sc_hd__nor2_1_67/A sky130_fd_sc_hd__o21a_1_5/A1
+ sky130_fd_sc_hd__a21oi_1_77/Y sky130_fd_sc_hd__nor2_1_67/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_88 sky130_fd_sc_hd__a211o_1_3/A1 sky130_fd_sc_hd__o21ai_1_104/Y
+ sky130_fd_sc_hd__a21oi_1_88/Y sky130_fd_sc_hd__a21oi_1_88/A2 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__fa_2_770 sky130_fd_sc_hd__fa_2_768/A sky130_fd_sc_hd__fa_2_766/B
+ sky130_fd_sc_hd__ha_2_143/A sky130_fd_sc_hd__ha_2_143/B sky130_fd_sc_hd__fa_2_758/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a21oi_1_99 sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__o21ai_1_114/Y
+ sky130_fd_sc_hd__a21oi_1_99/Y sky130_fd_sc_hd__fa_2_985/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__fa_2_781 sky130_fd_sc_hd__fa_2_780/A sky130_fd_sc_hd__fa_2_781/SUM
+ sky130_fd_sc_hd__ha_2_144/B sky130_fd_sc_hd__ha_2_144/A sky130_fd_sc_hd__fa_2_758/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_792 sky130_fd_sc_hd__fa_2_796/CIN sky130_fd_sc_hd__fa_2_790/B
+ sky130_fd_sc_hd__ha_2_138/A sky130_fd_sc_hd__ha_2_136/A sky130_fd_sc_hd__fa_2_792/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor3_1_3 sky130_fd_sc_hd__or2_0_0/B sky130_fd_sc_hd__nor3_1_3/Y
+ sky130_fd_sc_hd__nor3_1_3/A sky130_fd_sc_hd__nor3_1_4/A VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__clkinv_1_408 sky130_fd_sc_hd__nand2_1_216/B sky130_fd_sc_hd__nor4_1_6/D
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_408/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_419 sky130_fd_sc_hd__or3_1_0/C sky130_fd_sc_hd__dfxtp_1_498/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_419/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__bufinv_16_0 sky130_fd_sc_hd__bufinv_16_0/A sky130_fd_sc_hd__buf_12_79/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufinv_16
Xsky130_fd_sc_hd__buf_6_40 VDD VSS sky130_fd_sc_hd__buf_6_40/X sky130_fd_sc_hd__buf_6_40/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_51 VDD VSS sky130_fd_sc_hd__buf_6_51/X sky130_fd_sc_hd__buf_6_51/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_62 VDD VSS sky130_fd_sc_hd__buf_6_62/X sky130_fd_sc_hd__buf_6_62/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_73 VDD VSS sky130_fd_sc_hd__buf_6_73/X sky130_fd_sc_hd__buf_6_73/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_84 VDD VSS sky130_fd_sc_hd__buf_6_84/X sky130_fd_sc_hd__buf_6_84/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_20 sky130_fd_sc_hd__buf_2_123/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_305 sky130_fd_sc_hd__nor2_1_188/A sky130_fd_sc_hd__o21a_1_34/A1
+ sky130_fd_sc_hd__a21oi_1_305/Y sky130_fd_sc_hd__nor2_1_188/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_31 sky130_fd_sc_hd__buf_2_107/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_316 sky130_fd_sc_hd__nor2_1_199/A sky130_fd_sc_hd__nor2_1_199/Y
+ sky130_fd_sc_hd__a21oi_1_316/Y sky130_fd_sc_hd__nor2_1_199/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_42 sky130_fd_sc_hd__buf_2_105/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_327 sky130_fd_sc_hd__clkinv_1_902/Y sky130_fd_sc_hd__nor2_1_215/Y
+ sky130_fd_sc_hd__a21oi_1_327/Y sky130_fd_sc_hd__nor2b_2_3/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_53 sky130_fd_sc_hd__buf_2_109/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_338 sky130_fd_sc_hd__fa_2_1179/A sky130_fd_sc_hd__o22ai_1_305/Y
+ sky130_fd_sc_hd__a21oi_1_338/Y sky130_fd_sc_hd__nor3_1_39/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_64 sky130_fd_sc_hd__buf_2_103/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_349 sky130_fd_sc_hd__nand2_1_439/B sky130_fd_sc_hd__o22ai_1_312/Y
+ sky130_fd_sc_hd__a21oi_1_349/Y sky130_fd_sc_hd__o21ai_1_383/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_75 sky130_fd_sc_hd__clkbuf_4_83/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_86 sky130_fd_sc_hd__clkinv_2_8/Y VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_97 sky130_fd_sc_hd__clkbuf_1_535/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a222oi_1_8 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1125/A sky130_fd_sc_hd__nor2_2_15/Y
+ sky130_fd_sc_hd__nor3_1_38/A sky130_fd_sc_hd__fa_2_1127/A sky130_fd_sc_hd__nor3_1_38/B
+ sky130_fd_sc_hd__a222oi_1_8/Y sky130_fd_sc_hd__fa_2_1124/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2_1_310 sky130_fd_sc_hd__o21a_1_11/B1 sky130_fd_sc_hd__fa_2_1062/A
+ sky130_fd_sc_hd__o21a_1_11/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_321 sky130_fd_sc_hd__nand2_1_321/Y sky130_fd_sc_hd__xor2_1_87/A
+ sky130_fd_sc_hd__nand2_1_321/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_920 sky130_fd_sc_hd__o21ai_1_365/A2 sky130_fd_sc_hd__o21ai_1_376/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_920/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_332 sky130_fd_sc_hd__nand2_1_332/Y sky130_fd_sc_hd__nand2_1_333/B
+ sky130_fd_sc_hd__nand2_1_332/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_931 sky130_fd_sc_hd__nor2_1_225/B sky130_fd_sc_hd__o21ai_1_382/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_931/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_343 sky130_fd_sc_hd__o21a_1_18/B1 sky130_fd_sc_hd__fa_2_1136/A
+ sky130_fd_sc_hd__o21a_1_18/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_290 sky130_fd_sc_hd__nand2_1_412/Y sky130_fd_sc_hd__nand2_1_411/Y
+ sky130_fd_sc_hd__o22ai_1_290/Y sky130_fd_sc_hd__nand2_1_424/B sky130_fd_sc_hd__o21ai_1_336/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_942 sky130_fd_sc_hd__nor2_1_200/B sky130_fd_sc_hd__o21bai_1_3/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_942/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_354 sky130_fd_sc_hd__o21a_1_28/B1 sky130_fd_sc_hd__fa_2_1145/A
+ sky130_fd_sc_hd__o21a_1_28/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_953 sky130_fd_sc_hd__nor2_1_265/A sky130_fd_sc_hd__nor2b_2_4/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_953/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_365 sky130_fd_sc_hd__nand2_1_365/Y sky130_fd_sc_hd__mux2_2_99/S
+ sky130_fd_sc_hd__nand2_1_365/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_964 sky130_fd_sc_hd__nor2_1_246/B sky130_fd_sc_hd__xor2_1_230/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_964/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_376 sky130_fd_sc_hd__nand2_1_376/Y sky130_fd_sc_hd__nor2b_1_104/A
+ sky130_fd_sc_hd__xor2_1_164/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_975 sky130_fd_sc_hd__nor2_1_241/B sky130_fd_sc_hd__fa_2_1246/A
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_387 sky130_fd_sc_hd__nand2_1_387/Y sky130_fd_sc_hd__nand2_1_387/B
+ sky130_fd_sc_hd__o21ai_1_316/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_986 sky130_fd_sc_hd__clkinv_1_986/Y sky130_fd_sc_hd__nand2_1_480/Y
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_398 sky130_fd_sc_hd__o21a_1_34/B1 sky130_fd_sc_hd__fa_2_1181/A
+ sky130_fd_sc_hd__o21a_1_34/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_997 sky130_fd_sc_hd__nor2_1_231/B sky130_fd_sc_hd__fa_2_1231/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_997/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_150 VDD VSS sky130_fd_sc_hd__ha_2_37/A sky130_fd_sc_hd__dfxtp_1_155/CLK
+ sky130_fd_sc_hd__and2_0_31/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_161 VDD VSS sky130_fd_sc_hd__ha_2_48/A sky130_fd_sc_hd__dfxtp_1_170/CLK
+ sky130_fd_sc_hd__nor2b_1_18/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_172 VDD VSS sky130_fd_sc_hd__nor3_2_4/B sky130_fd_sc_hd__clkinv_4_9/Y
+ sky130_fd_sc_hd__ha_2_40/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_183 VDD VSS sky130_fd_sc_hd__ha_2_51/A sky130_fd_sc_hd__dfxtp_1_185/CLK
+ sky130_fd_sc_hd__and2_0_54/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_194 VDD VSS sky130_fd_sc_hd__ha_2_62/A sky130_fd_sc_hd__dfxtp_1_197/CLK
+ sky130_fd_sc_hd__nor2b_1_34/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a21boi_1_4 sky130_fd_sc_hd__a21boi_1_4/Y sky130_fd_sc_hd__nor2_2_16/Y
+ sky130_fd_sc_hd__a21oi_1_345/Y sky130_fd_sc_hd__fa_2_1204/A VDD VSS VDD VSS sky130_fd_sc_hd__a21boi_1
Xsky130_fd_sc_hd__o211ai_1_14 sky130_fd_sc_hd__a21oi_1_200/Y sky130_fd_sc_hd__nor2_1_127/A
+ sky130_fd_sc_hd__xor2_1_119/A sky130_fd_sc_hd__nand2_1_318/Y sky130_fd_sc_hd__nand2_1_320/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_25 sky130_fd_sc_hd__nor2_1_180/A sky130_fd_sc_hd__nor2_1_174/B
+ sky130_fd_sc_hd__xor2_1_172/A sky130_fd_sc_hd__nand2_1_375/Y sky130_fd_sc_hd__nand2_1_376/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_36 sky130_fd_sc_hd__nor2_1_222/A sky130_fd_sc_hd__nor2_1_214/B
+ sky130_fd_sc_hd__xor2_1_216/A sky130_fd_sc_hd__nand2_1_426/Y sky130_fd_sc_hd__nand2_1_428/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_47 sky130_fd_sc_hd__a21oi_1_354/Y sky130_fd_sc_hd__nor2_1_222/A
+ sky130_fd_sc_hd__xor2_1_203/A sky130_fd_sc_hd__a21oi_1_351/Y sky130_fd_sc_hd__nand2_1_441/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__fa_2_1260 sky130_fd_sc_hd__fa_2_1261/CIN sky130_fd_sc_hd__mux2_2_219/A1
+ sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1260/B sky130_fd_sc_hd__nor2_8_1/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o211ai_1_58 sky130_fd_sc_hd__nor2_1_267/A sky130_fd_sc_hd__a21oi_1_414/Y
+ sky130_fd_sc_hd__xor2_1_244/A sky130_fd_sc_hd__nand2_1_492/Y sky130_fd_sc_hd__a21oi_1_406/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__fa_2_1271 sky130_fd_sc_hd__fa_2_1272/CIN sky130_fd_sc_hd__mux2_2_196/A1
+ sky130_fd_sc_hd__fa_2_1271/A sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1271/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o211ai_1_69 sky130_fd_sc_hd__nor2_1_299/A sky130_fd_sc_hd__a222oi_1_40/Y
+ sky130_fd_sc_hd__xor2_1_288/A sky130_fd_sc_hd__nand2_1_543/Y sky130_fd_sc_hd__a21oi_1_464/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__fa_2_1282 sky130_fd_sc_hd__fa_2_1283/CIN sky130_fd_sc_hd__mux2_2_246/A1
+ sky130_fd_sc_hd__fa_2_1282/A sky130_fd_sc_hd__fa_2_1282/B sky130_fd_sc_hd__fa_2_1282/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1293 sky130_fd_sc_hd__fa_2_1294/CIN sky130_fd_sc_hd__and2_0_335/A
+ sky130_fd_sc_hd__nor2_4_20/Y sky130_fd_sc_hd__fa_2_1293/B sky130_fd_sc_hd__xor2_1_317/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1090 VDD VSS sky130_fd_sc_hd__fa_2_1209/B sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__mux2_2_171/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o2bb2ai_1_30 sky130_fd_sc_hd__a221o_1_0/B2 sky130_fd_sc_hd__o21ai_1_38/A2
+ sky130_fd_sc_hd__o21ai_1_38/A1 sky130_fd_sc_hd__o21ai_1_38/Y sky130_fd_sc_hd__xor2_1_30/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__clkinv_1_205 sky130_fd_sc_hd__clkinv_1_207/A sky130_fd_sc_hd__buf_2_162/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_205/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_216 sky130_fd_sc_hd__inv_2_111/A sky130_fd_sc_hd__a22o_1_18/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_216/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_227 sky130_fd_sc_hd__inv_2_119/A sky130_fd_sc_hd__buf_8_186/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_227/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_238 sky130_fd_sc_hd__clkinv_1_238/Y sky130_fd_sc_hd__clkinv_1_238/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_238/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_249 sky130_fd_sc_hd__clkinv_1_250/A sky130_fd_sc_hd__inv_2_122/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_249/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_102 sky130_fd_sc_hd__a21o_2_3/A2 sky130_fd_sc_hd__o22ai_1_107/Y
+ sky130_fd_sc_hd__a21oi_1_102/Y sky130_fd_sc_hd__fa_2_974/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_113 sky130_fd_sc_hd__a21o_2_3/A2 sky130_fd_sc_hd__o21ai_1_137/Y
+ sky130_fd_sc_hd__o22ai_1_92/A1 sky130_fd_sc_hd__fa_2_1013/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_124 sky130_fd_sc_hd__a21o_2_3/A2 sky130_fd_sc_hd__o21ai_1_149/Y
+ sky130_fd_sc_hd__a21oi_1_124/Y sky130_fd_sc_hd__fa_2_1002/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_135 sky130_fd_sc_hd__nor2_2_10/Y sky130_fd_sc_hd__o22ai_1_135/Y
+ sky130_fd_sc_hd__a21oi_1_135/Y sky130_fd_sc_hd__fa_2_1107/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_146 sky130_fd_sc_hd__nor2_2_10/Y sky130_fd_sc_hd__o22ai_1_146/Y
+ sky130_fd_sc_hd__a21oi_1_146/Y sky130_fd_sc_hd__fa_2_1118/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nor2_1_310 sky130_fd_sc_hd__nor2_1_310/B sky130_fd_sc_hd__nor2_1_310/Y
+ sky130_fd_sc_hd__nor2_1_310/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_321 sky130_fd_sc_hd__nor2_1_321/B sky130_fd_sc_hd__nor2_1_321/Y
+ sky130_fd_sc_hd__nor2_1_322/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a21oi_1_157 sky130_fd_sc_hd__nor2_2_11/Y sky130_fd_sc_hd__o22ai_1_156/Y
+ sky130_fd_sc_hd__a21oi_1_157/Y sky130_fd_sc_hd__fa_2_1114/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_168 sky130_fd_sc_hd__clkinv_1_669/Y sky130_fd_sc_hd__nor2_1_96/B
+ sky130_fd_sc_hd__xnor2_1_81/A sky130_fd_sc_hd__xnor2_1_79/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_179 sky130_fd_sc_hd__xnor2_1_62/B sky130_fd_sc_hd__nor2_1_92/A
+ sky130_fd_sc_hd__xnor2_1_64/A sky130_fd_sc_hd__nand2_1_301/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_8_109 sky130_fd_sc_hd__buf_8_109/A sky130_fd_sc_hd__buf_8_109/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__nand2_1_140 sky130_fd_sc_hd__nand2_1_140/Y sky130_fd_sc_hd__fa_2_713/SUM
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_151 sky130_fd_sc_hd__fa_2_62/A sky130_fd_sc_hd__fa_2_92/B
+ sky130_fd_sc_hd__fa_2_87/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_750 sky130_fd_sc_hd__nor2_1_121/B sky130_fd_sc_hd__nor2_1_139/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_750/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_162 sky130_fd_sc_hd__fa_2_239/A sky130_fd_sc_hd__fa_2_258/A
+ sky130_fd_sc_hd__fa_2_261/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_761 sky130_fd_sc_hd__ha_2_193/B sky130_fd_sc_hd__fa_2_1114/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_761/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_173 sky130_fd_sc_hd__fa_2_413/B sky130_fd_sc_hd__fa_2_424/B
+ sky130_fd_sc_hd__fa_2_286/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_772 sky130_fd_sc_hd__o22ai_1_206/B1 sky130_fd_sc_hd__nor2_4_13/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_772/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_184 sky130_fd_sc_hd__fa_2_462/A sky130_fd_sc_hd__fa_2_558/B
+ sky130_fd_sc_hd__ha_2_124/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_783 sky130_fd_sc_hd__o22ai_1_265/A2 sky130_fd_sc_hd__nor3_1_38/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_783/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_195 sky130_fd_sc_hd__fa_2_759/B sky130_fd_sc_hd__ha_2_136/A
+ sky130_fd_sc_hd__ha_2_141/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_794 sky130_fd_sc_hd__nor2_1_156/A sky130_fd_sc_hd__nor2_1_157/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_794/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor2_1_0 sky130_fd_sc_hd__xor2_1_0/B sky130_fd_sc_hd__xor2_1_0/X
+ sky130_fd_sc_hd__xor2_1_0/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand3_2_1 sky130_fd_sc_hd__nand3_2_2/A sky130_fd_sc_hd__buf_2_99/A
+ sky130_fd_sc_hd__ha_2_30/A sky130_fd_sc_hd__xor2_1_3/B VSS VDD VSS VDD sky130_fd_sc_hd__nand3_2
Xsky130_fd_sc_hd__xor2_1_15 sky130_fd_sc_hd__xor2_1_15/B sky130_fd_sc_hd__xor2_1_15/X
+ sky130_fd_sc_hd__xor2_1_15/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_26 sky130_fd_sc_hd__xor2_1_26/B sky130_fd_sc_hd__xor2_1_26/X
+ sky130_fd_sc_hd__xor2_1_26/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_37 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_990/B
+ sky130_fd_sc_hd__xor2_1_37/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_48 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_979/B
+ sky130_fd_sc_hd__xor2_1_48/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_59 sky130_fd_sc_hd__xor2_1_60/X sky130_fd_sc_hd__xor2_1_59/X
+ sky130_fd_sc_hd__nor2_4_9/B VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand2b_1_9 sky130_fd_sc_hd__nand2b_1_9/Y sky130_fd_sc_hd__nand2_1_223/A
+ sky130_fd_sc_hd__fa_2_966/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__a21o_2_5 sky130_fd_sc_hd__a21o_2_5/X sky130_fd_sc_hd__a21o_2_5/B1
+ sky130_fd_sc_hd__fa_2_1082/A sky130_fd_sc_hd__a21o_2_5/A2 VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__dfxtp_1_908 VDD VSS sky130_fd_sc_hd__fa_2_943/B sky130_fd_sc_hd__clkinv_4_22/Y
+ sky130_fd_sc_hd__o21a_1_17/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_919 VDD VSS sky130_fd_sc_hd__fa_2_1148/A sky130_fd_sc_hd__clkinv_8_73/Y
+ sky130_fd_sc_hd__mux2_2_98/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_1090 sky130_fd_sc_hd__fa_2_1091/CIN sky130_fd_sc_hd__mux2_2_42/A0
+ sky130_fd_sc_hd__fa_2_1090/A sky130_fd_sc_hd__fa_2_1090/B sky130_fd_sc_hd__fa_2_1090/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_506 VSS VDD sky130_fd_sc_hd__buf_8_198/A sky130_fd_sc_hd__clkbuf_1_515/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_517 VSS VDD sky130_fd_sc_hd__buf_8_212/A sky130_fd_sc_hd__buf_6_66/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_528 VSS VDD sky130_fd_sc_hd__buf_2_248/A sky130_fd_sc_hd__clkbuf_1_528/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_539 VSS VDD sky130_fd_sc_hd__clkbuf_1_539/X sky130_fd_sc_hd__clkbuf_1_539/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_107 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_107/A sky130_fd_sc_hd__fa_2_283/B
+ sky130_fd_sc_hd__fa_2_279/A sky130_fd_sc_hd__fa_2_5/A sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_118 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_121/B sky130_fd_sc_hd__maj3_1_107/C
+ sky130_fd_sc_hd__ha_2_118/SUM sky130_fd_sc_hd__ha_2_118/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_129 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_130/A sky130_fd_sc_hd__fa_2_591/CIN
+ sky130_fd_sc_hd__fa_2_588/A sky130_fd_sc_hd__ha_2_129/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_20 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_20/A sky130_fd_sc_hd__xor2_1_2/A
+ sky130_fd_sc_hd__ha_2_20/SUM sky130_fd_sc_hd__ha_2_20/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_31 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_31/A sky130_fd_sc_hd__ha_2_30/B
+ sky130_fd_sc_hd__ha_2_31/SUM sky130_fd_sc_hd__ha_2_31/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_42 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_42/A sky130_fd_sc_hd__ha_2_41/B
+ sky130_fd_sc_hd__ha_2_42/SUM sky130_fd_sc_hd__ha_2_42/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_53 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_53/A sky130_fd_sc_hd__ha_2_52/B
+ sky130_fd_sc_hd__ha_2_53/SUM sky130_fd_sc_hd__ha_2_53/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_64 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_64/A sky130_fd_sc_hd__ha_2_63/B
+ sky130_fd_sc_hd__ha_2_64/SUM sky130_fd_sc_hd__ha_2_64/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_75 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_75/A sky130_fd_sc_hd__ha_2_74/B
+ sky130_fd_sc_hd__ha_2_75/SUM sky130_fd_sc_hd__ha_2_75/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_86 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_86/A sky130_fd_sc_hd__ha_2_85/B
+ sky130_fd_sc_hd__ha_2_86/SUM sky130_fd_sc_hd__ha_2_86/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_97 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_97/A sky130_fd_sc_hd__fa_2_116/B
+ sky130_fd_sc_hd__ha_2_97/SUM sky130_fd_sc_hd__ha_2_97/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_5 VSS VDD sky130_fd_sc_hd__buf_4_4/A sky130_fd_sc_hd__clkbuf_1_5/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__sdlclkp_4_60 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__clkinv_8_61/Y
+ sky130_fd_sc_hd__dfxtp_1_520/CLK sky130_fd_sc_hd__nand2b_1_5/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_71 sky130_fd_sc_hd__conb_1_23/LO sky130_fd_sc_hd__clkinv_8_40/A
+ sky130_fd_sc_hd__dfxtp_1_627/CLK sky130_fd_sc_hd__or2_0_6/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_82 sky130_fd_sc_hd__conb_1_26/LO sky130_fd_sc_hd__clkinv_8_68/Y
+ sky130_fd_sc_hd__dfxtp_1_1038/CLK sky130_fd_sc_hd__or2_0_10/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_140 sky130_fd_sc_hd__nor2_1_140/B sky130_fd_sc_hd__nor2_1_140/Y
+ sky130_fd_sc_hd__or2_0_7/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_151 sky130_fd_sc_hd__nor2_1_151/B sky130_fd_sc_hd__o21a_1_24/A1
+ sky130_fd_sc_hd__o21a_1_25/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_1_5 sky130_fd_sc_hd__nor2_4_4/A sky130_fd_sc_hd__nand2_1_9/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_5/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_162 sky130_fd_sc_hd__or3_1_2/C sky130_fd_sc_hd__nor2_1_162/Y
+ sky130_fd_sc_hd__or3_1_2/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_173 sky130_fd_sc_hd__nor2_1_183/A sky130_fd_sc_hd__nor2_1_173/Y
+ sky130_fd_sc_hd__nor2_1_173/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_184 sky130_fd_sc_hd__nor2_1_218/A sky130_fd_sc_hd__o21a_1_30/A1
+ sky130_fd_sc_hd__o21a_1_31/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_60 sky130_fd_sc_hd__nor2_2_2/Y sky130_fd_sc_hd__a22oi_1_82/A1
+ sky130_fd_sc_hd__clkbuf_1_61/X sky130_fd_sc_hd__a22oi_1_60/A2 sky130_fd_sc_hd__nand4_1_9/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_195 sky130_fd_sc_hd__nor2_1_195/B sky130_fd_sc_hd__o21a_1_39/A1
+ sky130_fd_sc_hd__o21a_1_40/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_71 sky130_fd_sc_hd__a22oi_2_9/B1 sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__clkbuf_4_29/X sky130_fd_sc_hd__a22oi_1_71/A2 sky130_fd_sc_hd__a22oi_1_71/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_82 sky130_fd_sc_hd__nor2_2_2/Y sky130_fd_sc_hd__a22oi_1_82/A1
+ sky130_fd_sc_hd__clkbuf_1_55/X sky130_fd_sc_hd__clkbuf_1_51/X sky130_fd_sc_hd__nand4_1_15/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_93 sky130_fd_sc_hd__a22oi_1_97/B1 sky130_fd_sc_hd__a22oi_1_97/A1
+ sky130_fd_sc_hd__buf_2_63/X sky130_fd_sc_hd__clkbuf_4_87/X sky130_fd_sc_hd__nand4_1_18/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_380 sky130_fd_sc_hd__buf_12_380/A sky130_fd_sc_hd__buf_12_505/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_391 sky130_fd_sc_hd__buf_4_112/A sky130_fd_sc_hd__buf_12_490/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_250 sky130_fd_sc_hd__a22oi_2_25/B1 sky130_fd_sc_hd__a22oi_2_25/A1
+ sky130_fd_sc_hd__clkbuf_1_383/X sky130_fd_sc_hd__a22oi_1_250/A2 sky130_fd_sc_hd__buf_2_236/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_261 sky130_fd_sc_hd__clkbuf_4_165/X sky130_fd_sc_hd__clkinv_2_23/Y
+ sky130_fd_sc_hd__clkbuf_1_412/X sky130_fd_sc_hd__a22oi_1_261/A2 sky130_fd_sc_hd__a22oi_1_261/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_272 sky130_fd_sc_hd__clkbuf_1_376/X sky130_fd_sc_hd__nor2_2_5/Y
+ sky130_fd_sc_hd__buf_2_214/X sky130_fd_sc_hd__clkbuf_1_470/X sky130_fd_sc_hd__nand4_1_67/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_283 sky130_fd_sc_hd__nor2_2_4/Y sky130_fd_sc_hd__clkbuf_1_377/X
+ sky130_fd_sc_hd__a22oi_1_283/B2 sky130_fd_sc_hd__clkbuf_4_186/X sky130_fd_sc_hd__nand4_1_70/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_4_101 VDD VSS sky130_fd_sc_hd__buf_4_101/X sky130_fd_sc_hd__buf_4_101/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__a22oi_1_294 sky130_fd_sc_hd__clkbuf_1_378/X sky130_fd_sc_hd__clkbuf_1_379/X
+ sky130_fd_sc_hd__clkbuf_4_169/X sky130_fd_sc_hd__buf_2_193/X sky130_fd_sc_hd__nand4_1_73/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_4_112 VDD VSS sky130_fd_sc_hd__buf_6_81/A sky130_fd_sc_hd__buf_4_112/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_8_19 sky130_fd_sc_hd__buf_8_19/A sky130_fd_sc_hd__buf_8_19/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__clkinv_1_580 sky130_fd_sc_hd__o22ai_1_132/B2 sky130_fd_sc_hd__fa_2_1009/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_580/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_591 sky130_fd_sc_hd__nor2_1_71/B sky130_fd_sc_hd__nor2_1_89/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_591/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_4_60 sky130_fd_sc_hd__clkinv_4_60/A sky130_fd_sc_hd__clkinv_4_60/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_60/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_71 sky130_fd_sc_hd__clkinv_4_71/A sky130_fd_sc_hd__clkinv_4_73/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_71/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_1/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__o21ai_1_505 VSS VDD sky130_fd_sc_hd__nand2_1_566/A sky130_fd_sc_hd__o21ai_1_507/A1
+ sky130_fd_sc_hd__nand2_1_566/Y sky130_fd_sc_hd__and2_0_354/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_310 sky130_fd_sc_hd__nor2_4_20/Y sky130_fd_sc_hd__fa_2_1300/B
+ sky130_fd_sc_hd__xor2_1_310/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_705 VDD VSS sky130_fd_sc_hd__mux2_2_23/A1 sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__o21ai_1_45/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_716 VDD VSS sky130_fd_sc_hd__mux2_2_2/A1 sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__o21ai_1_56/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_727 VDD VSS sky130_fd_sc_hd__mux2_2_18/A1 sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__o21ai_1_64/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_738 VDD VSS sky130_fd_sc_hd__and2_0_179/A sky130_fd_sc_hd__dfxtp_1_747/CLK
+ sky130_fd_sc_hd__fa_2_1093/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_749 VDD VSS sky130_fd_sc_hd__and2_0_173/A sky130_fd_sc_hd__dfxtp_1_755/CLK
+ sky130_fd_sc_hd__fa_2_1104/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_303 VSS VDD sky130_fd_sc_hd__nand4_1_42/D sky130_fd_sc_hd__a22oi_1_187/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_314 VSS VDD sky130_fd_sc_hd__inv_2_74/A sky130_fd_sc_hd__a22o_1_10/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_325 VSS VDD sky130_fd_sc_hd__buf_8_154/A sky130_fd_sc_hd__buf_4_90/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_336 VSS VDD sky130_fd_sc_hd__clkbuf_1_336/X sky130_fd_sc_hd__clkbuf_1_336/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_347 VSS VDD sky130_fd_sc_hd__buf_8_162/A sky130_fd_sc_hd__buf_4_82/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_358 VSS VDD sky130_fd_sc_hd__clkbuf_1_359/A sky130_fd_sc_hd__buf_8_129/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_369 VSS VDD sky130_fd_sc_hd__buf_4_84/A sky130_fd_sc_hd__buf_8_164/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_40 VDD VSS sky130_fd_sc_hd__fa_2_911/CIN sky130_fd_sc_hd__clkinv_4_80/Y
+ sky130_fd_sc_hd__buf_2_288/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_51 VDD VSS sky130_fd_sc_hd__ha_2_122/B sky130_fd_sc_hd__dfxtp_1_61/CLK
+ sky130_fd_sc_hd__nand4_1_37/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_62 VDD VSS sky130_fd_sc_hd__ha_2_91/A sky130_fd_sc_hd__dfxtp_1_73/CLK
+ sky130_fd_sc_hd__dfxtp_1_62/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_73 VDD VSS sky130_fd_sc_hd__ha_2_97/B sky130_fd_sc_hd__dfxtp_1_73/CLK
+ sky130_fd_sc_hd__buf_2_287/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_84 VDD VSS sky130_fd_sc_hd__a22o_1_0/B2 sky130_fd_sc_hd__dfxtp_1_93/CLK
+ sky130_fd_sc_hd__dfxtp_1_84/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_95 VDD VSS sky130_fd_sc_hd__ha_2_9/A sky130_fd_sc_hd__dfxtp_1_95/CLK
+ sky130_fd_sc_hd__and2_0_13/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_4_130 sky130_fd_sc_hd__clkbuf_4_130/X sky130_fd_sc_hd__clkbuf_4_130/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_301 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_301/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_301/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_141 sky130_fd_sc_hd__nand4_1_44/B sky130_fd_sc_hd__a22oi_1_197/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_312 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_312/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_312/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_152 sky130_fd_sc_hd__nand4_1_33/B sky130_fd_sc_hd__a22oi_1_153/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_323 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_323/X sky130_fd_sc_hd__buf_2_263/A
+ sky130_fd_sc_hd__nor3_1_38/C sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_163 sky130_fd_sc_hd__clkbuf_4_163/X sky130_fd_sc_hd__buf_2_147/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_334 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_334/X sky130_fd_sc_hd__inv_2_140/Y
+ sky130_fd_sc_hd__and2_0_334/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_174 sky130_fd_sc_hd__clkbuf_4_174/X sky130_fd_sc_hd__clkbuf_4_174/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_345 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_345/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_345/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_185 sky130_fd_sc_hd__clkbuf_4_185/X sky130_fd_sc_hd__clkbuf_4_185/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_196 sky130_fd_sc_hd__nand4_1_76/D sky130_fd_sc_hd__a22oi_1_305/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__conb_1_9 sky130_fd_sc_hd__conb_1_9/LO sky130_fd_sc_hd__conb_1_9/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__inv_2_101 sky130_fd_sc_hd__inv_2_101/A sky130_fd_sc_hd__inv_2_101/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_112 sky130_fd_sc_hd__inv_2_112/A sky130_fd_sc_hd__inv_2_112/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__or2_0_3 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__or2_0_3/X sky130_fd_sc_hd__or2_0_3/B
+ VSS VDD VSS VDD sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__inv_2_123 sky130_fd_sc_hd__inv_2_123/A sky130_fd_sc_hd__inv_2_123/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_134 sky130_fd_sc_hd__buf_6_62/A sky130_fd_sc_hd__inv_2_134/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__o22ai_1_108 sky130_fd_sc_hd__o21a_1_8/A2 sky130_fd_sc_hd__nor2_1_66/B
+ sky130_fd_sc_hd__nor2_1_81/B sky130_fd_sc_hd__o22ai_1_117/A1 sky130_fd_sc_hd__o21ai_1_92/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__o22ai_1_119 sky130_fd_sc_hd__o22ai_1_132/B1 sky130_fd_sc_hd__nor2_1_67/B
+ sky130_fd_sc_hd__o22ai_1_119/Y sky130_fd_sc_hd__o22ai_1_119/A1 sky130_fd_sc_hd__o21ai_1_92/A1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nor2_2_19 sky130_fd_sc_hd__nor2_2_19/B sky130_fd_sc_hd__nor2_2_19/Y
+ sky130_fd_sc_hd__nor4_1_13/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__o211ai_1_9 sky130_fd_sc_hd__nor2_1_83/Y sky130_fd_sc_hd__nor2_1_77/A
+ sky130_fd_sc_hd__xor2_1_82/A sky130_fd_sc_hd__o211ai_1_9/C1 sky130_fd_sc_hd__o211ai_1_9/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__a211o_1_2 VSS VDD VSS VDD sky130_fd_sc_hd__a211o_1_2/X sky130_fd_sc_hd__o221ai_1_1/Y
+ sky130_fd_sc_hd__o22ai_1_59/Y sky130_fd_sc_hd__a31oi_1_1/A1 sky130_fd_sc_hd__a21oi_1_25/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o21ai_1_302 VSS VDD sky130_fd_sc_hd__nor2_1_180/A sky130_fd_sc_hd__a21oi_1_278/Y
+ sky130_fd_sc_hd__a211oi_1_12/Y sky130_fd_sc_hd__xor2_1_180/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_313 VSS VDD sky130_fd_sc_hd__a222oi_1_10/Y sky130_fd_sc_hd__nor2_1_180/A
+ sky130_fd_sc_hd__a21oi_1_281/Y sky130_fd_sc_hd__xor2_1_149/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_324 VSS VDD sky130_fd_sc_hd__nor2_1_180/A sky130_fd_sc_hd__a21oi_1_296/Y
+ sky130_fd_sc_hd__a211oi_1_15/Y sky130_fd_sc_hd__xor2_1_159/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_335 VSS VDD sky130_fd_sc_hd__nand2_1_423/B sky130_fd_sc_hd__nor2_1_212/Y
+ sky130_fd_sc_hd__nor2_1_211/B sky130_fd_sc_hd__o21ai_1_335/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_40 sky130_fd_sc_hd__o21a_1_40/X sky130_fd_sc_hd__o21a_1_40/A1
+ sky130_fd_sc_hd__o21a_1_40/B1 sky130_fd_sc_hd__fa_2_1199/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21ai_1_346 VSS VDD sky130_fd_sc_hd__nor2_1_217/B sky130_fd_sc_hd__nor2_1_224/A
+ sky130_fd_sc_hd__a21oi_1_323/Y sky130_fd_sc_hd__xor2_1_214/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_51 sky130_fd_sc_hd__o21a_1_51/X sky130_fd_sc_hd__o21a_1_51/A1
+ sky130_fd_sc_hd__o21a_1_51/B1 sky130_fd_sc_hd__fa_2_1254/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21ai_1_357 VSS VDD sky130_fd_sc_hd__a222oi_1_18/Y sky130_fd_sc_hd__nor2_1_224/A
+ sky130_fd_sc_hd__a22oi_1_383/Y sky130_fd_sc_hd__o21ai_1_357/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_62 sky130_fd_sc_hd__o21a_1_62/X sky130_fd_sc_hd__o21a_1_62/A1
+ sky130_fd_sc_hd__o21a_1_62/B1 sky130_fd_sc_hd__fa_2_1309/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__a211oi_1_18 sky130_fd_sc_hd__nor2_1_224/Y sky130_fd_sc_hd__nor2_1_214/Y
+ sky130_fd_sc_hd__nor2_1_215/Y sky130_fd_sc_hd__a211oi_1_18/Y sky130_fd_sc_hd__fa_2_1182/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_368 VSS VDD sky130_fd_sc_hd__o21a_1_42/X sky130_fd_sc_hd__nor2_1_224/A
+ sky130_fd_sc_hd__a21oi_1_342/Y sky130_fd_sc_hd__xor2_1_197/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a211oi_1_29 sky130_fd_sc_hd__nor2b_1_119/Y sky130_fd_sc_hd__nor2_1_264/Y
+ sky130_fd_sc_hd__o21ai_1_433/Y sky130_fd_sc_hd__a211oi_1_29/Y sky130_fd_sc_hd__o21ai_1_434/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_379 VSS VDD sky130_fd_sc_hd__a211oi_1_23/Y sky130_fd_sc_hd__nor2_1_225/A
+ sky130_fd_sc_hd__a22oi_1_386/Y sky130_fd_sc_hd__o21ai_1_379/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__mux2_2_15 VSS VDD sky130_fd_sc_hd__mux2_2_15/A1 sky130_fd_sc_hd__mux2_2_15/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_15/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_26 VSS VDD sky130_fd_sc_hd__mux2_2_26/A1 sky130_fd_sc_hd__mux2_2_26/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_26/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_37 VSS VDD sky130_fd_sc_hd__mux2_2_37/A1 sky130_fd_sc_hd__mux2_2_37/A0
+ sky130_fd_sc_hd__mux2_2_37/S sky130_fd_sc_hd__mux2_2_37/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_48 VSS VDD sky130_fd_sc_hd__mux2_2_48/A1 sky130_fd_sc_hd__mux2_2_48/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_48/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_59 VSS VDD sky130_fd_sc_hd__mux2_2_59/A1 sky130_fd_sc_hd__mux2_2_59/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_59/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__xor2_1_140 sky130_fd_sc_hd__xor2_1_185/B sky130_fd_sc_hd__xor2_1_140/X
+ sky130_fd_sc_hd__xor2_1_185/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_151 sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__fa_2_1132/B
+ sky130_fd_sc_hd__xor2_1_151/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_502 VDD VSS sky130_fd_sc_hd__dfxtp_1_502/Q sky130_fd_sc_hd__dfxtp_1_502/CLK
+ sky130_fd_sc_hd__nor2b_1_62/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_162 sky130_fd_sc_hd__xor2_1_162/B sky130_fd_sc_hd__xor2_1_162/X
+ sky130_fd_sc_hd__xor2_1_163/X VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_513 VDD VSS sky130_fd_sc_hd__nor4_1_11/B sky130_fd_sc_hd__dfxtp_1_520/CLK
+ sky130_fd_sc_hd__a22o_1_58/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_173 sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__fa_2_1149/B
+ sky130_fd_sc_hd__xor2_1_173/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_524 VDD VSS sky130_fd_sc_hd__fa_2_967/A sky130_fd_sc_hd__dfxtp_1_526/CLK
+ sky130_fd_sc_hd__and2_0_268/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_184 sky130_fd_sc_hd__fa_2_1172/B sky130_fd_sc_hd__xor2_1_184/X
+ sky130_fd_sc_hd__nor2_4_14/B VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_195 sky130_fd_sc_hd__fa_2_1173/A sky130_fd_sc_hd__fa_2_1184/B
+ sky130_fd_sc_hd__xor2_1_195/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_535 VDD VSS sky130_fd_sc_hd__fa_2_956/A sky130_fd_sc_hd__dfxtp_1_538/CLK
+ sky130_fd_sc_hd__a22o_1_50/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_546 VDD VSS sky130_fd_sc_hd__fa_2_945/A sky130_fd_sc_hd__dfxtp_1_548/CLK
+ sky130_fd_sc_hd__a22o_1_39/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_557 VDD VSS sky130_fd_sc_hd__and2_0_221/A sky130_fd_sc_hd__dfxtp_1_571/CLK
+ sky130_fd_sc_hd__dfxtp_1_558/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_568 VDD VSS sky130_fd_sc_hd__dfxtp_1_568/Q sky130_fd_sc_hd__dfxtp_1_595/CLK
+ sky130_fd_sc_hd__nor2_1_24/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_579 VDD VSS sky130_fd_sc_hd__nor4_1_7/A sky130_fd_sc_hd__dfxtp_1_591/CLK
+ sky130_fd_sc_hd__and2_0_254/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_100 VSS VDD sky130_fd_sc_hd__a22oi_1_81/B1 sky130_fd_sc_hd__nor3_1_6/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_111 VSS VDD sky130_fd_sc_hd__buf_8_48/A sky130_fd_sc_hd__inv_2_3/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_122 VSS VDD sky130_fd_sc_hd__clkbuf_1_122/X sky130_fd_sc_hd__buf_8_8/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_133 VSS VDD sky130_fd_sc_hd__clkbuf_1_193/A sky130_fd_sc_hd__ha_2_47/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_144 VSS VDD sky130_fd_sc_hd__clkbuf_1_144/X sky130_fd_sc_hd__clkbuf_1_144/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_155 VSS VDD sky130_fd_sc_hd__clkbuf_1_155/X sky130_fd_sc_hd__clkbuf_1_155/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_2 VDD VSS sky130_fd_sc_hd__dfxtp_1_2/Q sky130_fd_sc_hd__dfxtp_1_8/CLK
+ sky130_fd_sc_hd__o21a_1_0/A2 VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_166 VSS VDD sky130_fd_sc_hd__clkbuf_1_166/X sky130_fd_sc_hd__clkbuf_1_166/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_177 VSS VDD sky130_fd_sc_hd__nand4_1_29/B sky130_fd_sc_hd__a22oi_1_137/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_188 VSS VDD sky130_fd_sc_hd__nand4_1_17/B sky130_fd_sc_hd__a22oi_1_90/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_199 VSS VDD sky130_fd_sc_hd__buf_8_75/A sky130_fd_sc_hd__ha_2_49/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_407 sky130_fd_sc_hd__fa_2_410/B sky130_fd_sc_hd__fa_2_407/SUM
+ sky130_fd_sc_hd__fa_2_407/A sky130_fd_sc_hd__fa_2_407/B sky130_fd_sc_hd__o22ai_1_27/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_418 sky130_fd_sc_hd__fa_2_322/A sky130_fd_sc_hd__maj3_1_56/A
+ sky130_fd_sc_hd__fa_2_418/A sky130_fd_sc_hd__fa_2_418/B sky130_fd_sc_hd__fa_2_420/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_429 sky130_fd_sc_hd__fa_2_428/CIN sky130_fd_sc_hd__fa_2_429/SUM
+ sky130_fd_sc_hd__fa_2_429/A sky130_fd_sc_hd__fa_2_429/B sky130_fd_sc_hd__fa_2_429/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nand3_1_11 sky130_fd_sc_hd__nand3_1_11/Y sky130_fd_sc_hd__a22oi_2_0/Y
+ sky130_fd_sc_hd__nand3_1_11/C sky130_fd_sc_hd__nand3_1_11/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_22 sky130_fd_sc_hd__nand3_1_22/Y sky130_fd_sc_hd__nor2_4_3/Y
+ sky130_fd_sc_hd__nand3_2_0/B sky130_fd_sc_hd__xor2_1_2/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_33 sky130_fd_sc_hd__buf_2_132/A sky130_fd_sc_hd__and2_0_37/X
+ sky130_fd_sc_hd__nand3_2_4/C sky130_fd_sc_hd__nor2_4_2/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_44 sky130_fd_sc_hd__nand3_1_44/Y sky130_fd_sc_hd__or4_1_2/D
+ sky130_fd_sc_hd__nor3_1_31/B sky130_fd_sc_hd__nor3_1_32/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__dfxtp_1_1420 VDD VSS sky130_fd_sc_hd__mux2_2_250/A0 sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__dfxtp_1_435/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1431 VDD VSS sky130_fd_sc_hd__mux2_2_242/A0 sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__o22ai_1_402/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1442 VDD VSS sky130_fd_sc_hd__buf_6_87/A sky130_fd_sc_hd__clkinv_8_116/Y
+ sky130_fd_sc_hd__nor4_1_13/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1453 VDD VSS sky130_fd_sc_hd__buf_4_64/A sky130_fd_sc_hd__sdlclkp_1_6/GCLK
+ sky130_fd_sc_hd__and2_0_348/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1464 VDD VSS sky130_fd_sc_hd__buf_4_56/A sky130_fd_sc_hd__dfxtp_1_1464/CLK
+ sky130_fd_sc_hd__and2_0_340/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_120 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_120/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_919/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_131 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_131/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__fa_2_868/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_142 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_142/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_895/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_50 sky130_fd_sc_hd__inv_2_39/A sky130_fd_sc_hd__inv_2_25/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_50/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_153 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_153/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_845/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_61 sky130_fd_sc_hd__clkinv_1_61/Y sky130_fd_sc_hd__ha_2_49/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_61/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_164 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_164/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_164/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_72 sky130_fd_sc_hd__inv_2_46/A sky130_fd_sc_hd__dfxtp_1_256/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_72/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_175 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_175/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__xor2_1_14/X sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_83 sky130_fd_sc_hd__clkinv_1_95/A sky130_fd_sc_hd__clkinv_2_5/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_83/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_186 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_186/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__fa_2_929/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_94 sky130_fd_sc_hd__inv_2_58/A sky130_fd_sc_hd__buf_2_47/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_94/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_197 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_197/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__ha_2_163/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__fa_2_930 sky130_fd_sc_hd__fa_2_929/CIN sky130_fd_sc_hd__fa_2_930/SUM
+ sky130_fd_sc_hd__ha_2_119/A sky130_fd_sc_hd__fa_2_930/B sky130_fd_sc_hd__fa_2_930/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_941 sky130_fd_sc_hd__fa_2_917/A sky130_fd_sc_hd__fa_2_918/B
+ sky130_fd_sc_hd__fa_2_941/A sky130_fd_sc_hd__fa_2_941/B sky130_fd_sc_hd__fa_2_546/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_952 sky130_fd_sc_hd__fa_2_951/CIN sky130_fd_sc_hd__fa_2_952/SUM
+ sky130_fd_sc_hd__fa_2_952/A sky130_fd_sc_hd__fa_2_952/B sky130_fd_sc_hd__fa_2_952/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_963 sky130_fd_sc_hd__fa_2_962/CIN sky130_fd_sc_hd__fa_2_963/SUM
+ sky130_fd_sc_hd__fa_2_963/A sky130_fd_sc_hd__fa_2_963/B sky130_fd_sc_hd__fa_2_963/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_974 sky130_fd_sc_hd__fa_2_975/CIN sky130_fd_sc_hd__fa_2_974/SUM
+ sky130_fd_sc_hd__fa_2_974/A sky130_fd_sc_hd__fa_2_974/B sky130_fd_sc_hd__fa_2_974/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_985 sky130_fd_sc_hd__fa_2_986/CIN sky130_fd_sc_hd__mux2_2_17/A0
+ sky130_fd_sc_hd__fa_2_985/A sky130_fd_sc_hd__fa_2_985/B sky130_fd_sc_hd__fa_2_985/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_996 sky130_fd_sc_hd__fa_2_997/CIN sky130_fd_sc_hd__fa_2_996/SUM
+ sky130_fd_sc_hd__fa_2_996/A sky130_fd_sc_hd__fa_2_996/B sky130_fd_sc_hd__fa_2_996/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_1_3 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_72/A
+ sky130_fd_sc_hd__clkinv_2_40/A sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_1
Xsky130_fd_sc_hd__mux2_2_230 VSS VDD sky130_fd_sc_hd__mux2_2_230/A1 sky130_fd_sc_hd__mux2_2_230/A0
+ sky130_fd_sc_hd__nor2_8_2/A sky130_fd_sc_hd__mux2_2_230/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_241 VSS VDD sky130_fd_sc_hd__mux2_2_241/A1 sky130_fd_sc_hd__mux2_2_241/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_241/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_252 VSS VDD sky130_fd_sc_hd__mux2_2_252/A1 sky130_fd_sc_hd__mux2_2_252/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_252/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_263 VSS VDD sky130_fd_sc_hd__mux2_2_263/A1 sky130_fd_sc_hd__mux2_2_263/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_263/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__o21ai_1_110 VSS VDD sky130_fd_sc_hd__o21a_1_8/A2 sky130_fd_sc_hd__nor2_1_63/B
+ sky130_fd_sc_hd__a22oi_1_326/Y sky130_fd_sc_hd__o21ai_1_110/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_121 VSS VDD sky130_fd_sc_hd__nor2_1_68/B sky130_fd_sc_hd__o21a_1_8/A2
+ sky130_fd_sc_hd__a21oi_1_106/Y sky130_fd_sc_hd__a211o_1_5/A2 VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_132 VSS VDD sky130_fd_sc_hd__o21a_1_8/X sky130_fd_sc_hd__nor2_1_76/A
+ sky130_fd_sc_hd__nand2b_1_13/Y sky130_fd_sc_hd__o21ai_1_132/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_143 VSS VDD sky130_fd_sc_hd__o21a_1_8/A2 sky130_fd_sc_hd__o21ai_1_143/A1
+ sky130_fd_sc_hd__a22oi_1_337/Y sky130_fd_sc_hd__o21ai_1_143/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_154 VSS VDD sky130_fd_sc_hd__nor2_1_76/A sky130_fd_sc_hd__a21oi_1_134/Y
+ sky130_fd_sc_hd__a21oi_1_130/Y sky130_fd_sc_hd__xor2_1_57/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_165 VSS VDD sky130_fd_sc_hd__o21ai_1_171/A2 sky130_fd_sc_hd__xnor2_1_77/Y
+ sky130_fd_sc_hd__a21oi_1_142/Y sky130_fd_sc_hd__o21ai_1_165/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_176 VSS VDD sky130_fd_sc_hd__nand2_2_5/Y sky130_fd_sc_hd__xnor2_1_65/Y
+ sky130_fd_sc_hd__a21oi_1_151/Y sky130_fd_sc_hd__o21ai_1_176/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_187 VSS VDD sky130_fd_sc_hd__nand2_2_5/Y sky130_fd_sc_hd__xnor2_1_87/Y
+ sky130_fd_sc_hd__a21oi_1_162/Y sky130_fd_sc_hd__o21ai_1_187/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_198 VSS VDD sky130_fd_sc_hd__xnor2_1_65/A sky130_fd_sc_hd__o21ai_1_198/A1
+ sky130_fd_sc_hd__nand2_1_287/B sky130_fd_sc_hd__xnor2_1_67/B VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21bai_1_0 sky130_fd_sc_hd__buf_2_263/X sky130_fd_sc_hd__o21bai_1_0/Y
+ sky130_fd_sc_hd__buf_2_262/X sky130_fd_sc_hd__nor2_1_89/Y VDD VSS VDD VSS sky130_fd_sc_hd__o21bai_1
Xsky130_fd_sc_hd__maj3_1_60 sky130_fd_sc_hd__maj3_1_61/X sky130_fd_sc_hd__maj3_1_60/X
+ sky130_fd_sc_hd__maj3_1_60/B sky130_fd_sc_hd__maj3_1_60/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_503 sky130_fd_sc_hd__o21a_1_61/B1 sky130_fd_sc_hd__fa_2_1280/A
+ sky130_fd_sc_hd__o21a_1_61/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_71 sky130_fd_sc_hd__maj3_1_72/X sky130_fd_sc_hd__maj3_1_71/X
+ sky130_fd_sc_hd__maj3_1_71/B sky130_fd_sc_hd__maj3_1_71/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_514 sky130_fd_sc_hd__nand2_1_514/Y sky130_fd_sc_hd__nor2_1_288/B
+ sky130_fd_sc_hd__nor2_1_286/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_82 sky130_fd_sc_hd__maj3_1_83/X sky130_fd_sc_hd__maj3_1_82/X
+ sky130_fd_sc_hd__maj3_1_82/B sky130_fd_sc_hd__maj3_1_82/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_525 sky130_fd_sc_hd__nor2_1_294/B sky130_fd_sc_hd__nand2_1_525/B
+ sky130_fd_sc_hd__nor2_1_295/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_93 sky130_fd_sc_hd__maj3_1_94/X sky130_fd_sc_hd__maj3_1_93/X
+ sky130_fd_sc_hd__maj3_1_93/B sky130_fd_sc_hd__maj3_1_93/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_536 sky130_fd_sc_hd__nand2_1_536/Y sky130_fd_sc_hd__fa_2_1292/A
+ sky130_fd_sc_hd__nor3_1_41/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_547 sky130_fd_sc_hd__nor2_1_310/A sky130_fd_sc_hd__nor2b_2_5/A
+ sky130_fd_sc_hd__o32ai_1_11/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_558 sky130_fd_sc_hd__nand2_1_558/Y sky130_fd_sc_hd__buf_6_88/A
+ sky130_fd_sc_hd__nand2_1_558/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_569 sky130_fd_sc_hd__nand2_1_569/Y sky130_fd_sc_hd__nor2_1_320/Y
+ sky130_fd_sc_hd__nand2_1_569/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_5 sky130_fd_sc_hd__ha_2_29/SUM sky130_fd_sc_hd__nor2b_1_5/Y
+ sky130_fd_sc_hd__or2_0_1/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1105 sky130_fd_sc_hd__nor2_1_282/B sky130_fd_sc_hd__fa_2_1299/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1105/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1116 sky130_fd_sc_hd__nor2_1_315/B sky130_fd_sc_hd__nor2_1_314/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1116/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1127 sky130_fd_sc_hd__clkinv_2_43/A sky130_fd_sc_hd__buf_6_84/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1127/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_310 VDD VSS sky130_fd_sc_hd__a22o_1_39/A1 sky130_fd_sc_hd__dfxtp_1_313/CLK
+ sky130_fd_sc_hd__and2_0_88/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_321 VDD VSS sky130_fd_sc_hd__nor4_1_2/A sky130_fd_sc_hd__dfxtp_1_325/CLK
+ sky130_fd_sc_hd__and2_0_191/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_332 VDD VSS sky130_fd_sc_hd__a22o_1_31/B2 sky130_fd_sc_hd__clkinv_4_27/Y
+ sky130_fd_sc_hd__o21ai_1_24/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_343 VDD VSS sky130_fd_sc_hd__ha_2_156/A sky130_fd_sc_hd__dfxtp_1_347/CLK
+ sky130_fd_sc_hd__o2bb2ai_1_2/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_354 VDD VSS sky130_fd_sc_hd__a22o_1_18/B2 sky130_fd_sc_hd__dfxtp_1_354/CLK
+ sky130_fd_sc_hd__ha_2_150/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_365 VDD VSS sky130_fd_sc_hd__fa_2_1109/A sky130_fd_sc_hd__dfxtp_1_380/CLK
+ sky130_fd_sc_hd__and2_0_169/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_376 VDD VSS sky130_fd_sc_hd__fa_2_1120/A sky130_fd_sc_hd__clkinv_4_32/Y
+ sky130_fd_sc_hd__and2_0_109/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_387 VDD VSS sky130_fd_sc_hd__fa_2_1115/B sky130_fd_sc_hd__dfxtp_1_391/CLK
+ sky130_fd_sc_hd__and2_0_130/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_7 sky130_fd_sc_hd__nand3_1_7/C sky130_fd_sc_hd__nand2_1_7/B
+ sky130_fd_sc_hd__nand2_1_9/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_398 VDD VSS sky130_fd_sc_hd__nor2_1_57/A sky130_fd_sc_hd__dfxtp_1_411/CLK
+ sky130_fd_sc_hd__and2_0_162/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o31ai_1_10 sky130_fd_sc_hd__o31ai_1_10/Y sky130_fd_sc_hd__o31ai_1_9/A1
+ sky130_fd_sc_hd__nor2_1_245/A sky130_fd_sc_hd__o31ai_1_9/A3 sky130_fd_sc_hd__o31ai_1_10/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__o31ai_1
Xsky130_fd_sc_hd__fa_2_204 sky130_fd_sc_hd__fa_2_206/CIN sky130_fd_sc_hd__fa_2_201/A
+ sky130_fd_sc_hd__fa_2_204/A sky130_fd_sc_hd__fa_2_204/B sky130_fd_sc_hd__fa_2_204/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_215 sky130_fd_sc_hd__maj3_1_40/B sky130_fd_sc_hd__maj3_1_41/A
+ sky130_fd_sc_hd__fa_2_215/A sky130_fd_sc_hd__fa_2_215/B sky130_fd_sc_hd__fa_2_216/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_226 sky130_fd_sc_hd__maj3_1_38/B sky130_fd_sc_hd__maj3_1_39/A
+ sky130_fd_sc_hd__fa_2_226/A sky130_fd_sc_hd__fa_2_226/B sky130_fd_sc_hd__fa_2_227/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_237 sky130_fd_sc_hd__fa_2_240/B sky130_fd_sc_hd__fa_2_237/SUM
+ sky130_fd_sc_hd__fa_2_237/A sky130_fd_sc_hd__fa_2_237/B sky130_fd_sc_hd__fa_2_237/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_248 sky130_fd_sc_hd__fa_2_250/CIN sky130_fd_sc_hd__fa_2_241/B
+ sky130_fd_sc_hd__fa_2_5/A sky130_fd_sc_hd__ha_2_91/B sky130_fd_sc_hd__fa_2_144/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_259 sky130_fd_sc_hd__maj3_1_31/B sky130_fd_sc_hd__maj3_1_32/A
+ sky130_fd_sc_hd__fa_2_259/A sky130_fd_sc_hd__fa_2_259/B sky130_fd_sc_hd__fa_2_260/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_40 sky130_fd_sc_hd__fa_2_42/CIN sky130_fd_sc_hd__fa_2_38/B
+ sky130_fd_sc_hd__ha_2_96/B sky130_fd_sc_hd__fa_2_87/A sky130_fd_sc_hd__fa_2_91/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_8 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_8/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_3/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__diode_2_109 sky130_fd_sc_hd__buf_2_211/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__fa_2_51 sky130_fd_sc_hd__fa_2_54/A sky130_fd_sc_hd__fa_2_51/SUM
+ sky130_fd_sc_hd__fa_2_51/A sky130_fd_sc_hd__fa_2_51/B sky130_fd_sc_hd__fa_2_51/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_62 sky130_fd_sc_hd__fa_2_64/CIN sky130_fd_sc_hd__fa_2_59/A
+ sky130_fd_sc_hd__fa_2_62/A sky130_fd_sc_hd__fa_2_62/B sky130_fd_sc_hd__fa_2_62/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_73 sky130_fd_sc_hd__maj3_1_14/B sky130_fd_sc_hd__maj3_1_15/A
+ sky130_fd_sc_hd__fa_2_73/A sky130_fd_sc_hd__fa_2_73/B sky130_fd_sc_hd__fa_2_74/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_84 sky130_fd_sc_hd__maj3_1_12/B sky130_fd_sc_hd__maj3_1_13/A
+ sky130_fd_sc_hd__fa_2_84/A sky130_fd_sc_hd__fa_2_84/B sky130_fd_sc_hd__fa_2_85/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_95 sky130_fd_sc_hd__fa_2_98/B sky130_fd_sc_hd__fa_2_95/SUM
+ sky130_fd_sc_hd__fa_2_95/A sky130_fd_sc_hd__fa_2_95/B sky130_fd_sc_hd__fa_2_95/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_210 VDD VSS sky130_fd_sc_hd__buf_2_210/X sky130_fd_sc_hd__buf_2_210/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_221 VDD VSS sky130_fd_sc_hd__buf_2_221/X sky130_fd_sc_hd__buf_2_221/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_232 VDD VSS sky130_fd_sc_hd__buf_2_232/X sky130_fd_sc_hd__buf_2_232/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_243 VDD VSS sky130_fd_sc_hd__buf_2_243/X sky130_fd_sc_hd__a22o_2_8/X
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_254 VDD VSS sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__buf_2_254/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_265 VDD VSS sky130_fd_sc_hd__buf_2_265/X sky130_fd_sc_hd__buf_2_265/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_276 VDD VSS sky130_fd_sc_hd__inv_2_2/A debug_en VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_287 VDD VSS sky130_fd_sc_hd__buf_2_287/X sky130_fd_sc_hd__buf_2_287/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1250 VDD VSS sky130_fd_sc_hd__nor2_8_1/A sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__nor2b_1_124/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1261 VDD VSS sky130_fd_sc_hd__mux2_2_190/A0 sky130_fd_sc_hd__clkinv_8_75/Y
+ sky130_fd_sc_hd__o22ai_1_330/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1272 VDD VSS sky130_fd_sc_hd__mux2_2_217/A0 sky130_fd_sc_hd__clkinv_8_63/Y
+ sky130_fd_sc_hd__dfxtp_1_428/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1283 VDD VSS sky130_fd_sc_hd__nand2_1_468/B sky130_fd_sc_hd__clkinv_8_66/Y
+ sky130_fd_sc_hd__xnor2_1_99/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1294 VDD VSS sky130_fd_sc_hd__mux2_2_184/A0 sky130_fd_sc_hd__clkinv_8_116/Y
+ sky130_fd_sc_hd__o22ai_1_341/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a21oi_1_12 sky130_fd_sc_hd__o21ai_1_29/Y sky130_fd_sc_hd__nor2_1_12/Y
+ sky130_fd_sc_hd__a21oi_1_12/Y sky130_fd_sc_hd__nand2_1_49/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_23 sky130_fd_sc_hd__fa_2_954/A sky130_fd_sc_hd__nor3_1_35/C
+ sky130_fd_sc_hd__nand4_1_84/D sky130_fd_sc_hd__nor3_1_35/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_34 sky130_fd_sc_hd__nor2_1_41/Y sky130_fd_sc_hd__o22ai_1_67/Y
+ sky130_fd_sc_hd__a21oi_1_34/Y sky130_fd_sc_hd__fa_2_1037/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_45 sky130_fd_sc_hd__nor2_2_6/Y sky130_fd_sc_hd__o22ai_1_77/Y
+ sky130_fd_sc_hd__a21oi_1_45/Y sky130_fd_sc_hd__fa_2_1033/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__buf_12_209 sky130_fd_sc_hd__buf_12_209/A sky130_fd_sc_hd__buf_12_209/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a21oi_1_56 sky130_fd_sc_hd__nor2_2_6/Y sky130_fd_sc_hd__o22ai_1_88/Y
+ sky130_fd_sc_hd__a21oi_1_56/Y sky130_fd_sc_hd__fa_2_1044/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_67 sky130_fd_sc_hd__nand2_1_249/Y sky130_fd_sc_hd__nor2_1_50/Y
+ sky130_fd_sc_hd__xnor2_1_55/A sky130_fd_sc_hd__xnor2_1_53/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_78 sky130_fd_sc_hd__o21a_1_6/B1 sky130_fd_sc_hd__nor2_1_68/Y
+ sky130_fd_sc_hd__a21oi_1_78/Y sky130_fd_sc_hd__nor2_1_68/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__fa_2_760 sky130_fd_sc_hd__maj3_1_143/B sky130_fd_sc_hd__maj3_1_144/A
+ sky130_fd_sc_hd__fa_2_760/A sky130_fd_sc_hd__fa_2_760/B sky130_fd_sc_hd__fa_2_761/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a21oi_1_89 sky130_fd_sc_hd__a21oi_1_89/A1 sky130_fd_sc_hd__o21ai_1_106/Y
+ sky130_fd_sc_hd__a21oi_1_89/Y sky130_fd_sc_hd__a211o_1_6/A1 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__fa_2_771 sky130_fd_sc_hd__fa_2_773/B sky130_fd_sc_hd__fa_2_767/A
+ sky130_fd_sc_hd__fa_2_832/A sky130_fd_sc_hd__ha_2_136/A sky130_fd_sc_hd__fa_2_826/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_782 sky130_fd_sc_hd__fa_2_784/B sky130_fd_sc_hd__fa_2_779/A
+ sky130_fd_sc_hd__fa_2_832/A sky130_fd_sc_hd__ha_2_136/A sky130_fd_sc_hd__ha_2_138/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_793 sky130_fd_sc_hd__fa_2_792/CIN sky130_fd_sc_hd__fa_2_793/SUM
+ sky130_fd_sc_hd__fa_2_793/A sky130_fd_sc_hd__fa_2_801/B sky130_fd_sc_hd__ha_2_145/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor3_1_4 sky130_fd_sc_hd__or2_0_0/B sky130_fd_sc_hd__nor3_1_4/Y
+ sky130_fd_sc_hd__nor3_1_4/A sky130_fd_sc_hd__nor3_1_4/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__clkinv_1_409 sky130_fd_sc_hd__nand2_1_214/B sky130_fd_sc_hd__nor4_1_8/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_409/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__bufinv_16_1 sky130_fd_sc_hd__bufinv_8_2/A sky130_fd_sc_hd__buf_6_27/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufinv_16
Xsky130_fd_sc_hd__buf_6_30 VDD VSS sky130_fd_sc_hd__buf_6_30/X sky130_fd_sc_hd__buf_6_30/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_41 VDD VSS sky130_fd_sc_hd__buf_6_41/X sky130_fd_sc_hd__buf_6_41/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_52 VDD VSS sky130_fd_sc_hd__buf_6_52/X sky130_fd_sc_hd__buf_6_52/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_63 VDD VSS sky130_fd_sc_hd__buf_6_63/X sky130_fd_sc_hd__buf_6_63/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_74 VDD VSS sky130_fd_sc_hd__buf_6_74/X sky130_fd_sc_hd__buf_6_74/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_10 sky130_fd_sc_hd__clkbuf_1_247/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__buf_6_85 VDD VSS sky130_fd_sc_hd__buf_6_85/X sky130_fd_sc_hd__buf_6_85/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_21 sky130_fd_sc_hd__buf_2_123/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_306 sky130_fd_sc_hd__o21a_1_35/B1 sky130_fd_sc_hd__nor2_1_189/Y
+ sky130_fd_sc_hd__a21oi_1_306/Y sky130_fd_sc_hd__nor2_1_189/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_32 sky130_fd_sc_hd__buf_2_107/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_317 sky130_fd_sc_hd__nor3_1_39/B sky130_fd_sc_hd__nor2b_1_112/Y
+ sky130_fd_sc_hd__a21oi_1_317/Y sky130_fd_sc_hd__nor2b_2_3/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_43 sky130_fd_sc_hd__buf_2_105/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_328 sky130_fd_sc_hd__fa_2_1187/A sky130_fd_sc_hd__o22ai_1_300/Y
+ sky130_fd_sc_hd__a21oi_1_328/Y sky130_fd_sc_hd__clkinv_1_861/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_54 sky130_fd_sc_hd__buf_2_100/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_339 sky130_fd_sc_hd__nor3_1_39/A sky130_fd_sc_hd__o22ai_1_308/Y
+ sky130_fd_sc_hd__a21oi_1_339/Y sky130_fd_sc_hd__fa_2_1178/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_65 sky130_fd_sc_hd__buf_2_103/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_76 sky130_fd_sc_hd__clkbuf_4_64/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_87 sky130_fd_sc_hd__clkinv_2_8/Y VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_98 sky130_fd_sc_hd__clkbuf_1_525/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a222oi_1_9 VSS VDD VDD VSS sky130_fd_sc_hd__fa_2_1124/A sky130_fd_sc_hd__nor2_2_15/Y
+ sky130_fd_sc_hd__nor3_1_38/A sky130_fd_sc_hd__fa_2_1126/A sky130_fd_sc_hd__nor3_1_38/B
+ sky130_fd_sc_hd__a222oi_1_9/Y sky130_fd_sc_hd__fa_2_1123/A sky130_fd_sc_hd__a222oi_1
Xsky130_fd_sc_hd__nand2_1_300 sky130_fd_sc_hd__nand2_1_300/Y sky130_fd_sc_hd__nor2_1_106/B
+ sky130_fd_sc_hd__fa_2_1108/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_311 sky130_fd_sc_hd__o21a_1_12/B1 sky130_fd_sc_hd__fa_2_1060/A
+ sky130_fd_sc_hd__o21a_1_12/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_910 sky130_fd_sc_hd__o22ai_1_307/B1 sky130_fd_sc_hd__fa_2_1189/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_910/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_322 sky130_fd_sc_hd__nand2_1_322/Y sky130_fd_sc_hd__fa_2_1064/A
+ sky130_fd_sc_hd__nor2_4_12/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_921 sky130_fd_sc_hd__clkinv_1_921/Y sky130_fd_sc_hd__a21boi_1_4/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_921/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_333 sky130_fd_sc_hd__nand2_1_333/Y sky130_fd_sc_hd__nand2_1_333/B
+ sky130_fd_sc_hd__nand2_1_333/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_932 sky130_fd_sc_hd__nor2_1_223/A sky130_fd_sc_hd__fa_2_1207/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_932/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_280 sky130_fd_sc_hd__nand2_1_412/Y sky130_fd_sc_hd__o21ai_1_331/Y
+ sky130_fd_sc_hd__o22ai_1_280/Y sky130_fd_sc_hd__nand2_1_419/B sky130_fd_sc_hd__nand2_1_411/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_344 sky130_fd_sc_hd__o21a_1_19/B1 sky130_fd_sc_hd__fa_2_1134/A
+ sky130_fd_sc_hd__o21a_1_19/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_291 sky130_fd_sc_hd__nand2_1_412/Y sky130_fd_sc_hd__nand2_1_411/Y
+ sky130_fd_sc_hd__o22ai_1_291/Y sky130_fd_sc_hd__o22ai_1_291/A1 sky130_fd_sc_hd__a21o_2_17/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_943 sky130_fd_sc_hd__nor2_4_17/B sky130_fd_sc_hd__nor2_8_0/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_943/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_355 sky130_fd_sc_hd__nor2_1_157/A sky130_fd_sc_hd__fa_2_1142/A
+ sky130_fd_sc_hd__fa_2_1141/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_954 sky130_fd_sc_hd__o32ai_1_6/A3 sky130_fd_sc_hd__fa_2_1225/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_954/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_366 sky130_fd_sc_hd__nand2_1_366/Y sky130_fd_sc_hd__o31ai_1_6/A3
+ sky130_fd_sc_hd__o31ai_1_6/A2 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_965 sky130_fd_sc_hd__o22ai_1_338/A1 sky130_fd_sc_hd__nor2_1_251/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_965/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_377 sky130_fd_sc_hd__nand2_1_377/Y sky130_fd_sc_hd__nand2_1_387/B
+ sky130_fd_sc_hd__o21ai_1_308/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_976 sky130_fd_sc_hd__o32ai_1_6/B2 sky130_fd_sc_hd__fa_2_1226/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_976/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_388 sky130_fd_sc_hd__nand2_1_388/Y sky130_fd_sc_hd__nor2b_1_104/Y
+ sky130_fd_sc_hd__o21ai_1_323/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_987 sky130_fd_sc_hd__clkinv_1_987/Y sky130_fd_sc_hd__a21boi_1_5/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_987/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_399 sky130_fd_sc_hd__o21a_1_35/B1 sky130_fd_sc_hd__fa_2_1178/A
+ sky130_fd_sc_hd__o21a_1_35/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_998 sky130_fd_sc_hd__o22ai_1_365/A1 sky130_fd_sc_hd__fa_2_1232/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_998/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_140 VDD VSS sky130_fd_sc_hd__ha_2_22/A sky130_fd_sc_hd__dfxtp_1_140/CLK
+ sky130_fd_sc_hd__nor2b_1_8/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_151 VDD VSS sky130_fd_sc_hd__ha_2_36/A sky130_fd_sc_hd__dfxtp_1_155/CLK
+ sky130_fd_sc_hd__and2_0_28/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_162 VDD VSS sky130_fd_sc_hd__dfxtp_1_162/Q sky130_fd_sc_hd__clkinv_8_14/Y
+ sky130_fd_sc_hd__nor2b_1_23/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_173 VDD VSS sky130_fd_sc_hd__nor3_1_9/B sky130_fd_sc_hd__clkinv_4_9/Y
+ sky130_fd_sc_hd__xor2_1_4/B VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_184 VDD VSS sky130_fd_sc_hd__ha_2_50/A sky130_fd_sc_hd__dfxtp_1_185/CLK
+ sky130_fd_sc_hd__and2_0_57/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_195 VDD VSS sky130_fd_sc_hd__ha_2_61/A sky130_fd_sc_hd__dfxtp_1_195/CLK
+ sky130_fd_sc_hd__nor2b_1_29/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a21boi_1_5 sky130_fd_sc_hd__a21boi_1_5/Y sky130_fd_sc_hd__nor2_2_17/Y
+ sky130_fd_sc_hd__a21oi_1_388/Y sky130_fd_sc_hd__fa_2_1237/A VDD VSS VDD VSS sky130_fd_sc_hd__a21boi_1
Xsky130_fd_sc_hd__o211ai_1_15 sky130_fd_sc_hd__a21oi_1_202/Y sky130_fd_sc_hd__nand2_2_6/Y
+ sky130_fd_sc_hd__xor2_1_120/A sky130_fd_sc_hd__nand2_1_319/Y sky130_fd_sc_hd__nand2_1_320/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_26 sky130_fd_sc_hd__nor2_1_175/B sky130_fd_sc_hd__nor2_1_180/A
+ sky130_fd_sc_hd__xor2_1_173/A sky130_fd_sc_hd__nand2_1_377/Y sky130_fd_sc_hd__a21oi_1_265/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_37 sky130_fd_sc_hd__nor2_1_222/A sky130_fd_sc_hd__nor2_1_216/B
+ sky130_fd_sc_hd__xor2_1_217/A sky130_fd_sc_hd__nand2_1_427/Y sky130_fd_sc_hd__nand2_1_428/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__fa_2_1250 sky130_fd_sc_hd__fa_2_1251/CIN sky130_fd_sc_hd__mux2_2_194/A1
+ sky130_fd_sc_hd__fa_2_1250/A sky130_fd_sc_hd__fa_2_1250/B sky130_fd_sc_hd__fa_2_1250/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o211ai_1_48 sky130_fd_sc_hd__nor2_1_265/A sky130_fd_sc_hd__nor2_1_257/B
+ sky130_fd_sc_hd__xor2_1_261/A sky130_fd_sc_hd__nand2_1_478/Y sky130_fd_sc_hd__nand2_1_480/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__fa_2_1261 sky130_fd_sc_hd__fa_2_1262/CIN sky130_fd_sc_hd__mux2_2_218/A1
+ sky130_fd_sc_hd__fa_2_1261/A sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1261/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o211ai_1_59 sky130_fd_sc_hd__a21oi_1_414/Y sky130_fd_sc_hd__nor2_1_265/A
+ sky130_fd_sc_hd__xor2_1_248/A sky130_fd_sc_hd__a21oi_1_411/Y sky130_fd_sc_hd__nand2_1_493/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__fa_2_1272 sky130_fd_sc_hd__fa_2_1273/CIN sky130_fd_sc_hd__mux2_2_193/A1
+ sky130_fd_sc_hd__fa_2_1272/A sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1272/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1283 sky130_fd_sc_hd__fa_2_1284/CIN sky130_fd_sc_hd__mux2_2_243/A1
+ sky130_fd_sc_hd__fa_2_1283/A sky130_fd_sc_hd__fa_2_1283/B sky130_fd_sc_hd__fa_2_1283/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1294 sky130_fd_sc_hd__fa_2_1295/CIN sky130_fd_sc_hd__and2_0_336/A
+ sky130_fd_sc_hd__fa_2_1294/A sky130_fd_sc_hd__fa_2_1294/B sky130_fd_sc_hd__fa_2_1294/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1080 VDD VSS sky130_fd_sc_hd__fa_2_1182/A sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__mux2_2_144/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1091 VDD VSS sky130_fd_sc_hd__fa_2_1210/A sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__mux2_2_170/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o2bb2ai_1_20 sky130_fd_sc_hd__dfxtp_1_560/D sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__dfxtp_1_560/Q sky130_fd_sc_hd__nand2_1_210/Y sky130_fd_sc_hd__nand3_1_45/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__o2bb2ai_1_31 sky130_fd_sc_hd__o2bb2ai_1_31/Y sky130_fd_sc_hd__nor2_1_91/A
+ sky130_fd_sc_hd__nor2_1_91/B sky130_fd_sc_hd__nor2_1_91/B sky130_fd_sc_hd__nor2_1_91/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_590 sky130_fd_sc_hd__maj3_1_127/B sky130_fd_sc_hd__maj3_1_128/A
+ sky130_fd_sc_hd__fa_2_599/B sky130_fd_sc_hd__fa_2_590/B sky130_fd_sc_hd__fa_2_591/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_1_206 sky130_fd_sc_hd__inv_2_108/A sky130_fd_sc_hd__buf_2_162/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_206/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_217 sky130_fd_sc_hd__inv_2_112/A sky130_fd_sc_hd__a22o_1_19/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_217/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_228 sky130_fd_sc_hd__inv_2_120/A sky130_fd_sc_hd__buf_8_201/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_228/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_239 sky130_fd_sc_hd__clkinv_1_240/A sky130_fd_sc_hd__inv_2_123/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_239/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_103 sky130_fd_sc_hd__fa_2_982/A sky130_fd_sc_hd__o22ai_1_112/Y
+ sky130_fd_sc_hd__a21oi_1_103/Y sky130_fd_sc_hd__nor2_2_8/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_114 sky130_fd_sc_hd__a21o_2_3/A2 sky130_fd_sc_hd__o21ai_1_138/Y
+ sky130_fd_sc_hd__nor2_1_73/B sky130_fd_sc_hd__fa_2_1009/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_125 sky130_fd_sc_hd__clkinv_1_461/Y sky130_fd_sc_hd__o22ai_1_133/Y
+ sky130_fd_sc_hd__a21oi_1_125/Y sky130_fd_sc_hd__a211o_1_6/A1 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_136 sky130_fd_sc_hd__nor2_2_10/Y sky130_fd_sc_hd__o22ai_1_136/Y
+ sky130_fd_sc_hd__a21oi_1_136/Y sky130_fd_sc_hd__fa_2_1108/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nor2_1_300 sky130_fd_sc_hd__nor2_1_310/A sky130_fd_sc_hd__nor2_1_300/Y
+ sky130_fd_sc_hd__nor2_1_300/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a21oi_1_147 sky130_fd_sc_hd__nor2_2_10/Y sky130_fd_sc_hd__o22ai_1_147/Y
+ sky130_fd_sc_hd__a21oi_1_147/Y sky130_fd_sc_hd__fa_2_1119/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nor2_1_311 sky130_fd_sc_hd__nor4_1_13/D sky130_fd_sc_hd__nor2_1_311/Y
+ sky130_fd_sc_hd__nor2_1_311/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a21oi_1_158 sky130_fd_sc_hd__nor2_2_11/Y sky130_fd_sc_hd__o22ai_1_157/Y
+ sky130_fd_sc_hd__a21oi_1_158/Y sky130_fd_sc_hd__fa_2_1115/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nor2_1_322 sky130_fd_sc_hd__nor2_1_322/B sky130_fd_sc_hd__nor2_1_322/Y
+ sky130_fd_sc_hd__nor2_1_322/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a21oi_1_169 sky130_fd_sc_hd__clkinv_1_667/Y sky130_fd_sc_hd__nor2_1_95/B
+ sky130_fd_sc_hd__xnor2_1_77/A sky130_fd_sc_hd__xnor2_1_75/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nand2_1_130 sky130_fd_sc_hd__nand2_1_130/Y sky130_fd_sc_hd__fa_2_708/SUM
+ sky130_fd_sc_hd__and2_0_235/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_141 sky130_fd_sc_hd__nand2_1_141/Y sky130_fd_sc_hd__nand2_1_142/Y
+ sky130_fd_sc_hd__buf_2_264/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_740 sky130_fd_sc_hd__o21ai_1_265/A2 sky130_fd_sc_hd__fa_2_1075/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_740/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_152 sky130_fd_sc_hd__fa_2_77/A sky130_fd_sc_hd__fa_2_45/A
+ sky130_fd_sc_hd__fa_2_92/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_751 sky130_fd_sc_hd__nor2_2_13/A sky130_fd_sc_hd__nor2_4_13/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_751/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_163 sky130_fd_sc_hd__fa_2_262/B sky130_fd_sc_hd__fa_2_280/A
+ sky130_fd_sc_hd__fa_2_144/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_762 sky130_fd_sc_hd__ha_2_194/B sky130_fd_sc_hd__fa_2_1113/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_762/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_174 sky130_fd_sc_hd__fa_2_417/CIN sky130_fd_sc_hd__fa_2_389/B
+ sky130_fd_sc_hd__ha_2_108/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_773 sky130_fd_sc_hd__a21o_2_5/A2 sky130_fd_sc_hd__o21a_1_16/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_773/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_185 sky130_fd_sc_hd__fa_2_611/A sky130_fd_sc_hd__ha_2_130/A
+ sky130_fd_sc_hd__ha_2_135/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_784 sky130_fd_sc_hd__nor3_1_38/B sky130_fd_sc_hd__o32ai_1_2/A3
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_784/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_196 sky130_fd_sc_hd__fa_2_776/A sky130_fd_sc_hd__fa_2_817/B
+ sky130_fd_sc_hd__ha_2_138/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_795 sky130_fd_sc_hd__o31ai_1_5/B1 sky130_fd_sc_hd__a221oi_1_2/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_795/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor2_1_1 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__xor2_1_1/X
+ sky130_fd_sc_hd__xor2_1_1/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand3_2_2 sky130_fd_sc_hd__nand3_2_2/A sky130_fd_sc_hd__nand3_2_2/Y
+ sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__nand3_2_2/C VSS VDD VSS VDD sky130_fd_sc_hd__nand3_2
Xsky130_fd_sc_hd__xor2_1_16 sky130_fd_sc_hd__xor2_1_16/B sky130_fd_sc_hd__xor2_1_16/X
+ sky130_fd_sc_hd__ha_2_148/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_27 sky130_fd_sc_hd__xor2_1_27/B sky130_fd_sc_hd__xor2_1_27/X
+ sky130_fd_sc_hd__xor2_1_27/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_38 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_989/B
+ sky130_fd_sc_hd__xor2_1_38/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_49 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_978/B
+ sky130_fd_sc_hd__xor2_1_49/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nor3_1_40 sky130_fd_sc_hd__nor3_1_40/C sky130_fd_sc_hd__nor3_1_40/Y
+ sky130_fd_sc_hd__nor3_1_40/A sky130_fd_sc_hd__nor3_1_40/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__a21o_2_6 sky130_fd_sc_hd__a21o_2_6/X sky130_fd_sc_hd__a21o_2_6/B1
+ sky130_fd_sc_hd__a21o_2_6/A1 sky130_fd_sc_hd__a21o_2_6/A2 VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__dfxtp_1_909 VDD VSS sky130_fd_sc_hd__xor2_1_25/A sky130_fd_sc_hd__clkinv_4_22/Y
+ sky130_fd_sc_hd__xnor2_1_91/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_1080 sky130_fd_sc_hd__fa_2_1081/CIN sky130_fd_sc_hd__mux2_2_62/A0
+ sky130_fd_sc_hd__fa_2_1080/A sky130_fd_sc_hd__fa_2_1080/B sky130_fd_sc_hd__fa_2_1080/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1091 sky130_fd_sc_hd__xor2_1_112/B sky130_fd_sc_hd__mux2_2_39/A0
+ sky130_fd_sc_hd__fa_2_1091/A sky130_fd_sc_hd__fa_2_1091/B sky130_fd_sc_hd__fa_2_1091/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkbuf_1_507 VSS VDD sky130_fd_sc_hd__buf_8_205/A sky130_fd_sc_hd__a22o_1_22/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_518 VSS VDD sky130_fd_sc_hd__buf_4_116/A sky130_fd_sc_hd__buf_8_200/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_529 VSS VDD sky130_fd_sc_hd__clkbuf_4_189/A sky130_fd_sc_hd__clkbuf_1_529/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__ha_2_108 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_109/B sky130_fd_sc_hd__fa_2_312/B
+ sky130_fd_sc_hd__fa_2_316/A sky130_fd_sc_hd__ha_2_108/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_119 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_119/A sky130_fd_sc_hd__fa_2_484/CIN
+ sky130_fd_sc_hd__fa_2_480/B sky130_fd_sc_hd__ha_2_119/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_10 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_10/A sky130_fd_sc_hd__xor2_1_1/A
+ sky130_fd_sc_hd__and2_2_0/A sky130_fd_sc_hd__ha_2_10/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_21 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_21/A sky130_fd_sc_hd__ha_2_20/B
+ sky130_fd_sc_hd__ha_2_21/SUM sky130_fd_sc_hd__ha_2_21/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_32 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_32/A sky130_fd_sc_hd__ha_2_31/B
+ sky130_fd_sc_hd__ha_2_32/SUM sky130_fd_sc_hd__ha_2_32/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_43 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_43/A sky130_fd_sc_hd__ha_2_42/B
+ sky130_fd_sc_hd__ha_2_43/SUM sky130_fd_sc_hd__ha_2_43/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_54 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_54/A sky130_fd_sc_hd__ha_2_53/B
+ sky130_fd_sc_hd__ha_2_54/SUM sky130_fd_sc_hd__ha_2_54/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_65 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_65/A sky130_fd_sc_hd__ha_2_64/B
+ sky130_fd_sc_hd__ha_2_65/SUM sky130_fd_sc_hd__ha_2_65/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_76 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_76/A sky130_fd_sc_hd__ha_2_75/B
+ sky130_fd_sc_hd__ha_2_76/SUM sky130_fd_sc_hd__ha_2_76/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_87 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_87/A sky130_fd_sc_hd__ha_2_86/B
+ sky130_fd_sc_hd__ha_2_87/SUM sky130_fd_sc_hd__ha_2_87/B sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__ha_2_98 VSS VDD VSS VDD sky130_fd_sc_hd__ha_2_99/B sky130_fd_sc_hd__fa_2_141/B
+ sky130_fd_sc_hd__fa_2_137/A sky130_fd_sc_hd__fa_2_5/A sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkbuf_1_6 VSS VDD sky130_fd_sc_hd__buf_6_4/A sky130_fd_sc_hd__buf_6_3/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_16_10 sky130_fd_sc_hd__buf_4_120/A sky130_fd_sc_hd__buf_2_140/X
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__sdlclkp_4_50 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__clkinv_8_104/A
+ sky130_fd_sc_hd__dfxtp_1_457/CLK sky130_fd_sc_hd__clkbuf_4_211/X VSS VDD VDD VSS
+ sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_61 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__clkinv_8_61/Y
+ sky130_fd_sc_hd__dfxtp_1_595/CLK sky130_fd_sc_hd__nand2b_1_5/Y VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_72 sky130_fd_sc_hd__conb_1_23/LO sky130_fd_sc_hd__clkinv_8_53/A
+ sky130_fd_sc_hd__dfxtp_1_601/CLK sky130_fd_sc_hd__or2_0_6/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__sdlclkp_4_83 sky130_fd_sc_hd__conb_1_26/LO sky130_fd_sc_hd__clkinv_8_68/Y
+ sky130_fd_sc_hd__dfxtp_1_1050/CLK sky130_fd_sc_hd__or2_0_10/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_130 sky130_fd_sc_hd__nor2_1_130/B sky130_fd_sc_hd__nor2_1_130/Y
+ sky130_fd_sc_hd__nor2_1_130/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_141 sky130_fd_sc_hd__nor2_1_141/B sky130_fd_sc_hd__nor2_1_141/Y
+ sky130_fd_sc_hd__nor2_1_141/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_152 sky130_fd_sc_hd__o21a_1_29/A2 sky130_fd_sc_hd__o21a_1_25/A1
+ sky130_fd_sc_hd__o21a_1_26/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__clkinv_1_6 sky130_fd_sc_hd__nor3_1_0/A sky130_fd_sc_hd__nor3_2_0/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_6/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nor2_1_163 sky130_fd_sc_hd__nor2_1_163/B sky130_fd_sc_hd__nor2_1_163/Y
+ sky130_fd_sc_hd__nor2_1_163/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_50 sky130_fd_sc_hd__a22oi_1_81/B1 sky130_fd_sc_hd__clkbuf_1_99/X
+ sky130_fd_sc_hd__clkbuf_1_44/X sky130_fd_sc_hd__clkbuf_4_19/X sky130_fd_sc_hd__nand4_1_6/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_174 sky130_fd_sc_hd__nor2_1_174/B sky130_fd_sc_hd__nor2_1_174/Y
+ sky130_fd_sc_hd__nor2_1_183/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_185 sky130_fd_sc_hd__nor2_1_185/B sky130_fd_sc_hd__o21a_1_31/A1
+ sky130_fd_sc_hd__o21a_1_32/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_61 sky130_fd_sc_hd__clkbuf_4_8/X sky130_fd_sc_hd__clkbuf_4_9/X
+ sky130_fd_sc_hd__clkbuf_1_24/X sky130_fd_sc_hd__a22oi_1_61/A2 sky130_fd_sc_hd__a22oi_1_61/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__nor2_1_196 sky130_fd_sc_hd__nor2_1_196/B sky130_fd_sc_hd__o21a_1_40/A1
+ sky130_fd_sc_hd__nor2_1_196/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a22oi_1_72 sky130_fd_sc_hd__clkbuf_4_8/X sky130_fd_sc_hd__clkbuf_4_9/X
+ sky130_fd_sc_hd__clkbuf_1_21/X sky130_fd_sc_hd__a22oi_1_72/A2 sky130_fd_sc_hd__a22oi_1_72/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_83 sky130_fd_sc_hd__a22oi_2_9/B1 sky130_fd_sc_hd__nor2_4_5/Y
+ sky130_fd_sc_hd__clkbuf_4_26/X sky130_fd_sc_hd__a22oi_1_83/A2 sky130_fd_sc_hd__a22oi_1_83/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_94 sky130_fd_sc_hd__nor2_4_6/Y sky130_fd_sc_hd__a22oi_2_12/A1
+ sky130_fd_sc_hd__buf_2_79/X sky130_fd_sc_hd__a22oi_1_94/A2 sky130_fd_sc_hd__a22oi_1_94/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_370 sky130_fd_sc_hd__buf_12_370/A sky130_fd_sc_hd__buf_12_372/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__buf_12_381 sky130_fd_sc_hd__inv_2_119/Y sky130_fd_sc_hd__buf_12_381/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_240 sky130_fd_sc_hd__buf_2_164/X sky130_fd_sc_hd__nor2_4_8/Y
+ sky130_fd_sc_hd__clkbuf_1_418/X sky130_fd_sc_hd__buf_2_227/X sky130_fd_sc_hd__nand4_1_58/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_12_392 sky130_fd_sc_hd__buf_12_392/A sky130_fd_sc_hd__buf_12_419/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__a22oi_1_251 sky130_fd_sc_hd__buf_2_166/X sky130_fd_sc_hd__buf_2_167/X
+ sky130_fd_sc_hd__a22oi_1_251/B2 sky130_fd_sc_hd__buf_2_169/X sky130_fd_sc_hd__nand4_1_62/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_262 sky130_fd_sc_hd__clkbuf_1_378/X sky130_fd_sc_hd__clkbuf_1_379/X
+ sky130_fd_sc_hd__clkbuf_4_175/X sky130_fd_sc_hd__buf_2_201/X sky130_fd_sc_hd__nand4_1_65/C
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_273 sky130_fd_sc_hd__clkbuf_4_165/X sky130_fd_sc_hd__clkinv_2_23/Y
+ sky130_fd_sc_hd__clkbuf_1_409/X sky130_fd_sc_hd__a22oi_1_273/A2 sky130_fd_sc_hd__a22oi_1_273/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__a22oi_1_284 sky130_fd_sc_hd__clkbuf_1_376/X sky130_fd_sc_hd__nor2_2_5/Y
+ sky130_fd_sc_hd__buf_2_211/X sky130_fd_sc_hd__clkbuf_1_467/X sky130_fd_sc_hd__nand4_1_70/A
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_4_102 VDD VSS sky130_fd_sc_hd__buf_4_102/X sky130_fd_sc_hd__buf_4_102/A
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__a22oi_1_295 sky130_fd_sc_hd__nor2_2_4/Y sky130_fd_sc_hd__clkbuf_1_377/X
+ sky130_fd_sc_hd__a22oi_1_295/B2 sky130_fd_sc_hd__clkbuf_4_183/X sky130_fd_sc_hd__nand4_1_73/B
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__buf_4_113 VDD VSS sky130_fd_sc_hd__buf_4_113/X sky130_fd_sc_hd__buf_8_214/X
+ VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__xnor2_1_100 VSS VDD sky130_fd_sc_hd__o21a_1_56/B1 sky130_fd_sc_hd__xnor2_1_100/Y
+ sky130_fd_sc_hd__fa_2_1292/A VDD VSS sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__clkinv_1_570 sky130_fd_sc_hd__o21ai_1_135/A1 sky130_fd_sc_hd__a211o_1_4/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_570/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_581 sky130_fd_sc_hd__o21ai_1_152/A2 sky130_fd_sc_hd__fa_2_1001/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_581/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_592 sky130_fd_sc_hd__nor2_2_9/A sky130_fd_sc_hd__nor2_2_7/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_592/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_4_50 sky130_fd_sc_hd__clkinv_4_50/A sky130_fd_sc_hd__clkinv_4_50/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_50/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_61 sky130_fd_sc_hd__clkinv_8_7/A sky130_fd_sc_hd__clkinv_4_61/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_61/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_4_72 sky130_fd_sc_hd__clkinv_4_73/A sky130_fd_sc_hd__clkinv_4_72/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkinv_4_72/w_82_21# sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__inv_16_2/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__o21ai_1_506 VSS VDD sky130_fd_sc_hd__nand2_1_567/A sky130_fd_sc_hd__o21ai_1_507/A1
+ sky130_fd_sc_hd__nand2_1_567/Y sky130_fd_sc_hd__and2_0_347/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__xor2_1_300 sky130_fd_sc_hd__nor2_4_20/Y sky130_fd_sc_hd__fa_2_1310/B
+ sky130_fd_sc_hd__xor2_1_300/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_311 sky130_fd_sc_hd__nor2_4_20/Y sky130_fd_sc_hd__fa_2_1299/B
+ sky130_fd_sc_hd__xor2_1_311/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_706 VDD VSS sky130_fd_sc_hd__mux2_2_21/A1 sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__o21ai_1_46/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_717 VDD VSS sky130_fd_sc_hd__mux2_2_30/A1 sky130_fd_sc_hd__clkinv_8_43/Y
+ sky130_fd_sc_hd__a22o_1_68/A1 VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_728 VDD VSS sky130_fd_sc_hd__mux2_2_16/A1 sky130_fd_sc_hd__clkinv_8_42/Y
+ sky130_fd_sc_hd__o21ai_1_65/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_739 VDD VSS sky130_fd_sc_hd__and2_0_180/A sky130_fd_sc_hd__dfxtp_1_747/CLK
+ sky130_fd_sc_hd__fa_2_1094/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_304 VSS VDD sky130_fd_sc_hd__nand4_1_41/D sky130_fd_sc_hd__a22oi_1_183/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_315 VSS VDD sky130_fd_sc_hd__clkinv_2_15/A sky130_fd_sc_hd__a22o_1_10/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_326 VSS VDD sky130_fd_sc_hd__buf_12_277/A sky130_fd_sc_hd__clkbuf_1_362/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_337 VSS VDD sky130_fd_sc_hd__buf_8_132/A sky130_fd_sc_hd__and2_4_0/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_348 VSS VDD sky130_fd_sc_hd__buf_8_166/A sky130_fd_sc_hd__buf_4_93/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_359 VSS VDD sky130_fd_sc_hd__buf_8_143/A sky130_fd_sc_hd__clkbuf_1_359/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_30 VDD VSS sky130_fd_sc_hd__fa_2_902/A sky130_fd_sc_hd__clkinv_4_80/Y
+ sky130_fd_sc_hd__dfxtp_1_62/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_41 VDD VSS sky130_fd_sc_hd__fa_2_912/CIN sky130_fd_sc_hd__clkinv_4_80/Y
+ sky130_fd_sc_hd__buf_2_287/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_52 VDD VSS sky130_fd_sc_hd__ha_2_123/A sky130_fd_sc_hd__dfxtp_1_60/CLK
+ sky130_fd_sc_hd__nand4_1_38/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_63 VDD VSS sky130_fd_sc_hd__ha_2_93/A sky130_fd_sc_hd__dfxtp_1_77/CLK
+ sky130_fd_sc_hd__dfxtp_1_63/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_74 VDD VSS sky130_fd_sc_hd__fa_2_82/A sky130_fd_sc_hd__dfxtp_1_77/CLK
+ sky130_fd_sc_hd__buf_2_286/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_85 VDD VSS sky130_fd_sc_hd__a22o_1_1/B2 sky130_fd_sc_hd__dfxtp_1_93/CLK
+ sky130_fd_sc_hd__buf_6_57/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_96 VDD VSS sky130_fd_sc_hd__ha_2_8/A sky130_fd_sc_hd__dfxtp_1_99/CLK
+ sky130_fd_sc_hd__and2_0_3/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_4_120 sky130_fd_sc_hd__clkbuf_4_120/X sky130_fd_sc_hd__clkbuf_4_120/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_131 sky130_fd_sc_hd__clkbuf_4_131/X sky130_fd_sc_hd__clkbuf_4_131/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_302 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_302/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_302/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_142 sky130_fd_sc_hd__nand4_1_43/B sky130_fd_sc_hd__a22oi_1_193/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_313 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_313/X sky130_fd_sc_hd__mux2_2_75/S
+ sky130_fd_sc_hd__and2_0_313/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_153 sky130_fd_sc_hd__nand4_1_32/B sky130_fd_sc_hd__a22oi_1_149/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_324 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_324/X sky130_fd_sc_hd__mux2_2_171/S
+ sky130_fd_sc_hd__and2_0_324/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_164 sky130_fd_sc_hd__clkbuf_4_164/X sky130_fd_sc_hd__buf_2_148/X
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_335 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_335/X sky130_fd_sc_hd__inv_2_140/Y
+ sky130_fd_sc_hd__and2_0_335/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_175 sky130_fd_sc_hd__clkbuf_4_175/X sky130_fd_sc_hd__clkbuf_4_175/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__and2_0_346 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_346/X sky130_fd_sc_hd__buf_6_86/X
+ sky130_fd_sc_hd__and2_0_346/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkbuf_4_186 sky130_fd_sc_hd__clkbuf_4_186/X sky130_fd_sc_hd__clkbuf_4_186/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_197 sky130_fd_sc_hd__nand4_1_72/D sky130_fd_sc_hd__a22oi_1_289/Y
+ VSS VDD VDD VSS sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__inv_2_102 sky130_fd_sc_hd__inv_2_102/A sky130_fd_sc_hd__inv_2_102/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_113 sky130_fd_sc_hd__inv_2_113/A sky130_fd_sc_hd__inv_2_113/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__or2_0_4 sky130_fd_sc_hd__or2_0_4/A sky130_fd_sc_hd__or2_0_4/X sky130_fd_sc_hd__or2_0_4/B
+ VSS VDD VSS VDD sky130_fd_sc_hd__or2_0
Xsky130_fd_sc_hd__inv_2_124 sky130_fd_sc_hd__inv_2_124/A sky130_fd_sc_hd__inv_2_124/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_135 sky130_fd_sc_hd__inv_2_136/Y sky130_fd_sc_hd__inv_2_135/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__o22ai_1_109 sky130_fd_sc_hd__o22ai_1_130/B1 sky130_fd_sc_hd__nor2_1_67/B
+ sky130_fd_sc_hd__nor2_1_81/A sky130_fd_sc_hd__nor2_1_68/B sky130_fd_sc_hd__o22ai_1_132/B1
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__a211o_1_3 VSS VDD VSS VDD sky130_fd_sc_hd__xor2_1_55/A sky130_fd_sc_hd__a211o_1_4/A2
+ sky130_fd_sc_hd__nor2_1_72/Y sky130_fd_sc_hd__a211o_1_3/A1 sky130_fd_sc_hd__o22ai_1_91/Y
+ sky130_fd_sc_hd__a211o_1
Xsky130_fd_sc_hd__o21ai_1_303 VSS VDD sky130_fd_sc_hd__a222oi_1_8/Y sky130_fd_sc_hd__nor2_1_182/A
+ sky130_fd_sc_hd__a22oi_1_375/Y sky130_fd_sc_hd__o21ai_1_303/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_314 VSS VDD sky130_fd_sc_hd__o21a_1_29/X sky130_fd_sc_hd__nor2_1_182/A
+ sky130_fd_sc_hd__a21oi_1_282/Y sky130_fd_sc_hd__xor2_1_152/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_30 sky130_fd_sc_hd__o21a_1_30/X sky130_fd_sc_hd__o21a_1_30/A1
+ sky130_fd_sc_hd__xnor2_1_94/B sky130_fd_sc_hd__fa_2_1189/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21ai_1_325 VSS VDD sky130_fd_sc_hd__a211oi_1_16/Y sky130_fd_sc_hd__nor2_1_183/A
+ sky130_fd_sc_hd__a22oi_1_378/Y sky130_fd_sc_hd__o21ai_1_325/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_336 VSS VDD sky130_fd_sc_hd__nand2_1_424/B sky130_fd_sc_hd__nor2_1_213/Y
+ sky130_fd_sc_hd__nor2_1_212/B sky130_fd_sc_hd__o21ai_1_336/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_41 sky130_fd_sc_hd__o21a_1_41/X sky130_fd_sc_hd__o21a_1_41/A1
+ sky130_fd_sc_hd__o21a_1_41/B1 sky130_fd_sc_hd__fa_2_1196/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21a_1_52 sky130_fd_sc_hd__o21a_1_52/X sky130_fd_sc_hd__o21a_1_52/A1
+ sky130_fd_sc_hd__o21a_1_52/B1 sky130_fd_sc_hd__fa_2_1252/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__o21ai_1_347 VSS VDD sky130_fd_sc_hd__a222oi_1_16/Y sky130_fd_sc_hd__nor2_1_222/A
+ sky130_fd_sc_hd__a21oi_1_324/Y sky130_fd_sc_hd__xor2_1_215/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21a_1_63 sky130_fd_sc_hd__o21a_1_63/X sky130_fd_sc_hd__o21a_1_63/A1
+ sky130_fd_sc_hd__o21a_1_63/B1 sky130_fd_sc_hd__fa_2_1307/A VDD VSS VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__a211oi_1_19 sky130_fd_sc_hd__nor2b_1_112/Y sky130_fd_sc_hd__o21ai_1_357/Y
+ sky130_fd_sc_hd__nor2_1_216/Y sky130_fd_sc_hd__a211oi_1_19/Y sky130_fd_sc_hd__o21ai_1_359/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a211oi_1
Xsky130_fd_sc_hd__o21ai_1_358 VSS VDD sky130_fd_sc_hd__o21ai_1_358/A2 sky130_fd_sc_hd__o22ai_1_322/A2
+ sky130_fd_sc_hd__a22oi_1_384/Y sky130_fd_sc_hd__o21ai_1_358/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_369 VSS VDD sky130_fd_sc_hd__a21oi_1_350/Y sky130_fd_sc_hd__nor2_1_214/A
+ sky130_fd_sc_hd__o21ai_1_371/B1 sky130_fd_sc_hd__o21ai_1_369/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__mux2_2_16 VSS VDD sky130_fd_sc_hd__mux2_2_16/A1 sky130_fd_sc_hd__mux2_2_16/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_16/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_27 VSS VDD sky130_fd_sc_hd__mux2_2_27/A1 sky130_fd_sc_hd__mux2_2_27/A0
+ sky130_fd_sc_hd__or2_0_5/A sky130_fd_sc_hd__mux2_2_27/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_38 VSS VDD sky130_fd_sc_hd__mux2_2_38/A1 sky130_fd_sc_hd__xor2_1_112/X
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_38/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_49 VSS VDD sky130_fd_sc_hd__mux2_2_49/A1 sky130_fd_sc_hd__mux2_2_49/A0
+ sky130_fd_sc_hd__or2_0_7/A sky130_fd_sc_hd__mux2_2_49/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__xor2_1_130 sky130_fd_sc_hd__nor2_4_11/Y sky130_fd_sc_hd__fa_2_1076/B
+ sky130_fd_sc_hd__xor2_1_130/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_141 sky130_fd_sc_hd__xor2_1_141/B sky130_fd_sc_hd__xor2_1_141/X
+ sky130_fd_sc_hd__xor2_1_142/X VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_152 sky130_fd_sc_hd__nor2_4_14/Y sky130_fd_sc_hd__fa_2_1131/B
+ sky130_fd_sc_hd__xor2_1_152/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_503 VDD VSS sky130_fd_sc_hd__nor2_1_36/B sky130_fd_sc_hd__edfxtp_1_0/CLK
+ sky130_fd_sc_hd__nor2b_1_79/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_163 sky130_fd_sc_hd__xor2_1_164/X sky130_fd_sc_hd__xor2_1_163/X
+ sky130_fd_sc_hd__xor2_1_163/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_514 VDD VSS sky130_fd_sc_hd__nor4_1_9/B sky130_fd_sc_hd__dfxtp_1_520/CLK
+ sky130_fd_sc_hd__a22o_1_57/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_174 sky130_fd_sc_hd__nor2_4_15/Y sky130_fd_sc_hd__fa_2_1148/B
+ sky130_fd_sc_hd__xor2_1_174/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_185 sky130_fd_sc_hd__xor2_1_185/B sky130_fd_sc_hd__xor2_1_185/X
+ sky130_fd_sc_hd__xor2_1_185/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_525 VDD VSS sky130_fd_sc_hd__fa_2_966/A sky130_fd_sc_hd__dfxtp_1_526/CLK
+ sky130_fd_sc_hd__and2_0_264/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xor2_1_196 sky130_fd_sc_hd__fa_2_1173/A sky130_fd_sc_hd__fa_2_1183/B
+ sky130_fd_sc_hd__xor2_1_196/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__dfxtp_1_536 VDD VSS sky130_fd_sc_hd__fa_2_955/A sky130_fd_sc_hd__dfxtp_1_538/CLK
+ sky130_fd_sc_hd__a22o_1_49/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_547 VDD VSS sky130_fd_sc_hd__fa_2_944/A sky130_fd_sc_hd__dfxtp_1_548/CLK
+ sky130_fd_sc_hd__a22o_1_38/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_558 VDD VSS sky130_fd_sc_hd__dfxtp_1_558/Q sky130_fd_sc_hd__dfxtp_1_576/CLK
+ sky130_fd_sc_hd__dfxtp_1_558/D VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_569 VDD VSS sky130_fd_sc_hd__and2_0_216/A sky130_fd_sc_hd__dfxtp_1_571/CLK
+ sky130_fd_sc_hd__a22o_1_35/B1 VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_101 VSS VDD sky130_fd_sc_hd__a22oi_1_82/A1 sky130_fd_sc_hd__nor3_1_8/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_112 VSS VDD sky130_fd_sc_hd__buf_12_20/A sky130_fd_sc_hd__inv_2_44/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_123 VSS VDD sky130_fd_sc_hd__buf_6_6/A sky130_fd_sc_hd__buf_6_5/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_134 VSS VDD sky130_fd_sc_hd__a22oi_2_12/A1 sky130_fd_sc_hd__nor3_2_4/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_145 VSS VDD sky130_fd_sc_hd__clkbuf_1_145/X sky130_fd_sc_hd__clkbuf_1_145/A
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_156 VSS VDD sky130_fd_sc_hd__clkbuf_1_156/X sky130_fd_sc_hd__clkbuf_1_200/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__dfxtp_1_3 VDD VSS sky130_fd_sc_hd__dfxtp_1_3/Q sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__a22o_1_0/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkbuf_1_167 VSS VDD sky130_fd_sc_hd__clkbuf_1_167/X sky130_fd_sc_hd__clkbuf_1_247/X
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_178 VSS VDD sky130_fd_sc_hd__nand4_1_28/B sky130_fd_sc_hd__a22oi_1_133/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_189 VSS VDD sky130_fd_sc_hd__nand4_1_16/B sky130_fd_sc_hd__a22oi_1_86/Y
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__fa_2_408 sky130_fd_sc_hd__fa_2_409/CIN sky130_fd_sc_hd__fa_2_403/B
+ sky130_fd_sc_hd__ha_2_115/A sky130_fd_sc_hd__fa_2_417/B sky130_fd_sc_hd__fa_2_395/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_419 sky130_fd_sc_hd__fa_2_318/A sky130_fd_sc_hd__fa_2_322/B
+ sky130_fd_sc_hd__fa_2_419/A sky130_fd_sc_hd__fa_2_419/B sky130_fd_sc_hd__fa_2_423/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nand3_1_12 sky130_fd_sc_hd__nand3_1_12/Y sky130_fd_sc_hd__nand3_1_12/A
+ sky130_fd_sc_hd__nand3_1_12/C sky130_fd_sc_hd__nand3_1_12/B VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_23 sky130_fd_sc_hd__nand3_1_23/Y sky130_fd_sc_hd__ha_2_10/A
+ sky130_fd_sc_hd__nand3_1_25/C sky130_fd_sc_hd__nand3_2_2/A VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_34 sky130_fd_sc_hd__nand3_1_34/Y sky130_fd_sc_hd__nand3_4_0/B
+ sky130_fd_sc_hd__nand3_1_35/C sky130_fd_sc_hd__nand3_4_1/A VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__nand3_1_45 sky130_fd_sc_hd__nand3_1_45/Y sky130_fd_sc_hd__or4_1_2/B
+ sky130_fd_sc_hd__nand3_1_45/C sky130_fd_sc_hd__nor3_1_32/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__dfxtp_1_1410 VDD VSS sky130_fd_sc_hd__mux2_2_221/A1 sky130_fd_sc_hd__clkinv_8_77/Y
+ sky130_fd_sc_hd__a21oi_1_442/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1421 VDD VSS sky130_fd_sc_hd__mux2_2_247/A0 sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__dfxtp_1_436/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1432 VDD VSS sky130_fd_sc_hd__mux2_2_239/A0 sky130_fd_sc_hd__clkinv_8_50/Y
+ sky130_fd_sc_hd__o22ai_1_401/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1443 VDD VSS sky130_fd_sc_hd__buf_2_283/A sky130_fd_sc_hd__clkinv_8_132/Y
+ sky130_fd_sc_hd__buf_2_272/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1454 VDD VSS sky130_fd_sc_hd__buf_4_122/A sky130_fd_sc_hd__dfxtp_1_1461/CLK
+ sky130_fd_sc_hd__and2_0_355/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1465 VDD VSS sky130_fd_sc_hd__inv_2_1/A sky130_fd_sc_hd__clkinv_8_140/Y
+ sky130_fd_sc_hd__nor2b_1_138/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__and2_0_110 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_110/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_917/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_121 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_121/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__fa_2_866/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_132 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_132/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_893/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_40 sky130_fd_sc_hd__inv_2_29/A sky130_fd_sc_hd__buf_2_11/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_40/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_143 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_143/X sky130_fd_sc_hd__buf_2_256/X
+ sky130_fd_sc_hd__fa_2_857/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_51 sky130_fd_sc_hd__inv_2_40/A sky130_fd_sc_hd__inv_2_23/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_51/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_154 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_154/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__fa_2_859/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_62 sky130_fd_sc_hd__nor2_4_6/A sky130_fd_sc_hd__nor3_2_4/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_62/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_165 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_165/X sky130_fd_sc_hd__buf_2_257/X
+ sky130_fd_sc_hd__and2_0_165/A sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_73 sky130_fd_sc_hd__inv_2_47/A sky130_fd_sc_hd__dfxtp_1_257/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_73/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_176 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_176/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__fa_2_863/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_84 sky130_fd_sc_hd__clkinv_1_86/A sky130_fd_sc_hd__ha_2_41/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_84/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_187 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_187/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__fa_2_928/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_95 sky130_fd_sc_hd__inv_2_59/A sky130_fd_sc_hd__clkinv_1_95/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_95/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_198 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_198/X sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__ha_2_164/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__fa_2_920 sky130_fd_sc_hd__fa_2_919/CIN sky130_fd_sc_hd__fa_2_920/SUM
+ sky130_fd_sc_hd__fa_2_920/A sky130_fd_sc_hd__fa_2_920/B sky130_fd_sc_hd__fa_2_920/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_931 sky130_fd_sc_hd__fa_2_927/A sky130_fd_sc_hd__fa_2_928/B
+ sky130_fd_sc_hd__fa_2_931/A sky130_fd_sc_hd__fa_2_931/B sky130_fd_sc_hd__ha_2_118/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_942 sky130_fd_sc_hd__fa_2_916/A sky130_fd_sc_hd__fa_2_917/B
+ sky130_fd_sc_hd__fa_2_942/A sky130_fd_sc_hd__fa_2_942/B sky130_fd_sc_hd__ha_2_124/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_953 sky130_fd_sc_hd__fa_2_952/CIN sky130_fd_sc_hd__fa_2_953/SUM
+ sky130_fd_sc_hd__fa_2_953/A sky130_fd_sc_hd__fa_2_953/B sky130_fd_sc_hd__fa_2_953/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_964 sky130_fd_sc_hd__fa_2_963/CIN sky130_fd_sc_hd__fa_2_964/SUM
+ sky130_fd_sc_hd__fa_2_964/A sky130_fd_sc_hd__fa_2_964/B sky130_fd_sc_hd__fa_2_964/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_975 sky130_fd_sc_hd__fa_2_976/CIN sky130_fd_sc_hd__fa_2_975/SUM
+ sky130_fd_sc_hd__fa_2_975/A sky130_fd_sc_hd__fa_2_975/B sky130_fd_sc_hd__fa_2_975/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_986 sky130_fd_sc_hd__fa_2_987/CIN sky130_fd_sc_hd__mux2_2_15/A0
+ sky130_fd_sc_hd__fa_2_986/A sky130_fd_sc_hd__fa_2_986/B sky130_fd_sc_hd__fa_2_986/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_997 sky130_fd_sc_hd__fa_2_998/CIN sky130_fd_sc_hd__fa_2_997/SUM
+ sky130_fd_sc_hd__fa_2_997/A sky130_fd_sc_hd__fa_2_997/B sky130_fd_sc_hd__fa_2_997/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_1_4 sky130_fd_sc_hd__conb_1_25/LO sky130_fd_sc_hd__clkinv_4_60/A
+ sky130_fd_sc_hd__clkinv_2_32/A sky130_fd_sc_hd__or2_0_9/B VSS VDD VDD VSS sky130_fd_sc_hd__sdlclkp_1
Xsky130_fd_sc_hd__mux2_2_220 VSS VDD sky130_fd_sc_hd__mux2_2_220/A1 sky130_fd_sc_hd__xor2_1_297/X
+ sky130_fd_sc_hd__nor2_8_2/A sky130_fd_sc_hd__mux2_2_220/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_231 VSS VDD sky130_fd_sc_hd__mux2_2_231/A1 sky130_fd_sc_hd__mux2_2_231/A0
+ sky130_fd_sc_hd__nor2_8_2/A sky130_fd_sc_hd__mux2_2_231/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_242 VSS VDD sky130_fd_sc_hd__mux2_2_242/A1 sky130_fd_sc_hd__mux2_2_242/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_242/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_253 VSS VDD sky130_fd_sc_hd__mux2_2_253/A1 sky130_fd_sc_hd__mux2_2_253/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_253/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__mux2_2_264 VSS VDD sky130_fd_sc_hd__mux2_2_264/A1 sky130_fd_sc_hd__mux2_2_264/A0
+ sky130_fd_sc_hd__inv_2_140/Y sky130_fd_sc_hd__mux2_2_264/X VDD VSS sky130_fd_sc_hd__mux2_2
Xsky130_fd_sc_hd__o21ai_1_100 VSS VDD sky130_fd_sc_hd__a21oi_1_93/Y sky130_fd_sc_hd__nor2_1_76/A
+ sky130_fd_sc_hd__nand2_1_264/Y sky130_fd_sc_hd__o21ai_1_100/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_111 VSS VDD sky130_fd_sc_hd__o21ai_1_111/A2 sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__a21oi_1_96/Y sky130_fd_sc_hd__xor2_1_75/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_122 VSS VDD sky130_fd_sc_hd__o22ai_1_122/B1 sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__nand2_1_273/Y sky130_fd_sc_hd__xor2_1_35/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_133 VSS VDD sky130_fd_sc_hd__o21ai_1_133/A2 sky130_fd_sc_hd__nor2_1_74/A
+ sky130_fd_sc_hd__a21oi_1_111/Y sky130_fd_sc_hd__xor2_1_46/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_144 VSS VDD sky130_fd_sc_hd__nor2_1_77/A sky130_fd_sc_hd__a21oi_1_129/Y
+ sky130_fd_sc_hd__a21oi_1_120/Y sky130_fd_sc_hd__xor2_1_52/A VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_155 VSS VDD sky130_fd_sc_hd__o21a_1_8/A2 sky130_fd_sc_hd__o21ai_1_155/A1
+ sky130_fd_sc_hd__a22oi_1_344/Y sky130_fd_sc_hd__o21ai_1_155/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_166 VSS VDD sky130_fd_sc_hd__o21ai_1_171/A2 sky130_fd_sc_hd__xnor2_1_79/Y
+ sky130_fd_sc_hd__a21oi_1_143/Y sky130_fd_sc_hd__o21ai_1_166/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_177 VSS VDD sky130_fd_sc_hd__nand2_2_5/Y sky130_fd_sc_hd__xnor2_1_67/Y
+ sky130_fd_sc_hd__a21oi_1_152/Y sky130_fd_sc_hd__o21ai_1_177/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_188 VSS VDD sky130_fd_sc_hd__nand2_2_5/Y sky130_fd_sc_hd__xnor2_1_89/Y
+ sky130_fd_sc_hd__a21oi_1_163/Y sky130_fd_sc_hd__o21ai_1_188/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21ai_1_199 VSS VDD sky130_fd_sc_hd__xnor2_1_88/A sky130_fd_sc_hd__nor2_1_112/Y
+ sky130_fd_sc_hd__nand2_1_294/Y sky130_fd_sc_hd__o21ai_1_199/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__o21bai_1_1 sky130_fd_sc_hd__buf_2_263/A sky130_fd_sc_hd__o21bai_1_1/Y
+ sky130_fd_sc_hd__buf_2_262/X sky130_fd_sc_hd__nor2_1_139/Y VDD VSS VDD VSS sky130_fd_sc_hd__o21bai_1
Xsky130_fd_sc_hd__maj3_1_50 sky130_fd_sc_hd__maj3_1_51/X sky130_fd_sc_hd__maj3_1_50/X
+ sky130_fd_sc_hd__maj3_1_50/B sky130_fd_sc_hd__maj3_1_50/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__maj3_1_61 sky130_fd_sc_hd__maj3_1_62/X sky130_fd_sc_hd__maj3_1_61/X
+ sky130_fd_sc_hd__maj3_1_61/B sky130_fd_sc_hd__maj3_1_61/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_504 sky130_fd_sc_hd__nor2_1_276/A sky130_fd_sc_hd__fa_2_1277/A
+ sky130_fd_sc_hd__fa_2_1276/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_72 sky130_fd_sc_hd__maj3_1_73/X sky130_fd_sc_hd__maj3_1_72/X
+ sky130_fd_sc_hd__maj3_1_72/B sky130_fd_sc_hd__maj3_1_72/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_515 sky130_fd_sc_hd__nand2_1_515/Y sky130_fd_sc_hd__xor2_1_275/B
+ sky130_fd_sc_hd__nor2_1_287/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_83 sky130_fd_sc_hd__maj3_1_84/X sky130_fd_sc_hd__maj3_1_83/X
+ sky130_fd_sc_hd__maj3_1_83/B sky130_fd_sc_hd__maj3_1_83/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_526 sky130_fd_sc_hd__nor2_1_295/B sky130_fd_sc_hd__nand2_1_526/B
+ sky130_fd_sc_hd__nor2_1_296/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__maj3_1_94 sky130_fd_sc_hd__maj3_1_95/X sky130_fd_sc_hd__maj3_1_94/X
+ sky130_fd_sc_hd__maj3_1_94/B sky130_fd_sc_hd__maj3_1_94/A VDD VSS VSS VDD sky130_fd_sc_hd__maj3_1
Xsky130_fd_sc_hd__nand2_1_537 sky130_fd_sc_hd__nand2_1_537/Y sky130_fd_sc_hd__nor2b_1_126/Y
+ sky130_fd_sc_hd__o21ai_1_463/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_548 sky130_fd_sc_hd__nand3_1_51/A sky130_fd_sc_hd__nand3_1_1/Y
+ sky130_fd_sc_hd__nor2_1_314/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_559 sky130_fd_sc_hd__nand2_1_559/Y sky130_fd_sc_hd__buf_4_60/A
+ sky130_fd_sc_hd__nand2_1_559/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nor2b_1_6 sky130_fd_sc_hd__ha_2_27/SUM sky130_fd_sc_hd__nor2b_1_6/Y
+ sky130_fd_sc_hd__or2_0_1/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2b_1
Xsky130_fd_sc_hd__clkinv_1_1106 sky130_fd_sc_hd__o22ai_1_436/B1 sky130_fd_sc_hd__fa_2_1305/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1106/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1117 sky130_fd_sc_hd__nor2_1_323/B sky130_fd_sc_hd__nor2_1_319/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1117/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_1128 sky130_fd_sc_hd__clkinv_4_37/A sky130_fd_sc_hd__buf_4_122/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_1128/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_300 VDD VSS sky130_fd_sc_hd__a22o_1_49/A1 sky130_fd_sc_hd__dfxtp_1_304/CLK
+ sky130_fd_sc_hd__and2_0_98/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_311 VDD VSS sky130_fd_sc_hd__a22o_1_38/A1 sky130_fd_sc_hd__dfxtp_1_313/CLK
+ sky130_fd_sc_hd__and2_0_87/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_322 VDD VSS sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__dfxtp_1_325/CLK
+ sky130_fd_sc_hd__and2_0_190/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_333 VDD VSS sky130_fd_sc_hd__a22o_2_9/B2 sky130_fd_sc_hd__dfxtp_1_360/CLK
+ sky130_fd_sc_hd__o21ai_1_25/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_344 VDD VSS sky130_fd_sc_hd__a22o_1_20/B2 sky130_fd_sc_hd__dfxtp_1_360/CLK
+ sky130_fd_sc_hd__ha_2_155/A VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_355 VDD VSS sky130_fd_sc_hd__ha_2_150/A sky130_fd_sc_hd__dfxtp_1_361/CLK
+ sky130_fd_sc_hd__o2bb2ai_1_5/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_366 VDD VSS sky130_fd_sc_hd__fa_2_1110/A sky130_fd_sc_hd__dfxtp_1_393/CLK
+ sky130_fd_sc_hd__and2_0_161/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_377 VDD VSS sky130_fd_sc_hd__nor2_2_10/B sky130_fd_sc_hd__dfxtp_1_393/CLK
+ sky130_fd_sc_hd__and2_0_105/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_388 VDD VSS sky130_fd_sc_hd__fa_2_1116/B sky130_fd_sc_hd__dfxtp_1_391/CLK
+ sky130_fd_sc_hd__and2_0_125/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_8 sky130_fd_sc_hd__nand3_1_8/C sky130_fd_sc_hd__nand2_1_8/B
+ sky130_fd_sc_hd__nand2_1_9/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_399 VDD VSS sky130_fd_sc_hd__fa_2_1035/A sky130_fd_sc_hd__dfxtp_1_424/CLK
+ sky130_fd_sc_hd__and2_0_153/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o31ai_1_11 sky130_fd_sc_hd__o31ai_1_11/Y sky130_fd_sc_hd__nor2_1_286/A
+ sky130_fd_sc_hd__o31ai_1_12/A2 sky130_fd_sc_hd__o31ai_1_12/A3 sky130_fd_sc_hd__o31ai_1_11/B1
+ VDD VSS VDD VSS sky130_fd_sc_hd__o31ai_1
Xsky130_fd_sc_hd__fa_2_205 sky130_fd_sc_hd__maj3_1_42/B sky130_fd_sc_hd__maj3_1_43/A
+ sky130_fd_sc_hd__fa_2_205/A sky130_fd_sc_hd__fa_2_205/B sky130_fd_sc_hd__fa_2_206/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_216 sky130_fd_sc_hd__fa_2_220/B sky130_fd_sc_hd__fa_2_216/SUM
+ sky130_fd_sc_hd__fa_2_216/A sky130_fd_sc_hd__fa_2_216/B sky130_fd_sc_hd__fa_2_216/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_227 sky130_fd_sc_hd__fa_2_231/B sky130_fd_sc_hd__fa_2_227/SUM
+ sky130_fd_sc_hd__fa_2_227/A sky130_fd_sc_hd__fa_2_227/B sky130_fd_sc_hd__fa_2_227/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_238 sky130_fd_sc_hd__fa_2_237/B sky130_fd_sc_hd__fa_2_232/B
+ sky130_fd_sc_hd__fa_2_280/B sky130_fd_sc_hd__fa_2_238/B sky130_fd_sc_hd__fa_2_238/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_249 sky130_fd_sc_hd__fa_2_246/A sky130_fd_sc_hd__fa_2_241/A
+ sky130_fd_sc_hd__fa_2_5/B sky130_fd_sc_hd__fa_2_15/B sky130_fd_sc_hd__fa_2_280/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_30 sky130_fd_sc_hd__maj3_1_29/B sky130_fd_sc_hd__fa_2_30/SUM
+ sky130_fd_sc_hd__fa_2_67/B sky130_fd_sc_hd__ha_2_93/A sky130_fd_sc_hd__ha_2_99/A
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_41 sky130_fd_sc_hd__maj3_1_22/B sky130_fd_sc_hd__maj3_1_23/A
+ sky130_fd_sc_hd__fa_2_41/A sky130_fd_sc_hd__fa_2_41/B sky130_fd_sc_hd__fa_2_42/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__and2_0_9 VSS VDD VDD VSS sky130_fd_sc_hd__and2_0_9/X sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__ha_2_4/SUM sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__fa_2_52 sky130_fd_sc_hd__fa_2_55/CIN sky130_fd_sc_hd__fa_2_50/B
+ sky130_fd_sc_hd__ha_2_97/B sky130_fd_sc_hd__fa_2_52/B sky130_fd_sc_hd__fa_2_52/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_63 sky130_fd_sc_hd__maj3_1_16/B sky130_fd_sc_hd__maj3_1_17/A
+ sky130_fd_sc_hd__fa_2_63/A sky130_fd_sc_hd__fa_2_63/B sky130_fd_sc_hd__fa_2_64/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_74 sky130_fd_sc_hd__fa_2_78/B sky130_fd_sc_hd__fa_2_74/SUM
+ sky130_fd_sc_hd__fa_2_74/A sky130_fd_sc_hd__fa_2_74/B sky130_fd_sc_hd__fa_2_74/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_85 sky130_fd_sc_hd__fa_2_89/B sky130_fd_sc_hd__fa_2_85/SUM
+ sky130_fd_sc_hd__fa_2_85/A sky130_fd_sc_hd__fa_2_85/B sky130_fd_sc_hd__fa_2_85/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_96 sky130_fd_sc_hd__fa_2_95/B sky130_fd_sc_hd__fa_2_90/B sky130_fd_sc_hd__fa_2_96/A
+ sky130_fd_sc_hd__fa_2_9/A sky130_fd_sc_hd__fa_2_96/CIN VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__buf_2_200 VDD VSS sky130_fd_sc_hd__buf_2_200/X sky130_fd_sc_hd__buf_2_200/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_211 VDD VSS sky130_fd_sc_hd__buf_2_211/X sky130_fd_sc_hd__buf_2_211/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_222 VDD VSS sky130_fd_sc_hd__buf_2_222/X sky130_fd_sc_hd__buf_2_222/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_233 VDD VSS sky130_fd_sc_hd__buf_2_233/X sky130_fd_sc_hd__buf_2_233/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_244 VDD VSS sky130_fd_sc_hd__buf_2_244/X sky130_fd_sc_hd__buf_2_244/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_255 VDD VSS sky130_fd_sc_hd__fa_2_1172/B sky130_fd_sc_hd__nor2_4_14/Y
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_266 VDD VSS sky130_fd_sc_hd__buf_2_266/X sky130_fd_sc_hd__buf_2_266/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_277 VDD VSS sky130_fd_sc_hd__nor4_1_0/B sky130_fd_sc_hd__buf_2_277/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_288 VDD VSS sky130_fd_sc_hd__buf_2_288/X sky130_fd_sc_hd__buf_2_288/A
+ VDD VSS sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dfxtp_1_1240 VDD VSS sky130_fd_sc_hd__fa_2_1269/A sky130_fd_sc_hd__clkinv_8_105/Y
+ sky130_fd_sc_hd__mux2_2_202/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1251 VDD VSS sky130_fd_sc_hd__nor3_1_40/C sky130_fd_sc_hd__clkinv_8_74/Y
+ sky130_fd_sc_hd__o21bai_1_4/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1262 VDD VSS sky130_fd_sc_hd__mux2_2_187/A0 sky130_fd_sc_hd__clkinv_8_78/Y
+ sky130_fd_sc_hd__o22ai_1_329/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1273 VDD VSS sky130_fd_sc_hd__mux2_2_216/A0 sky130_fd_sc_hd__clkinv_8_102/Y
+ sky130_fd_sc_hd__dfxtp_1_429/Q VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1284 VDD VSS sky130_fd_sc_hd__mux2_2_212/A0 sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__nor2_1_244/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1295 VDD VSS sky130_fd_sc_hd__mux2_2_182/A1 sky130_fd_sc_hd__clkinv_8_116/Y
+ sky130_fd_sc_hd__o22ai_1_340/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a21oi_1_13 sky130_fd_sc_hd__a21oi_1_14/Y sky130_fd_sc_hd__nor2_1_13/Y
+ sky130_fd_sc_hd__maj3_1_3/A sky130_fd_sc_hd__ha_2_157/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_24 sky130_fd_sc_hd__fa_2_952/A sky130_fd_sc_hd__nor2b_1_86/Y
+ sky130_fd_sc_hd__nand4_1_84/C sky130_fd_sc_hd__a21oi_1_24/A2 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_35 sky130_fd_sc_hd__nor2_1_41/Y sky130_fd_sc_hd__o22ai_1_68/Y
+ sky130_fd_sc_hd__a21oi_1_35/Y sky130_fd_sc_hd__fa_2_1038/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_46 sky130_fd_sc_hd__nor2_2_6/Y sky130_fd_sc_hd__o22ai_1_78/Y
+ sky130_fd_sc_hd__a21oi_1_46/Y sky130_fd_sc_hd__fa_2_1034/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_57 sky130_fd_sc_hd__nor2_2_6/Y sky130_fd_sc_hd__o22ai_1_89/Y
+ sky130_fd_sc_hd__a21oi_1_57/Y sky130_fd_sc_hd__a22o_1_67/A2 VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_68 sky130_fd_sc_hd__nand2_1_248/Y sky130_fd_sc_hd__nor2_1_51/Y
+ sky130_fd_sc_hd__xnor2_1_51/A sky130_fd_sc_hd__xnor2_1_49/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__fa_2_750 sky130_fd_sc_hd__fa_2_753/B sky130_fd_sc_hd__fa_2_748/B
+ sky130_fd_sc_hd__fa_2_829/A sky130_fd_sc_hd__fa_2_823/B sky130_fd_sc_hd__fa_2_750/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a21oi_1_79 sky130_fd_sc_hd__o21a_1_7/B1 sky130_fd_sc_hd__o21a_1_6/A1
+ sky130_fd_sc_hd__a21oi_1_79/Y sky130_fd_sc_hd__nor2_1_69/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__fa_2_761 sky130_fd_sc_hd__fa_2_764/CIN sky130_fd_sc_hd__fa_2_761/SUM
+ sky130_fd_sc_hd__fa_2_761/A sky130_fd_sc_hd__fa_2_761/B sky130_fd_sc_hd__fa_2_761/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_772 sky130_fd_sc_hd__maj3_1_140/B sky130_fd_sc_hd__maj3_1_141/A
+ sky130_fd_sc_hd__fa_2_772/A sky130_fd_sc_hd__fa_2_772/B sky130_fd_sc_hd__fa_2_773/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_783 sky130_fd_sc_hd__maj3_1_137/B sky130_fd_sc_hd__maj3_1_138/A
+ sky130_fd_sc_hd__fa_2_783/A sky130_fd_sc_hd__fa_2_783/B sky130_fd_sc_hd__fa_2_784/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_794 sky130_fd_sc_hd__fa_2_716/A sky130_fd_sc_hd__maj3_1_135/A
+ sky130_fd_sc_hd__fa_2_794/A sky130_fd_sc_hd__fa_2_794/B sky130_fd_sc_hd__fa_2_796/SUM
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nor3_1_5 sky130_fd_sc_hd__nor3_2_2/B sky130_fd_sc_hd__nor3_1_5/Y
+ sky130_fd_sc_hd__nor3_2_3/A sky130_fd_sc_hd__nor3_2_3/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__bufinv_16_2 sky130_fd_sc_hd__bufinv_8_3/A sky130_fd_sc_hd__buf_12_183/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__bufinv_16
Xsky130_fd_sc_hd__buf_6_20 VDD VSS sky130_fd_sc_hd__buf_6_20/X sky130_fd_sc_hd__inv_2_53/Y
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_31 VDD VSS sky130_fd_sc_hd__buf_6_31/X sky130_fd_sc_hd__buf_6_31/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_42 VDD VSS sky130_fd_sc_hd__buf_6_42/X sky130_fd_sc_hd__buf_6_42/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_53 VDD VSS sky130_fd_sc_hd__buf_6_53/X sky130_fd_sc_hd__buf_6_53/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_64 VDD VSS sky130_fd_sc_hd__buf_6_64/X sky130_fd_sc_hd__buf_6_64/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_75 VDD VSS sky130_fd_sc_hd__buf_6_75/X sky130_fd_sc_hd__buf_6_75/A
+ VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__buf_6_86 VDD VSS sky130_fd_sc_hd__buf_6_86/X rst_n VDD VSS sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__diode_2_11 sky130_fd_sc_hd__clkbuf_1_247/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_22 sky130_fd_sc_hd__buf_2_123/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_307 sky130_fd_sc_hd__nor2_1_190/A sky130_fd_sc_hd__o21a_1_35/A1
+ sky130_fd_sc_hd__a21oi_1_307/Y sky130_fd_sc_hd__nor2_1_190/B VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_33 sky130_fd_sc_hd__nand4_1_23/A VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_318 sky130_fd_sc_hd__or3_1_3/C sky130_fd_sc_hd__o21ai_1_330/Y
+ sky130_fd_sc_hd__a21oi_1_318/Y sky130_fd_sc_hd__nor2_1_203/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_44 sky130_fd_sc_hd__buf_2_80/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__a21oi_1_329 sky130_fd_sc_hd__nor2b_2_3/Y sky130_fd_sc_hd__o21ai_1_350/Y
+ sky130_fd_sc_hd__a21oi_1_329/Y sky130_fd_sc_hd__o21ai_1_359/Y VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__diode_2_55 sky130_fd_sc_hd__buf_2_100/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_66 sky130_fd_sc_hd__buf_2_81/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_77 sky130_fd_sc_hd__buf_8_63/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_88 sky130_fd_sc_hd__clkbuf_1_535/X VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_99 sky130_fd_sc_hd__inv_2_135/Y VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__nand2_1_301 sky130_fd_sc_hd__nand2_1_301/Y sky130_fd_sc_hd__nor2_1_105/B
+ sky130_fd_sc_hd__fa_2_1107/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_900 sky130_fd_sc_hd__nand2_1_424/B sky130_fd_sc_hd__fa_2_306/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_900/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_312 sky130_fd_sc_hd__o21a_1_13/B1 sky130_fd_sc_hd__fa_2_1058/A
+ sky130_fd_sc_hd__o21a_1_13/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_911 sky130_fd_sc_hd__nor2_1_185/B sky130_fd_sc_hd__fa_2_1186/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_911/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_323 sky130_fd_sc_hd__nand2_1_323/Y sky130_fd_sc_hd__nor2_4_13/Y
+ sky130_fd_sc_hd__fa_2_1065/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_922 sky130_fd_sc_hd__o21ai_1_371/B1 sky130_fd_sc_hd__nor2_1_219/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_922/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_270 sky130_fd_sc_hd__nand2_1_410/Y sky130_fd_sc_hd__nand2_1_409/Y
+ sky130_fd_sc_hd__o22ai_1_270/Y sky130_fd_sc_hd__o22ai_1_283/A1 sky130_fd_sc_hd__a21o_2_13/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_334 sky130_fd_sc_hd__nand2_1_334/Y sky130_fd_sc_hd__nand2_1_339/B
+ sky130_fd_sc_hd__xor2_1_88/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_933 sky130_fd_sc_hd__nor2_1_193/B sky130_fd_sc_hd__fa_2_1204/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_933/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__o22ai_1_281 sky130_fd_sc_hd__nand2_1_412/Y sky130_fd_sc_hd__nand2_1_411/Y
+ sky130_fd_sc_hd__o22ai_1_281/Y sky130_fd_sc_hd__o22ai_1_281/A1 sky130_fd_sc_hd__a21o_2_12/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__nand2_1_345 sky130_fd_sc_hd__o21a_1_20/B1 sky130_fd_sc_hd__fa_2_1132/A
+ sky130_fd_sc_hd__o21a_1_20/A1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__o22ai_1_292 sky130_fd_sc_hd__nand2_1_412/Y sky130_fd_sc_hd__nand2_1_411/Y
+ sky130_fd_sc_hd__o22ai_1_292/Y sky130_fd_sc_hd__o22ai_1_292/A1 sky130_fd_sc_hd__o21ai_1_337/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkinv_1_944 sky130_fd_sc_hd__nor2_2_17/B sky130_fd_sc_hd__nor2_4_18/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_944/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_356 sky130_fd_sc_hd__o32ai_1_2/B1 sky130_fd_sc_hd__o32ai_1_2/A3
+ sky130_fd_sc_hd__o21bai_1_2/A2 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_955 sky130_fd_sc_hd__o32ai_1_6/A2 sky130_fd_sc_hd__fa_2_1224/B
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_955/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_367 sky130_fd_sc_hd__o31ai_1_6/A2 sky130_fd_sc_hd__nand2_1_367/B
+ sky130_fd_sc_hd__a21o_2_6/B1 VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_966 sky130_fd_sc_hd__o22ai_1_340/A1 sky130_fd_sc_hd__nor2_1_252/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_966/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_378 sky130_fd_sc_hd__nand2_1_378/Y sky130_fd_sc_hd__nand2_1_387/B
+ sky130_fd_sc_hd__o21ai_1_294/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_977 sky130_fd_sc_hd__nor2_1_233/B sky130_fd_sc_hd__fa_2_1228/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_977/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_389 sky130_fd_sc_hd__nand2_1_389/Y sky130_fd_sc_hd__nor2b_1_105/Y
+ sky130_fd_sc_hd__o21ai_1_323/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_988 sky130_fd_sc_hd__o22ai_1_358/A1 sky130_fd_sc_hd__o21ai_1_406/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_988/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_999 sky130_fd_sc_hd__nor2_1_232/B sky130_fd_sc_hd__fa_2_1230/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_999/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_130 VDD VSS sky130_fd_sc_hd__dfxtp_1_130/Q sky130_fd_sc_hd__clkinv_8_8/Y
+ sky130_fd_sc_hd__and2_2_0/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_141 VDD VSS sky130_fd_sc_hd__buf_2_33/A sky130_fd_sc_hd__dfxtp_1_143/CLK
+ sky130_fd_sc_hd__nor2b_1_9/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_152 VDD VSS sky130_fd_sc_hd__ha_2_35/A sky130_fd_sc_hd__dfxtp_1_155/CLK
+ sky130_fd_sc_hd__and2_0_26/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_163 VDD VSS sky130_fd_sc_hd__ha_2_46/A sky130_fd_sc_hd__clkinv_8_14/Y
+ sky130_fd_sc_hd__nor2b_1_17/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_174 VDD VSS sky130_fd_sc_hd__ha_2_59/B sky130_fd_sc_hd__dfxtp_1_185/CLK
+ sky130_fd_sc_hd__and2_0_61/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_185 VDD VSS sky130_fd_sc_hd__xor2_1_5/B sky130_fd_sc_hd__dfxtp_1_185/CLK
+ sky130_fd_sc_hd__and2_0_59/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_196 VDD VSS sky130_fd_sc_hd__ha_2_60/A sky130_fd_sc_hd__dfxtp_1_197/CLK
+ sky130_fd_sc_hd__nor2b_1_30/Y VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a21boi_1_6 sky130_fd_sc_hd__a21boi_1_6/Y sky130_fd_sc_hd__nor2_2_17/Y
+ sky130_fd_sc_hd__a21oi_1_405/Y sky130_fd_sc_hd__fa_2_1255/A VDD VSS VDD VSS sky130_fd_sc_hd__a21boi_1
Xsky130_fd_sc_hd__o211ai_1_16 sky130_fd_sc_hd__o21ai_1_225/A2 sky130_fd_sc_hd__o21a_1_16/A2
+ sky130_fd_sc_hd__o211ai_1_16/Y sky130_fd_sc_hd__nand2_1_322/Y sky130_fd_sc_hd__nand2_1_323/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__fa_2_1240 sky130_fd_sc_hd__fa_2_1241/CIN sky130_fd_sc_hd__mux2_2_177/A0
+ sky130_fd_sc_hd__fa_2_1240/A sky130_fd_sc_hd__fa_2_1240/B sky130_fd_sc_hd__fa_2_1240/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o211ai_1_27 sky130_fd_sc_hd__nor2_1_172/A sky130_fd_sc_hd__a222oi_1_6/Y
+ sky130_fd_sc_hd__xor2_1_174/A sky130_fd_sc_hd__nand2_1_378/Y sky130_fd_sc_hd__a21oi_1_267/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__o211ai_1_38 sky130_fd_sc_hd__nor2_1_217/B sky130_fd_sc_hd__nor2_1_222/A
+ sky130_fd_sc_hd__xor2_1_218/A sky130_fd_sc_hd__nand2_1_429/Y sky130_fd_sc_hd__a21oi_1_325/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__fa_2_1251 sky130_fd_sc_hd__fa_2_1252/CIN sky130_fd_sc_hd__mux2_2_191/A1
+ sky130_fd_sc_hd__fa_2_1251/A sky130_fd_sc_hd__fa_2_1251/B sky130_fd_sc_hd__fa_2_1251/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o211ai_1_49 sky130_fd_sc_hd__nor2_1_265/A sky130_fd_sc_hd__nor2_1_259/B
+ sky130_fd_sc_hd__xor2_1_262/A sky130_fd_sc_hd__nand2_1_479/Y sky130_fd_sc_hd__nand2_1_480/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o211ai_1
Xsky130_fd_sc_hd__fa_2_1262 sky130_fd_sc_hd__fa_2_1263/CIN sky130_fd_sc_hd__mux2_2_217/A1
+ sky130_fd_sc_hd__fa_2_1262/A sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1262/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1273 sky130_fd_sc_hd__fa_2_1274/CIN sky130_fd_sc_hd__nand2_1_466/A
+ sky130_fd_sc_hd__fa_2_1273/A sky130_fd_sc_hd__nor2_8_1/Y sky130_fd_sc_hd__fa_2_1273/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1284 sky130_fd_sc_hd__fa_2_1285/CIN sky130_fd_sc_hd__mux2_2_240/A1
+ sky130_fd_sc_hd__fa_2_1284/A sky130_fd_sc_hd__fa_2_1284/B sky130_fd_sc_hd__fa_2_1284/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1295 sky130_fd_sc_hd__fa_2_1296/CIN sky130_fd_sc_hd__mux2_2_260/A1
+ sky130_fd_sc_hd__fa_2_1295/A sky130_fd_sc_hd__fa_2_1295/B sky130_fd_sc_hd__fa_2_1295/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_1070 VDD VSS sky130_fd_sc_hd__xor2_1_208/A sky130_fd_sc_hd__clkinv_8_70/Y
+ sky130_fd_sc_hd__mux2_2_124/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_1081 VDD VSS sky130_fd_sc_hd__fa_2_1183/A sky130_fd_sc_hd__clkinv_8_48/Y
+ sky130_fd_sc_hd__mux2_2_142/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21ai_1_90 VSS VDD sky130_fd_sc_hd__nor2_1_89/A sky130_fd_sc_hd__o22ai_1_90/A1
+ sky130_fd_sc_hd__a21oi_1_81/Y sky130_fd_sc_hd__o21ai_1_90/Y VDD VSS sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__dfxtp_1_1092 VDD VSS sky130_fd_sc_hd__fa_2_1211/A sky130_fd_sc_hd__clkinv_8_67/Y
+ sky130_fd_sc_hd__mux2_2_169/X VDD VSS sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o2bb2ai_1_10 sky130_fd_sc_hd__dfxtp_1_361/D sky130_fd_sc_hd__nor2_1_18/Y
+ sky130_fd_sc_hd__xor2_1_12/X sky130_fd_sc_hd__o21ai_1_31/A1 sky130_fd_sc_hd__a21oi_2_0/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__o2bb2ai_1_21 sky130_fd_sc_hd__dfxtp_1_562/D sky130_fd_sc_hd__a21o_2_2/A2
+ sky130_fd_sc_hd__dfxtp_1_562/Q sky130_fd_sc_hd__nor4_1_5/C sky130_fd_sc_hd__nand3_1_46/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__o2bb2ai_1_32 sky130_fd_sc_hd__o2bb2ai_1_32/Y sky130_fd_sc_hd__nor2_1_141/A
+ sky130_fd_sc_hd__nor2_1_141/B sky130_fd_sc_hd__nor2_1_141/B sky130_fd_sc_hd__nor2_1_141/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2ai_1
Xsky130_fd_sc_hd__fa_2_580 sky130_fd_sc_hd__fa_2_579/CIN sky130_fd_sc_hd__and2_0_98/A
+ sky130_fd_sc_hd__fa_2_580/A sky130_fd_sc_hd__fa_2_580/B sky130_fd_sc_hd__fa_2_580/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_591 sky130_fd_sc_hd__fa_2_592/B sky130_fd_sc_hd__fa_2_591/SUM
+ sky130_fd_sc_hd__fa_2_689/B sky130_fd_sc_hd__ha_2_128/A sky130_fd_sc_hd__fa_2_591/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__clkinv_1_207 sky130_fd_sc_hd__buf_8_217/A sky130_fd_sc_hd__clkinv_1_207/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_207/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_218 sky130_fd_sc_hd__clkinv_1_219/A sky130_fd_sc_hd__a22o_1_23/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_218/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkinv_1_229 sky130_fd_sc_hd__inv_2_121/A sky130_fd_sc_hd__buf_2_160/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_229/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a21oi_1_104 sky130_fd_sc_hd__a21o_2_3/A2 sky130_fd_sc_hd__o22ai_1_113/Y
+ sky130_fd_sc_hd__a21oi_1_104/Y sky130_fd_sc_hd__fa_2_973/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_115 sky130_fd_sc_hd__nor2_2_8/Y sky130_fd_sc_hd__o22ai_1_123/Y
+ sky130_fd_sc_hd__a21oi_1_115/Y sky130_fd_sc_hd__fa_2_1006/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_126 sky130_fd_sc_hd__nor2_4_10/Y sky130_fd_sc_hd__a22o_1_69/X
+ sky130_fd_sc_hd__a21oi_1_126/Y sky130_fd_sc_hd__fa_2_994/A VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a21oi_1_137 sky130_fd_sc_hd__nor2_2_10/Y sky130_fd_sc_hd__o22ai_1_137/Y
+ sky130_fd_sc_hd__a21oi_1_137/Y sky130_fd_sc_hd__fa_2_1109/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nor2_1_301 sky130_fd_sc_hd__nor2_1_301/B sky130_fd_sc_hd__nor2_1_301/Y
+ sky130_fd_sc_hd__nor2_1_310/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a21oi_1_148 sky130_fd_sc_hd__nor2_2_10/Y sky130_fd_sc_hd__o22ai_1_148/Y
+ sky130_fd_sc_hd__a21oi_1_148/Y sky130_fd_sc_hd__fa_2_1120/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__nor2_1_312 sky130_fd_sc_hd__nor2_1_314/B sky130_fd_sc_hd__nor2_1_312/Y
+ sky130_fd_sc_hd__nor2_1_315/B VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_323 sky130_fd_sc_hd__nor2_1_323/B sky130_fd_sc_hd__or2_0_13/A
+ sky130_fd_sc_hd__nor2_1_323/A VDD VSS VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__a21oi_1_159 sky130_fd_sc_hd__nor2_2_11/Y sky130_fd_sc_hd__o22ai_1_158/Y
+ sky130_fd_sc_hd__a21oi_1_159/Y sky130_fd_sc_hd__fa_2_1116/SUM VDD VSS VDD VSS sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__a22oi_1_400 sky130_fd_sc_hd__a22oi_1_400/B1 sky130_fd_sc_hd__nor3_1_41/B
+ sky130_fd_sc_hd__fa_2_1291/A sky130_fd_sc_hd__fa_2_1292/A sky130_fd_sc_hd__a22oi_1_400/Y
+ VDD VSS VDD VSS sky130_fd_sc_hd__a22oi_1
Xsky130_fd_sc_hd__clkbuf_8_0 sky130_fd_sc_hd__clkbuf_8_0/X sky130_fd_sc_hd__buf_2_39/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkbuf_8
Xsky130_fd_sc_hd__nand2_1_120 sky130_fd_sc_hd__nand2_1_120/Y sky130_fd_sc_hd__fa_2_703/SUM
+ sky130_fd_sc_hd__and2_0_235/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_131 sky130_fd_sc_hd__nand2_1_131/Y sky130_fd_sc_hd__nand2_1_132/Y
+ sky130_fd_sc_hd__buf_2_264/X VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_730 sky130_fd_sc_hd__o22ai_1_196/B1 sky130_fd_sc_hd__o21ai_1_254/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_730/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_142 sky130_fd_sc_hd__nand2_1_142/Y sky130_fd_sc_hd__fa_2_714/SUM
+ sky130_fd_sc_hd__inv_4_1/Y VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_741 sky130_fd_sc_hd__o22ai_1_197/B2 sky130_fd_sc_hd__fa_2_1079/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_741/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_153 sky130_fd_sc_hd__fa_2_97/A sky130_fd_sc_hd__fa_2_76/B
+ sky130_fd_sc_hd__fa_2_80/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_752 sky130_fd_sc_hd__nor2_1_140/B sky130_fd_sc_hd__xor2_1_88/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_752/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_164 sky130_fd_sc_hd__fa_2_266/CIN sky130_fd_sc_hd__fa_2_238/B
+ sky130_fd_sc_hd__fa_2_5/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_763 sky130_fd_sc_hd__ha_2_195/B sky130_fd_sc_hd__fa_2_1112/SUM
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_763/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_175 sky130_fd_sc_hd__fa_2_320/A sky130_fd_sc_hd__fa_2_416/B
+ sky130_fd_sc_hd__ha_2_115/A VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_774 sky130_fd_sc_hd__nand2_1_333/B sky130_fd_sc_hd__nand2_2_6/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_774/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_186 sky130_fd_sc_hd__fa_2_621/B sky130_fd_sc_hd__ha_2_130/A
+ sky130_fd_sc_hd__ha_2_132/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_785 sky130_fd_sc_hd__nor2_1_172/A sky130_fd_sc_hd__nor2b_1_105/Y
+ VDD VSS VSS VDD VSS sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__nand2_1_197 sky130_fd_sc_hd__fa_2_787/A sky130_fd_sc_hd__fa_2_826/A
+ sky130_fd_sc_hd__fa_2_823/B VDD VSS VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_796 sky130_fd_sc_hd__o31ai_1_6/B1 sky130_fd_sc_hd__dfxtp_1_987/D
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_1_796/w_84_21# sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__xor2_1_2 sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__xor2_1_2/X
+ sky130_fd_sc_hd__xor2_1_2/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nand3_2_3 sky130_fd_sc_hd__nor2_4_2/Y sky130_fd_sc_hd__nand3_2_3/Y
+ sky130_fd_sc_hd__nand3_2_3/B sky130_fd_sc_hd__nand3_2_4/B VSS VDD VSS VDD sky130_fd_sc_hd__nand3_2
Xsky130_fd_sc_hd__clkinv_8_0 sky130_fd_sc_hd__clkinv_8_0/Y sky130_fd_sc_hd__clkinv_8_0/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_8_0/w_189_21# sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__xor2_1_17 sky130_fd_sc_hd__maj3_1_0/A sky130_fd_sc_hd__xor2_1_17/X
+ sky130_fd_sc_hd__xor2_1_17/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_28 sky130_fd_sc_hd__xor2_1_28/B sky130_fd_sc_hd__xor2_1_28/X
+ sky130_fd_sc_hd__or4_1_2/B VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_39 sky130_fd_sc_hd__fa_2_970/A sky130_fd_sc_hd__fa_2_988/B
+ sky130_fd_sc_hd__xor2_1_39/A VSS VDD VDD VSS sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__nor3_1_30 sky130_fd_sc_hd__nor3_1_31/C sky130_fd_sc_hd__nor3_1_30/Y
+ sky130_fd_sc_hd__or4_1_2/D sky130_fd_sc_hd__or4_1_2/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_41 sky130_fd_sc_hd__nor3_1_41/C sky130_fd_sc_hd__nor3_1_41/Y
+ sky130_fd_sc_hd__nor3_1_41/A sky130_fd_sc_hd__nor3_1_41/B VDD VSS VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__a21o_2_7 sky130_fd_sc_hd__a21o_2_7/X sky130_fd_sc_hd__a21o_2_7/B1
+ sky130_fd_sc_hd__a21o_2_7/A1 sky130_fd_sc_hd__a21o_2_7/A2 VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
Xsky130_fd_sc_hd__fa_2_1070 sky130_fd_sc_hd__fa_2_1071/CIN sky130_fd_sc_hd__and2_0_304/A
+ sky130_fd_sc_hd__fa_2_1070/A sky130_fd_sc_hd__fa_2_1070/B sky130_fd_sc_hd__fa_2_1070/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1081 sky130_fd_sc_hd__fa_2_1082/CIN sky130_fd_sc_hd__mux2_2_60/A0
+ sky130_fd_sc_hd__fa_2_1081/A sky130_fd_sc_hd__fa_2_1081/B sky130_fd_sc_hd__fa_2_1081/CIN
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_1092 sky130_fd_sc_hd__fa_2_1093/CIN sky130_fd_sc_hd__and2_0_294/A
+ sky130_fd_sc_hd__xor2_1_99/B sky130_fd_sc_hd__fa_2_1092/B sky130_fd_sc_hd__xor2_1_99/B
+ VSS VDD VDD VSS sky130_fd_sc_hd__fa_2
.ends

