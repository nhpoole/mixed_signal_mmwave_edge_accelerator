magic
tech sky130A
magscale 1 2
timestamp 1623661481
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 30 -17 64 17
<< locali >>
rect 103 333 169 493
rect 271 333 337 493
rect 471 333 537 493
rect 719 333 785 493
rect 103 289 785 333
rect 22 215 169 255
rect 214 215 340 255
rect 447 215 616 255
rect 674 211 785 289
rect 833 215 899 255
rect 719 127 785 211
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 18 299 69 527
rect 203 367 237 527
rect 371 367 437 527
rect 599 367 665 527
rect 819 289 885 527
rect 18 147 237 181
rect 18 51 85 147
rect 119 17 153 109
rect 187 93 237 147
rect 271 127 617 181
rect 651 93 685 177
rect 819 93 885 181
rect 187 51 425 93
rect 463 51 885 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 833 215 899 255 6 A
port 1 nsew signal input
rlabel locali s 447 215 616 255 6 B
port 2 nsew signal input
rlabel locali s 214 215 340 255 6 C
port 3 nsew signal input
rlabel locali s 22 215 169 255 6 D
port 4 nsew signal input
rlabel locali s 719 333 785 493 6 Y
port 5 nsew signal output
rlabel locali s 719 127 785 211 6 Y
port 5 nsew signal output
rlabel locali s 674 211 785 289 6 Y
port 5 nsew signal output
rlabel locali s 471 333 537 493 6 Y
port 5 nsew signal output
rlabel locali s 271 333 337 493 6 Y
port 5 nsew signal output
rlabel locali s 103 333 169 493 6 Y
port 5 nsew signal output
rlabel locali s 103 289 785 333 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 920 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 17 8 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 958 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
