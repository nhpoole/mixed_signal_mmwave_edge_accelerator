magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< pwell >>
rect -26 -26 392 362
<< scnmos >>
rect 60 0 90 336
rect 168 0 198 336
rect 276 0 306 336
<< ndiff >>
rect 0 0 60 336
rect 90 0 168 336
rect 198 0 276 336
rect 306 0 366 336
<< poly >>
rect 60 362 306 392
rect 60 336 90 362
rect 168 336 198 362
rect 276 336 306 362
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
<< locali >>
rect 112 235 358 269
rect 8 135 42 201
rect 112 168 146 235
rect 220 135 254 201
rect 324 168 358 235
use contact_11  contact_11_0
timestamp 1624494425
transform 1 0 316 0 1 135
box -26 -22 76 88
use contact_11  contact_11_1
timestamp 1624494425
transform 1 0 212 0 1 135
box -26 -22 76 88
use contact_11  contact_11_2
timestamp 1624494425
transform 1 0 104 0 1 135
box -26 -22 76 88
use contact_11  contact_11_3
timestamp 1624494425
transform 1 0 0 0 1 135
box -26 -22 76 88
<< labels >>
rlabel poly s 183 377 183 377 4 G
rlabel locali s 25 168 25 168 4 S
rlabel locali s 237 168 237 168 4 S
rlabel locali s 235 252 235 252 4 D
<< properties >>
string FIXED_BBOX -25 -26 391 392
<< end >>
