magic
tech sky130A
magscale 1 2
timestamp 1622760105
<< nwell >>
rect -398 -7578 12658 2958
<< pwell >>
rect -398 -10858 12658 -7742
<< nmos >>
rect 4956 -8860 5356 -8460
rect 5414 -8860 5814 -8460
rect 5872 -8860 6272 -8460
rect 6330 -8860 6730 -8460
rect 6788 -8860 7188 -8460
rect 7246 -8860 7646 -8460
rect 4956 -9660 5356 -9260
rect 5414 -9660 5814 -9260
rect 5872 -9660 6272 -9260
rect 6330 -9660 6730 -9260
rect 6788 -9660 7188 -9260
rect 7246 -9660 7646 -9260
<< pmos >>
rect 232 304 1032 1504
rect 1090 304 1890 1504
rect 1948 304 2748 1504
rect 2806 304 3606 1504
rect 3664 304 4464 1504
rect 4522 304 5322 1504
rect 5380 304 6180 1504
rect 6238 304 7038 1504
rect 7096 304 7896 1504
rect 7954 304 8754 1504
rect 8812 304 9612 1504
rect 9670 304 10470 1504
rect 10528 304 11328 1504
rect 11386 304 12186 1504
rect 232 -1436 1032 -236
rect 1090 -1436 1890 -236
rect 1948 -1436 2748 -236
rect 2806 -1436 3606 -236
rect 3664 -1436 4464 -236
rect 4522 -1436 5322 -236
rect 5380 -1436 6180 -236
rect 6238 -1436 7038 -236
rect 7096 -1436 7896 -236
rect 7954 -1436 8754 -236
rect 8812 -1436 9612 -236
rect 9670 -1436 10470 -236
rect 10528 -1436 11328 -236
rect 11386 -1436 12186 -236
rect 232 -3176 1032 -1976
rect 1090 -3176 1890 -1976
rect 1948 -3176 2748 -1976
rect 2806 -3176 3606 -1976
rect 3664 -3176 4464 -1976
rect 4522 -3176 5322 -1976
rect 5380 -3176 6180 -1976
rect 6238 -3176 7038 -1976
rect 7096 -3176 7896 -1976
rect 7954 -3176 8754 -1976
rect 8812 -3176 9612 -1976
rect 9670 -3176 10470 -1976
rect 10528 -3176 11328 -1976
rect 11386 -3176 12186 -1976
rect 232 -4916 1032 -3716
rect 1090 -4916 1890 -3716
rect 1948 -4916 2748 -3716
rect 2806 -4916 3606 -3716
rect 3664 -4916 4464 -3716
rect 4522 -4916 5322 -3716
rect 5380 -4916 6180 -3716
rect 6238 -4916 7038 -3716
rect 7096 -4916 7896 -3716
rect 7954 -4916 8754 -3716
rect 8812 -4916 9612 -3716
rect 9670 -4916 10470 -3716
rect 10528 -4916 11328 -3716
rect 11386 -4916 12186 -3716
rect 232 -6656 1032 -5456
rect 1090 -6656 1890 -5456
rect 1948 -6656 2748 -5456
rect 2806 -6656 3606 -5456
rect 3664 -6656 4464 -5456
rect 4522 -6656 5322 -5456
rect 5380 -6656 6180 -5456
rect 6238 -6656 7038 -5456
rect 7096 -6656 7896 -5456
rect 7954 -6656 8754 -5456
rect 8812 -6656 9612 -5456
rect 9670 -6656 10470 -5456
rect 10528 -6656 11328 -5456
rect 11386 -6656 12186 -5456
<< ndiff >>
rect 4898 -8472 4956 -8460
rect 4898 -8848 4910 -8472
rect 4944 -8848 4956 -8472
rect 4898 -8860 4956 -8848
rect 5356 -8472 5414 -8460
rect 5356 -8848 5368 -8472
rect 5402 -8848 5414 -8472
rect 5356 -8860 5414 -8848
rect 5814 -8472 5872 -8460
rect 5814 -8848 5826 -8472
rect 5860 -8848 5872 -8472
rect 5814 -8860 5872 -8848
rect 6272 -8472 6330 -8460
rect 6272 -8848 6284 -8472
rect 6318 -8848 6330 -8472
rect 6272 -8860 6330 -8848
rect 6730 -8472 6788 -8460
rect 6730 -8848 6742 -8472
rect 6776 -8848 6788 -8472
rect 6730 -8860 6788 -8848
rect 7188 -8472 7246 -8460
rect 7188 -8848 7200 -8472
rect 7234 -8848 7246 -8472
rect 7188 -8860 7246 -8848
rect 7646 -8472 7704 -8460
rect 7646 -8848 7658 -8472
rect 7692 -8848 7704 -8472
rect 7646 -8860 7704 -8848
rect 4898 -9272 4956 -9260
rect 4898 -9648 4910 -9272
rect 4944 -9648 4956 -9272
rect 4898 -9660 4956 -9648
rect 5356 -9272 5414 -9260
rect 5356 -9648 5368 -9272
rect 5402 -9648 5414 -9272
rect 5356 -9660 5414 -9648
rect 5814 -9272 5872 -9260
rect 5814 -9648 5826 -9272
rect 5860 -9648 5872 -9272
rect 5814 -9660 5872 -9648
rect 6272 -9272 6330 -9260
rect 6272 -9648 6284 -9272
rect 6318 -9648 6330 -9272
rect 6272 -9660 6330 -9648
rect 6730 -9272 6788 -9260
rect 6730 -9648 6742 -9272
rect 6776 -9648 6788 -9272
rect 6730 -9660 6788 -9648
rect 7188 -9272 7246 -9260
rect 7188 -9648 7200 -9272
rect 7234 -9648 7246 -9272
rect 7188 -9660 7246 -9648
rect 7646 -9272 7704 -9260
rect 7646 -9648 7658 -9272
rect 7692 -9648 7704 -9272
rect 7646 -9660 7704 -9648
<< pdiff >>
rect 174 1492 232 1504
rect 174 316 186 1492
rect 220 316 232 1492
rect 174 304 232 316
rect 1032 1492 1090 1504
rect 1032 316 1044 1492
rect 1078 316 1090 1492
rect 1032 304 1090 316
rect 1890 1492 1948 1504
rect 1890 316 1902 1492
rect 1936 316 1948 1492
rect 1890 304 1948 316
rect 2748 1492 2806 1504
rect 2748 316 2760 1492
rect 2794 316 2806 1492
rect 2748 304 2806 316
rect 3606 1492 3664 1504
rect 3606 316 3618 1492
rect 3652 316 3664 1492
rect 3606 304 3664 316
rect 4464 1492 4522 1504
rect 4464 316 4476 1492
rect 4510 316 4522 1492
rect 4464 304 4522 316
rect 5322 1492 5380 1504
rect 5322 316 5334 1492
rect 5368 316 5380 1492
rect 5322 304 5380 316
rect 6180 1492 6238 1504
rect 6180 316 6192 1492
rect 6226 316 6238 1492
rect 6180 304 6238 316
rect 7038 1492 7096 1504
rect 7038 316 7050 1492
rect 7084 316 7096 1492
rect 7038 304 7096 316
rect 7896 1492 7954 1504
rect 7896 316 7908 1492
rect 7942 316 7954 1492
rect 7896 304 7954 316
rect 8754 1492 8812 1504
rect 8754 316 8766 1492
rect 8800 316 8812 1492
rect 8754 304 8812 316
rect 9612 1492 9670 1504
rect 9612 316 9624 1492
rect 9658 316 9670 1492
rect 9612 304 9670 316
rect 10470 1492 10528 1504
rect 10470 316 10482 1492
rect 10516 316 10528 1492
rect 10470 304 10528 316
rect 11328 1492 11386 1504
rect 11328 316 11340 1492
rect 11374 316 11386 1492
rect 11328 304 11386 316
rect 12186 1492 12244 1504
rect 12186 316 12198 1492
rect 12232 316 12244 1492
rect 12186 304 12244 316
rect 174 -248 232 -236
rect 174 -1424 186 -248
rect 220 -1424 232 -248
rect 174 -1436 232 -1424
rect 1032 -248 1090 -236
rect 1032 -1424 1044 -248
rect 1078 -1424 1090 -248
rect 1032 -1436 1090 -1424
rect 1890 -248 1948 -236
rect 1890 -1424 1902 -248
rect 1936 -1424 1948 -248
rect 1890 -1436 1948 -1424
rect 2748 -248 2806 -236
rect 2748 -1424 2760 -248
rect 2794 -1424 2806 -248
rect 2748 -1436 2806 -1424
rect 3606 -248 3664 -236
rect 3606 -1424 3618 -248
rect 3652 -1424 3664 -248
rect 3606 -1436 3664 -1424
rect 4464 -248 4522 -236
rect 4464 -1424 4476 -248
rect 4510 -1424 4522 -248
rect 4464 -1436 4522 -1424
rect 5322 -248 5380 -236
rect 5322 -1424 5334 -248
rect 5368 -1424 5380 -248
rect 5322 -1436 5380 -1424
rect 6180 -248 6238 -236
rect 6180 -1424 6192 -248
rect 6226 -1424 6238 -248
rect 6180 -1436 6238 -1424
rect 7038 -248 7096 -236
rect 7038 -1424 7050 -248
rect 7084 -1424 7096 -248
rect 7038 -1436 7096 -1424
rect 7896 -248 7954 -236
rect 7896 -1424 7908 -248
rect 7942 -1424 7954 -248
rect 7896 -1436 7954 -1424
rect 8754 -248 8812 -236
rect 8754 -1424 8766 -248
rect 8800 -1424 8812 -248
rect 8754 -1436 8812 -1424
rect 9612 -248 9670 -236
rect 9612 -1424 9624 -248
rect 9658 -1424 9670 -248
rect 9612 -1436 9670 -1424
rect 10470 -248 10528 -236
rect 10470 -1424 10482 -248
rect 10516 -1424 10528 -248
rect 10470 -1436 10528 -1424
rect 11328 -248 11386 -236
rect 11328 -1424 11340 -248
rect 11374 -1424 11386 -248
rect 11328 -1436 11386 -1424
rect 12186 -248 12244 -236
rect 12186 -1424 12198 -248
rect 12232 -1424 12244 -248
rect 12186 -1436 12244 -1424
rect 174 -1988 232 -1976
rect 174 -3164 186 -1988
rect 220 -3164 232 -1988
rect 174 -3176 232 -3164
rect 1032 -1988 1090 -1976
rect 1032 -3164 1044 -1988
rect 1078 -3164 1090 -1988
rect 1032 -3176 1090 -3164
rect 1890 -1988 1948 -1976
rect 1890 -3164 1902 -1988
rect 1936 -3164 1948 -1988
rect 1890 -3176 1948 -3164
rect 2748 -1988 2806 -1976
rect 2748 -3164 2760 -1988
rect 2794 -3164 2806 -1988
rect 2748 -3176 2806 -3164
rect 3606 -1988 3664 -1976
rect 3606 -3164 3618 -1988
rect 3652 -3164 3664 -1988
rect 3606 -3176 3664 -3164
rect 4464 -1988 4522 -1976
rect 4464 -3164 4476 -1988
rect 4510 -3164 4522 -1988
rect 4464 -3176 4522 -3164
rect 5322 -1988 5380 -1976
rect 5322 -3164 5334 -1988
rect 5368 -3164 5380 -1988
rect 5322 -3176 5380 -3164
rect 6180 -1988 6238 -1976
rect 6180 -3164 6192 -1988
rect 6226 -3164 6238 -1988
rect 6180 -3176 6238 -3164
rect 7038 -1988 7096 -1976
rect 7038 -3164 7050 -1988
rect 7084 -3164 7096 -1988
rect 7038 -3176 7096 -3164
rect 7896 -1988 7954 -1976
rect 7896 -3164 7908 -1988
rect 7942 -3164 7954 -1988
rect 7896 -3176 7954 -3164
rect 8754 -1988 8812 -1976
rect 8754 -3164 8766 -1988
rect 8800 -3164 8812 -1988
rect 8754 -3176 8812 -3164
rect 9612 -1988 9670 -1976
rect 9612 -3164 9624 -1988
rect 9658 -3164 9670 -1988
rect 9612 -3176 9670 -3164
rect 10470 -1988 10528 -1976
rect 10470 -3164 10482 -1988
rect 10516 -3164 10528 -1988
rect 10470 -3176 10528 -3164
rect 11328 -1988 11386 -1976
rect 11328 -3164 11340 -1988
rect 11374 -3164 11386 -1988
rect 11328 -3176 11386 -3164
rect 12186 -1988 12244 -1976
rect 12186 -3164 12198 -1988
rect 12232 -3164 12244 -1988
rect 12186 -3176 12244 -3164
rect 174 -3728 232 -3716
rect 174 -4904 186 -3728
rect 220 -4904 232 -3728
rect 174 -4916 232 -4904
rect 1032 -3728 1090 -3716
rect 1032 -4904 1044 -3728
rect 1078 -4904 1090 -3728
rect 1032 -4916 1090 -4904
rect 1890 -3728 1948 -3716
rect 1890 -4904 1902 -3728
rect 1936 -4904 1948 -3728
rect 1890 -4916 1948 -4904
rect 2748 -3728 2806 -3716
rect 2748 -4904 2760 -3728
rect 2794 -4904 2806 -3728
rect 2748 -4916 2806 -4904
rect 3606 -3728 3664 -3716
rect 3606 -4904 3618 -3728
rect 3652 -4904 3664 -3728
rect 3606 -4916 3664 -4904
rect 4464 -3728 4522 -3716
rect 4464 -4904 4476 -3728
rect 4510 -4904 4522 -3728
rect 4464 -4916 4522 -4904
rect 5322 -3728 5380 -3716
rect 5322 -4904 5334 -3728
rect 5368 -4904 5380 -3728
rect 5322 -4916 5380 -4904
rect 6180 -3728 6238 -3716
rect 6180 -4904 6192 -3728
rect 6226 -4904 6238 -3728
rect 6180 -4916 6238 -4904
rect 7038 -3728 7096 -3716
rect 7038 -4904 7050 -3728
rect 7084 -4904 7096 -3728
rect 7038 -4916 7096 -4904
rect 7896 -3728 7954 -3716
rect 7896 -4904 7908 -3728
rect 7942 -4904 7954 -3728
rect 7896 -4916 7954 -4904
rect 8754 -3728 8812 -3716
rect 8754 -4904 8766 -3728
rect 8800 -4904 8812 -3728
rect 8754 -4916 8812 -4904
rect 9612 -3728 9670 -3716
rect 9612 -4904 9624 -3728
rect 9658 -4904 9670 -3728
rect 9612 -4916 9670 -4904
rect 10470 -3728 10528 -3716
rect 10470 -4904 10482 -3728
rect 10516 -4904 10528 -3728
rect 10470 -4916 10528 -4904
rect 11328 -3728 11386 -3716
rect 11328 -4904 11340 -3728
rect 11374 -4904 11386 -3728
rect 11328 -4916 11386 -4904
rect 12186 -3728 12244 -3716
rect 12186 -4904 12198 -3728
rect 12232 -4904 12244 -3728
rect 12186 -4916 12244 -4904
rect 174 -5468 232 -5456
rect 174 -6644 186 -5468
rect 220 -6644 232 -5468
rect 174 -6656 232 -6644
rect 1032 -5468 1090 -5456
rect 1032 -6644 1044 -5468
rect 1078 -6644 1090 -5468
rect 1032 -6656 1090 -6644
rect 1890 -5468 1948 -5456
rect 1890 -6644 1902 -5468
rect 1936 -6644 1948 -5468
rect 1890 -6656 1948 -6644
rect 2748 -5468 2806 -5456
rect 2748 -6644 2760 -5468
rect 2794 -6644 2806 -5468
rect 2748 -6656 2806 -6644
rect 3606 -5468 3664 -5456
rect 3606 -6644 3618 -5468
rect 3652 -6644 3664 -5468
rect 3606 -6656 3664 -6644
rect 4464 -5468 4522 -5456
rect 4464 -6644 4476 -5468
rect 4510 -6644 4522 -5468
rect 4464 -6656 4522 -6644
rect 5322 -5468 5380 -5456
rect 5322 -6644 5334 -5468
rect 5368 -6644 5380 -5468
rect 5322 -6656 5380 -6644
rect 6180 -5468 6238 -5456
rect 6180 -6644 6192 -5468
rect 6226 -6644 6238 -5468
rect 6180 -6656 6238 -6644
rect 7038 -5468 7096 -5456
rect 7038 -6644 7050 -5468
rect 7084 -6644 7096 -5468
rect 7038 -6656 7096 -6644
rect 7896 -5468 7954 -5456
rect 7896 -6644 7908 -5468
rect 7942 -6644 7954 -5468
rect 7896 -6656 7954 -6644
rect 8754 -5468 8812 -5456
rect 8754 -6644 8766 -5468
rect 8800 -6644 8812 -5468
rect 8754 -6656 8812 -6644
rect 9612 -5468 9670 -5456
rect 9612 -6644 9624 -5468
rect 9658 -6644 9670 -5468
rect 9612 -6656 9670 -6644
rect 10470 -5468 10528 -5456
rect 10470 -6644 10482 -5468
rect 10516 -6644 10528 -5468
rect 10470 -6656 10528 -6644
rect 11328 -5468 11386 -5456
rect 11328 -6644 11340 -5468
rect 11374 -6644 11386 -5468
rect 11328 -6656 11386 -6644
rect 12186 -5468 12244 -5456
rect 12186 -6644 12198 -5468
rect 12232 -6644 12244 -5468
rect 12186 -6656 12244 -6644
<< ndiffc >>
rect 4910 -8848 4944 -8472
rect 5368 -8848 5402 -8472
rect 5826 -8848 5860 -8472
rect 6284 -8848 6318 -8472
rect 6742 -8848 6776 -8472
rect 7200 -8848 7234 -8472
rect 7658 -8848 7692 -8472
rect 4910 -9648 4944 -9272
rect 5368 -9648 5402 -9272
rect 5826 -9648 5860 -9272
rect 6284 -9648 6318 -9272
rect 6742 -9648 6776 -9272
rect 7200 -9648 7234 -9272
rect 7658 -9648 7692 -9272
<< pdiffc >>
rect 186 316 220 1492
rect 1044 316 1078 1492
rect 1902 316 1936 1492
rect 2760 316 2794 1492
rect 3618 316 3652 1492
rect 4476 316 4510 1492
rect 5334 316 5368 1492
rect 6192 316 6226 1492
rect 7050 316 7084 1492
rect 7908 316 7942 1492
rect 8766 316 8800 1492
rect 9624 316 9658 1492
rect 10482 316 10516 1492
rect 11340 316 11374 1492
rect 12198 316 12232 1492
rect 186 -1424 220 -248
rect 1044 -1424 1078 -248
rect 1902 -1424 1936 -248
rect 2760 -1424 2794 -248
rect 3618 -1424 3652 -248
rect 4476 -1424 4510 -248
rect 5334 -1424 5368 -248
rect 6192 -1424 6226 -248
rect 7050 -1424 7084 -248
rect 7908 -1424 7942 -248
rect 8766 -1424 8800 -248
rect 9624 -1424 9658 -248
rect 10482 -1424 10516 -248
rect 11340 -1424 11374 -248
rect 12198 -1424 12232 -248
rect 186 -3164 220 -1988
rect 1044 -3164 1078 -1988
rect 1902 -3164 1936 -1988
rect 2760 -3164 2794 -1988
rect 3618 -3164 3652 -1988
rect 4476 -3164 4510 -1988
rect 5334 -3164 5368 -1988
rect 6192 -3164 6226 -1988
rect 7050 -3164 7084 -1988
rect 7908 -3164 7942 -1988
rect 8766 -3164 8800 -1988
rect 9624 -3164 9658 -1988
rect 10482 -3164 10516 -1988
rect 11340 -3164 11374 -1988
rect 12198 -3164 12232 -1988
rect 186 -4904 220 -3728
rect 1044 -4904 1078 -3728
rect 1902 -4904 1936 -3728
rect 2760 -4904 2794 -3728
rect 3618 -4904 3652 -3728
rect 4476 -4904 4510 -3728
rect 5334 -4904 5368 -3728
rect 6192 -4904 6226 -3728
rect 7050 -4904 7084 -3728
rect 7908 -4904 7942 -3728
rect 8766 -4904 8800 -3728
rect 9624 -4904 9658 -3728
rect 10482 -4904 10516 -3728
rect 11340 -4904 11374 -3728
rect 12198 -4904 12232 -3728
rect 186 -6644 220 -5468
rect 1044 -6644 1078 -5468
rect 1902 -6644 1936 -5468
rect 2760 -6644 2794 -5468
rect 3618 -6644 3652 -5468
rect 4476 -6644 4510 -5468
rect 5334 -6644 5368 -5468
rect 6192 -6644 6226 -5468
rect 7050 -6644 7084 -5468
rect 7908 -6644 7942 -5468
rect 8766 -6644 8800 -5468
rect 9624 -6644 9658 -5468
rect 10482 -6644 10516 -5468
rect 11340 -6644 11374 -5468
rect 12198 -6644 12232 -5468
<< psubdiff >>
rect -362 -7878 -200 -7778
rect 12460 -7878 12622 -7778
rect -362 -7940 -262 -7878
rect 12522 -7940 12622 -7878
rect -362 -10722 -262 -10660
rect 12522 -10722 12622 -10660
rect -362 -10822 -200 -10722
rect 12460 -10822 12622 -10722
<< nsubdiff >>
rect -362 2822 -200 2922
rect 12460 2822 12622 2922
rect -362 2760 -262 2822
rect 12522 2760 12622 2822
rect -362 -7442 -262 -7380
rect 12522 -7442 12622 -7380
rect -362 -7542 -200 -7442
rect 12460 -7542 12622 -7442
<< psubdiffcont >>
rect -200 -7878 12460 -7778
rect -362 -10660 -262 -7940
rect 12522 -10660 12622 -7940
rect -200 -10822 12460 -10722
<< nsubdiffcont >>
rect -200 2822 12460 2922
rect -362 -7380 -262 2760
rect 12522 -7380 12622 2760
rect -200 -7542 12460 -7442
<< poly >>
rect 386 1585 878 1601
rect 386 1568 402 1585
rect 232 1551 402 1568
rect 862 1568 878 1585
rect 1244 1585 1736 1601
rect 1244 1568 1260 1585
rect 862 1551 1032 1568
rect 232 1504 1032 1551
rect 1090 1551 1260 1568
rect 1720 1568 1736 1585
rect 2102 1585 2594 1601
rect 2102 1568 2118 1585
rect 1720 1551 1890 1568
rect 1090 1504 1890 1551
rect 1948 1551 2118 1568
rect 2578 1568 2594 1585
rect 2960 1585 3452 1601
rect 2960 1568 2976 1585
rect 2578 1551 2748 1568
rect 1948 1504 2748 1551
rect 2806 1551 2976 1568
rect 3436 1568 3452 1585
rect 3818 1585 4310 1601
rect 3818 1568 3834 1585
rect 3436 1551 3606 1568
rect 2806 1504 3606 1551
rect 3664 1551 3834 1568
rect 4294 1568 4310 1585
rect 4676 1585 5168 1601
rect 4676 1568 4692 1585
rect 4294 1551 4464 1568
rect 3664 1504 4464 1551
rect 4522 1551 4692 1568
rect 5152 1568 5168 1585
rect 5534 1585 6026 1601
rect 5534 1568 5550 1585
rect 5152 1551 5322 1568
rect 4522 1504 5322 1551
rect 5380 1551 5550 1568
rect 6010 1568 6026 1585
rect 6392 1585 6884 1601
rect 6392 1568 6408 1585
rect 6010 1551 6180 1568
rect 5380 1504 6180 1551
rect 6238 1551 6408 1568
rect 6868 1568 6884 1585
rect 7250 1585 7742 1601
rect 7250 1568 7266 1585
rect 6868 1551 7038 1568
rect 6238 1504 7038 1551
rect 7096 1551 7266 1568
rect 7726 1568 7742 1585
rect 8108 1585 8600 1601
rect 8108 1568 8124 1585
rect 7726 1551 7896 1568
rect 7096 1504 7896 1551
rect 7954 1551 8124 1568
rect 8584 1568 8600 1585
rect 8966 1585 9458 1601
rect 8966 1568 8982 1585
rect 8584 1551 8754 1568
rect 7954 1504 8754 1551
rect 8812 1551 8982 1568
rect 9442 1568 9458 1585
rect 9824 1585 10316 1601
rect 9824 1568 9840 1585
rect 9442 1551 9612 1568
rect 8812 1504 9612 1551
rect 9670 1551 9840 1568
rect 10300 1568 10316 1585
rect 10682 1585 11174 1601
rect 10682 1568 10698 1585
rect 10300 1551 10470 1568
rect 9670 1504 10470 1551
rect 10528 1551 10698 1568
rect 11158 1568 11174 1585
rect 11540 1585 12032 1601
rect 11540 1568 11556 1585
rect 11158 1551 11328 1568
rect 10528 1504 11328 1551
rect 11386 1551 11556 1568
rect 12016 1568 12032 1585
rect 12016 1551 12186 1568
rect 11386 1504 12186 1551
rect 232 257 1032 304
rect 232 240 402 257
rect 386 223 402 240
rect 862 240 1032 257
rect 1090 257 1890 304
rect 1090 240 1260 257
rect 862 223 878 240
rect 386 207 878 223
rect 1244 223 1260 240
rect 1720 240 1890 257
rect 1948 257 2748 304
rect 1948 240 2118 257
rect 1720 223 1736 240
rect 1244 207 1736 223
rect 2102 223 2118 240
rect 2578 240 2748 257
rect 2806 257 3606 304
rect 2806 240 2976 257
rect 2578 223 2594 240
rect 2102 207 2594 223
rect 2960 223 2976 240
rect 3436 240 3606 257
rect 3664 257 4464 304
rect 3664 240 3834 257
rect 3436 223 3452 240
rect 2960 207 3452 223
rect 3818 223 3834 240
rect 4294 240 4464 257
rect 4522 257 5322 304
rect 4522 240 4692 257
rect 4294 223 4310 240
rect 3818 207 4310 223
rect 4676 223 4692 240
rect 5152 240 5322 257
rect 5380 257 6180 304
rect 5380 240 5550 257
rect 5152 223 5168 240
rect 4676 207 5168 223
rect 5534 223 5550 240
rect 6010 240 6180 257
rect 6238 257 7038 304
rect 6238 240 6408 257
rect 6010 223 6026 240
rect 5534 207 6026 223
rect 6392 223 6408 240
rect 6868 240 7038 257
rect 7096 257 7896 304
rect 7096 240 7266 257
rect 6868 223 6884 240
rect 6392 207 6884 223
rect 7250 223 7266 240
rect 7726 240 7896 257
rect 7954 257 8754 304
rect 7954 240 8124 257
rect 7726 223 7742 240
rect 7250 207 7742 223
rect 8108 223 8124 240
rect 8584 240 8754 257
rect 8812 257 9612 304
rect 8812 240 8982 257
rect 8584 223 8600 240
rect 8108 207 8600 223
rect 8966 223 8982 240
rect 9442 240 9612 257
rect 9670 257 10470 304
rect 9670 240 9840 257
rect 9442 223 9458 240
rect 8966 207 9458 223
rect 9824 223 9840 240
rect 10300 240 10470 257
rect 10528 257 11328 304
rect 10528 240 10698 257
rect 10300 223 10316 240
rect 9824 207 10316 223
rect 10682 223 10698 240
rect 11158 240 11328 257
rect 11386 257 12186 304
rect 11386 240 11556 257
rect 11158 223 11174 240
rect 10682 207 11174 223
rect 11540 223 11556 240
rect 12016 240 12186 257
rect 12016 223 12032 240
rect 11540 207 12032 223
rect 386 -155 878 -139
rect 386 -172 402 -155
rect 232 -189 402 -172
rect 862 -172 878 -155
rect 1244 -155 1736 -139
rect 1244 -172 1260 -155
rect 862 -189 1032 -172
rect 232 -236 1032 -189
rect 1090 -189 1260 -172
rect 1720 -172 1736 -155
rect 2102 -155 2594 -139
rect 2102 -172 2118 -155
rect 1720 -189 1890 -172
rect 1090 -236 1890 -189
rect 1948 -189 2118 -172
rect 2578 -172 2594 -155
rect 2960 -155 3452 -139
rect 2960 -172 2976 -155
rect 2578 -189 2748 -172
rect 1948 -236 2748 -189
rect 2806 -189 2976 -172
rect 3436 -172 3452 -155
rect 3818 -155 4310 -139
rect 3818 -172 3834 -155
rect 3436 -189 3606 -172
rect 2806 -236 3606 -189
rect 3664 -189 3834 -172
rect 4294 -172 4310 -155
rect 4676 -155 5168 -139
rect 4676 -172 4692 -155
rect 4294 -189 4464 -172
rect 3664 -236 4464 -189
rect 4522 -189 4692 -172
rect 5152 -172 5168 -155
rect 5534 -155 6026 -139
rect 5534 -172 5550 -155
rect 5152 -189 5322 -172
rect 4522 -236 5322 -189
rect 5380 -189 5550 -172
rect 6010 -172 6026 -155
rect 6392 -155 6884 -139
rect 6392 -172 6408 -155
rect 6010 -189 6180 -172
rect 5380 -236 6180 -189
rect 6238 -189 6408 -172
rect 6868 -172 6884 -155
rect 7250 -155 7742 -139
rect 7250 -172 7266 -155
rect 6868 -189 7038 -172
rect 6238 -236 7038 -189
rect 7096 -189 7266 -172
rect 7726 -172 7742 -155
rect 8108 -155 8600 -139
rect 8108 -172 8124 -155
rect 7726 -189 7896 -172
rect 7096 -236 7896 -189
rect 7954 -189 8124 -172
rect 8584 -172 8600 -155
rect 8966 -155 9458 -139
rect 8966 -172 8982 -155
rect 8584 -189 8754 -172
rect 7954 -236 8754 -189
rect 8812 -189 8982 -172
rect 9442 -172 9458 -155
rect 9824 -155 10316 -139
rect 9824 -172 9840 -155
rect 9442 -189 9612 -172
rect 8812 -236 9612 -189
rect 9670 -189 9840 -172
rect 10300 -172 10316 -155
rect 10682 -155 11174 -139
rect 10682 -172 10698 -155
rect 10300 -189 10470 -172
rect 9670 -236 10470 -189
rect 10528 -189 10698 -172
rect 11158 -172 11174 -155
rect 11540 -155 12032 -139
rect 11540 -172 11556 -155
rect 11158 -189 11328 -172
rect 10528 -236 11328 -189
rect 11386 -189 11556 -172
rect 12016 -172 12032 -155
rect 12016 -189 12186 -172
rect 11386 -236 12186 -189
rect 232 -1483 1032 -1436
rect 232 -1500 402 -1483
rect 386 -1517 402 -1500
rect 862 -1500 1032 -1483
rect 1090 -1483 1890 -1436
rect 1090 -1500 1260 -1483
rect 862 -1517 878 -1500
rect 386 -1533 878 -1517
rect 1244 -1517 1260 -1500
rect 1720 -1500 1890 -1483
rect 1948 -1483 2748 -1436
rect 1948 -1500 2118 -1483
rect 1720 -1517 1736 -1500
rect 1244 -1533 1736 -1517
rect 2102 -1517 2118 -1500
rect 2578 -1500 2748 -1483
rect 2806 -1483 3606 -1436
rect 2806 -1500 2976 -1483
rect 2578 -1517 2594 -1500
rect 2102 -1533 2594 -1517
rect 2960 -1517 2976 -1500
rect 3436 -1500 3606 -1483
rect 3664 -1483 4464 -1436
rect 3664 -1500 3834 -1483
rect 3436 -1517 3452 -1500
rect 2960 -1533 3452 -1517
rect 3818 -1517 3834 -1500
rect 4294 -1500 4464 -1483
rect 4522 -1483 5322 -1436
rect 4522 -1500 4692 -1483
rect 4294 -1517 4310 -1500
rect 3818 -1533 4310 -1517
rect 4676 -1517 4692 -1500
rect 5152 -1500 5322 -1483
rect 5380 -1483 6180 -1436
rect 5380 -1500 5550 -1483
rect 5152 -1517 5168 -1500
rect 4676 -1533 5168 -1517
rect 5534 -1517 5550 -1500
rect 6010 -1500 6180 -1483
rect 6238 -1483 7038 -1436
rect 6238 -1500 6408 -1483
rect 6010 -1517 6026 -1500
rect 5534 -1533 6026 -1517
rect 6392 -1517 6408 -1500
rect 6868 -1500 7038 -1483
rect 7096 -1483 7896 -1436
rect 7096 -1500 7266 -1483
rect 6868 -1517 6884 -1500
rect 6392 -1533 6884 -1517
rect 7250 -1517 7266 -1500
rect 7726 -1500 7896 -1483
rect 7954 -1483 8754 -1436
rect 7954 -1500 8124 -1483
rect 7726 -1517 7742 -1500
rect 7250 -1533 7742 -1517
rect 8108 -1517 8124 -1500
rect 8584 -1500 8754 -1483
rect 8812 -1483 9612 -1436
rect 8812 -1500 8982 -1483
rect 8584 -1517 8600 -1500
rect 8108 -1533 8600 -1517
rect 8966 -1517 8982 -1500
rect 9442 -1500 9612 -1483
rect 9670 -1483 10470 -1436
rect 9670 -1500 9840 -1483
rect 9442 -1517 9458 -1500
rect 8966 -1533 9458 -1517
rect 9824 -1517 9840 -1500
rect 10300 -1500 10470 -1483
rect 10528 -1483 11328 -1436
rect 10528 -1500 10698 -1483
rect 10300 -1517 10316 -1500
rect 9824 -1533 10316 -1517
rect 10682 -1517 10698 -1500
rect 11158 -1500 11328 -1483
rect 11386 -1483 12186 -1436
rect 11386 -1500 11556 -1483
rect 11158 -1517 11174 -1500
rect 10682 -1533 11174 -1517
rect 11540 -1517 11556 -1500
rect 12016 -1500 12186 -1483
rect 12016 -1517 12032 -1500
rect 11540 -1533 12032 -1517
rect 386 -1895 878 -1879
rect 386 -1912 402 -1895
rect 232 -1929 402 -1912
rect 862 -1912 878 -1895
rect 1244 -1895 1736 -1879
rect 1244 -1912 1260 -1895
rect 862 -1929 1032 -1912
rect 232 -1976 1032 -1929
rect 1090 -1929 1260 -1912
rect 1720 -1912 1736 -1895
rect 2102 -1895 2594 -1879
rect 2102 -1912 2118 -1895
rect 1720 -1929 1890 -1912
rect 1090 -1976 1890 -1929
rect 1948 -1929 2118 -1912
rect 2578 -1912 2594 -1895
rect 2960 -1895 3452 -1879
rect 2960 -1912 2976 -1895
rect 2578 -1929 2748 -1912
rect 1948 -1976 2748 -1929
rect 2806 -1929 2976 -1912
rect 3436 -1912 3452 -1895
rect 3818 -1895 4310 -1879
rect 3818 -1912 3834 -1895
rect 3436 -1929 3606 -1912
rect 2806 -1976 3606 -1929
rect 3664 -1929 3834 -1912
rect 4294 -1912 4310 -1895
rect 4676 -1895 5168 -1879
rect 4676 -1912 4692 -1895
rect 4294 -1929 4464 -1912
rect 3664 -1976 4464 -1929
rect 4522 -1929 4692 -1912
rect 5152 -1912 5168 -1895
rect 5534 -1895 6026 -1879
rect 5534 -1912 5550 -1895
rect 5152 -1929 5322 -1912
rect 4522 -1976 5322 -1929
rect 5380 -1929 5550 -1912
rect 6010 -1912 6026 -1895
rect 6392 -1895 6884 -1879
rect 6392 -1912 6408 -1895
rect 6010 -1929 6180 -1912
rect 5380 -1976 6180 -1929
rect 6238 -1929 6408 -1912
rect 6868 -1912 6884 -1895
rect 7250 -1895 7742 -1879
rect 7250 -1912 7266 -1895
rect 6868 -1929 7038 -1912
rect 6238 -1976 7038 -1929
rect 7096 -1929 7266 -1912
rect 7726 -1912 7742 -1895
rect 8108 -1895 8600 -1879
rect 8108 -1912 8124 -1895
rect 7726 -1929 7896 -1912
rect 7096 -1976 7896 -1929
rect 7954 -1929 8124 -1912
rect 8584 -1912 8600 -1895
rect 8966 -1895 9458 -1879
rect 8966 -1912 8982 -1895
rect 8584 -1929 8754 -1912
rect 7954 -1976 8754 -1929
rect 8812 -1929 8982 -1912
rect 9442 -1912 9458 -1895
rect 9824 -1895 10316 -1879
rect 9824 -1912 9840 -1895
rect 9442 -1929 9612 -1912
rect 8812 -1976 9612 -1929
rect 9670 -1929 9840 -1912
rect 10300 -1912 10316 -1895
rect 10682 -1895 11174 -1879
rect 10682 -1912 10698 -1895
rect 10300 -1929 10470 -1912
rect 9670 -1976 10470 -1929
rect 10528 -1929 10698 -1912
rect 11158 -1912 11174 -1895
rect 11540 -1895 12032 -1879
rect 11540 -1912 11556 -1895
rect 11158 -1929 11328 -1912
rect 10528 -1976 11328 -1929
rect 11386 -1929 11556 -1912
rect 12016 -1912 12032 -1895
rect 12016 -1929 12186 -1912
rect 11386 -1976 12186 -1929
rect 232 -3223 1032 -3176
rect 232 -3240 402 -3223
rect 386 -3257 402 -3240
rect 862 -3240 1032 -3223
rect 1090 -3223 1890 -3176
rect 1090 -3240 1260 -3223
rect 862 -3257 878 -3240
rect 386 -3273 878 -3257
rect 1244 -3257 1260 -3240
rect 1720 -3240 1890 -3223
rect 1948 -3223 2748 -3176
rect 1948 -3240 2118 -3223
rect 1720 -3257 1736 -3240
rect 1244 -3273 1736 -3257
rect 2102 -3257 2118 -3240
rect 2578 -3240 2748 -3223
rect 2806 -3223 3606 -3176
rect 2806 -3240 2976 -3223
rect 2578 -3257 2594 -3240
rect 2102 -3273 2594 -3257
rect 2960 -3257 2976 -3240
rect 3436 -3240 3606 -3223
rect 3664 -3223 4464 -3176
rect 3664 -3240 3834 -3223
rect 3436 -3257 3452 -3240
rect 2960 -3273 3452 -3257
rect 3818 -3257 3834 -3240
rect 4294 -3240 4464 -3223
rect 4522 -3223 5322 -3176
rect 4522 -3240 4692 -3223
rect 4294 -3257 4310 -3240
rect 3818 -3273 4310 -3257
rect 4676 -3257 4692 -3240
rect 5152 -3240 5322 -3223
rect 5380 -3223 6180 -3176
rect 5380 -3240 5550 -3223
rect 5152 -3257 5168 -3240
rect 4676 -3273 5168 -3257
rect 5534 -3257 5550 -3240
rect 6010 -3240 6180 -3223
rect 6238 -3223 7038 -3176
rect 6238 -3240 6408 -3223
rect 6010 -3257 6026 -3240
rect 5534 -3273 6026 -3257
rect 6392 -3257 6408 -3240
rect 6868 -3240 7038 -3223
rect 7096 -3223 7896 -3176
rect 7096 -3240 7266 -3223
rect 6868 -3257 6884 -3240
rect 6392 -3273 6884 -3257
rect 7250 -3257 7266 -3240
rect 7726 -3240 7896 -3223
rect 7954 -3223 8754 -3176
rect 7954 -3240 8124 -3223
rect 7726 -3257 7742 -3240
rect 7250 -3273 7742 -3257
rect 8108 -3257 8124 -3240
rect 8584 -3240 8754 -3223
rect 8812 -3223 9612 -3176
rect 8812 -3240 8982 -3223
rect 8584 -3257 8600 -3240
rect 8108 -3273 8600 -3257
rect 8966 -3257 8982 -3240
rect 9442 -3240 9612 -3223
rect 9670 -3223 10470 -3176
rect 9670 -3240 9840 -3223
rect 9442 -3257 9458 -3240
rect 8966 -3273 9458 -3257
rect 9824 -3257 9840 -3240
rect 10300 -3240 10470 -3223
rect 10528 -3223 11328 -3176
rect 10528 -3240 10698 -3223
rect 10300 -3257 10316 -3240
rect 9824 -3273 10316 -3257
rect 10682 -3257 10698 -3240
rect 11158 -3240 11328 -3223
rect 11386 -3223 12186 -3176
rect 11386 -3240 11556 -3223
rect 11158 -3257 11174 -3240
rect 10682 -3273 11174 -3257
rect 11540 -3257 11556 -3240
rect 12016 -3240 12186 -3223
rect 12016 -3257 12032 -3240
rect 11540 -3273 12032 -3257
rect 386 -3635 878 -3619
rect 386 -3652 402 -3635
rect 232 -3669 402 -3652
rect 862 -3652 878 -3635
rect 1244 -3635 1736 -3619
rect 1244 -3652 1260 -3635
rect 862 -3669 1032 -3652
rect 232 -3716 1032 -3669
rect 1090 -3669 1260 -3652
rect 1720 -3652 1736 -3635
rect 2102 -3635 2594 -3619
rect 2102 -3652 2118 -3635
rect 1720 -3669 1890 -3652
rect 1090 -3716 1890 -3669
rect 1948 -3669 2118 -3652
rect 2578 -3652 2594 -3635
rect 2960 -3635 3452 -3619
rect 2960 -3652 2976 -3635
rect 2578 -3669 2748 -3652
rect 1948 -3716 2748 -3669
rect 2806 -3669 2976 -3652
rect 3436 -3652 3452 -3635
rect 3818 -3635 4310 -3619
rect 3818 -3652 3834 -3635
rect 3436 -3669 3606 -3652
rect 2806 -3716 3606 -3669
rect 3664 -3669 3834 -3652
rect 4294 -3652 4310 -3635
rect 4676 -3635 5168 -3619
rect 4676 -3652 4692 -3635
rect 4294 -3669 4464 -3652
rect 3664 -3716 4464 -3669
rect 4522 -3669 4692 -3652
rect 5152 -3652 5168 -3635
rect 5534 -3635 6026 -3619
rect 5534 -3652 5550 -3635
rect 5152 -3669 5322 -3652
rect 4522 -3716 5322 -3669
rect 5380 -3669 5550 -3652
rect 6010 -3652 6026 -3635
rect 6392 -3635 6884 -3619
rect 6392 -3652 6408 -3635
rect 6010 -3669 6180 -3652
rect 5380 -3716 6180 -3669
rect 6238 -3669 6408 -3652
rect 6868 -3652 6884 -3635
rect 7250 -3635 7742 -3619
rect 7250 -3652 7266 -3635
rect 6868 -3669 7038 -3652
rect 6238 -3716 7038 -3669
rect 7096 -3669 7266 -3652
rect 7726 -3652 7742 -3635
rect 8108 -3635 8600 -3619
rect 8108 -3652 8124 -3635
rect 7726 -3669 7896 -3652
rect 7096 -3716 7896 -3669
rect 7954 -3669 8124 -3652
rect 8584 -3652 8600 -3635
rect 8966 -3635 9458 -3619
rect 8966 -3652 8982 -3635
rect 8584 -3669 8754 -3652
rect 7954 -3716 8754 -3669
rect 8812 -3669 8982 -3652
rect 9442 -3652 9458 -3635
rect 9824 -3635 10316 -3619
rect 9824 -3652 9840 -3635
rect 9442 -3669 9612 -3652
rect 8812 -3716 9612 -3669
rect 9670 -3669 9840 -3652
rect 10300 -3652 10316 -3635
rect 10682 -3635 11174 -3619
rect 10682 -3652 10698 -3635
rect 10300 -3669 10470 -3652
rect 9670 -3716 10470 -3669
rect 10528 -3669 10698 -3652
rect 11158 -3652 11174 -3635
rect 11540 -3635 12032 -3619
rect 11540 -3652 11556 -3635
rect 11158 -3669 11328 -3652
rect 10528 -3716 11328 -3669
rect 11386 -3669 11556 -3652
rect 12016 -3652 12032 -3635
rect 12016 -3669 12186 -3652
rect 11386 -3716 12186 -3669
rect 232 -4963 1032 -4916
rect 232 -4980 402 -4963
rect 386 -4997 402 -4980
rect 862 -4980 1032 -4963
rect 1090 -4963 1890 -4916
rect 1090 -4980 1260 -4963
rect 862 -4997 878 -4980
rect 386 -5013 878 -4997
rect 1244 -4997 1260 -4980
rect 1720 -4980 1890 -4963
rect 1948 -4963 2748 -4916
rect 1948 -4980 2118 -4963
rect 1720 -4997 1736 -4980
rect 1244 -5013 1736 -4997
rect 2102 -4997 2118 -4980
rect 2578 -4980 2748 -4963
rect 2806 -4963 3606 -4916
rect 2806 -4980 2976 -4963
rect 2578 -4997 2594 -4980
rect 2102 -5013 2594 -4997
rect 2960 -4997 2976 -4980
rect 3436 -4980 3606 -4963
rect 3664 -4963 4464 -4916
rect 3664 -4980 3834 -4963
rect 3436 -4997 3452 -4980
rect 2960 -5013 3452 -4997
rect 3818 -4997 3834 -4980
rect 4294 -4980 4464 -4963
rect 4522 -4963 5322 -4916
rect 4522 -4980 4692 -4963
rect 4294 -4997 4310 -4980
rect 3818 -5013 4310 -4997
rect 4676 -4997 4692 -4980
rect 5152 -4980 5322 -4963
rect 5380 -4963 6180 -4916
rect 5380 -4980 5550 -4963
rect 5152 -4997 5168 -4980
rect 4676 -5013 5168 -4997
rect 5534 -4997 5550 -4980
rect 6010 -4980 6180 -4963
rect 6238 -4963 7038 -4916
rect 6238 -4980 6408 -4963
rect 6010 -4997 6026 -4980
rect 5534 -5013 6026 -4997
rect 6392 -4997 6408 -4980
rect 6868 -4980 7038 -4963
rect 7096 -4963 7896 -4916
rect 7096 -4980 7266 -4963
rect 6868 -4997 6884 -4980
rect 6392 -5013 6884 -4997
rect 7250 -4997 7266 -4980
rect 7726 -4980 7896 -4963
rect 7954 -4963 8754 -4916
rect 7954 -4980 8124 -4963
rect 7726 -4997 7742 -4980
rect 7250 -5013 7742 -4997
rect 8108 -4997 8124 -4980
rect 8584 -4980 8754 -4963
rect 8812 -4963 9612 -4916
rect 8812 -4980 8982 -4963
rect 8584 -4997 8600 -4980
rect 8108 -5013 8600 -4997
rect 8966 -4997 8982 -4980
rect 9442 -4980 9612 -4963
rect 9670 -4963 10470 -4916
rect 9670 -4980 9840 -4963
rect 9442 -4997 9458 -4980
rect 8966 -5013 9458 -4997
rect 9824 -4997 9840 -4980
rect 10300 -4980 10470 -4963
rect 10528 -4963 11328 -4916
rect 10528 -4980 10698 -4963
rect 10300 -4997 10316 -4980
rect 9824 -5013 10316 -4997
rect 10682 -4997 10698 -4980
rect 11158 -4980 11328 -4963
rect 11386 -4963 12186 -4916
rect 11386 -4980 11556 -4963
rect 11158 -4997 11174 -4980
rect 10682 -5013 11174 -4997
rect 11540 -4997 11556 -4980
rect 12016 -4980 12186 -4963
rect 12016 -4997 12032 -4980
rect 11540 -5013 12032 -4997
rect 386 -5375 878 -5359
rect 386 -5392 402 -5375
rect 232 -5409 402 -5392
rect 862 -5392 878 -5375
rect 1244 -5375 1736 -5359
rect 1244 -5392 1260 -5375
rect 862 -5409 1032 -5392
rect 232 -5456 1032 -5409
rect 1090 -5409 1260 -5392
rect 1720 -5392 1736 -5375
rect 2102 -5375 2594 -5359
rect 2102 -5392 2118 -5375
rect 1720 -5409 1890 -5392
rect 1090 -5456 1890 -5409
rect 1948 -5409 2118 -5392
rect 2578 -5392 2594 -5375
rect 2960 -5375 3452 -5359
rect 2960 -5392 2976 -5375
rect 2578 -5409 2748 -5392
rect 1948 -5456 2748 -5409
rect 2806 -5409 2976 -5392
rect 3436 -5392 3452 -5375
rect 3818 -5375 4310 -5359
rect 3818 -5392 3834 -5375
rect 3436 -5409 3606 -5392
rect 2806 -5456 3606 -5409
rect 3664 -5409 3834 -5392
rect 4294 -5392 4310 -5375
rect 4676 -5375 5168 -5359
rect 4676 -5392 4692 -5375
rect 4294 -5409 4464 -5392
rect 3664 -5456 4464 -5409
rect 4522 -5409 4692 -5392
rect 5152 -5392 5168 -5375
rect 5534 -5375 6026 -5359
rect 5534 -5392 5550 -5375
rect 5152 -5409 5322 -5392
rect 4522 -5456 5322 -5409
rect 5380 -5409 5550 -5392
rect 6010 -5392 6026 -5375
rect 6392 -5375 6884 -5359
rect 6392 -5392 6408 -5375
rect 6010 -5409 6180 -5392
rect 5380 -5456 6180 -5409
rect 6238 -5409 6408 -5392
rect 6868 -5392 6884 -5375
rect 7250 -5375 7742 -5359
rect 7250 -5392 7266 -5375
rect 6868 -5409 7038 -5392
rect 6238 -5456 7038 -5409
rect 7096 -5409 7266 -5392
rect 7726 -5392 7742 -5375
rect 8108 -5375 8600 -5359
rect 8108 -5392 8124 -5375
rect 7726 -5409 7896 -5392
rect 7096 -5456 7896 -5409
rect 7954 -5409 8124 -5392
rect 8584 -5392 8600 -5375
rect 8966 -5375 9458 -5359
rect 8966 -5392 8982 -5375
rect 8584 -5409 8754 -5392
rect 7954 -5456 8754 -5409
rect 8812 -5409 8982 -5392
rect 9442 -5392 9458 -5375
rect 9824 -5375 10316 -5359
rect 9824 -5392 9840 -5375
rect 9442 -5409 9612 -5392
rect 8812 -5456 9612 -5409
rect 9670 -5409 9840 -5392
rect 10300 -5392 10316 -5375
rect 10682 -5375 11174 -5359
rect 10682 -5392 10698 -5375
rect 10300 -5409 10470 -5392
rect 9670 -5456 10470 -5409
rect 10528 -5409 10698 -5392
rect 11158 -5392 11174 -5375
rect 11540 -5375 12032 -5359
rect 11540 -5392 11556 -5375
rect 11158 -5409 11328 -5392
rect 10528 -5456 11328 -5409
rect 11386 -5409 11556 -5392
rect 12016 -5392 12032 -5375
rect 12016 -5409 12186 -5392
rect 11386 -5456 12186 -5409
rect 232 -6703 1032 -6656
rect 232 -6720 402 -6703
rect 386 -6737 402 -6720
rect 862 -6720 1032 -6703
rect 1090 -6703 1890 -6656
rect 1090 -6720 1260 -6703
rect 862 -6737 878 -6720
rect 386 -6753 878 -6737
rect 1244 -6737 1260 -6720
rect 1720 -6720 1890 -6703
rect 1948 -6703 2748 -6656
rect 1948 -6720 2118 -6703
rect 1720 -6737 1736 -6720
rect 1244 -6753 1736 -6737
rect 2102 -6737 2118 -6720
rect 2578 -6720 2748 -6703
rect 2806 -6703 3606 -6656
rect 2806 -6720 2976 -6703
rect 2578 -6737 2594 -6720
rect 2102 -6753 2594 -6737
rect 2960 -6737 2976 -6720
rect 3436 -6720 3606 -6703
rect 3664 -6703 4464 -6656
rect 3664 -6720 3834 -6703
rect 3436 -6737 3452 -6720
rect 2960 -6753 3452 -6737
rect 3818 -6737 3834 -6720
rect 4294 -6720 4464 -6703
rect 4522 -6703 5322 -6656
rect 4522 -6720 4692 -6703
rect 4294 -6737 4310 -6720
rect 3818 -6753 4310 -6737
rect 4676 -6737 4692 -6720
rect 5152 -6720 5322 -6703
rect 5380 -6703 6180 -6656
rect 5380 -6720 5550 -6703
rect 5152 -6737 5168 -6720
rect 4676 -6753 5168 -6737
rect 5534 -6737 5550 -6720
rect 6010 -6720 6180 -6703
rect 6238 -6703 7038 -6656
rect 6238 -6720 6408 -6703
rect 6010 -6737 6026 -6720
rect 5534 -6753 6026 -6737
rect 6392 -6737 6408 -6720
rect 6868 -6720 7038 -6703
rect 7096 -6703 7896 -6656
rect 7096 -6720 7266 -6703
rect 6868 -6737 6884 -6720
rect 6392 -6753 6884 -6737
rect 7250 -6737 7266 -6720
rect 7726 -6720 7896 -6703
rect 7954 -6703 8754 -6656
rect 7954 -6720 8124 -6703
rect 7726 -6737 7742 -6720
rect 7250 -6753 7742 -6737
rect 8108 -6737 8124 -6720
rect 8584 -6720 8754 -6703
rect 8812 -6703 9612 -6656
rect 8812 -6720 8982 -6703
rect 8584 -6737 8600 -6720
rect 8108 -6753 8600 -6737
rect 8966 -6737 8982 -6720
rect 9442 -6720 9612 -6703
rect 9670 -6703 10470 -6656
rect 9670 -6720 9840 -6703
rect 9442 -6737 9458 -6720
rect 8966 -6753 9458 -6737
rect 9824 -6737 9840 -6720
rect 10300 -6720 10470 -6703
rect 10528 -6703 11328 -6656
rect 10528 -6720 10698 -6703
rect 10300 -6737 10316 -6720
rect 9824 -6753 10316 -6737
rect 10682 -6737 10698 -6720
rect 11158 -6720 11328 -6703
rect 11386 -6703 12186 -6656
rect 11386 -6720 11556 -6703
rect 11158 -6737 11174 -6720
rect 10682 -6753 11174 -6737
rect 11540 -6737 11556 -6720
rect 12016 -6720 12186 -6703
rect 12016 -6737 12032 -6720
rect 11540 -6753 12032 -6737
rect 5030 -8388 5282 -8372
rect 5030 -8405 5046 -8388
rect 4956 -8422 5046 -8405
rect 5266 -8405 5282 -8388
rect 5488 -8388 5740 -8372
rect 5488 -8405 5504 -8388
rect 5266 -8422 5356 -8405
rect 4956 -8460 5356 -8422
rect 5414 -8422 5504 -8405
rect 5724 -8405 5740 -8388
rect 5946 -8388 6198 -8372
rect 5946 -8405 5962 -8388
rect 5724 -8422 5814 -8405
rect 5414 -8460 5814 -8422
rect 5872 -8422 5962 -8405
rect 6182 -8405 6198 -8388
rect 6404 -8388 6656 -8372
rect 6404 -8405 6420 -8388
rect 6182 -8422 6272 -8405
rect 5872 -8460 6272 -8422
rect 6330 -8422 6420 -8405
rect 6640 -8405 6656 -8388
rect 6862 -8388 7114 -8372
rect 6862 -8405 6878 -8388
rect 6640 -8422 6730 -8405
rect 6330 -8460 6730 -8422
rect 6788 -8422 6878 -8405
rect 7098 -8405 7114 -8388
rect 7320 -8388 7572 -8372
rect 7320 -8405 7336 -8388
rect 7098 -8422 7188 -8405
rect 6788 -8460 7188 -8422
rect 7246 -8422 7336 -8405
rect 7556 -8405 7572 -8388
rect 7556 -8422 7646 -8405
rect 7246 -8460 7646 -8422
rect 4956 -8898 5356 -8860
rect 4956 -8915 5046 -8898
rect 5030 -8932 5046 -8915
rect 5266 -8915 5356 -8898
rect 5414 -8898 5814 -8860
rect 5414 -8915 5504 -8898
rect 5266 -8932 5282 -8915
rect 5030 -8948 5282 -8932
rect 5488 -8932 5504 -8915
rect 5724 -8915 5814 -8898
rect 5872 -8898 6272 -8860
rect 5872 -8915 5962 -8898
rect 5724 -8932 5740 -8915
rect 5488 -8948 5740 -8932
rect 5946 -8932 5962 -8915
rect 6182 -8915 6272 -8898
rect 6330 -8898 6730 -8860
rect 6330 -8915 6420 -8898
rect 6182 -8932 6198 -8915
rect 5946 -8948 6198 -8932
rect 6404 -8932 6420 -8915
rect 6640 -8915 6730 -8898
rect 6788 -8898 7188 -8860
rect 6788 -8915 6878 -8898
rect 6640 -8932 6656 -8915
rect 6404 -8948 6656 -8932
rect 6862 -8932 6878 -8915
rect 7098 -8915 7188 -8898
rect 7246 -8898 7646 -8860
rect 7246 -8915 7336 -8898
rect 7098 -8932 7114 -8915
rect 6862 -8948 7114 -8932
rect 7320 -8932 7336 -8915
rect 7556 -8915 7646 -8898
rect 7556 -8932 7572 -8915
rect 7320 -8948 7572 -8932
rect 5030 -9188 5282 -9172
rect 5030 -9205 5046 -9188
rect 4956 -9222 5046 -9205
rect 5266 -9205 5282 -9188
rect 5488 -9188 5740 -9172
rect 5488 -9205 5504 -9188
rect 5266 -9222 5356 -9205
rect 4956 -9260 5356 -9222
rect 5414 -9222 5504 -9205
rect 5724 -9205 5740 -9188
rect 5946 -9188 6198 -9172
rect 5946 -9205 5962 -9188
rect 5724 -9222 5814 -9205
rect 5414 -9260 5814 -9222
rect 5872 -9222 5962 -9205
rect 6182 -9205 6198 -9188
rect 6404 -9188 6656 -9172
rect 6404 -9205 6420 -9188
rect 6182 -9222 6272 -9205
rect 5872 -9260 6272 -9222
rect 6330 -9222 6420 -9205
rect 6640 -9205 6656 -9188
rect 6862 -9188 7114 -9172
rect 6862 -9205 6878 -9188
rect 6640 -9222 6730 -9205
rect 6330 -9260 6730 -9222
rect 6788 -9222 6878 -9205
rect 7098 -9205 7114 -9188
rect 7320 -9188 7572 -9172
rect 7320 -9205 7336 -9188
rect 7098 -9222 7188 -9205
rect 6788 -9260 7188 -9222
rect 7246 -9222 7336 -9205
rect 7556 -9205 7572 -9188
rect 7556 -9222 7646 -9205
rect 7246 -9260 7646 -9222
rect 4956 -9698 5356 -9660
rect 4956 -9715 5046 -9698
rect 5030 -9732 5046 -9715
rect 5266 -9715 5356 -9698
rect 5414 -9698 5814 -9660
rect 5414 -9715 5504 -9698
rect 5266 -9732 5282 -9715
rect 5030 -9748 5282 -9732
rect 5488 -9732 5504 -9715
rect 5724 -9715 5814 -9698
rect 5872 -9698 6272 -9660
rect 5872 -9715 5962 -9698
rect 5724 -9732 5740 -9715
rect 5488 -9748 5740 -9732
rect 5946 -9732 5962 -9715
rect 6182 -9715 6272 -9698
rect 6330 -9698 6730 -9660
rect 6330 -9715 6420 -9698
rect 6182 -9732 6198 -9715
rect 5946 -9748 6198 -9732
rect 6404 -9732 6420 -9715
rect 6640 -9715 6730 -9698
rect 6788 -9698 7188 -9660
rect 6788 -9715 6878 -9698
rect 6640 -9732 6656 -9715
rect 6404 -9748 6656 -9732
rect 6862 -9732 6878 -9715
rect 7098 -9715 7188 -9698
rect 7246 -9698 7646 -9660
rect 7246 -9715 7336 -9698
rect 7098 -9732 7114 -9715
rect 6862 -9748 7114 -9732
rect 7320 -9732 7336 -9715
rect 7556 -9715 7646 -9698
rect 7556 -9732 7572 -9715
rect 7320 -9748 7572 -9732
<< polycont >>
rect 402 1551 862 1585
rect 1260 1551 1720 1585
rect 2118 1551 2578 1585
rect 2976 1551 3436 1585
rect 3834 1551 4294 1585
rect 4692 1551 5152 1585
rect 5550 1551 6010 1585
rect 6408 1551 6868 1585
rect 7266 1551 7726 1585
rect 8124 1551 8584 1585
rect 8982 1551 9442 1585
rect 9840 1551 10300 1585
rect 10698 1551 11158 1585
rect 11556 1551 12016 1585
rect 402 223 862 257
rect 1260 223 1720 257
rect 2118 223 2578 257
rect 2976 223 3436 257
rect 3834 223 4294 257
rect 4692 223 5152 257
rect 5550 223 6010 257
rect 6408 223 6868 257
rect 7266 223 7726 257
rect 8124 223 8584 257
rect 8982 223 9442 257
rect 9840 223 10300 257
rect 10698 223 11158 257
rect 11556 223 12016 257
rect 402 -189 862 -155
rect 1260 -189 1720 -155
rect 2118 -189 2578 -155
rect 2976 -189 3436 -155
rect 3834 -189 4294 -155
rect 4692 -189 5152 -155
rect 5550 -189 6010 -155
rect 6408 -189 6868 -155
rect 7266 -189 7726 -155
rect 8124 -189 8584 -155
rect 8982 -189 9442 -155
rect 9840 -189 10300 -155
rect 10698 -189 11158 -155
rect 11556 -189 12016 -155
rect 402 -1517 862 -1483
rect 1260 -1517 1720 -1483
rect 2118 -1517 2578 -1483
rect 2976 -1517 3436 -1483
rect 3834 -1517 4294 -1483
rect 4692 -1517 5152 -1483
rect 5550 -1517 6010 -1483
rect 6408 -1517 6868 -1483
rect 7266 -1517 7726 -1483
rect 8124 -1517 8584 -1483
rect 8982 -1517 9442 -1483
rect 9840 -1517 10300 -1483
rect 10698 -1517 11158 -1483
rect 11556 -1517 12016 -1483
rect 402 -1929 862 -1895
rect 1260 -1929 1720 -1895
rect 2118 -1929 2578 -1895
rect 2976 -1929 3436 -1895
rect 3834 -1929 4294 -1895
rect 4692 -1929 5152 -1895
rect 5550 -1929 6010 -1895
rect 6408 -1929 6868 -1895
rect 7266 -1929 7726 -1895
rect 8124 -1929 8584 -1895
rect 8982 -1929 9442 -1895
rect 9840 -1929 10300 -1895
rect 10698 -1929 11158 -1895
rect 11556 -1929 12016 -1895
rect 402 -3257 862 -3223
rect 1260 -3257 1720 -3223
rect 2118 -3257 2578 -3223
rect 2976 -3257 3436 -3223
rect 3834 -3257 4294 -3223
rect 4692 -3257 5152 -3223
rect 5550 -3257 6010 -3223
rect 6408 -3257 6868 -3223
rect 7266 -3257 7726 -3223
rect 8124 -3257 8584 -3223
rect 8982 -3257 9442 -3223
rect 9840 -3257 10300 -3223
rect 10698 -3257 11158 -3223
rect 11556 -3257 12016 -3223
rect 402 -3669 862 -3635
rect 1260 -3669 1720 -3635
rect 2118 -3669 2578 -3635
rect 2976 -3669 3436 -3635
rect 3834 -3669 4294 -3635
rect 4692 -3669 5152 -3635
rect 5550 -3669 6010 -3635
rect 6408 -3669 6868 -3635
rect 7266 -3669 7726 -3635
rect 8124 -3669 8584 -3635
rect 8982 -3669 9442 -3635
rect 9840 -3669 10300 -3635
rect 10698 -3669 11158 -3635
rect 11556 -3669 12016 -3635
rect 402 -4997 862 -4963
rect 1260 -4997 1720 -4963
rect 2118 -4997 2578 -4963
rect 2976 -4997 3436 -4963
rect 3834 -4997 4294 -4963
rect 4692 -4997 5152 -4963
rect 5550 -4997 6010 -4963
rect 6408 -4997 6868 -4963
rect 7266 -4997 7726 -4963
rect 8124 -4997 8584 -4963
rect 8982 -4997 9442 -4963
rect 9840 -4997 10300 -4963
rect 10698 -4997 11158 -4963
rect 11556 -4997 12016 -4963
rect 402 -5409 862 -5375
rect 1260 -5409 1720 -5375
rect 2118 -5409 2578 -5375
rect 2976 -5409 3436 -5375
rect 3834 -5409 4294 -5375
rect 4692 -5409 5152 -5375
rect 5550 -5409 6010 -5375
rect 6408 -5409 6868 -5375
rect 7266 -5409 7726 -5375
rect 8124 -5409 8584 -5375
rect 8982 -5409 9442 -5375
rect 9840 -5409 10300 -5375
rect 10698 -5409 11158 -5375
rect 11556 -5409 12016 -5375
rect 402 -6737 862 -6703
rect 1260 -6737 1720 -6703
rect 2118 -6737 2578 -6703
rect 2976 -6737 3436 -6703
rect 3834 -6737 4294 -6703
rect 4692 -6737 5152 -6703
rect 5550 -6737 6010 -6703
rect 6408 -6737 6868 -6703
rect 7266 -6737 7726 -6703
rect 8124 -6737 8584 -6703
rect 8982 -6737 9442 -6703
rect 9840 -6737 10300 -6703
rect 10698 -6737 11158 -6703
rect 11556 -6737 12016 -6703
rect 5046 -8422 5266 -8388
rect 5504 -8422 5724 -8388
rect 5962 -8422 6182 -8388
rect 6420 -8422 6640 -8388
rect 6878 -8422 7098 -8388
rect 7336 -8422 7556 -8388
rect 5046 -8932 5266 -8898
rect 5504 -8932 5724 -8898
rect 5962 -8932 6182 -8898
rect 6420 -8932 6640 -8898
rect 6878 -8932 7098 -8898
rect 7336 -8932 7556 -8898
rect 5046 -9222 5266 -9188
rect 5504 -9222 5724 -9188
rect 5962 -9222 6182 -9188
rect 6420 -9222 6640 -9188
rect 6878 -9222 7098 -9188
rect 7336 -9222 7556 -9188
rect 5046 -9732 5266 -9698
rect 5504 -9732 5724 -9698
rect 5962 -9732 6182 -9698
rect 6420 -9732 6640 -9698
rect 6878 -9732 7098 -9698
rect 7336 -9732 7556 -9698
<< locali >>
rect -362 2760 -262 2922
rect 12522 2760 12622 2922
rect 386 1551 402 1585
rect 862 1551 878 1585
rect 1244 1551 1260 1585
rect 1720 1551 1736 1585
rect 2102 1551 2118 1585
rect 2578 1551 2594 1585
rect 2960 1551 2976 1585
rect 3436 1551 3452 1585
rect 3818 1551 3834 1585
rect 4294 1551 4310 1585
rect 4676 1551 4692 1585
rect 5152 1551 5168 1585
rect 5534 1551 5550 1585
rect 6010 1551 6026 1585
rect 6392 1551 6408 1585
rect 6868 1551 6884 1585
rect 7250 1551 7266 1585
rect 7726 1551 7742 1585
rect 8108 1551 8124 1585
rect 8584 1551 8600 1585
rect 8966 1551 8982 1585
rect 9442 1551 9458 1585
rect 9824 1551 9840 1585
rect 10300 1551 10316 1585
rect 10682 1551 10698 1585
rect 11158 1551 11174 1585
rect 11540 1551 11556 1585
rect 12016 1551 12032 1585
rect 186 1492 220 1508
rect 186 300 220 316
rect 1044 1492 1078 1508
rect 1044 300 1078 316
rect 1902 1492 1936 1508
rect 1902 300 1936 316
rect 2760 1492 2794 1508
rect 2760 300 2794 316
rect 3618 1492 3652 1508
rect 3618 300 3652 316
rect 4476 1492 4510 1508
rect 4476 300 4510 316
rect 5334 1492 5368 1508
rect 5334 300 5368 316
rect 6192 1492 6226 1508
rect 6192 300 6226 316
rect 7050 1492 7084 1508
rect 7050 300 7084 316
rect 7908 1492 7942 1508
rect 7908 300 7942 316
rect 8766 1492 8800 1508
rect 8766 300 8800 316
rect 9624 1492 9658 1508
rect 9624 300 9658 316
rect 10482 1492 10516 1508
rect 10482 300 10516 316
rect 11340 1492 11374 1508
rect 11340 300 11374 316
rect 12198 1492 12232 1508
rect 12198 300 12232 316
rect 386 223 402 257
rect 862 223 878 257
rect 1244 223 1260 257
rect 1720 223 1736 257
rect 2102 223 2118 257
rect 2578 223 2594 257
rect 2960 223 2976 257
rect 3436 223 3452 257
rect 3818 223 3834 257
rect 4294 223 4310 257
rect 4676 223 4692 257
rect 5152 223 5168 257
rect 5534 223 5550 257
rect 6010 223 6026 257
rect 6392 223 6408 257
rect 6868 223 6884 257
rect 7250 223 7266 257
rect 7726 223 7742 257
rect 8108 223 8124 257
rect 8584 223 8600 257
rect 8966 223 8982 257
rect 9442 223 9458 257
rect 9824 223 9840 257
rect 10300 223 10316 257
rect 10682 223 10698 257
rect 11158 223 11174 257
rect 11540 223 11556 257
rect 12016 223 12032 257
rect 386 -189 402 -155
rect 862 -189 878 -155
rect 1244 -189 1260 -155
rect 1720 -189 1736 -155
rect 2102 -189 2118 -155
rect 2578 -189 2594 -155
rect 2960 -189 2976 -155
rect 3436 -189 3452 -155
rect 3818 -189 3834 -155
rect 4294 -189 4310 -155
rect 4676 -189 4692 -155
rect 5152 -189 5168 -155
rect 5534 -189 5550 -155
rect 6010 -189 6026 -155
rect 6392 -189 6408 -155
rect 6868 -189 6884 -155
rect 7250 -189 7266 -155
rect 7726 -189 7742 -155
rect 8108 -189 8124 -155
rect 8584 -189 8600 -155
rect 8966 -189 8982 -155
rect 9442 -189 9458 -155
rect 9824 -189 9840 -155
rect 10300 -189 10316 -155
rect 10682 -189 10698 -155
rect 11158 -189 11174 -155
rect 11540 -189 11556 -155
rect 12016 -189 12032 -155
rect 186 -248 220 -232
rect 186 -1440 220 -1424
rect 1044 -248 1078 -232
rect 1044 -1440 1078 -1424
rect 1902 -248 1936 -232
rect 1902 -1440 1936 -1424
rect 2760 -248 2794 -232
rect 2760 -1440 2794 -1424
rect 3618 -248 3652 -232
rect 3618 -1440 3652 -1424
rect 4476 -248 4510 -232
rect 4476 -1440 4510 -1424
rect 5334 -248 5368 -232
rect 5334 -1440 5368 -1424
rect 6192 -248 6226 -232
rect 6192 -1440 6226 -1424
rect 7050 -248 7084 -232
rect 7050 -1440 7084 -1424
rect 7908 -248 7942 -232
rect 7908 -1440 7942 -1424
rect 8766 -248 8800 -232
rect 8766 -1440 8800 -1424
rect 9624 -248 9658 -232
rect 9624 -1440 9658 -1424
rect 10482 -248 10516 -232
rect 10482 -1440 10516 -1424
rect 11340 -248 11374 -232
rect 11340 -1440 11374 -1424
rect 12198 -248 12232 -232
rect 12198 -1440 12232 -1424
rect 386 -1517 402 -1483
rect 862 -1517 878 -1483
rect 1244 -1517 1260 -1483
rect 1720 -1517 1736 -1483
rect 2102 -1517 2118 -1483
rect 2578 -1517 2594 -1483
rect 2960 -1517 2976 -1483
rect 3436 -1517 3452 -1483
rect 3818 -1517 3834 -1483
rect 4294 -1517 4310 -1483
rect 4676 -1517 4692 -1483
rect 5152 -1517 5168 -1483
rect 5534 -1517 5550 -1483
rect 6010 -1517 6026 -1483
rect 6392 -1517 6408 -1483
rect 6868 -1517 6884 -1483
rect 7250 -1517 7266 -1483
rect 7726 -1517 7742 -1483
rect 8108 -1517 8124 -1483
rect 8584 -1517 8600 -1483
rect 8966 -1517 8982 -1483
rect 9442 -1517 9458 -1483
rect 9824 -1517 9840 -1483
rect 10300 -1517 10316 -1483
rect 10682 -1517 10698 -1483
rect 11158 -1517 11174 -1483
rect 11540 -1517 11556 -1483
rect 12016 -1517 12032 -1483
rect 386 -1929 402 -1895
rect 862 -1929 878 -1895
rect 1244 -1929 1260 -1895
rect 1720 -1929 1736 -1895
rect 2102 -1929 2118 -1895
rect 2578 -1929 2594 -1895
rect 2960 -1929 2976 -1895
rect 3436 -1929 3452 -1895
rect 3818 -1929 3834 -1895
rect 4294 -1929 4310 -1895
rect 4676 -1929 4692 -1895
rect 5152 -1929 5168 -1895
rect 5534 -1929 5550 -1895
rect 6010 -1929 6026 -1895
rect 6392 -1929 6408 -1895
rect 6868 -1929 6884 -1895
rect 7250 -1929 7266 -1895
rect 7726 -1929 7742 -1895
rect 8108 -1929 8124 -1895
rect 8584 -1929 8600 -1895
rect 8966 -1929 8982 -1895
rect 9442 -1929 9458 -1895
rect 9824 -1929 9840 -1895
rect 10300 -1929 10316 -1895
rect 10682 -1929 10698 -1895
rect 11158 -1929 11174 -1895
rect 11540 -1929 11556 -1895
rect 12016 -1929 12032 -1895
rect 186 -1988 220 -1972
rect 186 -3180 220 -3164
rect 1044 -1988 1078 -1972
rect 1044 -3180 1078 -3164
rect 1902 -1988 1936 -1972
rect 1902 -3180 1936 -3164
rect 2760 -1988 2794 -1972
rect 2760 -3180 2794 -3164
rect 3618 -1988 3652 -1972
rect 3618 -3180 3652 -3164
rect 4476 -1988 4510 -1972
rect 4476 -3180 4510 -3164
rect 5334 -1988 5368 -1972
rect 5334 -3180 5368 -3164
rect 6192 -1988 6226 -1972
rect 6192 -3180 6226 -3164
rect 7050 -1988 7084 -1972
rect 7050 -3180 7084 -3164
rect 7908 -1988 7942 -1972
rect 7908 -3180 7942 -3164
rect 8766 -1988 8800 -1972
rect 8766 -3180 8800 -3164
rect 9624 -1988 9658 -1972
rect 9624 -3180 9658 -3164
rect 10482 -1988 10516 -1972
rect 10482 -3180 10516 -3164
rect 11340 -1988 11374 -1972
rect 11340 -3180 11374 -3164
rect 12198 -1988 12232 -1972
rect 12198 -3180 12232 -3164
rect 386 -3257 402 -3223
rect 862 -3257 878 -3223
rect 1244 -3257 1260 -3223
rect 1720 -3257 1736 -3223
rect 2102 -3257 2118 -3223
rect 2578 -3257 2594 -3223
rect 2960 -3257 2976 -3223
rect 3436 -3257 3452 -3223
rect 3818 -3257 3834 -3223
rect 4294 -3257 4310 -3223
rect 4676 -3257 4692 -3223
rect 5152 -3257 5168 -3223
rect 5534 -3257 5550 -3223
rect 6010 -3257 6026 -3223
rect 6392 -3257 6408 -3223
rect 6868 -3257 6884 -3223
rect 7250 -3257 7266 -3223
rect 7726 -3257 7742 -3223
rect 8108 -3257 8124 -3223
rect 8584 -3257 8600 -3223
rect 8966 -3257 8982 -3223
rect 9442 -3257 9458 -3223
rect 9824 -3257 9840 -3223
rect 10300 -3257 10316 -3223
rect 10682 -3257 10698 -3223
rect 11158 -3257 11174 -3223
rect 11540 -3257 11556 -3223
rect 12016 -3257 12032 -3223
rect 386 -3669 402 -3635
rect 862 -3669 878 -3635
rect 1244 -3669 1260 -3635
rect 1720 -3669 1736 -3635
rect 2102 -3669 2118 -3635
rect 2578 -3669 2594 -3635
rect 2960 -3669 2976 -3635
rect 3436 -3669 3452 -3635
rect 3818 -3669 3834 -3635
rect 4294 -3669 4310 -3635
rect 4676 -3669 4692 -3635
rect 5152 -3669 5168 -3635
rect 5534 -3669 5550 -3635
rect 6010 -3669 6026 -3635
rect 6392 -3669 6408 -3635
rect 6868 -3669 6884 -3635
rect 7250 -3669 7266 -3635
rect 7726 -3669 7742 -3635
rect 8108 -3669 8124 -3635
rect 8584 -3669 8600 -3635
rect 8966 -3669 8982 -3635
rect 9442 -3669 9458 -3635
rect 9824 -3669 9840 -3635
rect 10300 -3669 10316 -3635
rect 10682 -3669 10698 -3635
rect 11158 -3669 11174 -3635
rect 11540 -3669 11556 -3635
rect 12016 -3669 12032 -3635
rect 186 -3728 220 -3712
rect 186 -4920 220 -4904
rect 1044 -3728 1078 -3712
rect 1044 -4920 1078 -4904
rect 1902 -3728 1936 -3712
rect 1902 -4920 1936 -4904
rect 2760 -3728 2794 -3712
rect 2760 -4920 2794 -4904
rect 3618 -3728 3652 -3712
rect 3618 -4920 3652 -4904
rect 4476 -3728 4510 -3712
rect 4476 -4920 4510 -4904
rect 5334 -3728 5368 -3712
rect 5334 -4920 5368 -4904
rect 6192 -3728 6226 -3712
rect 6192 -4920 6226 -4904
rect 7050 -3728 7084 -3712
rect 7050 -4920 7084 -4904
rect 7908 -3728 7942 -3712
rect 7908 -4920 7942 -4904
rect 8766 -3728 8800 -3712
rect 8766 -4920 8800 -4904
rect 9624 -3728 9658 -3712
rect 9624 -4920 9658 -4904
rect 10482 -3728 10516 -3712
rect 10482 -4920 10516 -4904
rect 11340 -3728 11374 -3712
rect 11340 -4920 11374 -4904
rect 12198 -3728 12232 -3712
rect 12198 -4920 12232 -4904
rect 386 -4997 402 -4963
rect 862 -4997 878 -4963
rect 1244 -4997 1260 -4963
rect 1720 -4997 1736 -4963
rect 2102 -4997 2118 -4963
rect 2578 -4997 2594 -4963
rect 2960 -4997 2976 -4963
rect 3436 -4997 3452 -4963
rect 3818 -4997 3834 -4963
rect 4294 -4997 4310 -4963
rect 4676 -4997 4692 -4963
rect 5152 -4997 5168 -4963
rect 5534 -4997 5550 -4963
rect 6010 -4997 6026 -4963
rect 6392 -4997 6408 -4963
rect 6868 -4997 6884 -4963
rect 7250 -4997 7266 -4963
rect 7726 -4997 7742 -4963
rect 8108 -4997 8124 -4963
rect 8584 -4997 8600 -4963
rect 8966 -4997 8982 -4963
rect 9442 -4997 9458 -4963
rect 9824 -4997 9840 -4963
rect 10300 -4997 10316 -4963
rect 10682 -4997 10698 -4963
rect 11158 -4997 11174 -4963
rect 11540 -4997 11556 -4963
rect 12016 -4997 12032 -4963
rect 386 -5409 402 -5375
rect 862 -5409 878 -5375
rect 1244 -5409 1260 -5375
rect 1720 -5409 1736 -5375
rect 2102 -5409 2118 -5375
rect 2578 -5409 2594 -5375
rect 2960 -5409 2976 -5375
rect 3436 -5409 3452 -5375
rect 3818 -5409 3834 -5375
rect 4294 -5409 4310 -5375
rect 4676 -5409 4692 -5375
rect 5152 -5409 5168 -5375
rect 5534 -5409 5550 -5375
rect 6010 -5409 6026 -5375
rect 6392 -5409 6408 -5375
rect 6868 -5409 6884 -5375
rect 7250 -5409 7266 -5375
rect 7726 -5409 7742 -5375
rect 8108 -5409 8124 -5375
rect 8584 -5409 8600 -5375
rect 8966 -5409 8982 -5375
rect 9442 -5409 9458 -5375
rect 9824 -5409 9840 -5375
rect 10300 -5409 10316 -5375
rect 10682 -5409 10698 -5375
rect 11158 -5409 11174 -5375
rect 11540 -5409 11556 -5375
rect 12016 -5409 12032 -5375
rect 186 -5468 220 -5452
rect 186 -6660 220 -6644
rect 1044 -5468 1078 -5452
rect 1044 -6660 1078 -6644
rect 1902 -5468 1936 -5452
rect 1902 -6660 1936 -6644
rect 2760 -5468 2794 -5452
rect 2760 -6660 2794 -6644
rect 3618 -5468 3652 -5452
rect 3618 -6660 3652 -6644
rect 4476 -5468 4510 -5452
rect 4476 -6660 4510 -6644
rect 5334 -5468 5368 -5452
rect 5334 -6660 5368 -6644
rect 6192 -5468 6226 -5452
rect 6192 -6660 6226 -6644
rect 7050 -5468 7084 -5452
rect 7050 -6660 7084 -6644
rect 7908 -5468 7942 -5452
rect 7908 -6660 7942 -6644
rect 8766 -5468 8800 -5452
rect 8766 -6660 8800 -6644
rect 9624 -5468 9658 -5452
rect 9624 -6660 9658 -6644
rect 10482 -5468 10516 -5452
rect 10482 -6660 10516 -6644
rect 11340 -5468 11374 -5452
rect 11340 -6660 11374 -6644
rect 12198 -5468 12232 -5452
rect 12198 -6660 12232 -6644
rect 386 -6737 402 -6703
rect 862 -6737 878 -6703
rect 1244 -6737 1260 -6703
rect 1720 -6737 1736 -6703
rect 2102 -6737 2118 -6703
rect 2578 -6737 2594 -6703
rect 2960 -6737 2976 -6703
rect 3436 -6737 3452 -6703
rect 3818 -6737 3834 -6703
rect 4294 -6737 4310 -6703
rect 4676 -6737 4692 -6703
rect 5152 -6737 5168 -6703
rect 5534 -6737 5550 -6703
rect 6010 -6737 6026 -6703
rect 6392 -6737 6408 -6703
rect 6868 -6737 6884 -6703
rect 7250 -6737 7266 -6703
rect 7726 -6737 7742 -6703
rect 8108 -6737 8124 -6703
rect 8584 -6737 8600 -6703
rect 8966 -6737 8982 -6703
rect 9442 -6737 9458 -6703
rect 9824 -6737 9840 -6703
rect 10300 -6737 10316 -6703
rect 10682 -6737 10698 -6703
rect 11158 -6737 11174 -6703
rect 11540 -6737 11556 -6703
rect 12016 -6737 12032 -6703
rect -362 -7542 -262 -7380
rect 12522 -7542 12622 -7380
rect -362 -7940 -262 -7778
rect 12522 -7940 12622 -7778
rect 5030 -8422 5046 -8388
rect 5266 -8422 5282 -8388
rect 5488 -8422 5504 -8388
rect 5724 -8422 5740 -8388
rect 5946 -8422 5962 -8388
rect 6182 -8422 6198 -8388
rect 6404 -8422 6420 -8388
rect 6640 -8422 6656 -8388
rect 6862 -8422 6878 -8388
rect 7098 -8422 7114 -8388
rect 7320 -8422 7336 -8388
rect 7556 -8422 7572 -8388
rect 4910 -8472 4944 -8456
rect 4910 -8864 4944 -8848
rect 5368 -8472 5402 -8456
rect 5368 -8864 5402 -8848
rect 5826 -8472 5860 -8456
rect 5826 -8864 5860 -8848
rect 6284 -8472 6318 -8456
rect 6284 -8864 6318 -8848
rect 6742 -8472 6776 -8456
rect 6742 -8864 6776 -8848
rect 7200 -8472 7234 -8456
rect 7200 -8864 7234 -8848
rect 7658 -8472 7692 -8456
rect 7658 -8864 7692 -8848
rect 5030 -8932 5046 -8898
rect 5266 -8932 5282 -8898
rect 5488 -8932 5504 -8898
rect 5724 -8932 5740 -8898
rect 5946 -8932 5962 -8898
rect 6182 -8932 6198 -8898
rect 6404 -8932 6420 -8898
rect 6640 -8932 6656 -8898
rect 6862 -8932 6878 -8898
rect 7098 -8932 7114 -8898
rect 7320 -8932 7336 -8898
rect 7556 -8932 7572 -8898
rect 5030 -9222 5046 -9188
rect 5266 -9222 5282 -9188
rect 5488 -9222 5504 -9188
rect 5724 -9222 5740 -9188
rect 5946 -9222 5962 -9188
rect 6182 -9222 6198 -9188
rect 6404 -9222 6420 -9188
rect 6640 -9222 6656 -9188
rect 6862 -9222 6878 -9188
rect 7098 -9222 7114 -9188
rect 7320 -9222 7336 -9188
rect 7556 -9222 7572 -9188
rect 4910 -9272 4944 -9256
rect 4910 -9664 4944 -9648
rect 5368 -9272 5402 -9256
rect 5368 -9664 5402 -9648
rect 5826 -9272 5860 -9256
rect 5826 -9664 5860 -9648
rect 6284 -9272 6318 -9256
rect 6284 -9664 6318 -9648
rect 6742 -9272 6776 -9256
rect 6742 -9664 6776 -9648
rect 7200 -9272 7234 -9256
rect 7200 -9664 7234 -9648
rect 7658 -9272 7692 -9256
rect 7658 -9664 7692 -9648
rect 5030 -9732 5046 -9698
rect 5266 -9732 5282 -9698
rect 5488 -9732 5504 -9698
rect 5724 -9732 5740 -9698
rect 5946 -9732 5962 -9698
rect 6182 -9732 6198 -9698
rect 6404 -9732 6420 -9698
rect 6640 -9732 6656 -9698
rect 6862 -9732 6878 -9698
rect 7098 -9732 7114 -9698
rect 7320 -9732 7336 -9698
rect 7556 -9732 7572 -9698
rect -362 -10822 -262 -10660
rect 12522 -10822 12622 -10660
<< viali >>
rect -262 2822 -200 2922
rect -200 2822 12460 2922
rect 12460 2822 12522 2922
rect -362 -7119 -262 2299
rect 440 1551 824 1585
rect 1298 1551 1682 1585
rect 2156 1551 2540 1585
rect 3014 1551 3398 1585
rect 3872 1551 4256 1585
rect 4730 1551 5114 1585
rect 5588 1551 5972 1585
rect 6446 1551 6830 1585
rect 7304 1551 7688 1585
rect 8162 1551 8546 1585
rect 9020 1551 9404 1585
rect 9878 1551 10262 1585
rect 10736 1551 11120 1585
rect 11594 1551 11978 1585
rect 186 316 220 1492
rect 1044 316 1078 1492
rect 1902 316 1936 1492
rect 2760 316 2794 1492
rect 3618 316 3652 1492
rect 4476 316 4510 1492
rect 5334 316 5368 1492
rect 6192 316 6226 1492
rect 7050 316 7084 1492
rect 7908 316 7942 1492
rect 8766 316 8800 1492
rect 9624 316 9658 1492
rect 10482 316 10516 1492
rect 11340 316 11374 1492
rect 12198 316 12232 1492
rect 440 223 824 257
rect 1298 223 1682 257
rect 2156 223 2540 257
rect 3014 223 3398 257
rect 3872 223 4256 257
rect 4730 223 5114 257
rect 5588 223 5972 257
rect 6446 223 6830 257
rect 7304 223 7688 257
rect 8162 223 8546 257
rect 9020 223 9404 257
rect 9878 223 10262 257
rect 10736 223 11120 257
rect 11594 223 11978 257
rect 440 -189 824 -155
rect 1298 -189 1682 -155
rect 2156 -189 2540 -155
rect 3014 -189 3398 -155
rect 3872 -189 4256 -155
rect 4730 -189 5114 -155
rect 5588 -189 5972 -155
rect 6446 -189 6830 -155
rect 7304 -189 7688 -155
rect 8162 -189 8546 -155
rect 9020 -189 9404 -155
rect 9878 -189 10262 -155
rect 10736 -189 11120 -155
rect 11594 -189 11978 -155
rect 186 -1424 220 -248
rect 1044 -1424 1078 -248
rect 1902 -1424 1936 -248
rect 2760 -1424 2794 -248
rect 3618 -1424 3652 -248
rect 4476 -1424 4510 -248
rect 5334 -1424 5368 -248
rect 6192 -1424 6226 -248
rect 7050 -1424 7084 -248
rect 7908 -1424 7942 -248
rect 8766 -1424 8800 -248
rect 9624 -1424 9658 -248
rect 10482 -1424 10516 -248
rect 11340 -1424 11374 -248
rect 12198 -1424 12232 -248
rect 440 -1517 824 -1483
rect 1298 -1517 1682 -1483
rect 2156 -1517 2540 -1483
rect 3014 -1517 3398 -1483
rect 3872 -1517 4256 -1483
rect 4730 -1517 5114 -1483
rect 5588 -1517 5972 -1483
rect 6446 -1517 6830 -1483
rect 7304 -1517 7688 -1483
rect 8162 -1517 8546 -1483
rect 9020 -1517 9404 -1483
rect 9878 -1517 10262 -1483
rect 10736 -1517 11120 -1483
rect 11594 -1517 11978 -1483
rect 440 -1929 824 -1895
rect 1298 -1929 1682 -1895
rect 2156 -1929 2540 -1895
rect 3014 -1929 3398 -1895
rect 3872 -1929 4256 -1895
rect 4730 -1929 5114 -1895
rect 5588 -1929 5972 -1895
rect 6446 -1929 6830 -1895
rect 7304 -1929 7688 -1895
rect 8162 -1929 8546 -1895
rect 9020 -1929 9404 -1895
rect 9878 -1929 10262 -1895
rect 10736 -1929 11120 -1895
rect 11594 -1929 11978 -1895
rect 186 -3164 220 -1988
rect 1044 -3164 1078 -1988
rect 1902 -3164 1936 -1988
rect 2760 -3164 2794 -1988
rect 3618 -3164 3652 -1988
rect 4476 -3164 4510 -1988
rect 5334 -3164 5368 -1988
rect 6192 -3164 6226 -1988
rect 7050 -3164 7084 -1988
rect 7908 -3164 7942 -1988
rect 8766 -3164 8800 -1988
rect 9624 -3164 9658 -1988
rect 10482 -3164 10516 -1988
rect 11340 -3164 11374 -1988
rect 12198 -3164 12232 -1988
rect 440 -3257 824 -3223
rect 1298 -3257 1682 -3223
rect 2156 -3257 2540 -3223
rect 3014 -3257 3398 -3223
rect 3872 -3257 4256 -3223
rect 4730 -3257 5114 -3223
rect 5588 -3257 5972 -3223
rect 6446 -3257 6830 -3223
rect 7304 -3257 7688 -3223
rect 8162 -3257 8546 -3223
rect 9020 -3257 9404 -3223
rect 9878 -3257 10262 -3223
rect 10736 -3257 11120 -3223
rect 11594 -3257 11978 -3223
rect 440 -3669 824 -3635
rect 1298 -3669 1682 -3635
rect 2156 -3669 2540 -3635
rect 3014 -3669 3398 -3635
rect 3872 -3669 4256 -3635
rect 4730 -3669 5114 -3635
rect 5588 -3669 5972 -3635
rect 6446 -3669 6830 -3635
rect 7304 -3669 7688 -3635
rect 8162 -3669 8546 -3635
rect 9020 -3669 9404 -3635
rect 9878 -3669 10262 -3635
rect 10736 -3669 11120 -3635
rect 11594 -3669 11978 -3635
rect 186 -4904 220 -3728
rect 1044 -4904 1078 -3728
rect 1902 -4904 1936 -3728
rect 2760 -4904 2794 -3728
rect 3618 -4904 3652 -3728
rect 4476 -4904 4510 -3728
rect 5334 -4904 5368 -3728
rect 6192 -4904 6226 -3728
rect 7050 -4904 7084 -3728
rect 7908 -4904 7942 -3728
rect 8766 -4904 8800 -3728
rect 9624 -4904 9658 -3728
rect 10482 -4904 10516 -3728
rect 11340 -4904 11374 -3728
rect 12198 -4904 12232 -3728
rect 440 -4997 824 -4963
rect 1298 -4997 1682 -4963
rect 2156 -4997 2540 -4963
rect 3014 -4997 3398 -4963
rect 3872 -4997 4256 -4963
rect 4730 -4997 5114 -4963
rect 5588 -4997 5972 -4963
rect 6446 -4997 6830 -4963
rect 7304 -4997 7688 -4963
rect 8162 -4997 8546 -4963
rect 9020 -4997 9404 -4963
rect 9878 -4997 10262 -4963
rect 10736 -4997 11120 -4963
rect 11594 -4997 11978 -4963
rect 440 -5409 824 -5375
rect 1298 -5409 1682 -5375
rect 2156 -5409 2540 -5375
rect 3014 -5409 3398 -5375
rect 3872 -5409 4256 -5375
rect 4730 -5409 5114 -5375
rect 5588 -5409 5972 -5375
rect 6446 -5409 6830 -5375
rect 7304 -5409 7688 -5375
rect 8162 -5409 8546 -5375
rect 9020 -5409 9404 -5375
rect 9878 -5409 10262 -5375
rect 10736 -5409 11120 -5375
rect 11594 -5409 11978 -5375
rect 186 -6644 220 -5468
rect 1044 -6644 1078 -5468
rect 1902 -6644 1936 -5468
rect 2760 -6644 2794 -5468
rect 3618 -6644 3652 -5468
rect 4476 -6644 4510 -5468
rect 5334 -6644 5368 -5468
rect 6192 -6644 6226 -5468
rect 7050 -6644 7084 -5468
rect 7908 -6644 7942 -5468
rect 8766 -6644 8800 -5468
rect 9624 -6644 9658 -5468
rect 10482 -6644 10516 -5468
rect 11340 -6644 11374 -5468
rect 12198 -6644 12232 -5468
rect 440 -6737 824 -6703
rect 1298 -6737 1682 -6703
rect 2156 -6737 2540 -6703
rect 3014 -6737 3398 -6703
rect 3872 -6737 4256 -6703
rect 4730 -6737 5114 -6703
rect 5588 -6737 5972 -6703
rect 6446 -6737 6830 -6703
rect 7304 -6737 7688 -6703
rect 8162 -6737 8546 -6703
rect 9020 -6737 9404 -6703
rect 9878 -6737 10262 -6703
rect 10736 -6737 11120 -6703
rect 11594 -6737 11978 -6703
rect 12522 -7119 12622 2299
rect -262 -7542 -200 -7442
rect -200 -7542 12460 -7442
rect 12460 -7542 12522 -7442
rect -262 -7878 -200 -7778
rect -200 -7878 12460 -7778
rect 12460 -7878 12522 -7778
rect -362 -10570 -262 -7982
rect 5064 -8422 5248 -8388
rect 5522 -8422 5706 -8388
rect 5980 -8422 6164 -8388
rect 6438 -8422 6622 -8388
rect 6896 -8422 7080 -8388
rect 7354 -8422 7538 -8388
rect 4910 -8848 4944 -8472
rect 5368 -8848 5402 -8472
rect 5826 -8848 5860 -8472
rect 6284 -8848 6318 -8472
rect 6742 -8848 6776 -8472
rect 7200 -8848 7234 -8472
rect 7658 -8848 7692 -8472
rect 5064 -8932 5248 -8898
rect 5522 -8932 5706 -8898
rect 5980 -8932 6164 -8898
rect 6438 -8932 6622 -8898
rect 6896 -8932 7080 -8898
rect 7354 -8932 7538 -8898
rect 5064 -9222 5248 -9188
rect 5522 -9222 5706 -9188
rect 5980 -9222 6164 -9188
rect 6438 -9222 6622 -9188
rect 6896 -9222 7080 -9188
rect 7354 -9222 7538 -9188
rect 4910 -9648 4944 -9272
rect 5368 -9648 5402 -9272
rect 5826 -9648 5860 -9272
rect 6284 -9648 6318 -9272
rect 6742 -9648 6776 -9272
rect 7200 -9648 7234 -9272
rect 7658 -9648 7692 -9272
rect 5064 -9732 5248 -9698
rect 5522 -9732 5706 -9698
rect 5980 -9732 6164 -9698
rect 6438 -9732 6622 -9698
rect 6896 -9732 7080 -9698
rect 7354 -9732 7538 -9698
rect 12522 -10570 12622 -7982
rect -262 -10822 -200 -10722
rect -200 -10822 12460 -10722
rect 12460 -10822 12522 -10722
<< metal1 >>
rect -368 2922 12628 2928
rect -368 2822 -262 2922
rect 12522 2822 12628 2922
rect -368 2816 12628 2822
rect -368 2299 -256 2816
rect 344 2516 354 2816
rect 11906 2516 11916 2816
rect -368 -7119 -362 2299
rect -262 2108 -256 2299
rect 110 2396 12310 2438
rect 110 2232 158 2396
rect 12268 2232 12310 2396
rect 110 2192 12310 2232
rect 12516 2299 12628 2816
rect 172 2110 232 2192
rect 596 2110 656 2192
rect 1032 2110 1092 2192
rect 2746 2110 2806 2192
rect 4466 2110 4526 2192
rect 6174 2110 6234 2192
rect 7894 2110 7954 2192
rect 9608 2110 9668 2192
rect 11326 2110 11386 2192
rect 11754 2110 11814 2192
rect 12186 2110 12246 2192
rect 166 2108 172 2110
rect -262 2050 172 2108
rect 232 2050 238 2110
rect 590 2050 596 2110
rect 656 2050 662 2110
rect 1026 2050 1032 2110
rect 1092 2050 1098 2110
rect 2740 2050 2746 2110
rect 2806 2050 2812 2110
rect 4460 2050 4466 2110
rect 4526 2050 4532 2110
rect 6168 2050 6174 2110
rect 6234 2050 6240 2110
rect 7888 2050 7894 2110
rect 7954 2050 7960 2110
rect 9602 2050 9608 2110
rect 9668 2050 9674 2110
rect 11320 2050 11326 2110
rect 11386 2050 11392 2110
rect 11748 2050 11754 2110
rect 11814 2050 11820 2110
rect 12180 2050 12186 2110
rect 12246 2108 12252 2110
rect 12516 2108 12522 2299
rect 12246 2050 12522 2108
rect -262 2048 232 2050
rect -262 -5150 -256 2048
rect -98 1786 -92 1846
rect -32 1786 -26 1846
rect -92 -50 -32 1786
rect 44 1658 50 1718
rect 110 1658 116 1718
rect 50 56 110 1658
rect 172 1492 232 2048
rect 596 1591 656 2050
rect 428 1585 836 1591
rect 428 1551 440 1585
rect 824 1551 836 1585
rect 428 1545 836 1551
rect 172 1414 186 1492
rect 180 394 186 1414
rect 170 316 186 394
rect 220 1414 232 1492
rect 1032 1492 1092 2050
rect 1452 1922 1458 1982
rect 1518 1922 1524 1982
rect 2306 1922 2312 1982
rect 2372 1922 2378 1982
rect 1458 1591 1518 1922
rect 2312 1591 2372 1922
rect 1286 1585 1694 1591
rect 1286 1551 1298 1585
rect 1682 1551 1694 1585
rect 1286 1545 1694 1551
rect 2144 1585 2552 1591
rect 2144 1551 2156 1585
rect 2540 1551 2552 1585
rect 2144 1545 2552 1551
rect 1032 1414 1044 1492
rect 220 394 226 1414
rect 1038 396 1044 1414
rect 220 316 230 394
rect 170 62 230 316
rect 1030 316 1044 396
rect 1078 1414 1092 1492
rect 1896 1492 1942 1504
rect 1078 396 1084 1414
rect 1896 454 1902 1492
rect 1078 316 1090 396
rect 428 257 836 263
rect 428 223 440 257
rect 824 223 836 257
rect 428 217 836 223
rect 600 62 660 217
rect 1030 62 1090 316
rect 1888 316 1902 454
rect 1936 454 1942 1492
rect 2746 1492 2806 2050
rect 3166 1922 3172 1982
rect 3232 1922 3238 1982
rect 4026 1922 4032 1982
rect 4092 1922 4098 1982
rect 3172 1591 3232 1922
rect 4032 1591 4092 1922
rect 3002 1585 3410 1591
rect 3002 1551 3014 1585
rect 3398 1551 3410 1585
rect 3002 1545 3410 1551
rect 3860 1585 4268 1591
rect 3860 1551 3872 1585
rect 4256 1551 4268 1585
rect 3860 1545 4268 1551
rect 2746 1422 2760 1492
rect 1936 316 1948 454
rect 2754 388 2760 1422
rect 1286 257 1694 263
rect 1286 223 1298 257
rect 1682 223 1694 257
rect 1286 217 1694 223
rect 44 -4 50 56
rect 110 -4 116 56
rect 170 -6 1090 62
rect -98 -110 -92 -50
rect -32 -110 -26 -50
rect 170 -248 230 -6
rect 600 -149 660 -6
rect 428 -155 836 -149
rect 428 -189 440 -155
rect 824 -189 836 -155
rect 428 -195 836 -189
rect 170 -1424 186 -248
rect 220 -1424 230 -248
rect -98 -1640 -92 -1580
rect -32 -1640 -26 -1580
rect -92 -3530 -32 -1640
rect 170 -1682 230 -1424
rect 1030 -248 1090 -6
rect 1460 -149 1520 217
rect 1888 156 1948 316
rect 2748 316 2760 388
rect 2794 1422 2806 1492
rect 3612 1492 3658 1504
rect 2794 388 2800 1422
rect 2794 316 2808 388
rect 3612 360 3618 1492
rect 2144 257 2552 263
rect 2144 223 2156 257
rect 2540 223 2552 257
rect 2144 217 2552 223
rect 1882 96 1888 156
rect 1948 96 1954 156
rect 1884 -110 1890 -50
rect 1950 -110 1956 -50
rect 1286 -155 1694 -149
rect 1286 -189 1298 -155
rect 1682 -189 1694 -155
rect 1286 -195 1694 -189
rect 1030 -1424 1044 -248
rect 1078 -1424 1090 -248
rect 1890 -248 1950 -110
rect 2320 -149 2380 217
rect 2144 -155 2552 -149
rect 2144 -189 2156 -155
rect 2540 -189 2552 -155
rect 2144 -195 2552 -189
rect 1890 -298 1902 -248
rect 428 -1483 836 -1477
rect 428 -1517 440 -1483
rect 824 -1517 836 -1483
rect 428 -1523 836 -1517
rect 600 -1682 660 -1523
rect 1030 -1682 1090 -1424
rect 1896 -1424 1902 -298
rect 1936 -298 1950 -248
rect 2748 -248 2808 316
rect 3604 316 3618 360
rect 3652 360 3658 1492
rect 4466 1492 4526 2050
rect 4886 1922 4892 1982
rect 4952 1922 4958 1982
rect 5746 1922 5752 1982
rect 5812 1922 5818 1982
rect 4892 1591 4952 1922
rect 5752 1591 5812 1922
rect 4718 1585 5126 1591
rect 4718 1551 4730 1585
rect 5114 1551 5126 1585
rect 4718 1545 5126 1551
rect 5576 1585 5984 1591
rect 5576 1551 5588 1585
rect 5972 1551 5984 1585
rect 5576 1545 5984 1551
rect 4466 1436 4476 1492
rect 4470 386 4476 1436
rect 3652 316 3664 360
rect 3002 257 3410 263
rect 3002 223 3014 257
rect 3398 223 3410 257
rect 3002 217 3410 223
rect 3180 -149 3240 217
rect 3464 -4 3470 56
rect 3530 -4 3536 56
rect 3604 54 3664 316
rect 4462 316 4476 386
rect 4510 1436 4526 1492
rect 5328 1492 5374 1504
rect 4510 386 4516 1436
rect 5328 420 5334 1492
rect 4510 316 4522 386
rect 3860 257 4268 263
rect 3860 223 3872 257
rect 4256 223 4268 257
rect 3860 217 4268 223
rect 3470 -48 3530 -4
rect 3598 -6 3604 54
rect 3664 -6 3670 54
rect 3470 -108 3664 -48
rect 3002 -155 3410 -149
rect 3002 -189 3014 -155
rect 3398 -189 3410 -155
rect 3002 -195 3410 -189
rect 1936 -1424 1942 -298
rect 1896 -1436 1942 -1424
rect 2748 -1424 2760 -248
rect 2794 -1424 2808 -248
rect 3604 -248 3664 -108
rect 4040 -149 4100 217
rect 3860 -155 4268 -149
rect 3860 -189 3872 -155
rect 4256 -189 4268 -155
rect 3860 -195 4268 -189
rect 3604 -312 3618 -248
rect 1286 -1483 1694 -1477
rect 1286 -1517 1298 -1483
rect 1682 -1517 1694 -1483
rect 1286 -1523 1694 -1517
rect 2144 -1483 2552 -1477
rect 2144 -1517 2156 -1483
rect 2540 -1517 2552 -1483
rect 2144 -1523 2552 -1517
rect 1460 -1678 1520 -1523
rect 170 -1742 1090 -1682
rect 44 -1846 50 -1786
rect 110 -1846 116 -1786
rect 50 -3424 110 -1846
rect 170 -1988 230 -1742
rect 600 -1889 660 -1742
rect 428 -1895 836 -1889
rect 428 -1929 440 -1895
rect 824 -1929 836 -1895
rect 428 -1935 836 -1929
rect 170 -3164 186 -1988
rect 220 -3164 230 -1988
rect 170 -3424 230 -3164
rect 1030 -1988 1090 -1742
rect 1458 -1684 1520 -1678
rect 1518 -1744 1520 -1684
rect 1458 -1750 1520 -1744
rect 1460 -1889 1520 -1750
rect 2320 -1684 2380 -1523
rect 2320 -1889 2380 -1744
rect 1286 -1895 1694 -1889
rect 1286 -1929 1298 -1895
rect 1682 -1929 1694 -1895
rect 1286 -1935 1694 -1929
rect 2144 -1895 2552 -1889
rect 2144 -1929 2156 -1895
rect 2540 -1929 2552 -1895
rect 2144 -1935 2552 -1929
rect 1030 -3164 1044 -1988
rect 1078 -3164 1090 -1988
rect 1896 -1988 1942 -1976
rect 1896 -3026 1902 -1988
rect 428 -3223 836 -3217
rect 428 -3257 440 -3223
rect 824 -3257 836 -3223
rect 428 -3263 836 -3257
rect 600 -3424 660 -3263
rect 1030 -3424 1090 -3164
rect 1888 -3164 1902 -3026
rect 1936 -3026 1942 -1988
rect 2748 -1988 2808 -1424
rect 3612 -1424 3618 -312
rect 3652 -312 3664 -248
rect 4462 -248 4522 316
rect 5318 316 5334 420
rect 5368 420 5374 1492
rect 6174 1492 6234 2050
rect 6606 1922 6612 1982
rect 6672 1922 6678 1982
rect 7466 1922 7472 1982
rect 7532 1922 7538 1982
rect 6612 1591 6672 1922
rect 7472 1591 7532 1922
rect 6434 1585 6842 1591
rect 6434 1551 6446 1585
rect 6830 1551 6842 1585
rect 6434 1545 6842 1551
rect 7292 1585 7700 1591
rect 7292 1551 7304 1585
rect 7688 1551 7700 1585
rect 7292 1545 7700 1551
rect 6174 1436 6192 1492
rect 5368 316 5378 420
rect 4718 257 5126 263
rect 4718 223 4730 257
rect 5114 223 5126 257
rect 4718 217 5126 223
rect 4900 -149 4960 217
rect 5318 54 5378 316
rect 6186 316 6192 1436
rect 6226 1436 6234 1492
rect 7044 1492 7090 1504
rect 6226 316 6232 1436
rect 7044 368 7050 1492
rect 6186 304 6232 316
rect 7038 316 7050 368
rect 7084 368 7090 1492
rect 7894 1492 7954 2050
rect 8326 1922 8332 1982
rect 8392 1922 8398 1982
rect 9166 1922 9172 1982
rect 9232 1922 9238 1982
rect 8332 1591 8392 1922
rect 8746 1658 8752 1718
rect 8812 1658 8818 1718
rect 8150 1585 8558 1591
rect 8150 1551 8162 1585
rect 8546 1551 8558 1585
rect 8150 1545 8558 1551
rect 7894 1416 7908 1492
rect 7902 384 7908 1416
rect 7084 316 7098 368
rect 5576 257 5984 263
rect 5576 223 5588 257
rect 5972 223 5984 257
rect 5576 217 5984 223
rect 6434 257 6842 263
rect 6434 223 6446 257
rect 6830 223 6842 257
rect 6434 217 6842 223
rect 7038 156 7098 316
rect 7894 316 7908 384
rect 7942 1416 7954 1492
rect 8752 1492 8812 1658
rect 9172 1591 9232 1922
rect 9008 1585 9416 1591
rect 9008 1551 9020 1585
rect 9404 1551 9416 1585
rect 9008 1545 9416 1551
rect 7942 384 7948 1416
rect 8752 1342 8766 1492
rect 7942 316 7954 384
rect 7292 257 7700 263
rect 7292 223 7304 257
rect 7688 223 7700 257
rect 7292 217 7700 223
rect 7038 96 7226 156
rect 5318 -6 7096 54
rect 5314 -110 5320 -50
rect 5380 -110 5386 -50
rect 4718 -155 5126 -149
rect 4718 -189 4730 -155
rect 5114 -189 5126 -155
rect 4718 -195 5126 -189
rect 3652 -1424 3658 -312
rect 3612 -1436 3658 -1424
rect 4462 -1424 4476 -248
rect 4510 -1424 4522 -248
rect 5320 -248 5380 -110
rect 7036 -112 7096 -6
rect 7166 -50 7226 96
rect 7160 -110 7166 -50
rect 7226 -110 7232 -50
rect 5576 -155 5984 -149
rect 5576 -189 5588 -155
rect 5972 -189 5984 -155
rect 5576 -195 5984 -189
rect 6434 -155 6842 -149
rect 6434 -189 6446 -155
rect 6830 -189 6842 -155
rect 6434 -195 6842 -189
rect 5320 -406 5334 -248
rect 3002 -1483 3410 -1477
rect 3002 -1517 3014 -1483
rect 3398 -1517 3410 -1483
rect 3002 -1523 3410 -1517
rect 3860 -1483 4268 -1477
rect 3860 -1517 3872 -1483
rect 4256 -1517 4268 -1483
rect 3860 -1523 4268 -1517
rect 3180 -1678 3240 -1523
rect 3180 -1684 3242 -1678
rect 3180 -1744 3182 -1684
rect 3180 -1750 3242 -1744
rect 4040 -1684 4100 -1523
rect 3180 -1889 3240 -1750
rect 4040 -1889 4100 -1744
rect 3002 -1895 3410 -1889
rect 3002 -1929 3014 -1895
rect 3398 -1929 3410 -1895
rect 3002 -1935 3410 -1929
rect 3860 -1895 4268 -1889
rect 3860 -1929 3872 -1895
rect 4256 -1929 4268 -1895
rect 3860 -1935 4268 -1929
rect 1936 -3164 1948 -3026
rect 1286 -3223 1694 -3217
rect 1286 -3257 1298 -3223
rect 1682 -3257 1694 -3223
rect 1286 -3263 1694 -3257
rect 44 -3484 50 -3424
rect 110 -3484 116 -3424
rect 170 -3484 1090 -3424
rect -98 -3590 -92 -3530
rect -32 -3590 -26 -3530
rect 170 -3728 230 -3484
rect 600 -3629 660 -3484
rect 428 -3635 836 -3629
rect 428 -3669 440 -3635
rect 824 -3669 836 -3635
rect 428 -3675 836 -3669
rect 170 -4904 186 -3728
rect 220 -4904 230 -3728
rect 170 -5150 230 -4904
rect 1030 -3728 1090 -3484
rect 1460 -3629 1520 -3263
rect 1888 -3324 1948 -3164
rect 2748 -3164 2760 -1988
rect 2794 -3164 2808 -1988
rect 3612 -1988 3658 -1976
rect 3612 -3120 3618 -1988
rect 2144 -3223 2552 -3217
rect 2144 -3257 2156 -3223
rect 2540 -3257 2552 -3223
rect 2144 -3263 2552 -3257
rect 1882 -3384 1888 -3324
rect 1948 -3384 1954 -3324
rect 1884 -3590 1890 -3530
rect 1950 -3590 1956 -3530
rect 1286 -3635 1694 -3629
rect 1286 -3669 1298 -3635
rect 1682 -3669 1694 -3635
rect 1286 -3675 1694 -3669
rect 1030 -4904 1044 -3728
rect 1078 -4904 1090 -3728
rect 1890 -3728 1950 -3590
rect 2320 -3629 2380 -3263
rect 2144 -3635 2552 -3629
rect 2144 -3669 2156 -3635
rect 2540 -3669 2552 -3635
rect 2144 -3675 2552 -3669
rect 1890 -3778 1902 -3728
rect 428 -4963 836 -4957
rect 428 -4997 440 -4963
rect 824 -4997 836 -4963
rect 428 -5003 836 -4997
rect 600 -5150 660 -5003
rect 1030 -5150 1090 -4904
rect 1896 -4904 1902 -3778
rect 1936 -3778 1950 -3728
rect 2748 -3728 2808 -3164
rect 3604 -3164 3618 -3120
rect 3652 -3120 3658 -1988
rect 4462 -1988 4522 -1424
rect 5328 -1424 5334 -406
rect 5368 -406 5380 -248
rect 6186 -248 6232 -236
rect 6186 -332 6192 -248
rect 5368 -1424 5374 -406
rect 5328 -1436 5374 -1424
rect 6180 -1424 6192 -332
rect 6226 -332 6232 -248
rect 7036 -248 7098 -112
rect 7480 -149 7540 217
rect 7292 -155 7700 -149
rect 7292 -189 7304 -155
rect 7688 -189 7700 -155
rect 7292 -195 7700 -189
rect 7036 -280 7050 -248
rect 7038 -294 7050 -280
rect 6226 -1424 6240 -332
rect 4718 -1483 5126 -1477
rect 4718 -1517 4730 -1483
rect 5114 -1517 5126 -1483
rect 4718 -1523 5126 -1517
rect 5576 -1483 5984 -1477
rect 5576 -1517 5588 -1483
rect 5972 -1517 5984 -1483
rect 5576 -1523 5984 -1517
rect 4900 -1684 4960 -1523
rect 4900 -1889 4960 -1744
rect 5744 -1684 5804 -1523
rect 5744 -1889 5804 -1744
rect 4718 -1895 5126 -1889
rect 4718 -1929 4730 -1895
rect 5114 -1929 5126 -1895
rect 4718 -1935 5126 -1929
rect 5576 -1895 5984 -1889
rect 5576 -1929 5588 -1895
rect 5972 -1929 5984 -1895
rect 5576 -1935 5984 -1929
rect 5744 -1936 5804 -1935
rect 3652 -3164 3664 -3120
rect 3002 -3223 3410 -3217
rect 3002 -3257 3014 -3223
rect 3398 -3257 3410 -3223
rect 3002 -3263 3410 -3257
rect 3180 -3629 3240 -3263
rect 3464 -3484 3470 -3424
rect 3530 -3484 3536 -3424
rect 3604 -3426 3664 -3164
rect 4462 -3164 4476 -1988
rect 4510 -3164 4522 -1988
rect 5328 -1988 5374 -1976
rect 5328 -3060 5334 -1988
rect 3860 -3223 4268 -3217
rect 3860 -3257 3872 -3223
rect 4256 -3257 4268 -3223
rect 3860 -3263 4268 -3257
rect 3470 -3528 3530 -3484
rect 3598 -3486 3604 -3426
rect 3664 -3486 3670 -3426
rect 3470 -3588 3664 -3528
rect 3002 -3635 3410 -3629
rect 3002 -3669 3014 -3635
rect 3398 -3669 3410 -3635
rect 3002 -3675 3410 -3669
rect 1936 -4904 1942 -3778
rect 1896 -4916 1942 -4904
rect 2748 -4904 2760 -3728
rect 2794 -4904 2808 -3728
rect 3604 -3728 3664 -3588
rect 4040 -3629 4100 -3263
rect 4462 -3532 4522 -3164
rect 5318 -3164 5334 -3060
rect 5368 -3060 5374 -1988
rect 6180 -1988 6240 -1424
rect 7044 -1424 7050 -294
rect 7084 -294 7098 -248
rect 7894 -248 7954 316
rect 8760 316 8766 1342
rect 8800 1342 8812 1492
rect 9608 1492 9668 2050
rect 10024 1922 10030 1982
rect 10090 1922 10096 1982
rect 10886 1922 10892 1982
rect 10952 1922 10958 1982
rect 10030 1591 10090 1922
rect 10462 1786 10468 1846
rect 10528 1786 10534 1846
rect 9866 1585 10274 1591
rect 9866 1551 9878 1585
rect 10262 1551 10274 1585
rect 9866 1545 10274 1551
rect 9608 1414 9624 1492
rect 8800 316 8806 1342
rect 9618 390 9624 1414
rect 8760 304 8806 316
rect 9608 316 9624 390
rect 9658 1414 9668 1492
rect 10468 1492 10528 1786
rect 10892 1591 10952 1922
rect 10724 1585 11132 1591
rect 10724 1551 10736 1585
rect 11120 1551 11132 1585
rect 10724 1545 11132 1551
rect 9658 390 9664 1414
rect 10468 1356 10482 1492
rect 9658 316 9668 390
rect 8150 257 8558 263
rect 8150 223 8162 257
rect 8546 223 8558 257
rect 8150 217 8558 223
rect 9008 257 9416 263
rect 9008 223 9020 257
rect 9404 223 9416 257
rect 9008 217 9416 223
rect 8336 -149 8396 217
rect 8750 -6 8756 54
rect 8816 -6 8822 54
rect 8150 -155 8558 -149
rect 8150 -189 8162 -155
rect 8546 -189 8558 -155
rect 8150 -195 8558 -189
rect 7084 -1424 7090 -294
rect 7044 -1436 7090 -1424
rect 7894 -1424 7908 -248
rect 7942 -1424 7954 -248
rect 8756 -248 8816 -6
rect 9192 -149 9252 217
rect 9008 -155 9416 -149
rect 9008 -189 9020 -155
rect 9404 -189 9416 -155
rect 9008 -195 9416 -189
rect 8756 -340 8766 -248
rect 6434 -1483 6842 -1477
rect 6434 -1517 6446 -1483
rect 6830 -1517 6842 -1483
rect 6434 -1523 6842 -1517
rect 7292 -1483 7700 -1477
rect 7292 -1517 7304 -1483
rect 7688 -1517 7700 -1483
rect 7292 -1523 7700 -1517
rect 6614 -1684 6674 -1523
rect 6614 -1889 6674 -1744
rect 7480 -1684 7540 -1523
rect 7480 -1889 7540 -1744
rect 6434 -1895 6842 -1889
rect 6434 -1929 6446 -1895
rect 6830 -1929 6842 -1895
rect 6434 -1935 6842 -1929
rect 7292 -1895 7700 -1889
rect 7292 -1929 7304 -1895
rect 7688 -1929 7700 -1895
rect 7292 -1935 7700 -1929
rect 5368 -3164 5378 -3060
rect 4718 -3223 5126 -3217
rect 4718 -3257 4730 -3223
rect 5114 -3257 5126 -3223
rect 4718 -3263 5126 -3257
rect 3860 -3635 4268 -3629
rect 3860 -3669 3872 -3635
rect 4256 -3669 4268 -3635
rect 3860 -3675 4268 -3669
rect 3604 -3792 3618 -3728
rect 1286 -4963 1694 -4957
rect 1286 -4997 1298 -4963
rect 1682 -4997 1694 -4963
rect 1286 -5003 1694 -4997
rect 2144 -4963 2552 -4957
rect 2144 -4997 2156 -4963
rect 2540 -4997 2552 -4963
rect 2144 -5003 2552 -4997
rect 1460 -5050 1520 -5003
rect 2320 -5050 2380 -5003
rect 1454 -5110 1460 -5050
rect 1520 -5110 1526 -5050
rect -262 -5210 1090 -5150
rect -262 -7076 -256 -5210
rect 170 -5468 230 -5210
rect 600 -5369 660 -5210
rect 428 -5375 836 -5369
rect 428 -5409 440 -5375
rect 824 -5409 836 -5375
rect 428 -5415 836 -5409
rect 170 -6644 186 -5468
rect 220 -6644 230 -5468
rect 1030 -5468 1090 -5210
rect 1460 -5369 1520 -5110
rect 1882 -5328 1888 -5268
rect 1948 -5328 1954 -5268
rect 1286 -5375 1694 -5369
rect 1286 -5409 1298 -5375
rect 1682 -5409 1694 -5375
rect 1286 -5415 1694 -5409
rect 1030 -5542 1044 -5468
rect 1038 -6548 1044 -5542
rect 170 -7070 230 -6644
rect 1030 -6644 1044 -6548
rect 1078 -5542 1090 -5468
rect 1888 -5468 1948 -5328
rect 2320 -5369 2380 -5110
rect 2144 -5375 2552 -5369
rect 2144 -5409 2156 -5375
rect 2540 -5409 2552 -5375
rect 2144 -5415 2552 -5409
rect 1078 -6548 1084 -5542
rect 1888 -5580 1902 -5468
rect 1078 -6644 1090 -6548
rect 428 -6703 836 -6697
rect 428 -6737 440 -6703
rect 824 -6737 836 -6703
rect 428 -6743 836 -6737
rect 590 -7070 650 -6743
rect 1030 -7070 1090 -6644
rect 1896 -6644 1902 -5580
rect 1936 -5580 1948 -5468
rect 2748 -5468 2808 -4904
rect 3612 -4904 3618 -3792
rect 3652 -3792 3664 -3728
rect 4462 -3728 4522 -3592
rect 4900 -3629 4960 -3263
rect 5318 -3426 5378 -3164
rect 6180 -3164 6192 -1988
rect 6226 -3164 6240 -1988
rect 7044 -1988 7090 -1976
rect 7044 -3112 7050 -1988
rect 6180 -3196 6240 -3164
rect 5576 -3223 5984 -3217
rect 5576 -3257 5588 -3223
rect 5972 -3257 5984 -3223
rect 5576 -3263 5984 -3257
rect 7038 -3164 7050 -3112
rect 7084 -3112 7090 -1988
rect 7894 -1988 7954 -1424
rect 8760 -1424 8766 -340
rect 8800 -340 8816 -248
rect 9608 -248 9668 316
rect 10476 316 10482 1356
rect 10516 1356 10528 1492
rect 11326 1492 11386 2050
rect 11754 1591 11814 2050
rect 12186 2048 12522 2050
rect 11582 1585 11990 1591
rect 11582 1551 11594 1585
rect 11978 1551 11990 1585
rect 11582 1545 11990 1551
rect 11754 1544 11814 1545
rect 11326 1432 11340 1492
rect 10516 316 10522 1356
rect 11334 406 11340 1432
rect 10476 304 10522 316
rect 11326 316 11340 406
rect 11374 1432 11386 1492
rect 12186 1492 12246 2048
rect 11374 406 11380 1432
rect 12186 1418 12198 1492
rect 11374 316 11386 406
rect 12192 394 12198 1418
rect 9866 257 10274 263
rect 9866 223 9878 257
rect 10262 223 10274 257
rect 9866 217 10274 223
rect 10724 257 11132 263
rect 10724 223 10736 257
rect 11120 223 11132 257
rect 10724 217 11132 223
rect 10048 -149 10108 217
rect 10464 96 10470 156
rect 10530 96 10536 156
rect 9866 -155 10274 -149
rect 9866 -189 9878 -155
rect 10262 -189 10274 -155
rect 9866 -195 10274 -189
rect 8800 -1424 8806 -340
rect 8760 -1436 8806 -1424
rect 9608 -1424 9624 -248
rect 9658 -1424 9668 -248
rect 10470 -248 10530 96
rect 10904 -149 10964 217
rect 11326 66 11386 316
rect 12184 316 12198 394
rect 12232 1418 12246 1492
rect 12232 394 12238 1418
rect 12232 316 12244 394
rect 11582 257 11990 263
rect 11582 223 11594 257
rect 11978 223 11990 257
rect 11582 217 11990 223
rect 11750 66 11810 217
rect 12184 66 12244 316
rect 12516 66 12522 2048
rect 11326 6 12522 66
rect 10724 -155 11132 -149
rect 10724 -189 10736 -155
rect 11120 -189 11132 -155
rect 10724 -195 11132 -189
rect 10470 -304 10482 -248
rect 8150 -1483 8558 -1477
rect 8150 -1517 8162 -1483
rect 8546 -1517 8558 -1483
rect 8150 -1523 8558 -1517
rect 9008 -1483 9416 -1477
rect 9008 -1517 9020 -1483
rect 9404 -1517 9416 -1483
rect 9008 -1523 9416 -1517
rect 8336 -1684 8396 -1523
rect 8336 -1889 8396 -1744
rect 9192 -1684 9252 -1523
rect 8746 -1846 8752 -1786
rect 8812 -1846 8818 -1786
rect 8150 -1895 8558 -1889
rect 8150 -1929 8162 -1895
rect 8546 -1929 8558 -1895
rect 8150 -1935 8558 -1929
rect 7084 -3164 7098 -3112
rect 6180 -3262 6240 -3256
rect 6434 -3223 6842 -3217
rect 6434 -3257 6446 -3223
rect 6830 -3257 6842 -3223
rect 6434 -3263 6842 -3257
rect 7038 -3324 7098 -3164
rect 7894 -3164 7908 -1988
rect 7942 -3164 7954 -1988
rect 8752 -1988 8812 -1846
rect 9192 -1889 9252 -1744
rect 9008 -1895 9416 -1889
rect 9008 -1929 9020 -1895
rect 9404 -1929 9416 -1895
rect 9008 -1935 9416 -1929
rect 8752 -2138 8766 -1988
rect 7292 -3223 7700 -3217
rect 7292 -3257 7304 -3223
rect 7688 -3257 7700 -3223
rect 7292 -3263 7700 -3257
rect 7038 -3384 7226 -3324
rect 5318 -3486 7096 -3426
rect 5314 -3590 5320 -3530
rect 5380 -3590 5386 -3530
rect 4718 -3635 5126 -3629
rect 4718 -3669 4730 -3635
rect 5114 -3669 5126 -3635
rect 4718 -3675 5126 -3669
rect 3652 -4904 3658 -3792
rect 3612 -4916 3658 -4904
rect 4462 -4904 4476 -3728
rect 4510 -4904 4522 -3728
rect 5320 -3728 5380 -3590
rect 7036 -3592 7096 -3486
rect 7166 -3530 7226 -3384
rect 7160 -3590 7166 -3530
rect 7226 -3590 7232 -3530
rect 5576 -3635 5984 -3629
rect 5576 -3669 5588 -3635
rect 5972 -3669 5984 -3635
rect 5576 -3675 5984 -3669
rect 6434 -3635 6842 -3629
rect 6434 -3669 6446 -3635
rect 6830 -3669 6842 -3635
rect 6434 -3675 6842 -3669
rect 5320 -3886 5334 -3728
rect 3002 -4963 3410 -4957
rect 3002 -4997 3014 -4963
rect 3398 -4997 3410 -4963
rect 3002 -5003 3410 -4997
rect 3860 -4963 4268 -4957
rect 3860 -4997 3872 -4963
rect 4256 -4997 4268 -4963
rect 3860 -5003 4268 -4997
rect 3180 -5044 3240 -5003
rect 3176 -5050 3240 -5044
rect 3236 -5110 3240 -5050
rect 3176 -5116 3240 -5110
rect 3180 -5369 3240 -5116
rect 4040 -5044 4100 -5003
rect 4040 -5050 4102 -5044
rect 4040 -5110 4042 -5050
rect 4040 -5116 4102 -5110
rect 3600 -5214 3606 -5154
rect 3666 -5214 3672 -5154
rect 3002 -5375 3410 -5369
rect 3002 -5409 3014 -5375
rect 3398 -5409 3410 -5375
rect 3002 -5415 3410 -5409
rect 1936 -6644 1942 -5580
rect 1896 -6656 1942 -6644
rect 2748 -6644 2760 -5468
rect 2794 -6644 2808 -5468
rect 3606 -5468 3666 -5214
rect 4040 -5369 4100 -5116
rect 3860 -5375 4268 -5369
rect 3860 -5409 3872 -5375
rect 4256 -5409 4268 -5375
rect 3860 -5415 4268 -5409
rect 3606 -5520 3618 -5468
rect 1286 -6703 1694 -6697
rect 1286 -6737 1298 -6703
rect 1682 -6737 1694 -6703
rect 1286 -6743 1694 -6737
rect 2144 -6703 2552 -6697
rect 2144 -6737 2156 -6703
rect 2540 -6737 2552 -6703
rect 2144 -6743 2552 -6737
rect 1456 -6926 1516 -6743
rect 2326 -6926 2386 -6743
rect 1450 -6986 1456 -6926
rect 1516 -6986 1522 -6926
rect 2320 -6986 2326 -6926
rect 2386 -6986 2392 -6926
rect 2748 -7070 2808 -6644
rect 3612 -6644 3618 -5520
rect 3652 -5520 3666 -5468
rect 4462 -5468 4522 -4904
rect 5328 -4904 5334 -3886
rect 5368 -3886 5380 -3728
rect 6186 -3728 6232 -3716
rect 6186 -3788 6192 -3728
rect 5368 -4904 5374 -3886
rect 5328 -4916 5374 -4904
rect 6180 -4904 6192 -3788
rect 6226 -3788 6232 -3728
rect 7036 -3728 7098 -3592
rect 7480 -3629 7540 -3263
rect 7894 -3530 7954 -3164
rect 8760 -3164 8766 -2138
rect 8800 -2138 8812 -1988
rect 9608 -1988 9668 -1424
rect 10476 -1424 10482 -304
rect 10516 -304 10530 -248
rect 11326 -248 11386 6
rect 11750 -149 11810 6
rect 11582 -155 11990 -149
rect 11582 -189 11594 -155
rect 11978 -189 11990 -155
rect 11582 -195 11990 -189
rect 11750 -196 11810 -195
rect 10516 -1424 10522 -304
rect 10476 -1436 10522 -1424
rect 11326 -1424 11340 -248
rect 11374 -1424 11386 -248
rect 9866 -1483 10274 -1477
rect 9866 -1517 9878 -1483
rect 10262 -1517 10274 -1483
rect 9866 -1523 10274 -1517
rect 10724 -1483 11132 -1477
rect 10724 -1517 10736 -1483
rect 11120 -1517 11132 -1483
rect 10724 -1523 11132 -1517
rect 10048 -1678 10108 -1523
rect 10462 -1640 10468 -1580
rect 10528 -1640 10534 -1580
rect 10046 -1684 10108 -1678
rect 10106 -1744 10108 -1684
rect 10046 -1750 10108 -1744
rect 10048 -1889 10108 -1750
rect 9866 -1895 10274 -1889
rect 9866 -1929 9878 -1895
rect 10262 -1929 10274 -1895
rect 9866 -1935 10274 -1929
rect 8800 -3164 8806 -2138
rect 8760 -3176 8806 -3164
rect 9608 -3164 9624 -1988
rect 9658 -3164 9668 -1988
rect 10468 -1988 10528 -1640
rect 10904 -1684 10964 -1523
rect 11326 -1680 11386 -1424
rect 12184 -248 12244 6
rect 12184 -1424 12198 -248
rect 12232 -1424 12244 -248
rect 11582 -1483 11990 -1477
rect 11582 -1517 11594 -1483
rect 11978 -1517 11990 -1483
rect 11582 -1523 11990 -1517
rect 11754 -1680 11814 -1523
rect 12184 -1680 12244 -1424
rect 12516 -1680 12522 6
rect 10898 -1744 10904 -1684
rect 10964 -1744 10970 -1684
rect 11326 -1740 12522 -1680
rect 10904 -1889 10964 -1744
rect 10724 -1895 11132 -1889
rect 10724 -1929 10736 -1895
rect 11120 -1929 11132 -1895
rect 10724 -1935 11132 -1929
rect 10468 -2124 10482 -1988
rect 8150 -3223 8558 -3217
rect 8150 -3257 8162 -3223
rect 8546 -3257 8558 -3223
rect 8150 -3263 8558 -3257
rect 9008 -3223 9416 -3217
rect 9008 -3257 9020 -3223
rect 9404 -3257 9416 -3223
rect 9008 -3263 9416 -3257
rect 7292 -3635 7700 -3629
rect 7292 -3669 7304 -3635
rect 7688 -3669 7700 -3635
rect 7292 -3675 7700 -3669
rect 7036 -3760 7050 -3728
rect 7038 -3774 7050 -3760
rect 6226 -4904 6240 -3788
rect 4718 -4963 5126 -4957
rect 4718 -4997 4730 -4963
rect 5114 -4997 5126 -4963
rect 4718 -5003 5126 -4997
rect 5576 -4963 5984 -4957
rect 5576 -4997 5588 -4963
rect 5972 -4997 5984 -4963
rect 5576 -5003 5984 -4997
rect 4900 -5044 4960 -5003
rect 4898 -5050 4960 -5044
rect 4958 -5110 4960 -5050
rect 4898 -5116 4960 -5110
rect 4900 -5369 4960 -5116
rect 5742 -5044 5802 -5003
rect 5742 -5050 5806 -5044
rect 5742 -5110 5746 -5050
rect 5742 -5116 5806 -5110
rect 5742 -5369 5802 -5116
rect 4718 -5375 5126 -5369
rect 4718 -5409 4730 -5375
rect 5114 -5409 5126 -5375
rect 4718 -5415 5126 -5409
rect 5576 -5375 5984 -5369
rect 5576 -5409 5588 -5375
rect 5972 -5409 5984 -5375
rect 5576 -5415 5984 -5409
rect 5742 -5418 5802 -5415
rect 3652 -6644 3658 -5520
rect 3612 -6656 3658 -6644
rect 4462 -6644 4476 -5468
rect 4510 -6644 4522 -5468
rect 5328 -5468 5374 -5456
rect 5328 -6540 5334 -5468
rect 3002 -6703 3410 -6697
rect 3002 -6737 3014 -6703
rect 3398 -6737 3410 -6703
rect 3002 -6743 3410 -6737
rect 3860 -6703 4268 -6697
rect 3860 -6737 3872 -6703
rect 4256 -6737 4268 -6703
rect 3860 -6743 4268 -6737
rect 3184 -6926 3244 -6743
rect 4042 -6926 4102 -6743
rect 3178 -6986 3184 -6926
rect 3244 -6986 3250 -6926
rect 4036 -6986 4042 -6926
rect 4102 -6986 4108 -6926
rect 4462 -7070 4522 -6644
rect 5320 -6644 5334 -6540
rect 5368 -6540 5374 -5468
rect 6180 -5468 6240 -4904
rect 7044 -4904 7050 -3774
rect 7084 -3774 7098 -3728
rect 7894 -3728 7954 -3590
rect 8336 -3629 8396 -3263
rect 8750 -3486 8756 -3426
rect 8816 -3486 8822 -3426
rect 8150 -3635 8558 -3629
rect 8150 -3669 8162 -3635
rect 8546 -3669 8558 -3635
rect 8150 -3675 8558 -3669
rect 7084 -4904 7090 -3774
rect 7044 -4916 7090 -4904
rect 7894 -4904 7908 -3728
rect 7942 -4904 7954 -3728
rect 8756 -3728 8816 -3486
rect 9192 -3629 9252 -3263
rect 9008 -3635 9416 -3629
rect 9008 -3669 9020 -3635
rect 9404 -3669 9416 -3635
rect 9008 -3675 9416 -3669
rect 8756 -3820 8766 -3728
rect 6434 -4963 6842 -4957
rect 6434 -4997 6446 -4963
rect 6830 -4997 6842 -4963
rect 6434 -5003 6842 -4997
rect 7292 -4963 7700 -4957
rect 7292 -4997 7304 -4963
rect 7688 -4997 7700 -4963
rect 7292 -5003 7700 -4997
rect 6602 -5044 6662 -5003
rect 6600 -5050 6662 -5044
rect 6660 -5110 6662 -5050
rect 6600 -5116 6662 -5110
rect 6602 -5369 6662 -5116
rect 7480 -5050 7540 -5003
rect 7480 -5369 7540 -5110
rect 6434 -5375 6842 -5369
rect 6434 -5409 6446 -5375
rect 6830 -5409 6842 -5375
rect 6434 -5415 6842 -5409
rect 7292 -5375 7700 -5369
rect 7292 -5409 7304 -5375
rect 7688 -5409 7700 -5375
rect 7292 -5415 7700 -5409
rect 5368 -6644 5380 -6540
rect 4718 -6703 5126 -6697
rect 4718 -6737 4730 -6703
rect 5114 -6737 5126 -6703
rect 4718 -6743 5126 -6737
rect 4900 -6926 4960 -6743
rect 5320 -6800 5380 -6644
rect 6180 -6644 6192 -5468
rect 6226 -6644 6240 -5468
rect 7044 -5468 7090 -5456
rect 7044 -6602 7050 -5468
rect 5576 -6703 5984 -6697
rect 5576 -6737 5588 -6703
rect 5972 -6737 5984 -6703
rect 5576 -6743 5984 -6737
rect 5314 -6860 5320 -6800
rect 5380 -6860 5386 -6800
rect 5758 -6926 5818 -6743
rect 4894 -6986 4900 -6926
rect 4960 -6986 4966 -6926
rect 5752 -6986 5758 -6926
rect 5818 -6986 5824 -6926
rect 6180 -7070 6240 -6644
rect 7038 -6644 7050 -6602
rect 7084 -6602 7090 -5468
rect 7894 -5468 7954 -4904
rect 8760 -4904 8766 -3820
rect 8800 -3820 8816 -3728
rect 9608 -3728 9668 -3164
rect 10476 -3164 10482 -2124
rect 10516 -2124 10528 -1988
rect 11326 -1988 11386 -1740
rect 11754 -1889 11814 -1740
rect 11582 -1895 11990 -1889
rect 11582 -1929 11594 -1895
rect 11978 -1929 11990 -1895
rect 11582 -1935 11990 -1929
rect 10516 -3164 10522 -2124
rect 10476 -3176 10522 -3164
rect 11326 -3164 11340 -1988
rect 11374 -3164 11386 -1988
rect 9866 -3223 10274 -3217
rect 9866 -3257 9878 -3223
rect 10262 -3257 10274 -3223
rect 9866 -3263 10274 -3257
rect 10724 -3223 11132 -3217
rect 10724 -3257 10736 -3223
rect 11120 -3257 11132 -3223
rect 10724 -3263 11132 -3257
rect 10048 -3629 10108 -3263
rect 10464 -3384 10470 -3324
rect 10530 -3384 10536 -3324
rect 9866 -3635 10274 -3629
rect 9866 -3669 9878 -3635
rect 10262 -3669 10274 -3635
rect 9866 -3675 10274 -3669
rect 8800 -4904 8806 -3820
rect 8760 -4916 8806 -4904
rect 9608 -4904 9624 -3728
rect 9658 -4904 9668 -3728
rect 10470 -3728 10530 -3384
rect 10904 -3629 10964 -3263
rect 11326 -3412 11386 -3164
rect 12184 -1988 12244 -1740
rect 12184 -3164 12198 -1988
rect 12232 -3164 12244 -1988
rect 11582 -3223 11990 -3217
rect 11582 -3257 11594 -3223
rect 11978 -3257 11990 -3223
rect 11582 -3263 11990 -3257
rect 11750 -3412 11810 -3263
rect 12184 -3412 12244 -3164
rect 12516 -3412 12522 -1740
rect 11326 -3472 12522 -3412
rect 10724 -3635 11132 -3629
rect 10724 -3669 10736 -3635
rect 11120 -3669 11132 -3635
rect 10724 -3675 11132 -3669
rect 10470 -3784 10482 -3728
rect 8150 -4963 8558 -4957
rect 8150 -4997 8162 -4963
rect 8546 -4997 8558 -4963
rect 8150 -5003 8558 -4997
rect 9008 -4963 9416 -4957
rect 9008 -4997 9020 -4963
rect 9404 -4997 9416 -4963
rect 9008 -5003 9416 -4997
rect 8336 -5044 8396 -5003
rect 8334 -5050 8396 -5044
rect 8394 -5110 8396 -5050
rect 8334 -5116 8396 -5110
rect 8336 -5369 8396 -5116
rect 9192 -5054 9252 -5003
rect 8746 -5214 8752 -5154
rect 8812 -5214 8818 -5154
rect 8150 -5375 8558 -5369
rect 8150 -5409 8162 -5375
rect 8546 -5409 8558 -5375
rect 8150 -5415 8558 -5409
rect 7084 -6644 7098 -6602
rect 6434 -6703 6842 -6697
rect 6434 -6737 6446 -6703
rect 6830 -6737 6842 -6703
rect 6434 -6743 6842 -6737
rect 6616 -6926 6676 -6743
rect 7038 -6800 7098 -6644
rect 7894 -6644 7908 -5468
rect 7942 -6644 7954 -5468
rect 8752 -5468 8812 -5214
rect 9192 -5369 9252 -5114
rect 9008 -5375 9416 -5369
rect 9008 -5409 9020 -5375
rect 9404 -5409 9416 -5375
rect 9008 -5415 9416 -5409
rect 8752 -5518 8766 -5468
rect 7292 -6703 7700 -6697
rect 7292 -6737 7304 -6703
rect 7688 -6737 7700 -6703
rect 7292 -6743 7700 -6737
rect 7032 -6860 7038 -6800
rect 7098 -6860 7104 -6800
rect 7474 -6926 7534 -6743
rect 6610 -6986 6616 -6926
rect 6676 -6986 6682 -6926
rect 7468 -6986 7474 -6926
rect 7534 -6986 7540 -6926
rect 7894 -7070 7954 -6644
rect 8760 -6644 8766 -5518
rect 8800 -5518 8812 -5468
rect 9608 -5468 9668 -4904
rect 10476 -4904 10482 -3784
rect 10516 -3784 10530 -3728
rect 11326 -3728 11386 -3472
rect 11750 -3629 11810 -3472
rect 11582 -3635 11990 -3629
rect 11582 -3669 11594 -3635
rect 11978 -3669 11990 -3635
rect 11582 -3675 11990 -3669
rect 10516 -4904 10522 -3784
rect 10476 -4916 10522 -4904
rect 11326 -4904 11340 -3728
rect 11374 -4904 11386 -3728
rect 9866 -4963 10274 -4957
rect 9866 -4997 9878 -4963
rect 10262 -4997 10274 -4963
rect 9866 -5003 10274 -4997
rect 10724 -4963 11132 -4957
rect 10724 -4997 10736 -4963
rect 11120 -4997 11132 -4963
rect 10724 -5003 11132 -4997
rect 10048 -5050 10108 -5003
rect 10048 -5369 10108 -5110
rect 10904 -5044 10964 -5003
rect 10904 -5050 10966 -5044
rect 10904 -5110 10906 -5050
rect 10904 -5116 10966 -5110
rect 10464 -5328 10470 -5268
rect 10530 -5328 10536 -5268
rect 9866 -5375 10274 -5369
rect 9866 -5409 9878 -5375
rect 10262 -5409 10274 -5375
rect 9866 -5415 10274 -5409
rect 8800 -6644 8806 -5518
rect 8760 -6656 8806 -6644
rect 9608 -6644 9624 -5468
rect 9658 -6644 9668 -5468
rect 10470 -5468 10530 -5328
rect 10904 -5369 10964 -5116
rect 11326 -5154 11386 -4904
rect 12184 -3728 12244 -3472
rect 12184 -4904 12198 -3728
rect 12232 -4904 12244 -3728
rect 11582 -4963 11990 -4957
rect 11582 -4997 11594 -4963
rect 11978 -4997 11990 -4963
rect 11582 -5003 11990 -4997
rect 11754 -5154 11814 -5003
rect 12184 -5154 12244 -4904
rect 12516 -5154 12522 -3472
rect 11326 -5214 12522 -5154
rect 10724 -5375 11132 -5369
rect 10724 -5409 10736 -5375
rect 11120 -5409 11132 -5375
rect 10724 -5415 11132 -5409
rect 10470 -5518 10482 -5468
rect 8150 -6703 8558 -6697
rect 8150 -6737 8162 -6703
rect 8546 -6737 8558 -6703
rect 8150 -6743 8558 -6737
rect 9008 -6703 9416 -6697
rect 9008 -6737 9020 -6703
rect 9404 -6737 9416 -6703
rect 9008 -6743 9416 -6737
rect 8332 -6926 8392 -6743
rect 9190 -6926 9250 -6743
rect 8326 -6986 8332 -6926
rect 8392 -6986 8398 -6926
rect 9184 -6986 9190 -6926
rect 9250 -6986 9256 -6926
rect 9608 -7070 9668 -6644
rect 10476 -6644 10482 -5518
rect 10516 -5518 10530 -5468
rect 11326 -5468 11386 -5214
rect 11754 -5369 11814 -5214
rect 11582 -5375 11990 -5369
rect 11582 -5409 11594 -5375
rect 11978 -5409 11990 -5375
rect 11582 -5415 11990 -5409
rect 10516 -6644 10522 -5518
rect 11326 -5572 11340 -5468
rect 11334 -6594 11340 -5572
rect 10476 -6656 10522 -6644
rect 11324 -6644 11340 -6594
rect 11374 -5572 11386 -5468
rect 12184 -5468 12244 -5214
rect 12184 -5568 12198 -5468
rect 11374 -6594 11380 -5572
rect 12192 -6588 12198 -5568
rect 11374 -6644 11384 -6594
rect 9866 -6703 10274 -6697
rect 9866 -6737 9878 -6703
rect 10262 -6737 10274 -6703
rect 9866 -6743 10274 -6737
rect 10724 -6703 11132 -6697
rect 10724 -6737 10736 -6703
rect 11120 -6737 11132 -6703
rect 10724 -6743 11132 -6737
rect 10048 -6926 10108 -6743
rect 10904 -6926 10964 -6743
rect 10042 -6986 10048 -6926
rect 10108 -6986 10114 -6926
rect 10898 -6986 10904 -6926
rect 10964 -6986 10970 -6926
rect 11324 -7070 11384 -6644
rect 12184 -6644 12198 -6588
rect 12232 -5568 12244 -5468
rect 12232 -6588 12238 -5568
rect 12232 -6644 12244 -6588
rect 11582 -6703 11990 -6697
rect 11582 -6737 11594 -6703
rect 11978 -6737 11990 -6703
rect 11582 -6743 11990 -6737
rect 11750 -7070 11810 -6743
rect 12184 -7070 12244 -6644
rect 164 -7076 170 -7070
rect -262 -7119 170 -7076
rect -368 -7130 170 -7119
rect 230 -7130 236 -7070
rect 584 -7130 590 -7070
rect 650 -7130 656 -7070
rect 1024 -7130 1030 -7070
rect 1090 -7130 1096 -7070
rect 2742 -7130 2748 -7070
rect 2808 -7130 2814 -7070
rect 4456 -7130 4462 -7070
rect 4522 -7130 4528 -7070
rect 6174 -7130 6180 -7070
rect 6240 -7130 6246 -7070
rect 7888 -7130 7894 -7070
rect 7954 -7130 7960 -7070
rect 9602 -7130 9608 -7070
rect 9668 -7130 9674 -7070
rect 11318 -7130 11324 -7070
rect 11384 -7130 11390 -7070
rect 11744 -7130 11750 -7070
rect 11810 -7130 11816 -7070
rect 12178 -7130 12184 -7070
rect 12244 -7072 12250 -7070
rect 12516 -7072 12522 -5214
rect 12244 -7119 12522 -7072
rect 12622 -7119 12628 2299
rect 12244 -7130 12628 -7119
rect -368 -7136 230 -7130
rect -368 -7436 -256 -7136
rect 170 -7436 230 -7136
rect 590 -7436 650 -7130
rect 1030 -7436 1090 -7130
rect 2748 -7436 2808 -7130
rect 4462 -7436 4522 -7130
rect 6180 -7436 6240 -7130
rect 7894 -7436 7954 -7130
rect 9608 -7436 9668 -7130
rect 11324 -7436 11384 -7130
rect 11750 -7436 11810 -7130
rect 12184 -7132 12628 -7130
rect 12184 -7436 12244 -7132
rect 12516 -7436 12628 -7132
rect -368 -7442 12628 -7436
rect -368 -7542 -262 -7442
rect 12522 -7542 12628 -7442
rect -368 -7548 12628 -7542
rect -368 -7778 12628 -7772
rect -368 -7878 -262 -7778
rect 12522 -7878 12628 -7778
rect -368 -7884 12628 -7878
rect -368 -7982 -256 -7884
rect -368 -10570 -362 -7982
rect -262 -10570 -256 -7982
rect 4792 -8222 4798 -8162
rect 4858 -8222 4864 -8162
rect 4798 -9092 4858 -8222
rect 4896 -8272 4956 -7884
rect 5124 -8272 5184 -7884
rect 4896 -8332 5184 -8272
rect 5576 -8330 5582 -8270
rect 5642 -8330 5648 -8270
rect 4896 -8472 4956 -8332
rect 5124 -8382 5184 -8332
rect 5582 -8382 5642 -8330
rect 5052 -8388 5260 -8382
rect 5052 -8422 5064 -8388
rect 5248 -8422 5260 -8388
rect 5052 -8428 5260 -8422
rect 5510 -8388 5718 -8382
rect 5510 -8422 5522 -8388
rect 5706 -8422 5718 -8388
rect 5510 -8428 5718 -8422
rect 4896 -8848 4910 -8472
rect 4944 -8848 4956 -8472
rect 5362 -8472 5408 -8460
rect 5362 -8826 5368 -8472
rect 4896 -9032 4956 -8848
rect 5356 -8848 5368 -8826
rect 5402 -8826 5408 -8472
rect 5814 -8472 5874 -7884
rect 6264 -8222 6270 -8162
rect 6330 -8222 6336 -8162
rect 6036 -8330 6042 -8270
rect 6102 -8330 6108 -8270
rect 6042 -8382 6102 -8330
rect 5968 -8388 6176 -8382
rect 5968 -8422 5980 -8388
rect 6164 -8422 6176 -8388
rect 5968 -8428 6176 -8422
rect 5402 -8848 5416 -8826
rect 5052 -8898 5260 -8892
rect 5052 -8932 5064 -8898
rect 5248 -8932 5260 -8898
rect 5052 -8938 5260 -8932
rect 5124 -9032 5184 -8938
rect 5356 -8978 5416 -8848
rect 5814 -8848 5826 -8472
rect 5860 -8848 5874 -8472
rect 6270 -8472 6330 -8222
rect 6498 -8330 6504 -8270
rect 6564 -8330 6570 -8270
rect 6504 -8382 6564 -8330
rect 6426 -8388 6634 -8382
rect 6426 -8422 6438 -8388
rect 6622 -8422 6634 -8388
rect 6426 -8428 6634 -8422
rect 6270 -8494 6284 -8472
rect 5510 -8898 5718 -8892
rect 5510 -8932 5522 -8898
rect 5706 -8932 5718 -8898
rect 5510 -8938 5718 -8932
rect 4896 -9092 5184 -9032
rect 5350 -9038 5356 -8978
rect 5416 -9038 5422 -8978
rect 4792 -9152 4798 -9092
rect 4858 -9152 4864 -9092
rect 4896 -9272 4956 -9092
rect 5124 -9182 5184 -9092
rect 5350 -9152 5356 -9092
rect 5416 -9152 5422 -9092
rect 5052 -9188 5260 -9182
rect 5052 -9222 5064 -9188
rect 5248 -9222 5260 -9188
rect 5052 -9228 5260 -9222
rect 4896 -9648 4910 -9272
rect 4944 -9648 4956 -9272
rect 5356 -9272 5416 -9152
rect 5584 -9182 5644 -8938
rect 5510 -9188 5718 -9182
rect 5510 -9222 5522 -9188
rect 5706 -9222 5718 -9188
rect 5510 -9228 5718 -9222
rect 5356 -9316 5368 -9272
rect 4896 -9794 4956 -9648
rect 5362 -9648 5368 -9316
rect 5402 -9316 5416 -9272
rect 5814 -9272 5874 -8848
rect 6278 -8848 6284 -8494
rect 6318 -8494 6330 -8472
rect 6728 -8472 6788 -7884
rect 7422 -8268 7482 -7884
rect 7646 -8268 7706 -7884
rect 6954 -8330 6960 -8270
rect 7020 -8330 7026 -8270
rect 7422 -8328 7706 -8268
rect 6960 -8382 7020 -8330
rect 7422 -8382 7482 -8328
rect 6884 -8388 7092 -8382
rect 6884 -8422 6896 -8388
rect 7080 -8422 7092 -8388
rect 6884 -8428 7092 -8422
rect 7342 -8388 7550 -8382
rect 7342 -8422 7354 -8388
rect 7538 -8422 7550 -8388
rect 7342 -8428 7550 -8422
rect 6318 -8848 6324 -8494
rect 6278 -8860 6324 -8848
rect 6728 -8848 6742 -8472
rect 6776 -8848 6788 -8472
rect 7194 -8472 7240 -8460
rect 7194 -8804 7200 -8472
rect 5968 -8898 6176 -8892
rect 5968 -8932 5980 -8898
rect 6164 -8932 6176 -8898
rect 5968 -8938 6176 -8932
rect 6426 -8898 6634 -8892
rect 6426 -8932 6438 -8898
rect 6622 -8932 6634 -8898
rect 6426 -8938 6634 -8932
rect 6044 -9182 6104 -8938
rect 6264 -9038 6270 -8978
rect 6330 -9038 6336 -8978
rect 5968 -9188 6176 -9182
rect 5968 -9222 5980 -9188
rect 6164 -9222 6176 -9188
rect 5968 -9228 6176 -9222
rect 5402 -9648 5408 -9316
rect 5362 -9660 5408 -9648
rect 5814 -9648 5826 -9272
rect 5860 -9648 5874 -9272
rect 6270 -9272 6330 -9038
rect 6504 -9182 6564 -8938
rect 6426 -9188 6634 -9182
rect 6426 -9222 6438 -9188
rect 6622 -9222 6634 -9188
rect 6426 -9228 6634 -9222
rect 6270 -9324 6284 -9272
rect 5584 -9692 5644 -9690
rect 5052 -9698 5260 -9692
rect 5052 -9732 5064 -9698
rect 5248 -9732 5260 -9698
rect 5052 -9738 5260 -9732
rect 5510 -9698 5718 -9692
rect 5510 -9732 5522 -9698
rect 5706 -9732 5718 -9698
rect 5510 -9738 5718 -9732
rect 5124 -9794 5184 -9738
rect 5584 -9792 5644 -9738
rect 4896 -9854 5184 -9794
rect 5578 -9852 5584 -9792
rect 5644 -9852 5650 -9792
rect 4896 -10100 4956 -9854
rect 5124 -10100 5184 -9854
rect 5814 -9918 5874 -9648
rect 6278 -9648 6284 -9324
rect 6318 -9324 6330 -9272
rect 6728 -9272 6788 -8848
rect 7186 -8848 7200 -8804
rect 7234 -8804 7240 -8472
rect 7646 -8472 7706 -8328
rect 7234 -8848 7246 -8804
rect 6884 -8898 7092 -8892
rect 6884 -8932 6896 -8898
rect 7080 -8932 7092 -8898
rect 6884 -8938 7092 -8932
rect 6964 -9182 7024 -8938
rect 7186 -8978 7246 -8848
rect 7646 -8848 7658 -8472
rect 7692 -8848 7706 -8472
rect 7342 -8898 7550 -8892
rect 7342 -8932 7354 -8898
rect 7538 -8932 7550 -8898
rect 7342 -8938 7550 -8932
rect 7180 -9038 7186 -8978
rect 7246 -9038 7252 -8978
rect 7424 -9034 7484 -8938
rect 7646 -9034 7706 -8848
rect 7180 -9152 7186 -9092
rect 7246 -9152 7252 -9092
rect 7424 -9094 7706 -9034
rect 6884 -9188 7092 -9182
rect 6884 -9222 6896 -9188
rect 7080 -9222 7092 -9188
rect 6884 -9228 7092 -9222
rect 6318 -9648 6324 -9324
rect 6278 -9660 6324 -9648
rect 6728 -9648 6742 -9272
rect 6776 -9648 6788 -9272
rect 7186 -9272 7246 -9152
rect 7424 -9182 7484 -9094
rect 7342 -9188 7550 -9182
rect 7342 -9222 7354 -9188
rect 7538 -9222 7550 -9188
rect 7342 -9228 7550 -9222
rect 7186 -9314 7200 -9272
rect 5968 -9698 6176 -9692
rect 5968 -9732 5980 -9698
rect 6164 -9732 6176 -9698
rect 5968 -9738 6176 -9732
rect 6426 -9698 6634 -9692
rect 6426 -9732 6438 -9698
rect 6622 -9732 6634 -9698
rect 6426 -9738 6634 -9732
rect 6044 -9792 6104 -9738
rect 6504 -9792 6564 -9738
rect 6038 -9852 6044 -9792
rect 6104 -9852 6110 -9792
rect 6498 -9852 6504 -9792
rect 6564 -9852 6570 -9792
rect 6728 -9918 6788 -9648
rect 7194 -9648 7200 -9314
rect 7234 -9314 7246 -9272
rect 7646 -9272 7706 -9094
rect 7234 -9648 7240 -9314
rect 7194 -9660 7240 -9648
rect 7646 -9648 7658 -9272
rect 7692 -9648 7706 -9272
rect 6884 -9698 7092 -9692
rect 6884 -9732 6896 -9698
rect 7080 -9732 7092 -9698
rect 6884 -9738 7092 -9732
rect 7342 -9698 7550 -9692
rect 7342 -9732 7354 -9698
rect 7538 -9732 7550 -9698
rect 7342 -9738 7550 -9732
rect 6958 -9792 7018 -9738
rect 7422 -9790 7482 -9738
rect 7646 -9790 7706 -9648
rect 6952 -9852 6958 -9792
rect 7018 -9852 7024 -9792
rect 7422 -9850 7706 -9790
rect 5808 -9978 5814 -9918
rect 5874 -9978 5880 -9918
rect 6722 -9978 6728 -9918
rect 6788 -9978 6794 -9918
rect 5814 -10100 5874 -9978
rect 6728 -10100 6788 -9978
rect 7422 -10100 7482 -9850
rect 7646 -10100 7706 -9850
rect 12516 -7982 12628 -7884
rect 4664 -10168 7854 -10100
rect -368 -10716 -256 -10570
rect 344 -10716 354 -10416
rect 4664 -10594 4734 -10168
rect 7798 -10594 7854 -10168
rect 4664 -10646 7854 -10594
rect 11906 -10716 11916 -10416
rect 12516 -10570 12522 -7982
rect 12622 -10570 12628 -7982
rect 12516 -10716 12628 -10570
rect -368 -10722 12628 -10716
rect -368 -10822 -262 -10722
rect 12522 -10822 12628 -10722
rect -368 -10828 12628 -10822
<< via1 >>
rect -256 2516 344 2816
rect 11916 2516 12516 2816
rect 158 2232 12268 2396
rect 172 2050 232 2110
rect 596 2050 656 2110
rect 1032 2050 1092 2110
rect 2746 2050 2806 2110
rect 4466 2050 4526 2110
rect 6174 2050 6234 2110
rect 7894 2050 7954 2110
rect 9608 2050 9668 2110
rect 11326 2050 11386 2110
rect 11754 2050 11814 2110
rect 12186 2050 12246 2110
rect -92 1786 -32 1846
rect 50 1658 110 1718
rect 1458 1922 1518 1982
rect 2312 1922 2372 1982
rect 3172 1922 3232 1982
rect 4032 1922 4092 1982
rect 50 -4 110 56
rect -92 -110 -32 -50
rect -92 -1640 -32 -1580
rect 1888 96 1948 156
rect 1890 -110 1950 -50
rect 4892 1922 4952 1982
rect 5752 1922 5812 1982
rect 3470 -4 3530 56
rect 3604 -6 3664 54
rect 50 -1846 110 -1786
rect 1458 -1744 1518 -1684
rect 2320 -1744 2380 -1684
rect 6612 1922 6672 1982
rect 7472 1922 7532 1982
rect 8332 1922 8392 1982
rect 9172 1922 9232 1982
rect 8752 1658 8812 1718
rect 5320 -110 5380 -50
rect 7166 -110 7226 -50
rect 3182 -1744 3242 -1684
rect 4040 -1744 4100 -1684
rect 50 -3484 110 -3424
rect -92 -3590 -32 -3530
rect 1888 -3384 1948 -3324
rect 1890 -3590 1950 -3530
rect 4900 -1744 4960 -1684
rect 5744 -1744 5804 -1684
rect 3470 -3484 3530 -3424
rect 3604 -3486 3664 -3426
rect 10030 1922 10090 1982
rect 10892 1922 10952 1982
rect 10468 1786 10528 1846
rect 8756 -6 8816 54
rect 6614 -1744 6674 -1684
rect 7480 -1744 7540 -1684
rect 4462 -3592 4522 -3532
rect 1460 -5110 1520 -5050
rect 2320 -5110 2380 -5050
rect 1888 -5328 1948 -5268
rect 6180 -3256 6240 -3196
rect 10470 96 10530 156
rect 8336 -1744 8396 -1684
rect 9192 -1744 9252 -1684
rect 8752 -1846 8812 -1786
rect 5320 -3590 5380 -3530
rect 7166 -3590 7226 -3530
rect 3176 -5110 3236 -5050
rect 4042 -5110 4102 -5050
rect 3606 -5214 3666 -5154
rect 1456 -6986 1516 -6926
rect 2326 -6986 2386 -6926
rect 10468 -1640 10528 -1580
rect 10046 -1744 10106 -1684
rect 10904 -1744 10964 -1684
rect 7894 -3590 7954 -3530
rect 4898 -5110 4958 -5050
rect 5746 -5110 5806 -5050
rect 3184 -6986 3244 -6926
rect 4042 -6986 4102 -6926
rect 8756 -3486 8816 -3426
rect 6600 -5110 6660 -5050
rect 7480 -5110 7540 -5050
rect 5320 -6860 5380 -6800
rect 4900 -6986 4960 -6926
rect 5758 -6986 5818 -6926
rect 10470 -3384 10530 -3324
rect 8334 -5110 8394 -5050
rect 9192 -5114 9252 -5054
rect 8752 -5214 8812 -5154
rect 7038 -6860 7098 -6800
rect 6616 -6986 6676 -6926
rect 7474 -6986 7534 -6926
rect 10048 -5110 10108 -5050
rect 10906 -5110 10966 -5050
rect 10470 -5328 10530 -5268
rect 8332 -6986 8392 -6926
rect 9190 -6986 9250 -6926
rect 10048 -6986 10108 -6926
rect 10904 -6986 10964 -6926
rect 170 -7130 230 -7070
rect 590 -7130 650 -7070
rect 1030 -7130 1090 -7070
rect 2748 -7130 2808 -7070
rect 4462 -7130 4522 -7070
rect 6180 -7130 6240 -7070
rect 7894 -7130 7954 -7070
rect 9608 -7130 9668 -7070
rect 11324 -7130 11384 -7070
rect 11750 -7130 11810 -7070
rect 12184 -7130 12244 -7070
rect 4798 -8222 4858 -8162
rect 5582 -8330 5642 -8270
rect 6270 -8222 6330 -8162
rect 6042 -8330 6102 -8270
rect 6504 -8330 6564 -8270
rect 5356 -9038 5416 -8978
rect 4798 -9152 4858 -9092
rect 5356 -9152 5416 -9092
rect 6960 -8330 7020 -8270
rect 6270 -9038 6330 -8978
rect 5584 -9852 5644 -9792
rect 7186 -9038 7246 -8978
rect 7186 -9152 7246 -9092
rect 6044 -9852 6104 -9792
rect 6504 -9852 6564 -9792
rect 6958 -9852 7018 -9792
rect 5814 -9978 5874 -9918
rect 6728 -9978 6788 -9918
rect -256 -10716 344 -10416
rect 4734 -10594 7798 -10168
rect 11916 -10716 12516 -10416
<< metal2 >>
rect -256 2816 344 2826
rect -256 2506 344 2516
rect 11916 2816 12516 2826
rect 11916 2506 12516 2516
rect 110 2396 12310 2438
rect 110 2232 158 2396
rect 12268 2232 12310 2396
rect 110 2192 12310 2232
rect 172 2110 232 2116
rect 596 2110 656 2116
rect 1032 2110 1092 2116
rect 2746 2110 2806 2116
rect 4466 2110 4526 2116
rect 6174 2110 6234 2116
rect 7894 2110 7954 2116
rect 9608 2110 9668 2116
rect 11326 2110 11386 2116
rect 11754 2110 11814 2116
rect 12186 2110 12246 2116
rect 232 2050 596 2110
rect 656 2050 1032 2110
rect 1092 2050 2746 2110
rect 2806 2050 4466 2110
rect 4526 2050 6174 2110
rect 6234 2050 7894 2110
rect 7954 2050 9608 2110
rect 9668 2050 11326 2110
rect 11386 2050 11754 2110
rect 11814 2050 12186 2110
rect 172 2044 232 2050
rect 596 2044 656 2050
rect 1032 2044 1092 2050
rect 2746 2044 2806 2050
rect 4466 2044 4526 2050
rect 6174 2044 6234 2050
rect 7894 2044 7954 2050
rect 9608 2044 9668 2050
rect 11326 2044 11386 2050
rect 11754 2044 11814 2050
rect 12186 2044 12246 2050
rect 1458 1982 1518 1988
rect 2312 1982 2372 1988
rect 3172 1982 3232 1988
rect 4032 1982 4092 1988
rect 4892 1982 4952 1988
rect 5752 1982 5812 1988
rect 6612 1982 6672 1988
rect 7472 1982 7532 1988
rect 8332 1982 8392 1988
rect 9172 1982 9232 1988
rect 10030 1982 10090 1988
rect 10892 1982 10952 1988
rect 1518 1922 2312 1982
rect 2372 1922 3172 1982
rect 3232 1922 4032 1982
rect 4092 1922 4892 1982
rect 4952 1922 5752 1982
rect 5812 1922 6612 1982
rect 6672 1922 7472 1982
rect 7532 1922 8332 1982
rect 8392 1922 9172 1982
rect 9232 1922 10030 1982
rect 10090 1922 10892 1982
rect 1458 1916 1518 1922
rect 2312 1916 2372 1922
rect 3172 1916 3232 1922
rect 4032 1916 4092 1922
rect 4892 1916 4952 1922
rect 5752 1916 5812 1922
rect 6612 1916 6672 1922
rect 7472 1916 7532 1922
rect 8332 1916 8392 1922
rect 9172 1916 9232 1922
rect 10030 1916 10090 1922
rect 10892 1916 10952 1922
rect -92 1846 -32 1852
rect 10468 1846 10528 1852
rect -32 1786 10468 1846
rect -92 1780 -32 1786
rect 10468 1780 10528 1786
rect 50 1718 110 1724
rect 8752 1718 8812 1724
rect 110 1658 8752 1718
rect 50 1652 110 1658
rect 8752 1652 8812 1658
rect 1888 156 1948 162
rect 10470 156 10530 162
rect 1948 96 10470 156
rect 1888 90 1948 96
rect 10470 90 10530 96
rect 50 56 110 62
rect 3470 56 3530 62
rect 110 -4 3470 56
rect 50 -10 110 -4
rect 3470 -10 3530 -4
rect 3604 54 3664 60
rect 8756 54 8816 60
rect 3664 -6 8756 54
rect 3604 -12 3664 -6
rect 8756 -12 8816 -6
rect -92 -50 -32 -44
rect 1890 -50 1950 -44
rect -32 -110 1890 -50
rect -92 -116 -32 -110
rect 1890 -116 1950 -110
rect 5320 -50 5380 -44
rect 7166 -50 7226 -44
rect 5380 -110 7166 -50
rect 5320 -116 5380 -110
rect 7166 -116 7226 -110
rect -92 -1580 -32 -1574
rect 10468 -1580 10528 -1574
rect -32 -1640 10468 -1580
rect -92 -1646 -32 -1640
rect 10468 -1646 10528 -1640
rect 10904 -1684 10964 -1678
rect 1452 -1744 1458 -1684
rect 1518 -1744 2320 -1684
rect 2380 -1744 3182 -1684
rect 3242 -1744 4040 -1684
rect 4100 -1744 4900 -1684
rect 4960 -1744 5744 -1684
rect 5804 -1744 6614 -1684
rect 6674 -1744 7480 -1684
rect 7540 -1744 8336 -1684
rect 8396 -1744 9192 -1684
rect 9252 -1744 10046 -1684
rect 10106 -1744 10904 -1684
rect 10904 -1750 10964 -1744
rect 50 -1786 110 -1780
rect 8752 -1786 8812 -1780
rect 110 -1846 8752 -1786
rect 50 -1852 110 -1846
rect 8752 -1852 8812 -1846
rect 6180 -3196 6240 -3187
rect 6174 -3256 6180 -3196
rect 6240 -3256 6246 -3196
rect 6180 -3265 6240 -3256
rect 1888 -3324 1948 -3318
rect 10470 -3324 10530 -3318
rect 1948 -3384 10470 -3324
rect 1888 -3390 1948 -3384
rect 10470 -3390 10530 -3384
rect 50 -3424 110 -3418
rect 3470 -3424 3530 -3418
rect 110 -3484 3470 -3424
rect 50 -3490 110 -3484
rect 3470 -3490 3530 -3484
rect 3604 -3426 3664 -3420
rect 8756 -3426 8816 -3420
rect 3664 -3486 8756 -3426
rect 3604 -3492 3664 -3486
rect 8756 -3492 8816 -3486
rect -92 -3530 -32 -3524
rect 1890 -3530 1950 -3524
rect -32 -3590 1890 -3530
rect 4462 -3532 4522 -3523
rect 5320 -3530 5380 -3524
rect 7166 -3530 7226 -3524
rect 7894 -3530 7954 -3521
rect -92 -3596 -32 -3590
rect 1890 -3596 1950 -3590
rect 4456 -3592 4462 -3532
rect 4522 -3592 4528 -3532
rect 5380 -3590 7166 -3530
rect 7888 -3590 7894 -3530
rect 7954 -3590 7960 -3530
rect 4462 -3601 4522 -3592
rect 5320 -3596 5380 -3590
rect 7166 -3596 7226 -3590
rect 7894 -3599 7954 -3590
rect 1460 -5050 1520 -5044
rect 1520 -5110 2320 -5050
rect 2380 -5110 3176 -5050
rect 3236 -5110 4042 -5050
rect 4102 -5110 4898 -5050
rect 4958 -5110 5746 -5050
rect 5806 -5110 6600 -5050
rect 6660 -5110 7480 -5050
rect 7540 -5110 8334 -5050
rect 8394 -5054 10048 -5050
rect 8394 -5110 9192 -5054
rect 1460 -5116 1520 -5110
rect 9186 -5114 9192 -5110
rect 9252 -5110 10048 -5054
rect 10108 -5110 10906 -5050
rect 10966 -5110 10972 -5050
rect 9252 -5114 9258 -5110
rect 3606 -5154 3666 -5148
rect 8752 -5154 8812 -5148
rect 3666 -5214 8752 -5154
rect 3606 -5220 3666 -5214
rect 8752 -5220 8812 -5214
rect 1888 -5268 1948 -5262
rect 10470 -5268 10530 -5262
rect 1948 -5328 10470 -5268
rect 1888 -5334 1948 -5328
rect 10470 -5334 10530 -5328
rect 5320 -6800 5380 -6794
rect 7038 -6800 7098 -6794
rect 5380 -6860 7038 -6800
rect 5320 -6866 5380 -6860
rect 7038 -6866 7098 -6860
rect 1456 -6926 1516 -6920
rect 2326 -6926 2386 -6920
rect 3184 -6926 3244 -6920
rect 4042 -6926 4102 -6920
rect 4900 -6926 4960 -6920
rect 5758 -6926 5818 -6920
rect 6616 -6926 6676 -6920
rect 7474 -6926 7534 -6920
rect 8332 -6926 8392 -6920
rect 9190 -6926 9250 -6920
rect 10048 -6926 10108 -6920
rect 10904 -6926 10964 -6920
rect 1516 -6986 2326 -6926
rect 2386 -6986 3184 -6926
rect 3244 -6986 4042 -6926
rect 4102 -6986 4900 -6926
rect 4960 -6986 5758 -6926
rect 5818 -6986 6616 -6926
rect 6676 -6986 7474 -6926
rect 7534 -6986 8332 -6926
rect 8392 -6986 9190 -6926
rect 9250 -6986 10048 -6926
rect 10108 -6986 10904 -6926
rect 1456 -6992 1516 -6986
rect 2326 -6992 2386 -6986
rect 3184 -6992 3244 -6986
rect 4042 -6992 4102 -6986
rect 4900 -6992 4960 -6986
rect 5758 -6992 5818 -6986
rect 6616 -6992 6676 -6986
rect 7474 -6992 7534 -6986
rect 8332 -6992 8392 -6986
rect 9190 -6992 9250 -6986
rect 10048 -6992 10108 -6986
rect 10904 -6992 10964 -6986
rect 170 -7070 230 -7064
rect 590 -7070 650 -7064
rect 1030 -7070 1090 -7064
rect 2748 -7070 2808 -7064
rect 4462 -7070 4522 -7064
rect 6180 -7070 6240 -7064
rect 7894 -7070 7954 -7064
rect 9608 -7070 9668 -7064
rect 11324 -7070 11384 -7064
rect 11750 -7070 11810 -7064
rect 12184 -7070 12244 -7064
rect 230 -7130 590 -7070
rect 650 -7130 1030 -7070
rect 1090 -7130 2748 -7070
rect 2808 -7130 4462 -7070
rect 4522 -7130 6180 -7070
rect 6240 -7130 7894 -7070
rect 7954 -7130 9608 -7070
rect 9668 -7130 11324 -7070
rect 11384 -7130 11750 -7070
rect 11810 -7130 12184 -7070
rect 170 -7136 230 -7130
rect 590 -7136 650 -7130
rect 1030 -7136 1090 -7130
rect 2748 -7136 2808 -7130
rect 4462 -7136 4522 -7130
rect 6180 -7136 6240 -7130
rect 7894 -7136 7954 -7130
rect 9608 -7136 9668 -7130
rect 11324 -7136 11384 -7130
rect 11750 -7136 11810 -7130
rect 12184 -7136 12244 -7130
rect 4798 -8162 4858 -8156
rect 6270 -8162 6330 -8156
rect 4858 -8222 6270 -8162
rect 4798 -8228 4858 -8222
rect 6270 -8228 6330 -8222
rect 5582 -8270 5642 -8264
rect 6042 -8270 6102 -8264
rect 6504 -8270 6564 -8264
rect 6960 -8270 7020 -8264
rect 5642 -8330 6042 -8270
rect 6102 -8330 6504 -8270
rect 6564 -8330 6960 -8270
rect 5582 -8336 5642 -8330
rect 6042 -8336 6102 -8330
rect 6504 -8336 6564 -8330
rect 6960 -8336 7020 -8330
rect 5356 -8978 5416 -8972
rect 6270 -8978 6330 -8972
rect 7186 -8978 7246 -8972
rect 5416 -9038 6270 -8978
rect 6330 -9038 7186 -8978
rect 5356 -9044 5416 -9038
rect 6270 -9044 6330 -9038
rect 7186 -9044 7246 -9038
rect 4798 -9092 4858 -9086
rect 5356 -9092 5416 -9086
rect 7186 -9092 7246 -9086
rect 4858 -9152 5356 -9092
rect 5416 -9152 7186 -9092
rect 4798 -9158 4858 -9152
rect 5356 -9158 5416 -9152
rect 7186 -9158 7246 -9152
rect 5584 -9792 5644 -9786
rect 6044 -9792 6104 -9786
rect 6504 -9792 6564 -9786
rect 6958 -9792 7018 -9786
rect 5644 -9852 6044 -9792
rect 6104 -9852 6504 -9792
rect 6564 -9852 6958 -9792
rect 5584 -9858 5644 -9852
rect 6044 -9858 6104 -9852
rect 6504 -9858 6564 -9852
rect 6958 -9858 7018 -9852
rect 5814 -9918 5874 -9912
rect 6728 -9918 6788 -9912
rect 5874 -9978 6728 -9918
rect 5814 -9984 5874 -9978
rect 6728 -9984 6788 -9978
rect 4664 -10168 7854 -10100
rect -256 -10416 344 -10406
rect 4664 -10594 4734 -10168
rect 7798 -10594 7854 -10168
rect 4664 -10646 7854 -10594
rect 11916 -10416 12516 -10406
rect -256 -10726 344 -10716
rect 11916 -10726 12516 -10716
<< via2 >>
rect -256 2516 344 2816
rect 11916 2516 12516 2816
rect 158 2232 12268 2396
rect 6180 -3256 6240 -3196
rect 4462 -3592 4522 -3532
rect 7894 -3590 7954 -3530
rect -256 -10716 344 -10416
rect 4734 -10594 7798 -10168
rect 11916 -10716 12516 -10416
<< metal3 >>
rect -266 2816 354 2821
rect -266 2516 -256 2816
rect 344 2516 354 2816
rect -266 2511 354 2516
rect 11906 2816 12526 2821
rect 11906 2516 11916 2816
rect 12516 2516 12526 2816
rect 11906 2511 12526 2516
rect 110 2396 12310 2438
rect 110 2232 158 2396
rect 12268 2232 12310 2396
rect 110 2192 12310 2232
rect 6158 -3196 6258 -3176
rect 6158 -3256 6180 -3196
rect 6240 -3256 6258 -3196
rect 6158 -3512 6258 -3256
rect 4434 -3530 7988 -3512
rect 4434 -3532 7894 -3530
rect 4434 -3592 4462 -3532
rect 4522 -3590 7894 -3532
rect 7954 -3590 7988 -3530
rect 4522 -3592 7988 -3590
rect 4434 -3612 7988 -3592
rect 4664 -10168 7854 -10100
rect -266 -10416 354 -10411
rect -266 -10716 -256 -10416
rect 344 -10716 354 -10416
rect 4664 -10594 4734 -10168
rect 7798 -10594 7854 -10168
rect 4664 -10646 7854 -10594
rect 11906 -10416 12526 -10411
rect -266 -10721 354 -10716
rect 11906 -10716 11916 -10416
rect 12516 -10716 12526 -10416
rect 11906 -10721 12526 -10716
<< via3 >>
rect -256 2516 344 2816
rect 11916 2516 12516 2816
rect 158 2232 12268 2396
rect -256 -10716 344 -10416
rect 4734 -10594 7798 -10168
rect 11916 -10716 12516 -10416
<< metal4 >>
rect -440 2816 12700 3000
rect -440 2516 -256 2816
rect 344 2516 11916 2816
rect 12516 2516 12700 2816
rect -440 2396 12700 2516
rect -440 2232 158 2396
rect 12268 2232 12700 2396
rect -440 2200 12700 2232
rect -440 -10168 12700 -10100
rect -440 -10416 4734 -10168
rect -440 -10716 -256 -10416
rect 344 -10594 4734 -10416
rect 7798 -10416 12700 -10168
rect 7798 -10594 11916 -10416
rect 344 -10716 11916 -10594
rect 12516 -10716 12700 -10416
rect -440 -10900 12700 -10716
<< labels >>
flabel metal2 2170 120 2190 138 1 FreeSans 480 0 0 0 low_freq_pll_ibiasn
port 18 n
flabel metal2 1436 -74 1454 -64 1 FreeSans 480 0 0 0 comparator_ibiasn
port 13 n
flabel metal2 3796 12 3814 26 1 FreeSans 480 0 0 0 biquad_gm_c_filter_ibiasn4
port 17 n
flabel metal1 5340 180 5354 186 1 FreeSans 480 0 0 0 biquad_gm_c_filter_ibiasn3
port 16 n
flabel metal2 5890 -90 5904 -74 1 FreeSans 480 0 0 0 biquad_gm_c_filter_ibiasn2
port 15 n
flabel metal2 2212 16 2228 34 1 FreeSans 480 0 0 0 biquad_gm_c_filter_ibiasn1
port 14 n
flabel metal2 1210 -3580 1234 -3554 1 FreeSans 480 0 0 0 sample_and_hold_ibiasn_A
port 9 n
flabel metal2 1524 -3460 1542 -3444 1 FreeSans 480 0 0 0 peak_detector_ibiasn2
port 8 n
flabel metal2 6342 -3576 6354 -3558 1 FreeSans 480 0 0 0 peak_detector_ibiasn1
port 7 n
flabel metal1 5342 -3304 5356 -3294 1 FreeSans 480 0 0 0 diff_to_se_converter_ibiasn
port 6 n
flabel metal2 3948 -3460 3954 -3444 1 FreeSans 480 0 0 0 input_amplifier_ibiasn2
port 5 n
flabel metal2 3240 -3356 3256 -3342 1 FreeSans 480 0 0 0 input_amplifier_ibiasn1
port 4 n
flabel metal2 6058 -6832 6082 -6816 1 FreeSans 480 0 0 0 dac_8bit_ibiasn_B
port 12 n
flabel metal2 4048 -5194 4060 -5174 1 FreeSans 480 0 0 0 sample_and_hold_ibiasn_B
port 11 n
flabel metal2 2324 -5298 2344 -5282 1 FreeSans 480 0 0 0 dac_8bit_ibiasn_A
port 10 n
flabel metal2 3562 -6966 3574 -6948 1 FreeSans 480 0 0 0 vbiasp
port 3 n
flabel metal4 -414 2968 -398 2984 1 FreeSans 480 0 0 0 VDD
port 1 n power bidirectional
flabel metal2 6620 -9826 6626 -9814 1 FreeSans 480 0 0 0 vbiasn
port 19 n
flabel metal2 5934 -9020 5950 -9006 1 FreeSans 480 0 0 0 dac_8bit_ibiasp_A
port 20 n
flabel metal2 5264 -9132 5274 -9118 1 FreeSans 480 0 0 0 dac_8bit_ibiasp_B
port 21 n
flabel metal4 -398 -10890 -382 -10872 1 FreeSans 480 0 0 0 VSS
port 2 n ground bidirectional
<< end >>
