* Stimulus file.

.include ../layouts/continuous_time_comparator/comparator_pex.spice
.include comparator_lvs.spice

.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8/sky130_fd_pr__nfet_01v8__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8/sky130_fd_pr__pfet_01v8__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_05v0_nvt/sky130_fd_pr__nfet_05v0_nvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_nfet_01v8/sky130_fd_pr__esd_nfet_01v8__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_lvt/sky130_fd_pr__pfet_01v8_lvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_pfet_g5v0d10v5/sky130_fd_pr__esd_pfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d16v0/sky130_fd_pr__pfet_g5v0d16v0__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d10v5/sky130_fd_pr__nfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d16v0/sky130_fd_pr__nfet_g5v0d16v0__tt_discrete.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_nfet_g5v0d10v5/sky130_fd_pr__esd_nfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/nonfet.spice
* Mismatch parameters
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8/sky130_fd_pr__nfet_01v8__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8/sky130_fd_pr__pfet_01v8__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_lvt/sky130_fd_pr__pfet_01v8_lvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d10v5/sky130_fd_pr__nfet_g5v0d10v5__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_05v0_nvt/sky130_fd_pr__nfet_05v0_nvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__mismatch.corner.spice
* Resistor~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/Capacitor
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/r+c/res_typical__cap_typical.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/r+c/res_typical__cap_typical__lin.spice
* Special cells
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/specialized_cells.spice
* All models
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/all.spice
* Corner
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/rf.spice

.param Ibias_comp=10u vincm_comp=0.9 vsig=0 vdd=1.8 Wp_comp=4 Wn_comp=2

x0 vip vim vo ibiasn VDD VSS comparator_flat
*x1 vip vim vo ibiasn VDD VSS comparator_lvs
vdd VDD VSS 'vdd'
vss VSS 0 0
i1 VDD ibiasn 10u
*vip vip VSS pwl(0 'vincm_comp' 10n 'vincm_comp' 10.1n 'vincm_comp+5m' 50n 'vincm_comp+5m' 50.1n 'vincm_comp-5m' 110n 'vincm_comp-5m' 110.1n 'vincm_comp+5m' 200n 'vincm_comp+5m')
*vim vim VSS pwl(0 'vincm_comp' 10n 'vincm_comp' 10.1n 'vincm_comp-5m' 50n 'vincm_comp-5m' 50.1n 'vincm_comp+5m' 110n 'vincm_comp+5m' 110.1n 'vincm_comp-5m' 200n 'vincm_comp-5m')
vip vip VSS sin('vdd/2' '0.1*vdd/2' 50 0 0 0)
vim vim VSS sin('vdd/2' '0.1*vdd/2' 50 0 0 180)
*vip vip VSS dc 'vincm_comp+vsig' ac 0.5 0
*vim vim VSS dc 'vincm_comp-vsig' ac 0.5 180

.control
options savecurrents
save all
+ @m.xm1.msky130_fd_pr__nfet_01v8_lvt[id]
+ @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @m.xm2.msky130_fd_pr__nfet_01v8[gm]
+ @m.xm2.msky130_fd_pr__nfet_01v8[id]
+ @m.xm2.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm3.msky130_fd_pr__pfet_01v8[id]
+ @m.xm3.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm4.msky130_fd_pr__nfet_01v8_lvt[id]
+ @m.xm4.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @m.xm5.msky130_fd_pr__pfet_01v8[id]
+ @m.xm5.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm6.msky130_fd_pr__pfet_01v8[id]
+ @m.xm6.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm7.msky130_fd_pr__pfet_01v8[id]
+ @m.xm7.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm8.msky130_fd_pr__pfet_01v8[id]
+ @m.xm8.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm9.msky130_fd_pr__nfet_01v8[id]
+ @m.xm9.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm10.msky130_fd_pr__pfet_01v8[id]
+ @m.xm10.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm11.msky130_fd_pr__nfet_01v8[id]
+ @m.xm11.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm12.msky130_fd_pr__nfet_01v8[id]
+ @m.xm12.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm13.msky130_fd_pr__nfet_01v8[id]
+ @m.xm13.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm14.msky130_fd_pr__nfet_01v8[id]
+ @m.xm14.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm15.msky130_fd_pr__pfet_01v8_hvt[id]
+ @m.xm15.msky130_fd_pr__pfet_01v8_hvt[vth]

op
run
print all
*write comparator_lvs_op.raw

*tran 0.1n 200n
tran 10u 200m
run
write comparator_lvs_tran.raw

*dc vip 0.8999 0.9001 1e-7
*run
*write comparator_lvs_dc.raw

*ac dec 100 0.1 1g
*run
*write comparator_lvs_ac.raw
quit
.endc
