magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -1335 -1309 13042 19691
<< locali >>
rect 8998 8467 11698 8501
rect 8998 7053 11698 7087
rect 3573 6790 3792 6824
rect 3758 6308 3792 6790
rect 5908 5639 11698 5673
rect 4620 4225 11698 4259
rect 4620 2811 11698 2845
rect 3555 2541 3740 2575
rect 3555 2176 3589 2541
rect 3422 2142 3589 2176
rect 4988 1397 11698 1431
<< metal1 >>
rect 11666 8458 11730 8510
rect 2736 7801 3307 7829
rect 7502 7751 7566 7803
rect 11666 7044 11730 7096
rect 7970 6337 8034 6389
rect 2652 6160 3455 6188
rect 2820 5912 3355 5940
rect 11666 5630 11730 5682
rect 2652 5372 3322 5400
rect 2736 5248 3455 5276
rect 3072 5124 3588 5152
rect 4736 4923 4800 4975
rect 1553 4308 2652 4336
rect 11666 4216 11730 4268
rect 383 4148 2904 4176
rect 4094 3493 4158 3545
rect 3072 3332 3455 3360
rect 2904 3084 3355 3112
rect 11666 2802 11730 2854
rect 3791 2284 3855 2336
rect 2904 2145 3307 2173
rect 4462 2111 4526 2163
rect 11666 1388 11730 1440
rect 3275 643 3339 695
rect 9336 681 9400 733
rect 11666 -26 11730 26
<< metal2 >>
rect -57 17699 -29 17727
rect 1539 4322 1567 6401
rect 369 1414 397 4162
rect 137 538 203 590
rect 2554 0 2582 8524
rect 2638 0 2666 8524
rect 2722 0 2750 8524
rect 2806 0 2834 8524
rect 2890 0 2918 8524
rect 2974 0 3002 8524
rect 3058 0 3086 8524
rect 11670 8460 11726 8508
rect 7534 7763 11782 7791
rect 11670 7046 11726 7094
rect 8002 6349 11782 6377
rect 11670 5632 11726 5680
rect 4768 4935 11782 4963
rect 11670 4218 11726 4266
rect 4098 3495 4154 3543
rect 11670 2804 11726 2852
rect 3795 2286 3851 2334
rect 4480 1571 4508 2137
rect 11670 1390 11726 1438
rect 9368 707 11782 721
rect 9354 693 11782 707
rect 3293 655 3321 683
rect 9354 141 9382 693
rect 11670 -24 11726 24
<< metal3 >>
rect 607 18333 705 18431
rect 1343 18333 1441 18431
rect 607 16919 705 17017
rect 1343 16919 1441 17017
rect 607 15505 705 15603
rect 1343 15505 1441 15603
rect 607 14091 705 14189
rect 1343 14091 1441 14189
rect 607 12677 705 12775
rect 1343 12677 1441 12775
rect 607 11263 705 11361
rect 1343 11263 1441 11361
rect 607 9849 705 9947
rect 1343 9849 1441 9947
rect 607 8435 705 8533
rect 1343 8435 1441 8533
rect 11649 8435 11747 8533
rect 607 7021 705 7119
rect 1343 7021 1441 7119
rect 11649 7021 11747 7119
rect 607 5607 705 5705
rect 1343 5607 1441 5705
rect 11649 5607 11747 5705
rect 11649 4193 11747 4291
rect 2820 3489 4126 3549
rect 11649 2779 11747 2877
rect 3072 2280 3823 2340
rect 2736 1541 4494 1601
rect -49 1365 49 1463
rect 11649 1365 11747 1463
rect 1872 855 3072 915
rect 2378 473 2988 533
rect 2904 111 9368 171
rect -49 -49 49 49
rect 11649 -49 11747 49
use sky130_sram_2kbyte_1rw1r_32x512_8_dff_buf_array_0  sky130_sram_2kbyte_1rw1r_32x512_8_dff_buf_array_0_0
timestamp 1626486988
transform 1 0 0 0 1 0
box -49 -49 2590 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_16
timestamp 1626486988
transform 1 0 1839 0 1 848
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_15
timestamp 1626486988
transform 1 0 2345 0 1 466
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_pand2_1  sky130_sram_2kbyte_1rw1r_32x512_8_pand2_1_1
timestamp 1626486988
transform 1 0 3594 0 -1 2828
box -36 -17 1430 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_pinv_1  sky130_sram_2kbyte_1rw1r_32x512_8_pinv_1_0
timestamp 1626486988
transform 1 0 3226 0 -1 2828
box -36 -17 404 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_7
timestamp 1626486988
transform 1 0 3039 0 1 848
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_6
timestamp 1626486988
transform 1 0 2955 0 1 466
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_5
timestamp 1626486988
transform 1 0 2871 0 1 104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_24
timestamp 1626486988
transform 1 0 3275 0 1 637
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_24
timestamp 1626486988
transform 1 0 3278 0 1 636
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_0
timestamp 1626486988
transform 1 0 9335 0 1 104
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_15
timestamp 1626486988
transform 1 0 9336 0 1 675
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_14
timestamp 1626486988
transform 1 0 9336 0 1 675
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_15
timestamp 1626486988
transform 1 0 9339 0 1 674
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_14
timestamp 1626486988
transform 1 0 9339 0 1 674
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_11
timestamp 1626486988
transform 1 0 11665 0 1 1377
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_10
timestamp 1626486988
transform 1 0 11665 0 1 -37
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_9
timestamp 1626486988
transform 1 0 11665 0 1 1377
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_11
timestamp 1626486988
transform 1 0 11666 0 1 1382
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_10
timestamp 1626486988
transform 1 0 11666 0 1 -32
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_9
timestamp 1626486988
transform 1 0 11666 0 1 1382
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_11
timestamp 1626486988
transform 1 0 11669 0 1 1381
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_10
timestamp 1626486988
transform 1 0 11669 0 1 -33
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_9
timestamp 1626486988
transform 1 0 11669 0 1 1381
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_pdriver_6  sky130_sram_2kbyte_1rw1r_32x512_8_pdriver_6_0
timestamp 1626486988
transform 1 0 3226 0 1 0
box -36 -17 8508 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_2
timestamp 1626486988
transform 1 0 2703 0 1 1534
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_23
timestamp 1626486988
transform 1 0 2872 0 1 2127
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_23
timestamp 1626486988
transform 1 0 3278 0 1 2126
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_4
timestamp 1626486988
transform 1 0 3039 0 1 2273
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_14
timestamp 1626486988
transform 1 0 3790 0 1 2273
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_13
timestamp 1626486988
transform 1 0 3790 0 1 2273
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_22
timestamp 1626486988
transform 1 0 3791 0 1 2278
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_21
timestamp 1626486988
transform 1 0 3791 0 1 2278
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_22
timestamp 1626486988
transform 1 0 3794 0 1 2277
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_21
timestamp 1626486988
transform 1 0 3794 0 1 2277
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_pand2_1  sky130_sram_2kbyte_1rw1r_32x512_8_pand2_1_0
timestamp 1626486988
transform 1 0 3226 0 1 2828
box -36 -17 1430 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_20
timestamp 1626486988
transform 1 0 4465 0 1 2104
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_20
timestamp 1626486988
transform 1 0 4462 0 1 2105
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_3
timestamp 1626486988
transform 1 0 4461 0 1 1534
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_6
timestamp 1626486988
transform 1 0 11669 0 1 2795
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_8
timestamp 1626486988
transform 1 0 11669 0 1 2795
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_6
timestamp 1626486988
transform 1 0 11666 0 1 2796
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_8
timestamp 1626486988
transform 1 0 11666 0 1 2796
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_6
timestamp 1626486988
transform 1 0 11665 0 1 2791
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_8
timestamp 1626486988
transform 1 0 11665 0 1 2791
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_27
timestamp 1626486988
transform 1 0 2620 0 1 4290
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_28
timestamp 1626486988
transform 1 0 1521 0 1 4290
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_35
timestamp 1626486988
transform 1 0 351 0 1 4130
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_19
timestamp 1626486988
transform 1 0 2872 0 1 3066
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_1
timestamp 1626486988
transform 1 0 2787 0 1 3482
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_18
timestamp 1626486988
transform 1 0 3040 0 1 3314
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_18
timestamp 1626486988
transform 1 0 3426 0 1 3313
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_19
timestamp 1626486988
transform 1 0 3326 0 1 3065
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_16
timestamp 1626486988
transform 1 0 4097 0 1 3486
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_17
timestamp 1626486988
transform 1 0 4097 0 1 3486
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_16
timestamp 1626486988
transform 1 0 4094 0 1 3487
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_17
timestamp 1626486988
transform 1 0 4094 0 1 3487
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_12
timestamp 1626486988
transform 1 0 4093 0 1 3482
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_34
timestamp 1626486988
transform 1 0 2872 0 1 4130
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_pand3_0  sky130_sram_2kbyte_1rw1r_32x512_8_pand3_0_0
timestamp 1626486988
transform 1 0 3226 0 -1 5656
box -36 -17 2718 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_5
timestamp 1626486988
transform 1 0 11669 0 1 4209
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_7
timestamp 1626486988
transform 1 0 11669 0 1 4209
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_5
timestamp 1626486988
transform 1 0 11666 0 1 4210
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_7
timestamp 1626486988
transform 1 0 11666 0 1 4210
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_5
timestamp 1626486988
transform 1 0 11665 0 1 4205
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_7
timestamp 1626486988
transform 1 0 11665 0 1 4205
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_32
timestamp 1626486988
transform 1 0 2620 0 1 5354
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_31
timestamp 1626486988
transform 1 0 2704 0 1 5230
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_26
timestamp 1626486988
transform 1 0 2788 0 1 5894
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_pnand2_1  sky130_sram_2kbyte_1rw1r_32x512_8_pnand2_1_0
timestamp 1626486988
transform 1 0 3226 0 1 5656
box -36 -17 504 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_30
timestamp 1626486988
transform 1 0 3040 0 1 5106
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_29
timestamp 1626486988
transform 1 0 4736 0 1 4917
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_30
timestamp 1626486988
transform 1 0 3293 0 1 5353
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_29
timestamp 1626486988
transform 1 0 3426 0 1 5229
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_28
timestamp 1626486988
transform 1 0 3559 0 1 5105
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_27
timestamp 1626486988
transform 1 0 4739 0 1 4916
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_26
timestamp 1626486988
transform 1 0 3326 0 1 5893
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_pdriver_3  sky130_sram_2kbyte_1rw1r_32x512_8_pdriver_3_0
timestamp 1626486988
transform 1 0 3694 0 1 5656
box -36 -17 5808 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_2
timestamp 1626486988
transform 1 0 11669 0 1 5623
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_4
timestamp 1626486988
transform 1 0 11669 0 1 5623
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_2
timestamp 1626486988
transform 1 0 11666 0 1 5624
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_4
timestamp 1626486988
transform 1 0 11666 0 1 5624
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_2
timestamp 1626486988
transform 1 0 11665 0 1 5619
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_4
timestamp 1626486988
transform 1 0 11665 0 1 5619
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_25
timestamp 1626486988
transform 1 0 3426 0 1 6141
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_25
timestamp 1626486988
transform 1 0 2620 0 1 6142
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_pdriver_3  sky130_sram_2kbyte_1rw1r_32x512_8_pdriver_3_1
timestamp 1626486988
transform 1 0 3226 0 -1 8484
box -36 -17 5808 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_12
timestamp 1626486988
transform 1 0 7973 0 1 6330
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_13
timestamp 1626486988
transform 1 0 7970 0 1 6331
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1
timestamp 1626486988
transform 1 0 11669 0 1 7037
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_3
timestamp 1626486988
transform 1 0 11669 0 1 7037
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_1
timestamp 1626486988
transform 1 0 11666 0 1 7038
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_3
timestamp 1626486988
transform 1 0 11666 0 1 7038
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_1
timestamp 1626486988
transform 1 0 11665 0 1 7033
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_3
timestamp 1626486988
transform 1 0 11665 0 1 7033
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_0
timestamp 1626486988
transform 1 0 11665 0 1 8447
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_33
timestamp 1626486988
transform 1 0 2704 0 1 7783
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_12
timestamp 1626486988
transform 1 0 7502 0 1 7745
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_0
timestamp 1626486988
transform 1 0 11666 0 1 8452
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_31
timestamp 1626486988
transform 1 0 3278 0 1 7782
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_13
timestamp 1626486988
transform 1 0 7505 0 1 7744
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_0
timestamp 1626486988
transform 1 0 11669 0 1 8451
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_delay_chain  sky130_sram_2kbyte_1rw1r_32x512_8_delay_chain_0
timestamp 1626486988
transform 1 0 0 0 -1 18382
box -75 -49 1876 12783
<< labels >>
rlabel metal3 s 1343 11263 1441 11361 4 vdd
rlabel metal3 s 607 8435 705 8533 4 vdd
rlabel metal3 s 11649 1365 11747 1463 4 vdd
rlabel metal3 s 11649 4193 11747 4291 4 vdd
rlabel metal3 s 1343 5607 1441 5705 4 vdd
rlabel metal3 s 607 11263 705 11361 4 vdd
rlabel metal3 s 607 5607 705 5705 4 vdd
rlabel metal3 s 1343 16919 1441 17017 4 vdd
rlabel metal3 s 1343 14091 1441 14189 4 vdd
rlabel metal3 s -49 1365 49 1463 4 vdd
rlabel metal3 s 607 14091 705 14189 4 vdd
rlabel metal3 s 11649 7021 11747 7119 4 vdd
rlabel metal3 s 607 16919 705 17017 4 vdd
rlabel metal3 s 1343 8435 1441 8533 4 vdd
rlabel metal3 s 11649 -49 11747 49 4 gnd
rlabel metal3 s 1343 7021 1441 7119 4 gnd
rlabel metal3 s 607 15505 705 15603 4 gnd
rlabel metal3 s 11649 2779 11747 2877 4 gnd
rlabel metal3 s 1343 9849 1441 9947 4 gnd
rlabel metal3 s 1343 12677 1441 12775 4 gnd
rlabel metal3 s 11649 5607 11747 5705 4 gnd
rlabel metal3 s 1343 18333 1441 18431 4 gnd
rlabel metal3 s 11649 8435 11747 8533 4 gnd
rlabel metal3 s 607 9849 705 9947 4 gnd
rlabel metal3 s 607 18333 705 18431 4 gnd
rlabel metal3 s 607 7021 705 7119 4 gnd
rlabel metal3 s -49 -49 49 49 4 gnd
rlabel metal3 s 1343 15505 1441 15603 4 gnd
rlabel metal3 s 607 12677 705 12775 4 gnd
rlabel metal2 s 137 538 203 590 4 csb
rlabel metal2 s 7534 7763 11782 7791 4 wl_en
rlabel metal2 s 4768 4935 11782 4963 4 s_en
rlabel metal2 s -57 17699 -29 17727 4 rbl_bl
rlabel metal2 s 8002 6349 11782 6377 4 p_en_bar
rlabel metal2 s 3293 655 3321 683 4 clk
rlabel metal2 s 9368 693 11782 721 4 clk_buf
<< properties >>
string FIXED_BBOX 0 0 11782 18542
<< end >>
