magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -2810 -1560 2809 1560
<< metal3 >>
rect -1550 193 1549 300
rect -1550 129 1465 193
rect 1529 129 1549 193
rect -1550 113 1549 129
rect -1550 49 1465 113
rect 1529 49 1549 113
rect -1550 33 1549 49
rect -1550 -31 1465 33
rect 1529 -31 1549 33
rect -1550 -47 1549 -31
rect -1550 -111 1465 -47
rect 1529 -111 1549 -47
rect -1550 -127 1549 -111
rect -1550 -191 1465 -127
rect 1529 -191 1549 -127
rect -1550 -207 1549 -191
rect -1550 -271 1465 -207
rect 1529 -271 1549 -207
rect -1550 -300 1549 -271
<< via3 >>
rect 1465 129 1529 193
rect 1465 49 1529 113
rect 1465 -31 1529 33
rect 1465 -111 1529 -47
rect 1465 -191 1529 -127
rect 1465 -271 1529 -207
<< mimcap >>
rect -1450 152 1350 200
rect -1450 -152 -1402 152
rect 1302 -152 1350 152
rect -1450 -200 1350 -152
<< mimcapcontact >>
rect -1402 -152 1302 152
<< metal4 >>
rect 1449 193 1545 234
rect -1411 152 1311 161
rect -1411 -152 -1402 152
rect 1302 -152 1311 152
rect -1411 -161 1311 -152
rect 1449 129 1465 193
rect 1529 129 1545 193
rect 1449 113 1545 129
rect 1449 49 1465 113
rect 1529 49 1545 113
rect 1449 33 1545 49
rect 1449 -31 1465 33
rect 1529 -31 1545 33
rect 1449 -47 1545 -31
rect 1449 -111 1465 -47
rect 1529 -111 1545 -47
rect 1449 -127 1545 -111
rect 1449 -191 1465 -127
rect 1529 -191 1545 -127
rect 1449 -207 1545 -191
rect 1449 -271 1465 -207
rect 1529 -271 1545 -207
rect 1449 -288 1545 -271
<< properties >>
string FIXED_BBOX -1550 -300 1450 300
<< end >>
