magic
tech sky130A
timestamp 1620271567
<< nmoslvt >>
rect -805 -150 -685 150
rect -656 -150 -536 150
rect -507 -150 -387 150
rect -358 -150 -238 150
rect -209 -150 -89 150
rect -60 -150 60 150
rect 89 -150 209 150
rect 238 -150 358 150
rect 387 -150 507 150
rect 536 -150 656 150
rect 685 -150 805 150
<< ndiff >>
rect -834 144 -805 150
rect -834 -144 -828 144
rect -811 -144 -805 144
rect -834 -150 -805 -144
rect -685 144 -656 150
rect -685 -144 -679 144
rect -662 -144 -656 144
rect -685 -150 -656 -144
rect -536 144 -507 150
rect -536 -144 -530 144
rect -513 -144 -507 144
rect -536 -150 -507 -144
rect -387 144 -358 150
rect -387 -144 -381 144
rect -364 -144 -358 144
rect -387 -150 -358 -144
rect -238 144 -209 150
rect -238 -144 -232 144
rect -215 -144 -209 144
rect -238 -150 -209 -144
rect -89 144 -60 150
rect -89 -144 -83 144
rect -66 -144 -60 144
rect -89 -150 -60 -144
rect 60 144 89 150
rect 60 -144 66 144
rect 83 -144 89 144
rect 60 -150 89 -144
rect 209 144 238 150
rect 209 -144 215 144
rect 232 -144 238 144
rect 209 -150 238 -144
rect 358 144 387 150
rect 358 -144 364 144
rect 381 -144 387 144
rect 358 -150 387 -144
rect 507 144 536 150
rect 507 -144 513 144
rect 530 -144 536 144
rect 507 -150 536 -144
rect 656 144 685 150
rect 656 -144 662 144
rect 679 -144 685 144
rect 656 -150 685 -144
rect 805 144 834 150
rect 805 -144 811 144
rect 828 -144 834 144
rect 805 -150 834 -144
<< ndiffc >>
rect -828 -144 -811 144
rect -679 -144 -662 144
rect -530 -144 -513 144
rect -381 -144 -364 144
rect -232 -144 -215 144
rect -83 -144 -66 144
rect 66 -144 83 144
rect 215 -144 232 144
rect 364 -144 381 144
rect 513 -144 530 144
rect 662 -144 679 144
rect 811 -144 828 144
<< poly >>
rect -805 186 -685 194
rect -805 169 -797 186
rect -693 169 -685 186
rect -805 150 -685 169
rect -656 186 -536 194
rect -656 169 -648 186
rect -544 169 -536 186
rect -656 150 -536 169
rect -507 186 -387 194
rect -507 169 -499 186
rect -395 169 -387 186
rect -507 150 -387 169
rect -358 186 -238 194
rect -358 169 -350 186
rect -246 169 -238 186
rect -358 150 -238 169
rect -209 186 -89 194
rect -209 169 -201 186
rect -97 169 -89 186
rect -209 150 -89 169
rect -60 186 60 194
rect -60 169 -52 186
rect 52 169 60 186
rect -60 150 60 169
rect 89 186 209 194
rect 89 169 97 186
rect 201 169 209 186
rect 89 150 209 169
rect 238 186 358 194
rect 238 169 246 186
rect 350 169 358 186
rect 238 150 358 169
rect 387 186 507 194
rect 387 169 395 186
rect 499 169 507 186
rect 387 150 507 169
rect 536 186 656 194
rect 536 169 544 186
rect 648 169 656 186
rect 536 150 656 169
rect 685 186 805 194
rect 685 169 693 186
rect 797 169 805 186
rect 685 150 805 169
rect -805 -169 -685 -150
rect -805 -186 -797 -169
rect -693 -186 -685 -169
rect -805 -194 -685 -186
rect -656 -169 -536 -150
rect -656 -186 -648 -169
rect -544 -186 -536 -169
rect -656 -194 -536 -186
rect -507 -169 -387 -150
rect -507 -186 -499 -169
rect -395 -186 -387 -169
rect -507 -194 -387 -186
rect -358 -169 -238 -150
rect -358 -186 -350 -169
rect -246 -186 -238 -169
rect -358 -194 -238 -186
rect -209 -169 -89 -150
rect -209 -186 -201 -169
rect -97 -186 -89 -169
rect -209 -194 -89 -186
rect -60 -169 60 -150
rect -60 -186 -52 -169
rect 52 -186 60 -169
rect -60 -194 60 -186
rect 89 -169 209 -150
rect 89 -186 97 -169
rect 201 -186 209 -169
rect 89 -194 209 -186
rect 238 -169 358 -150
rect 238 -186 246 -169
rect 350 -186 358 -169
rect 238 -194 358 -186
rect 387 -169 507 -150
rect 387 -186 395 -169
rect 499 -186 507 -169
rect 387 -194 507 -186
rect 536 -169 656 -150
rect 536 -186 544 -169
rect 648 -186 656 -169
rect 536 -194 656 -186
rect 685 -169 805 -150
rect 685 -186 693 -169
rect 797 -186 805 -169
rect 685 -194 805 -186
<< polycont >>
rect -797 169 -693 186
rect -648 169 -544 186
rect -499 169 -395 186
rect -350 169 -246 186
rect -201 169 -97 186
rect -52 169 52 186
rect 97 169 201 186
rect 246 169 350 186
rect 395 169 499 186
rect 544 169 648 186
rect 693 169 797 186
rect -797 -186 -693 -169
rect -648 -186 -544 -169
rect -499 -186 -395 -169
rect -350 -186 -246 -169
rect -201 -186 -97 -169
rect -52 -186 52 -169
rect 97 -186 201 -169
rect 246 -186 350 -169
rect 395 -186 499 -169
rect 544 -186 648 -169
rect 693 -186 797 -169
<< locali >>
rect -805 169 -797 186
rect -693 169 -685 186
rect -656 169 -648 186
rect -544 169 -536 186
rect -507 169 -499 186
rect -395 169 -387 186
rect -358 169 -350 186
rect -246 169 -238 186
rect -209 169 -201 186
rect -97 169 -89 186
rect -60 169 -52 186
rect 52 169 60 186
rect 89 169 97 186
rect 201 169 209 186
rect 238 169 246 186
rect 350 169 358 186
rect 387 169 395 186
rect 499 169 507 186
rect 536 169 544 186
rect 648 169 656 186
rect 685 169 693 186
rect 797 169 805 186
rect -828 144 -811 152
rect -828 -152 -811 -144
rect -679 144 -662 152
rect -679 -152 -662 -144
rect -530 144 -513 152
rect -530 -152 -513 -144
rect -381 144 -364 152
rect -381 -152 -364 -144
rect -232 144 -215 152
rect -232 -152 -215 -144
rect -83 144 -66 152
rect -83 -152 -66 -144
rect 66 144 83 152
rect 66 -152 83 -144
rect 215 144 232 152
rect 215 -152 232 -144
rect 364 144 381 152
rect 364 -152 381 -144
rect 513 144 530 152
rect 513 -152 530 -144
rect 662 144 679 152
rect 662 -152 679 -144
rect 811 144 828 152
rect 811 -152 828 -144
rect -805 -186 -797 -169
rect -693 -186 -685 -169
rect -656 -186 -648 -169
rect -544 -186 -536 -169
rect -507 -186 -499 -169
rect -395 -186 -387 -169
rect -358 -186 -350 -169
rect -246 -186 -238 -169
rect -209 -186 -201 -169
rect -97 -186 -89 -169
rect -60 -186 -52 -169
rect 52 -186 60 -169
rect 89 -186 97 -169
rect 201 -186 209 -169
rect 238 -186 246 -169
rect 350 -186 358 -169
rect 387 -186 395 -169
rect 499 -186 507 -169
rect 536 -186 544 -169
rect 648 -186 656 -169
rect 685 -186 693 -169
rect 797 -186 805 -169
<< viali >>
rect -797 169 -693 186
rect -648 169 -544 186
rect -499 169 -395 186
rect -350 169 -246 186
rect -201 169 -97 186
rect -52 169 52 186
rect 97 169 201 186
rect 246 169 350 186
rect 395 169 499 186
rect 544 169 648 186
rect 693 169 797 186
rect -828 -144 -811 144
rect -679 -144 -662 144
rect -530 -144 -513 144
rect -381 -144 -364 144
rect -232 -144 -215 144
rect -83 -144 -66 144
rect 66 -144 83 144
rect 215 -144 232 144
rect 364 -144 381 144
rect 513 -144 530 144
rect 662 -144 679 144
rect 811 -144 828 144
rect -797 -186 -693 -169
rect -648 -186 -544 -169
rect -499 -186 -395 -169
rect -350 -186 -246 -169
rect -201 -186 -97 -169
rect -52 -186 52 -169
rect 97 -186 201 -169
rect 246 -186 350 -169
rect 395 -186 499 -169
rect 544 -186 648 -169
rect 693 -186 797 -169
<< metal1 >>
rect -803 186 -687 189
rect -803 169 -797 186
rect -693 169 -687 186
rect -803 166 -687 169
rect -654 186 -538 189
rect -654 169 -648 186
rect -544 169 -538 186
rect -654 166 -538 169
rect -505 186 -389 189
rect -505 169 -499 186
rect -395 169 -389 186
rect -505 166 -389 169
rect -356 186 -240 189
rect -356 169 -350 186
rect -246 169 -240 186
rect -356 166 -240 169
rect -207 186 -91 189
rect -207 169 -201 186
rect -97 169 -91 186
rect -207 166 -91 169
rect -58 186 58 189
rect -58 169 -52 186
rect 52 169 58 186
rect -58 166 58 169
rect 91 186 207 189
rect 91 169 97 186
rect 201 169 207 186
rect 91 166 207 169
rect 240 186 356 189
rect 240 169 246 186
rect 350 169 356 186
rect 240 166 356 169
rect 389 186 505 189
rect 389 169 395 186
rect 499 169 505 186
rect 389 166 505 169
rect 538 186 654 189
rect 538 169 544 186
rect 648 169 654 186
rect 538 166 654 169
rect 687 186 803 189
rect 687 169 693 186
rect 797 169 803 186
rect 687 166 803 169
rect -831 144 -808 150
rect -831 -144 -828 144
rect -811 -144 -808 144
rect -831 -150 -808 -144
rect -682 144 -659 150
rect -682 -144 -679 144
rect -662 -144 -659 144
rect -682 -150 -659 -144
rect -533 144 -510 150
rect -533 -144 -530 144
rect -513 -144 -510 144
rect -533 -150 -510 -144
rect -384 144 -361 150
rect -384 -144 -381 144
rect -364 -144 -361 144
rect -384 -150 -361 -144
rect -235 144 -212 150
rect -235 -144 -232 144
rect -215 -144 -212 144
rect -235 -150 -212 -144
rect -86 144 -63 150
rect -86 -144 -83 144
rect -66 -144 -63 144
rect -86 -150 -63 -144
rect 63 144 86 150
rect 63 -144 66 144
rect 83 -144 86 144
rect 63 -150 86 -144
rect 212 144 235 150
rect 212 -144 215 144
rect 232 -144 235 144
rect 212 -150 235 -144
rect 361 144 384 150
rect 361 -144 364 144
rect 381 -144 384 144
rect 361 -150 384 -144
rect 510 144 533 150
rect 510 -144 513 144
rect 530 -144 533 144
rect 510 -150 533 -144
rect 659 144 682 150
rect 659 -144 662 144
rect 679 -144 682 144
rect 659 -150 682 -144
rect 808 144 831 150
rect 808 -144 811 144
rect 828 -144 831 144
rect 808 -150 831 -144
rect -803 -169 -687 -166
rect -803 -186 -797 -169
rect -693 -186 -687 -169
rect -803 -189 -687 -186
rect -654 -169 -538 -166
rect -654 -186 -648 -169
rect -544 -186 -538 -169
rect -654 -189 -538 -186
rect -505 -169 -389 -166
rect -505 -186 -499 -169
rect -395 -186 -389 -169
rect -505 -189 -389 -186
rect -356 -169 -240 -166
rect -356 -186 -350 -169
rect -246 -186 -240 -169
rect -356 -189 -240 -186
rect -207 -169 -91 -166
rect -207 -186 -201 -169
rect -97 -186 -91 -169
rect -207 -189 -91 -186
rect -58 -169 58 -166
rect -58 -186 -52 -169
rect 52 -186 58 -169
rect -58 -189 58 -186
rect 91 -169 207 -166
rect 91 -186 97 -169
rect 201 -186 207 -169
rect 91 -189 207 -186
rect 240 -169 356 -166
rect 240 -186 246 -169
rect 350 -186 356 -169
rect 240 -189 356 -186
rect 389 -169 505 -166
rect 389 -186 395 -169
rect 499 -186 505 -169
rect 389 -189 505 -186
rect 538 -169 654 -166
rect 538 -186 544 -169
rect 648 -186 654 -169
rect 538 -189 654 -186
rect 687 -169 803 -166
rect 687 -186 693 -169
rect 797 -186 803 -169
rect 687 -189 803 -186
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string parameters w 3 l 1.2 m 1 nf 11 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
