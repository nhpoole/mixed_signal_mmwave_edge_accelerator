magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -6463 -1448 6463 1448
<< pwell >>
rect -5203 -126 5203 126
<< nmos >>
rect -5119 -100 -4319 100
rect -4261 -100 -3461 100
rect -3403 -100 -2603 100
rect -2545 -100 -1745 100
rect -1687 -100 -887 100
rect -829 -100 -29 100
rect 29 -100 829 100
rect 887 -100 1687 100
rect 1745 -100 2545 100
rect 2603 -100 3403 100
rect 3461 -100 4261 100
rect 4319 -100 5119 100
<< ndiff >>
rect -5177 85 -5119 100
rect -5177 51 -5165 85
rect -5131 51 -5119 85
rect -5177 17 -5119 51
rect -5177 -17 -5165 17
rect -5131 -17 -5119 17
rect -5177 -51 -5119 -17
rect -5177 -85 -5165 -51
rect -5131 -85 -5119 -51
rect -5177 -100 -5119 -85
rect -4319 85 -4261 100
rect -4319 51 -4307 85
rect -4273 51 -4261 85
rect -4319 17 -4261 51
rect -4319 -17 -4307 17
rect -4273 -17 -4261 17
rect -4319 -51 -4261 -17
rect -4319 -85 -4307 -51
rect -4273 -85 -4261 -51
rect -4319 -100 -4261 -85
rect -3461 85 -3403 100
rect -3461 51 -3449 85
rect -3415 51 -3403 85
rect -3461 17 -3403 51
rect -3461 -17 -3449 17
rect -3415 -17 -3403 17
rect -3461 -51 -3403 -17
rect -3461 -85 -3449 -51
rect -3415 -85 -3403 -51
rect -3461 -100 -3403 -85
rect -2603 85 -2545 100
rect -2603 51 -2591 85
rect -2557 51 -2545 85
rect -2603 17 -2545 51
rect -2603 -17 -2591 17
rect -2557 -17 -2545 17
rect -2603 -51 -2545 -17
rect -2603 -85 -2591 -51
rect -2557 -85 -2545 -51
rect -2603 -100 -2545 -85
rect -1745 85 -1687 100
rect -1745 51 -1733 85
rect -1699 51 -1687 85
rect -1745 17 -1687 51
rect -1745 -17 -1733 17
rect -1699 -17 -1687 17
rect -1745 -51 -1687 -17
rect -1745 -85 -1733 -51
rect -1699 -85 -1687 -51
rect -1745 -100 -1687 -85
rect -887 85 -829 100
rect -887 51 -875 85
rect -841 51 -829 85
rect -887 17 -829 51
rect -887 -17 -875 17
rect -841 -17 -829 17
rect -887 -51 -829 -17
rect -887 -85 -875 -51
rect -841 -85 -829 -51
rect -887 -100 -829 -85
rect -29 85 29 100
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -100 29 -85
rect 829 85 887 100
rect 829 51 841 85
rect 875 51 887 85
rect 829 17 887 51
rect 829 -17 841 17
rect 875 -17 887 17
rect 829 -51 887 -17
rect 829 -85 841 -51
rect 875 -85 887 -51
rect 829 -100 887 -85
rect 1687 85 1745 100
rect 1687 51 1699 85
rect 1733 51 1745 85
rect 1687 17 1745 51
rect 1687 -17 1699 17
rect 1733 -17 1745 17
rect 1687 -51 1745 -17
rect 1687 -85 1699 -51
rect 1733 -85 1745 -51
rect 1687 -100 1745 -85
rect 2545 85 2603 100
rect 2545 51 2557 85
rect 2591 51 2603 85
rect 2545 17 2603 51
rect 2545 -17 2557 17
rect 2591 -17 2603 17
rect 2545 -51 2603 -17
rect 2545 -85 2557 -51
rect 2591 -85 2603 -51
rect 2545 -100 2603 -85
rect 3403 85 3461 100
rect 3403 51 3415 85
rect 3449 51 3461 85
rect 3403 17 3461 51
rect 3403 -17 3415 17
rect 3449 -17 3461 17
rect 3403 -51 3461 -17
rect 3403 -85 3415 -51
rect 3449 -85 3461 -51
rect 3403 -100 3461 -85
rect 4261 85 4319 100
rect 4261 51 4273 85
rect 4307 51 4319 85
rect 4261 17 4319 51
rect 4261 -17 4273 17
rect 4307 -17 4319 17
rect 4261 -51 4319 -17
rect 4261 -85 4273 -51
rect 4307 -85 4319 -51
rect 4261 -100 4319 -85
rect 5119 85 5177 100
rect 5119 51 5131 85
rect 5165 51 5177 85
rect 5119 17 5177 51
rect 5119 -17 5131 17
rect 5165 -17 5177 17
rect 5119 -51 5177 -17
rect 5119 -85 5131 -51
rect 5165 -85 5177 -51
rect 5119 -100 5177 -85
<< ndiffc >>
rect -5165 51 -5131 85
rect -5165 -17 -5131 17
rect -5165 -85 -5131 -51
rect -4307 51 -4273 85
rect -4307 -17 -4273 17
rect -4307 -85 -4273 -51
rect -3449 51 -3415 85
rect -3449 -17 -3415 17
rect -3449 -85 -3415 -51
rect -2591 51 -2557 85
rect -2591 -17 -2557 17
rect -2591 -85 -2557 -51
rect -1733 51 -1699 85
rect -1733 -17 -1699 17
rect -1733 -85 -1699 -51
rect -875 51 -841 85
rect -875 -17 -841 17
rect -875 -85 -841 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 841 51 875 85
rect 841 -17 875 17
rect 841 -85 875 -51
rect 1699 51 1733 85
rect 1699 -17 1733 17
rect 1699 -85 1733 -51
rect 2557 51 2591 85
rect 2557 -17 2591 17
rect 2557 -85 2591 -51
rect 3415 51 3449 85
rect 3415 -17 3449 17
rect 3415 -85 3449 -51
rect 4273 51 4307 85
rect 4273 -17 4307 17
rect 4273 -85 4307 -51
rect 5131 51 5165 85
rect 5131 -17 5165 17
rect 5131 -85 5165 -51
<< poly >>
rect -4965 172 -4473 188
rect -4965 155 -4940 172
rect -5119 138 -4940 155
rect -4906 138 -4872 172
rect -4838 138 -4804 172
rect -4770 138 -4736 172
rect -4702 138 -4668 172
rect -4634 138 -4600 172
rect -4566 138 -4532 172
rect -4498 155 -4473 172
rect -4107 172 -3615 188
rect -4107 155 -4082 172
rect -4498 138 -4319 155
rect -5119 100 -4319 138
rect -4261 138 -4082 155
rect -4048 138 -4014 172
rect -3980 138 -3946 172
rect -3912 138 -3878 172
rect -3844 138 -3810 172
rect -3776 138 -3742 172
rect -3708 138 -3674 172
rect -3640 155 -3615 172
rect -3249 172 -2757 188
rect -3249 155 -3224 172
rect -3640 138 -3461 155
rect -4261 100 -3461 138
rect -3403 138 -3224 155
rect -3190 138 -3156 172
rect -3122 138 -3088 172
rect -3054 138 -3020 172
rect -2986 138 -2952 172
rect -2918 138 -2884 172
rect -2850 138 -2816 172
rect -2782 155 -2757 172
rect -2391 172 -1899 188
rect -2391 155 -2366 172
rect -2782 138 -2603 155
rect -3403 100 -2603 138
rect -2545 138 -2366 155
rect -2332 138 -2298 172
rect -2264 138 -2230 172
rect -2196 138 -2162 172
rect -2128 138 -2094 172
rect -2060 138 -2026 172
rect -1992 138 -1958 172
rect -1924 155 -1899 172
rect -1533 172 -1041 188
rect -1533 155 -1508 172
rect -1924 138 -1745 155
rect -2545 100 -1745 138
rect -1687 138 -1508 155
rect -1474 138 -1440 172
rect -1406 138 -1372 172
rect -1338 138 -1304 172
rect -1270 138 -1236 172
rect -1202 138 -1168 172
rect -1134 138 -1100 172
rect -1066 155 -1041 172
rect -675 172 -183 188
rect -675 155 -650 172
rect -1066 138 -887 155
rect -1687 100 -887 138
rect -829 138 -650 155
rect -616 138 -582 172
rect -548 138 -514 172
rect -480 138 -446 172
rect -412 138 -378 172
rect -344 138 -310 172
rect -276 138 -242 172
rect -208 155 -183 172
rect 183 172 675 188
rect 183 155 208 172
rect -208 138 -29 155
rect -829 100 -29 138
rect 29 138 208 155
rect 242 138 276 172
rect 310 138 344 172
rect 378 138 412 172
rect 446 138 480 172
rect 514 138 548 172
rect 582 138 616 172
rect 650 155 675 172
rect 1041 172 1533 188
rect 1041 155 1066 172
rect 650 138 829 155
rect 29 100 829 138
rect 887 138 1066 155
rect 1100 138 1134 172
rect 1168 138 1202 172
rect 1236 138 1270 172
rect 1304 138 1338 172
rect 1372 138 1406 172
rect 1440 138 1474 172
rect 1508 155 1533 172
rect 1899 172 2391 188
rect 1899 155 1924 172
rect 1508 138 1687 155
rect 887 100 1687 138
rect 1745 138 1924 155
rect 1958 138 1992 172
rect 2026 138 2060 172
rect 2094 138 2128 172
rect 2162 138 2196 172
rect 2230 138 2264 172
rect 2298 138 2332 172
rect 2366 155 2391 172
rect 2757 172 3249 188
rect 2757 155 2782 172
rect 2366 138 2545 155
rect 1745 100 2545 138
rect 2603 138 2782 155
rect 2816 138 2850 172
rect 2884 138 2918 172
rect 2952 138 2986 172
rect 3020 138 3054 172
rect 3088 138 3122 172
rect 3156 138 3190 172
rect 3224 155 3249 172
rect 3615 172 4107 188
rect 3615 155 3640 172
rect 3224 138 3403 155
rect 2603 100 3403 138
rect 3461 138 3640 155
rect 3674 138 3708 172
rect 3742 138 3776 172
rect 3810 138 3844 172
rect 3878 138 3912 172
rect 3946 138 3980 172
rect 4014 138 4048 172
rect 4082 155 4107 172
rect 4473 172 4965 188
rect 4473 155 4498 172
rect 4082 138 4261 155
rect 3461 100 4261 138
rect 4319 138 4498 155
rect 4532 138 4566 172
rect 4600 138 4634 172
rect 4668 138 4702 172
rect 4736 138 4770 172
rect 4804 138 4838 172
rect 4872 138 4906 172
rect 4940 155 4965 172
rect 4940 138 5119 155
rect 4319 100 5119 138
rect -5119 -138 -4319 -100
rect -5119 -155 -4940 -138
rect -4965 -172 -4940 -155
rect -4906 -172 -4872 -138
rect -4838 -172 -4804 -138
rect -4770 -172 -4736 -138
rect -4702 -172 -4668 -138
rect -4634 -172 -4600 -138
rect -4566 -172 -4532 -138
rect -4498 -155 -4319 -138
rect -4261 -138 -3461 -100
rect -4261 -155 -4082 -138
rect -4498 -172 -4473 -155
rect -4965 -188 -4473 -172
rect -4107 -172 -4082 -155
rect -4048 -172 -4014 -138
rect -3980 -172 -3946 -138
rect -3912 -172 -3878 -138
rect -3844 -172 -3810 -138
rect -3776 -172 -3742 -138
rect -3708 -172 -3674 -138
rect -3640 -155 -3461 -138
rect -3403 -138 -2603 -100
rect -3403 -155 -3224 -138
rect -3640 -172 -3615 -155
rect -4107 -188 -3615 -172
rect -3249 -172 -3224 -155
rect -3190 -172 -3156 -138
rect -3122 -172 -3088 -138
rect -3054 -172 -3020 -138
rect -2986 -172 -2952 -138
rect -2918 -172 -2884 -138
rect -2850 -172 -2816 -138
rect -2782 -155 -2603 -138
rect -2545 -138 -1745 -100
rect -2545 -155 -2366 -138
rect -2782 -172 -2757 -155
rect -3249 -188 -2757 -172
rect -2391 -172 -2366 -155
rect -2332 -172 -2298 -138
rect -2264 -172 -2230 -138
rect -2196 -172 -2162 -138
rect -2128 -172 -2094 -138
rect -2060 -172 -2026 -138
rect -1992 -172 -1958 -138
rect -1924 -155 -1745 -138
rect -1687 -138 -887 -100
rect -1687 -155 -1508 -138
rect -1924 -172 -1899 -155
rect -2391 -188 -1899 -172
rect -1533 -172 -1508 -155
rect -1474 -172 -1440 -138
rect -1406 -172 -1372 -138
rect -1338 -172 -1304 -138
rect -1270 -172 -1236 -138
rect -1202 -172 -1168 -138
rect -1134 -172 -1100 -138
rect -1066 -155 -887 -138
rect -829 -138 -29 -100
rect -829 -155 -650 -138
rect -1066 -172 -1041 -155
rect -1533 -188 -1041 -172
rect -675 -172 -650 -155
rect -616 -172 -582 -138
rect -548 -172 -514 -138
rect -480 -172 -446 -138
rect -412 -172 -378 -138
rect -344 -172 -310 -138
rect -276 -172 -242 -138
rect -208 -155 -29 -138
rect 29 -138 829 -100
rect 29 -155 208 -138
rect -208 -172 -183 -155
rect -675 -188 -183 -172
rect 183 -172 208 -155
rect 242 -172 276 -138
rect 310 -172 344 -138
rect 378 -172 412 -138
rect 446 -172 480 -138
rect 514 -172 548 -138
rect 582 -172 616 -138
rect 650 -155 829 -138
rect 887 -138 1687 -100
rect 887 -155 1066 -138
rect 650 -172 675 -155
rect 183 -188 675 -172
rect 1041 -172 1066 -155
rect 1100 -172 1134 -138
rect 1168 -172 1202 -138
rect 1236 -172 1270 -138
rect 1304 -172 1338 -138
rect 1372 -172 1406 -138
rect 1440 -172 1474 -138
rect 1508 -155 1687 -138
rect 1745 -138 2545 -100
rect 1745 -155 1924 -138
rect 1508 -172 1533 -155
rect 1041 -188 1533 -172
rect 1899 -172 1924 -155
rect 1958 -172 1992 -138
rect 2026 -172 2060 -138
rect 2094 -172 2128 -138
rect 2162 -172 2196 -138
rect 2230 -172 2264 -138
rect 2298 -172 2332 -138
rect 2366 -155 2545 -138
rect 2603 -138 3403 -100
rect 2603 -155 2782 -138
rect 2366 -172 2391 -155
rect 1899 -188 2391 -172
rect 2757 -172 2782 -155
rect 2816 -172 2850 -138
rect 2884 -172 2918 -138
rect 2952 -172 2986 -138
rect 3020 -172 3054 -138
rect 3088 -172 3122 -138
rect 3156 -172 3190 -138
rect 3224 -155 3403 -138
rect 3461 -138 4261 -100
rect 3461 -155 3640 -138
rect 3224 -172 3249 -155
rect 2757 -188 3249 -172
rect 3615 -172 3640 -155
rect 3674 -172 3708 -138
rect 3742 -172 3776 -138
rect 3810 -172 3844 -138
rect 3878 -172 3912 -138
rect 3946 -172 3980 -138
rect 4014 -172 4048 -138
rect 4082 -155 4261 -138
rect 4319 -138 5119 -100
rect 4319 -155 4498 -138
rect 4082 -172 4107 -155
rect 3615 -188 4107 -172
rect 4473 -172 4498 -155
rect 4532 -172 4566 -138
rect 4600 -172 4634 -138
rect 4668 -172 4702 -138
rect 4736 -172 4770 -138
rect 4804 -172 4838 -138
rect 4872 -172 4906 -138
rect 4940 -155 5119 -138
rect 4940 -172 4965 -155
rect 4473 -188 4965 -172
<< polycont >>
rect -4940 138 -4906 172
rect -4872 138 -4838 172
rect -4804 138 -4770 172
rect -4736 138 -4702 172
rect -4668 138 -4634 172
rect -4600 138 -4566 172
rect -4532 138 -4498 172
rect -4082 138 -4048 172
rect -4014 138 -3980 172
rect -3946 138 -3912 172
rect -3878 138 -3844 172
rect -3810 138 -3776 172
rect -3742 138 -3708 172
rect -3674 138 -3640 172
rect -3224 138 -3190 172
rect -3156 138 -3122 172
rect -3088 138 -3054 172
rect -3020 138 -2986 172
rect -2952 138 -2918 172
rect -2884 138 -2850 172
rect -2816 138 -2782 172
rect -2366 138 -2332 172
rect -2298 138 -2264 172
rect -2230 138 -2196 172
rect -2162 138 -2128 172
rect -2094 138 -2060 172
rect -2026 138 -1992 172
rect -1958 138 -1924 172
rect -1508 138 -1474 172
rect -1440 138 -1406 172
rect -1372 138 -1338 172
rect -1304 138 -1270 172
rect -1236 138 -1202 172
rect -1168 138 -1134 172
rect -1100 138 -1066 172
rect -650 138 -616 172
rect -582 138 -548 172
rect -514 138 -480 172
rect -446 138 -412 172
rect -378 138 -344 172
rect -310 138 -276 172
rect -242 138 -208 172
rect 208 138 242 172
rect 276 138 310 172
rect 344 138 378 172
rect 412 138 446 172
rect 480 138 514 172
rect 548 138 582 172
rect 616 138 650 172
rect 1066 138 1100 172
rect 1134 138 1168 172
rect 1202 138 1236 172
rect 1270 138 1304 172
rect 1338 138 1372 172
rect 1406 138 1440 172
rect 1474 138 1508 172
rect 1924 138 1958 172
rect 1992 138 2026 172
rect 2060 138 2094 172
rect 2128 138 2162 172
rect 2196 138 2230 172
rect 2264 138 2298 172
rect 2332 138 2366 172
rect 2782 138 2816 172
rect 2850 138 2884 172
rect 2918 138 2952 172
rect 2986 138 3020 172
rect 3054 138 3088 172
rect 3122 138 3156 172
rect 3190 138 3224 172
rect 3640 138 3674 172
rect 3708 138 3742 172
rect 3776 138 3810 172
rect 3844 138 3878 172
rect 3912 138 3946 172
rect 3980 138 4014 172
rect 4048 138 4082 172
rect 4498 138 4532 172
rect 4566 138 4600 172
rect 4634 138 4668 172
rect 4702 138 4736 172
rect 4770 138 4804 172
rect 4838 138 4872 172
rect 4906 138 4940 172
rect -4940 -172 -4906 -138
rect -4872 -172 -4838 -138
rect -4804 -172 -4770 -138
rect -4736 -172 -4702 -138
rect -4668 -172 -4634 -138
rect -4600 -172 -4566 -138
rect -4532 -172 -4498 -138
rect -4082 -172 -4048 -138
rect -4014 -172 -3980 -138
rect -3946 -172 -3912 -138
rect -3878 -172 -3844 -138
rect -3810 -172 -3776 -138
rect -3742 -172 -3708 -138
rect -3674 -172 -3640 -138
rect -3224 -172 -3190 -138
rect -3156 -172 -3122 -138
rect -3088 -172 -3054 -138
rect -3020 -172 -2986 -138
rect -2952 -172 -2918 -138
rect -2884 -172 -2850 -138
rect -2816 -172 -2782 -138
rect -2366 -172 -2332 -138
rect -2298 -172 -2264 -138
rect -2230 -172 -2196 -138
rect -2162 -172 -2128 -138
rect -2094 -172 -2060 -138
rect -2026 -172 -1992 -138
rect -1958 -172 -1924 -138
rect -1508 -172 -1474 -138
rect -1440 -172 -1406 -138
rect -1372 -172 -1338 -138
rect -1304 -172 -1270 -138
rect -1236 -172 -1202 -138
rect -1168 -172 -1134 -138
rect -1100 -172 -1066 -138
rect -650 -172 -616 -138
rect -582 -172 -548 -138
rect -514 -172 -480 -138
rect -446 -172 -412 -138
rect -378 -172 -344 -138
rect -310 -172 -276 -138
rect -242 -172 -208 -138
rect 208 -172 242 -138
rect 276 -172 310 -138
rect 344 -172 378 -138
rect 412 -172 446 -138
rect 480 -172 514 -138
rect 548 -172 582 -138
rect 616 -172 650 -138
rect 1066 -172 1100 -138
rect 1134 -172 1168 -138
rect 1202 -172 1236 -138
rect 1270 -172 1304 -138
rect 1338 -172 1372 -138
rect 1406 -172 1440 -138
rect 1474 -172 1508 -138
rect 1924 -172 1958 -138
rect 1992 -172 2026 -138
rect 2060 -172 2094 -138
rect 2128 -172 2162 -138
rect 2196 -172 2230 -138
rect 2264 -172 2298 -138
rect 2332 -172 2366 -138
rect 2782 -172 2816 -138
rect 2850 -172 2884 -138
rect 2918 -172 2952 -138
rect 2986 -172 3020 -138
rect 3054 -172 3088 -138
rect 3122 -172 3156 -138
rect 3190 -172 3224 -138
rect 3640 -172 3674 -138
rect 3708 -172 3742 -138
rect 3776 -172 3810 -138
rect 3844 -172 3878 -138
rect 3912 -172 3946 -138
rect 3980 -172 4014 -138
rect 4048 -172 4082 -138
rect 4498 -172 4532 -138
rect 4566 -172 4600 -138
rect 4634 -172 4668 -138
rect 4702 -172 4736 -138
rect 4770 -172 4804 -138
rect 4838 -172 4872 -138
rect 4906 -172 4940 -138
<< locali >>
rect -4965 138 -4940 172
rect -4906 138 -4880 172
rect -4838 138 -4808 172
rect -4770 138 -4736 172
rect -4702 138 -4668 172
rect -4630 138 -4600 172
rect -4558 138 -4532 172
rect -4498 138 -4473 172
rect -4107 138 -4082 172
rect -4048 138 -4022 172
rect -3980 138 -3950 172
rect -3912 138 -3878 172
rect -3844 138 -3810 172
rect -3772 138 -3742 172
rect -3700 138 -3674 172
rect -3640 138 -3615 172
rect -3249 138 -3224 172
rect -3190 138 -3164 172
rect -3122 138 -3092 172
rect -3054 138 -3020 172
rect -2986 138 -2952 172
rect -2914 138 -2884 172
rect -2842 138 -2816 172
rect -2782 138 -2757 172
rect -2391 138 -2366 172
rect -2332 138 -2306 172
rect -2264 138 -2234 172
rect -2196 138 -2162 172
rect -2128 138 -2094 172
rect -2056 138 -2026 172
rect -1984 138 -1958 172
rect -1924 138 -1899 172
rect -1533 138 -1508 172
rect -1474 138 -1448 172
rect -1406 138 -1376 172
rect -1338 138 -1304 172
rect -1270 138 -1236 172
rect -1198 138 -1168 172
rect -1126 138 -1100 172
rect -1066 138 -1041 172
rect -675 138 -650 172
rect -616 138 -590 172
rect -548 138 -518 172
rect -480 138 -446 172
rect -412 138 -378 172
rect -340 138 -310 172
rect -268 138 -242 172
rect -208 138 -183 172
rect 183 138 208 172
rect 242 138 268 172
rect 310 138 340 172
rect 378 138 412 172
rect 446 138 480 172
rect 518 138 548 172
rect 590 138 616 172
rect 650 138 675 172
rect 1041 138 1066 172
rect 1100 138 1126 172
rect 1168 138 1198 172
rect 1236 138 1270 172
rect 1304 138 1338 172
rect 1376 138 1406 172
rect 1448 138 1474 172
rect 1508 138 1533 172
rect 1899 138 1924 172
rect 1958 138 1984 172
rect 2026 138 2056 172
rect 2094 138 2128 172
rect 2162 138 2196 172
rect 2234 138 2264 172
rect 2306 138 2332 172
rect 2366 138 2391 172
rect 2757 138 2782 172
rect 2816 138 2842 172
rect 2884 138 2914 172
rect 2952 138 2986 172
rect 3020 138 3054 172
rect 3092 138 3122 172
rect 3164 138 3190 172
rect 3224 138 3249 172
rect 3615 138 3640 172
rect 3674 138 3700 172
rect 3742 138 3772 172
rect 3810 138 3844 172
rect 3878 138 3912 172
rect 3950 138 3980 172
rect 4022 138 4048 172
rect 4082 138 4107 172
rect 4473 138 4498 172
rect 4532 138 4558 172
rect 4600 138 4630 172
rect 4668 138 4702 172
rect 4736 138 4770 172
rect 4808 138 4838 172
rect 4880 138 4906 172
rect 4940 138 4965 172
rect -5165 85 -5131 104
rect -5165 17 -5131 19
rect -5165 -19 -5131 -17
rect -5165 -104 -5131 -85
rect -4307 85 -4273 104
rect -4307 17 -4273 19
rect -4307 -19 -4273 -17
rect -4307 -104 -4273 -85
rect -3449 85 -3415 104
rect -3449 17 -3415 19
rect -3449 -19 -3415 -17
rect -3449 -104 -3415 -85
rect -2591 85 -2557 104
rect -2591 17 -2557 19
rect -2591 -19 -2557 -17
rect -2591 -104 -2557 -85
rect -1733 85 -1699 104
rect -1733 17 -1699 19
rect -1733 -19 -1699 -17
rect -1733 -104 -1699 -85
rect -875 85 -841 104
rect -875 17 -841 19
rect -875 -19 -841 -17
rect -875 -104 -841 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 841 85 875 104
rect 841 17 875 19
rect 841 -19 875 -17
rect 841 -104 875 -85
rect 1699 85 1733 104
rect 1699 17 1733 19
rect 1699 -19 1733 -17
rect 1699 -104 1733 -85
rect 2557 85 2591 104
rect 2557 17 2591 19
rect 2557 -19 2591 -17
rect 2557 -104 2591 -85
rect 3415 85 3449 104
rect 3415 17 3449 19
rect 3415 -19 3449 -17
rect 3415 -104 3449 -85
rect 4273 85 4307 104
rect 4273 17 4307 19
rect 4273 -19 4307 -17
rect 4273 -104 4307 -85
rect 5131 85 5165 104
rect 5131 17 5165 19
rect 5131 -19 5165 -17
rect 5131 -104 5165 -85
rect -4965 -172 -4940 -138
rect -4906 -172 -4880 -138
rect -4838 -172 -4808 -138
rect -4770 -172 -4736 -138
rect -4702 -172 -4668 -138
rect -4630 -172 -4600 -138
rect -4558 -172 -4532 -138
rect -4498 -172 -4473 -138
rect -4107 -172 -4082 -138
rect -4048 -172 -4022 -138
rect -3980 -172 -3950 -138
rect -3912 -172 -3878 -138
rect -3844 -172 -3810 -138
rect -3772 -172 -3742 -138
rect -3700 -172 -3674 -138
rect -3640 -172 -3615 -138
rect -3249 -172 -3224 -138
rect -3190 -172 -3164 -138
rect -3122 -172 -3092 -138
rect -3054 -172 -3020 -138
rect -2986 -172 -2952 -138
rect -2914 -172 -2884 -138
rect -2842 -172 -2816 -138
rect -2782 -172 -2757 -138
rect -2391 -172 -2366 -138
rect -2332 -172 -2306 -138
rect -2264 -172 -2234 -138
rect -2196 -172 -2162 -138
rect -2128 -172 -2094 -138
rect -2056 -172 -2026 -138
rect -1984 -172 -1958 -138
rect -1924 -172 -1899 -138
rect -1533 -172 -1508 -138
rect -1474 -172 -1448 -138
rect -1406 -172 -1376 -138
rect -1338 -172 -1304 -138
rect -1270 -172 -1236 -138
rect -1198 -172 -1168 -138
rect -1126 -172 -1100 -138
rect -1066 -172 -1041 -138
rect -675 -172 -650 -138
rect -616 -172 -590 -138
rect -548 -172 -518 -138
rect -480 -172 -446 -138
rect -412 -172 -378 -138
rect -340 -172 -310 -138
rect -268 -172 -242 -138
rect -208 -172 -183 -138
rect 183 -172 208 -138
rect 242 -172 268 -138
rect 310 -172 340 -138
rect 378 -172 412 -138
rect 446 -172 480 -138
rect 518 -172 548 -138
rect 590 -172 616 -138
rect 650 -172 675 -138
rect 1041 -172 1066 -138
rect 1100 -172 1126 -138
rect 1168 -172 1198 -138
rect 1236 -172 1270 -138
rect 1304 -172 1338 -138
rect 1376 -172 1406 -138
rect 1448 -172 1474 -138
rect 1508 -172 1533 -138
rect 1899 -172 1924 -138
rect 1958 -172 1984 -138
rect 2026 -172 2056 -138
rect 2094 -172 2128 -138
rect 2162 -172 2196 -138
rect 2234 -172 2264 -138
rect 2306 -172 2332 -138
rect 2366 -172 2391 -138
rect 2757 -172 2782 -138
rect 2816 -172 2842 -138
rect 2884 -172 2914 -138
rect 2952 -172 2986 -138
rect 3020 -172 3054 -138
rect 3092 -172 3122 -138
rect 3164 -172 3190 -138
rect 3224 -172 3249 -138
rect 3615 -172 3640 -138
rect 3674 -172 3700 -138
rect 3742 -172 3772 -138
rect 3810 -172 3844 -138
rect 3878 -172 3912 -138
rect 3950 -172 3980 -138
rect 4022 -172 4048 -138
rect 4082 -172 4107 -138
rect 4473 -172 4498 -138
rect 4532 -172 4558 -138
rect 4600 -172 4630 -138
rect 4668 -172 4702 -138
rect 4736 -172 4770 -138
rect 4808 -172 4838 -138
rect 4880 -172 4906 -138
rect 4940 -172 4965 -138
<< viali >>
rect -4880 138 -4872 172
rect -4872 138 -4846 172
rect -4808 138 -4804 172
rect -4804 138 -4774 172
rect -4736 138 -4702 172
rect -4664 138 -4634 172
rect -4634 138 -4630 172
rect -4592 138 -4566 172
rect -4566 138 -4558 172
rect -4022 138 -4014 172
rect -4014 138 -3988 172
rect -3950 138 -3946 172
rect -3946 138 -3916 172
rect -3878 138 -3844 172
rect -3806 138 -3776 172
rect -3776 138 -3772 172
rect -3734 138 -3708 172
rect -3708 138 -3700 172
rect -3164 138 -3156 172
rect -3156 138 -3130 172
rect -3092 138 -3088 172
rect -3088 138 -3058 172
rect -3020 138 -2986 172
rect -2948 138 -2918 172
rect -2918 138 -2914 172
rect -2876 138 -2850 172
rect -2850 138 -2842 172
rect -2306 138 -2298 172
rect -2298 138 -2272 172
rect -2234 138 -2230 172
rect -2230 138 -2200 172
rect -2162 138 -2128 172
rect -2090 138 -2060 172
rect -2060 138 -2056 172
rect -2018 138 -1992 172
rect -1992 138 -1984 172
rect -1448 138 -1440 172
rect -1440 138 -1414 172
rect -1376 138 -1372 172
rect -1372 138 -1342 172
rect -1304 138 -1270 172
rect -1232 138 -1202 172
rect -1202 138 -1198 172
rect -1160 138 -1134 172
rect -1134 138 -1126 172
rect -590 138 -582 172
rect -582 138 -556 172
rect -518 138 -514 172
rect -514 138 -484 172
rect -446 138 -412 172
rect -374 138 -344 172
rect -344 138 -340 172
rect -302 138 -276 172
rect -276 138 -268 172
rect 268 138 276 172
rect 276 138 302 172
rect 340 138 344 172
rect 344 138 374 172
rect 412 138 446 172
rect 484 138 514 172
rect 514 138 518 172
rect 556 138 582 172
rect 582 138 590 172
rect 1126 138 1134 172
rect 1134 138 1160 172
rect 1198 138 1202 172
rect 1202 138 1232 172
rect 1270 138 1304 172
rect 1342 138 1372 172
rect 1372 138 1376 172
rect 1414 138 1440 172
rect 1440 138 1448 172
rect 1984 138 1992 172
rect 1992 138 2018 172
rect 2056 138 2060 172
rect 2060 138 2090 172
rect 2128 138 2162 172
rect 2200 138 2230 172
rect 2230 138 2234 172
rect 2272 138 2298 172
rect 2298 138 2306 172
rect 2842 138 2850 172
rect 2850 138 2876 172
rect 2914 138 2918 172
rect 2918 138 2948 172
rect 2986 138 3020 172
rect 3058 138 3088 172
rect 3088 138 3092 172
rect 3130 138 3156 172
rect 3156 138 3164 172
rect 3700 138 3708 172
rect 3708 138 3734 172
rect 3772 138 3776 172
rect 3776 138 3806 172
rect 3844 138 3878 172
rect 3916 138 3946 172
rect 3946 138 3950 172
rect 3988 138 4014 172
rect 4014 138 4022 172
rect 4558 138 4566 172
rect 4566 138 4592 172
rect 4630 138 4634 172
rect 4634 138 4664 172
rect 4702 138 4736 172
rect 4774 138 4804 172
rect 4804 138 4808 172
rect 4846 138 4872 172
rect 4872 138 4880 172
rect -5165 51 -5131 53
rect -5165 19 -5131 51
rect -5165 -51 -5131 -19
rect -5165 -53 -5131 -51
rect -4307 51 -4273 53
rect -4307 19 -4273 51
rect -4307 -51 -4273 -19
rect -4307 -53 -4273 -51
rect -3449 51 -3415 53
rect -3449 19 -3415 51
rect -3449 -51 -3415 -19
rect -3449 -53 -3415 -51
rect -2591 51 -2557 53
rect -2591 19 -2557 51
rect -2591 -51 -2557 -19
rect -2591 -53 -2557 -51
rect -1733 51 -1699 53
rect -1733 19 -1699 51
rect -1733 -51 -1699 -19
rect -1733 -53 -1699 -51
rect -875 51 -841 53
rect -875 19 -841 51
rect -875 -51 -841 -19
rect -875 -53 -841 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 841 51 875 53
rect 841 19 875 51
rect 841 -51 875 -19
rect 841 -53 875 -51
rect 1699 51 1733 53
rect 1699 19 1733 51
rect 1699 -51 1733 -19
rect 1699 -53 1733 -51
rect 2557 51 2591 53
rect 2557 19 2591 51
rect 2557 -51 2591 -19
rect 2557 -53 2591 -51
rect 3415 51 3449 53
rect 3415 19 3449 51
rect 3415 -51 3449 -19
rect 3415 -53 3449 -51
rect 4273 51 4307 53
rect 4273 19 4307 51
rect 4273 -51 4307 -19
rect 4273 -53 4307 -51
rect 5131 51 5165 53
rect 5131 19 5165 51
rect 5131 -51 5165 -19
rect 5131 -53 5165 -51
rect -4880 -172 -4872 -138
rect -4872 -172 -4846 -138
rect -4808 -172 -4804 -138
rect -4804 -172 -4774 -138
rect -4736 -172 -4702 -138
rect -4664 -172 -4634 -138
rect -4634 -172 -4630 -138
rect -4592 -172 -4566 -138
rect -4566 -172 -4558 -138
rect -4022 -172 -4014 -138
rect -4014 -172 -3988 -138
rect -3950 -172 -3946 -138
rect -3946 -172 -3916 -138
rect -3878 -172 -3844 -138
rect -3806 -172 -3776 -138
rect -3776 -172 -3772 -138
rect -3734 -172 -3708 -138
rect -3708 -172 -3700 -138
rect -3164 -172 -3156 -138
rect -3156 -172 -3130 -138
rect -3092 -172 -3088 -138
rect -3088 -172 -3058 -138
rect -3020 -172 -2986 -138
rect -2948 -172 -2918 -138
rect -2918 -172 -2914 -138
rect -2876 -172 -2850 -138
rect -2850 -172 -2842 -138
rect -2306 -172 -2298 -138
rect -2298 -172 -2272 -138
rect -2234 -172 -2230 -138
rect -2230 -172 -2200 -138
rect -2162 -172 -2128 -138
rect -2090 -172 -2060 -138
rect -2060 -172 -2056 -138
rect -2018 -172 -1992 -138
rect -1992 -172 -1984 -138
rect -1448 -172 -1440 -138
rect -1440 -172 -1414 -138
rect -1376 -172 -1372 -138
rect -1372 -172 -1342 -138
rect -1304 -172 -1270 -138
rect -1232 -172 -1202 -138
rect -1202 -172 -1198 -138
rect -1160 -172 -1134 -138
rect -1134 -172 -1126 -138
rect -590 -172 -582 -138
rect -582 -172 -556 -138
rect -518 -172 -514 -138
rect -514 -172 -484 -138
rect -446 -172 -412 -138
rect -374 -172 -344 -138
rect -344 -172 -340 -138
rect -302 -172 -276 -138
rect -276 -172 -268 -138
rect 268 -172 276 -138
rect 276 -172 302 -138
rect 340 -172 344 -138
rect 344 -172 374 -138
rect 412 -172 446 -138
rect 484 -172 514 -138
rect 514 -172 518 -138
rect 556 -172 582 -138
rect 582 -172 590 -138
rect 1126 -172 1134 -138
rect 1134 -172 1160 -138
rect 1198 -172 1202 -138
rect 1202 -172 1232 -138
rect 1270 -172 1304 -138
rect 1342 -172 1372 -138
rect 1372 -172 1376 -138
rect 1414 -172 1440 -138
rect 1440 -172 1448 -138
rect 1984 -172 1992 -138
rect 1992 -172 2018 -138
rect 2056 -172 2060 -138
rect 2060 -172 2090 -138
rect 2128 -172 2162 -138
rect 2200 -172 2230 -138
rect 2230 -172 2234 -138
rect 2272 -172 2298 -138
rect 2298 -172 2306 -138
rect 2842 -172 2850 -138
rect 2850 -172 2876 -138
rect 2914 -172 2918 -138
rect 2918 -172 2948 -138
rect 2986 -172 3020 -138
rect 3058 -172 3088 -138
rect 3088 -172 3092 -138
rect 3130 -172 3156 -138
rect 3156 -172 3164 -138
rect 3700 -172 3708 -138
rect 3708 -172 3734 -138
rect 3772 -172 3776 -138
rect 3776 -172 3806 -138
rect 3844 -172 3878 -138
rect 3916 -172 3946 -138
rect 3946 -172 3950 -138
rect 3988 -172 4014 -138
rect 4014 -172 4022 -138
rect 4558 -172 4566 -138
rect 4566 -172 4592 -138
rect 4630 -172 4634 -138
rect 4634 -172 4664 -138
rect 4702 -172 4736 -138
rect 4774 -172 4804 -138
rect 4804 -172 4808 -138
rect 4846 -172 4872 -138
rect 4872 -172 4880 -138
<< metal1 >>
rect -4923 172 -4515 178
rect -4923 138 -4880 172
rect -4846 138 -4808 172
rect -4774 138 -4736 172
rect -4702 138 -4664 172
rect -4630 138 -4592 172
rect -4558 138 -4515 172
rect -4923 132 -4515 138
rect -4065 172 -3657 178
rect -4065 138 -4022 172
rect -3988 138 -3950 172
rect -3916 138 -3878 172
rect -3844 138 -3806 172
rect -3772 138 -3734 172
rect -3700 138 -3657 172
rect -4065 132 -3657 138
rect -3207 172 -2799 178
rect -3207 138 -3164 172
rect -3130 138 -3092 172
rect -3058 138 -3020 172
rect -2986 138 -2948 172
rect -2914 138 -2876 172
rect -2842 138 -2799 172
rect -3207 132 -2799 138
rect -2349 172 -1941 178
rect -2349 138 -2306 172
rect -2272 138 -2234 172
rect -2200 138 -2162 172
rect -2128 138 -2090 172
rect -2056 138 -2018 172
rect -1984 138 -1941 172
rect -2349 132 -1941 138
rect -1491 172 -1083 178
rect -1491 138 -1448 172
rect -1414 138 -1376 172
rect -1342 138 -1304 172
rect -1270 138 -1232 172
rect -1198 138 -1160 172
rect -1126 138 -1083 172
rect -1491 132 -1083 138
rect -633 172 -225 178
rect -633 138 -590 172
rect -556 138 -518 172
rect -484 138 -446 172
rect -412 138 -374 172
rect -340 138 -302 172
rect -268 138 -225 172
rect -633 132 -225 138
rect 225 172 633 178
rect 225 138 268 172
rect 302 138 340 172
rect 374 138 412 172
rect 446 138 484 172
rect 518 138 556 172
rect 590 138 633 172
rect 225 132 633 138
rect 1083 172 1491 178
rect 1083 138 1126 172
rect 1160 138 1198 172
rect 1232 138 1270 172
rect 1304 138 1342 172
rect 1376 138 1414 172
rect 1448 138 1491 172
rect 1083 132 1491 138
rect 1941 172 2349 178
rect 1941 138 1984 172
rect 2018 138 2056 172
rect 2090 138 2128 172
rect 2162 138 2200 172
rect 2234 138 2272 172
rect 2306 138 2349 172
rect 1941 132 2349 138
rect 2799 172 3207 178
rect 2799 138 2842 172
rect 2876 138 2914 172
rect 2948 138 2986 172
rect 3020 138 3058 172
rect 3092 138 3130 172
rect 3164 138 3207 172
rect 2799 132 3207 138
rect 3657 172 4065 178
rect 3657 138 3700 172
rect 3734 138 3772 172
rect 3806 138 3844 172
rect 3878 138 3916 172
rect 3950 138 3988 172
rect 4022 138 4065 172
rect 3657 132 4065 138
rect 4515 172 4923 178
rect 4515 138 4558 172
rect 4592 138 4630 172
rect 4664 138 4702 172
rect 4736 138 4774 172
rect 4808 138 4846 172
rect 4880 138 4923 172
rect 4515 132 4923 138
rect -5171 53 -5125 100
rect -5171 19 -5165 53
rect -5131 19 -5125 53
rect -5171 -19 -5125 19
rect -5171 -53 -5165 -19
rect -5131 -53 -5125 -19
rect -5171 -100 -5125 -53
rect -4313 53 -4267 100
rect -4313 19 -4307 53
rect -4273 19 -4267 53
rect -4313 -19 -4267 19
rect -4313 -53 -4307 -19
rect -4273 -53 -4267 -19
rect -4313 -100 -4267 -53
rect -3455 53 -3409 100
rect -3455 19 -3449 53
rect -3415 19 -3409 53
rect -3455 -19 -3409 19
rect -3455 -53 -3449 -19
rect -3415 -53 -3409 -19
rect -3455 -100 -3409 -53
rect -2597 53 -2551 100
rect -2597 19 -2591 53
rect -2557 19 -2551 53
rect -2597 -19 -2551 19
rect -2597 -53 -2591 -19
rect -2557 -53 -2551 -19
rect -2597 -100 -2551 -53
rect -1739 53 -1693 100
rect -1739 19 -1733 53
rect -1699 19 -1693 53
rect -1739 -19 -1693 19
rect -1739 -53 -1733 -19
rect -1699 -53 -1693 -19
rect -1739 -100 -1693 -53
rect -881 53 -835 100
rect -881 19 -875 53
rect -841 19 -835 53
rect -881 -19 -835 19
rect -881 -53 -875 -19
rect -841 -53 -835 -19
rect -881 -100 -835 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 835 53 881 100
rect 835 19 841 53
rect 875 19 881 53
rect 835 -19 881 19
rect 835 -53 841 -19
rect 875 -53 881 -19
rect 835 -100 881 -53
rect 1693 53 1739 100
rect 1693 19 1699 53
rect 1733 19 1739 53
rect 1693 -19 1739 19
rect 1693 -53 1699 -19
rect 1733 -53 1739 -19
rect 1693 -100 1739 -53
rect 2551 53 2597 100
rect 2551 19 2557 53
rect 2591 19 2597 53
rect 2551 -19 2597 19
rect 2551 -53 2557 -19
rect 2591 -53 2597 -19
rect 2551 -100 2597 -53
rect 3409 53 3455 100
rect 3409 19 3415 53
rect 3449 19 3455 53
rect 3409 -19 3455 19
rect 3409 -53 3415 -19
rect 3449 -53 3455 -19
rect 3409 -100 3455 -53
rect 4267 53 4313 100
rect 4267 19 4273 53
rect 4307 19 4313 53
rect 4267 -19 4313 19
rect 4267 -53 4273 -19
rect 4307 -53 4313 -19
rect 4267 -100 4313 -53
rect 5125 53 5171 100
rect 5125 19 5131 53
rect 5165 19 5171 53
rect 5125 -19 5171 19
rect 5125 -53 5131 -19
rect 5165 -53 5171 -19
rect 5125 -100 5171 -53
rect -4923 -138 -4515 -132
rect -4923 -172 -4880 -138
rect -4846 -172 -4808 -138
rect -4774 -172 -4736 -138
rect -4702 -172 -4664 -138
rect -4630 -172 -4592 -138
rect -4558 -172 -4515 -138
rect -4923 -178 -4515 -172
rect -4065 -138 -3657 -132
rect -4065 -172 -4022 -138
rect -3988 -172 -3950 -138
rect -3916 -172 -3878 -138
rect -3844 -172 -3806 -138
rect -3772 -172 -3734 -138
rect -3700 -172 -3657 -138
rect -4065 -178 -3657 -172
rect -3207 -138 -2799 -132
rect -3207 -172 -3164 -138
rect -3130 -172 -3092 -138
rect -3058 -172 -3020 -138
rect -2986 -172 -2948 -138
rect -2914 -172 -2876 -138
rect -2842 -172 -2799 -138
rect -3207 -178 -2799 -172
rect -2349 -138 -1941 -132
rect -2349 -172 -2306 -138
rect -2272 -172 -2234 -138
rect -2200 -172 -2162 -138
rect -2128 -172 -2090 -138
rect -2056 -172 -2018 -138
rect -1984 -172 -1941 -138
rect -2349 -178 -1941 -172
rect -1491 -138 -1083 -132
rect -1491 -172 -1448 -138
rect -1414 -172 -1376 -138
rect -1342 -172 -1304 -138
rect -1270 -172 -1232 -138
rect -1198 -172 -1160 -138
rect -1126 -172 -1083 -138
rect -1491 -178 -1083 -172
rect -633 -138 -225 -132
rect -633 -172 -590 -138
rect -556 -172 -518 -138
rect -484 -172 -446 -138
rect -412 -172 -374 -138
rect -340 -172 -302 -138
rect -268 -172 -225 -138
rect -633 -178 -225 -172
rect 225 -138 633 -132
rect 225 -172 268 -138
rect 302 -172 340 -138
rect 374 -172 412 -138
rect 446 -172 484 -138
rect 518 -172 556 -138
rect 590 -172 633 -138
rect 225 -178 633 -172
rect 1083 -138 1491 -132
rect 1083 -172 1126 -138
rect 1160 -172 1198 -138
rect 1232 -172 1270 -138
rect 1304 -172 1342 -138
rect 1376 -172 1414 -138
rect 1448 -172 1491 -138
rect 1083 -178 1491 -172
rect 1941 -138 2349 -132
rect 1941 -172 1984 -138
rect 2018 -172 2056 -138
rect 2090 -172 2128 -138
rect 2162 -172 2200 -138
rect 2234 -172 2272 -138
rect 2306 -172 2349 -138
rect 1941 -178 2349 -172
rect 2799 -138 3207 -132
rect 2799 -172 2842 -138
rect 2876 -172 2914 -138
rect 2948 -172 2986 -138
rect 3020 -172 3058 -138
rect 3092 -172 3130 -138
rect 3164 -172 3207 -138
rect 2799 -178 3207 -172
rect 3657 -138 4065 -132
rect 3657 -172 3700 -138
rect 3734 -172 3772 -138
rect 3806 -172 3844 -138
rect 3878 -172 3916 -138
rect 3950 -172 3988 -138
rect 4022 -172 4065 -138
rect 3657 -178 4065 -172
rect 4515 -138 4923 -132
rect 4515 -172 4558 -138
rect 4592 -172 4630 -138
rect 4664 -172 4702 -138
rect 4736 -172 4774 -138
rect 4808 -172 4846 -138
rect 4880 -172 4923 -138
rect 4515 -178 4923 -172
<< end >>
