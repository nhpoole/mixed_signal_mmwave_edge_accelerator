magic
tech sky130A
magscale 1 2
timestamp 1622084140
<< nwell >>
rect 356 -11 780 310
<< pwell >>
rect 436 -251 622 -69
rect 653 -234 739 -77
rect 436 -255 457 -251
rect 423 -289 457 -255
<< scnmos >>
rect 514 -225 544 -95
<< scpmoshvt >>
rect 514 25 544 225
<< ndiff >>
rect 462 -107 514 -95
rect 462 -141 470 -107
rect 504 -141 514 -107
rect 462 -175 514 -141
rect 462 -209 470 -175
rect 504 -209 514 -175
rect 462 -225 514 -209
rect 544 -107 596 -95
rect 544 -141 554 -107
rect 588 -141 596 -107
rect 544 -175 596 -141
rect 544 -209 554 -175
rect 588 -209 596 -175
rect 544 -225 596 -209
<< pdiff >>
rect 462 213 514 225
rect 462 179 470 213
rect 504 179 514 213
rect 462 145 514 179
rect 462 111 470 145
rect 504 111 514 145
rect 462 77 514 111
rect 462 43 470 77
rect 504 43 514 77
rect 462 25 514 43
rect 544 213 596 225
rect 544 179 554 213
rect 588 179 596 213
rect 544 145 596 179
rect 544 111 554 145
rect 588 111 596 145
rect 544 77 596 111
rect 544 43 554 77
rect 588 43 596 77
rect 544 25 596 43
<< ndiffc >>
rect 470 -141 504 -107
rect 470 -209 504 -175
rect 554 -141 588 -107
rect 554 -209 588 -175
<< pdiffc >>
rect 470 179 504 213
rect 470 111 504 145
rect 470 43 504 77
rect 554 179 588 213
rect 554 111 588 145
rect 554 43 588 77
<< psubdiff >>
rect 679 -127 713 -103
rect 679 -208 713 -161
<< nsubdiff >>
rect 679 184 713 208
rect 679 91 713 150
rect 679 33 713 57
<< psubdiffcont >>
rect 679 -161 713 -127
<< nsubdiffcont >>
rect 679 150 713 184
rect 679 57 713 91
<< poly >>
rect 514 225 544 251
rect 514 -7 544 25
rect 458 -23 544 -7
rect 458 -57 474 -23
rect 508 -57 544 -23
rect 458 -73 544 -57
rect 514 -95 544 -73
rect 514 -251 544 -225
<< polycont >>
rect 474 -57 508 -23
<< locali >>
rect 394 255 423 289
rect 457 255 515 289
rect 549 255 607 289
rect 641 255 679 289
rect 713 255 742 289
rect 462 213 504 255
rect 462 179 470 213
rect 462 145 504 179
rect 462 111 470 145
rect 462 77 504 111
rect 462 43 470 77
rect 462 27 504 43
rect 538 213 604 221
rect 538 179 554 213
rect 588 179 604 213
rect 538 145 604 179
rect 538 111 554 145
rect 588 111 604 145
rect 538 77 604 111
rect 538 43 554 77
rect 588 43 604 77
rect 538 25 604 43
rect 458 -10 524 -9
rect 458 -56 464 -10
rect 512 -56 524 -10
rect 458 -57 474 -56
rect 508 -57 524 -56
rect 558 -10 604 25
rect 667 184 725 255
rect 667 150 679 184
rect 713 150 725 184
rect 667 91 725 150
rect 667 57 679 91
rect 713 57 725 91
rect 667 22 725 57
rect 558 -58 564 -10
rect 458 -107 504 -91
rect 558 -95 604 -58
rect 458 -141 470 -107
rect 458 -175 504 -141
rect 458 -209 470 -175
rect 458 -255 504 -209
rect 538 -107 604 -95
rect 538 -141 554 -107
rect 588 -141 604 -107
rect 538 -175 604 -141
rect 538 -209 554 -175
rect 588 -209 604 -175
rect 538 -221 604 -209
rect 667 -127 725 -110
rect 667 -161 679 -127
rect 713 -161 725 -127
rect 667 -255 725 -161
rect 394 -289 423 -255
rect 457 -289 515 -255
rect 549 -289 607 -255
rect 641 -289 679 -255
rect 713 -289 742 -255
<< viali >>
rect 423 255 457 289
rect 515 255 549 289
rect 607 255 641 289
rect 679 255 713 289
rect 464 -23 512 -10
rect 464 -56 474 -23
rect 474 -56 508 -23
rect 508 -56 512 -23
rect 564 -58 612 -10
rect 423 -289 457 -255
rect 515 -289 549 -255
rect 607 -289 641 -255
rect 679 -289 713 -255
<< metal1 >>
rect 260 289 742 320
rect 260 255 423 289
rect 457 255 515 289
rect 549 255 607 289
rect 641 255 679 289
rect 713 255 742 289
rect 260 224 742 255
rect 304 -10 524 -4
rect 304 -56 464 -10
rect 512 -56 524 -10
rect 304 -64 524 -56
rect 552 -10 718 -4
rect 552 -58 564 -10
rect 612 -58 718 -10
rect 552 -64 718 -58
rect 182 -255 742 -224
rect 182 -289 423 -255
rect 457 -289 515 -255
rect 549 -289 607 -255
rect 641 -289 679 -255
rect 713 -289 742 -255
rect 182 -320 742 -289
<< labels >>
flabel metal1 286 270 290 272 1 FreeSans 480 0 0 0 VDD
port 3 n power bidirectional
flabel metal1 278 -274 284 -270 1 FreeSans 480 0 0 0 VSS
port 4 n ground bidirectional
flabel metal1 332 -38 338 -32 1 FreeSans 480 0 0 0 A
port 1 n
flabel metal1 672 -34 676 -30 1 FreeSans 480 0 0 0 Y
port 2 n
flabel metal1 672 252 725 281 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VPWR
flabel metal1 671 -290 722 -252 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VGND
rlabel comment 650 -272 650 -272 4 sky130_fd_sc_hd__tapvpwrvgnd_1_0/tapvpwrvgnd_1
flabel locali 558 17 592 51 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali 558 -51 592 -17 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali 466 -51 500 -17 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/A
flabel nwell 423 255 457 289 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell 423 -289 457 -255 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 423 -289 457 -255 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 423 255 457 289 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment 394 -272 394 -272 4 sky130_fd_sc_hd__inv_1_0/inv_1
<< end >>
