magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -2228 -1560 2228 1560
<< nwell >>
rect -968 -300 968 300
<< pmos >>
rect -874 -200 -674 200
rect -616 -200 -416 200
rect -358 -200 -158 200
rect -100 -200 100 200
rect 158 -200 358 200
rect 416 -200 616 200
rect 674 -200 874 200
<< pdiff >>
rect -932 187 -874 200
rect -932 153 -920 187
rect -886 153 -874 187
rect -932 119 -874 153
rect -932 85 -920 119
rect -886 85 -874 119
rect -932 51 -874 85
rect -932 17 -920 51
rect -886 17 -874 51
rect -932 -17 -874 17
rect -932 -51 -920 -17
rect -886 -51 -874 -17
rect -932 -85 -874 -51
rect -932 -119 -920 -85
rect -886 -119 -874 -85
rect -932 -153 -874 -119
rect -932 -187 -920 -153
rect -886 -187 -874 -153
rect -932 -200 -874 -187
rect -674 187 -616 200
rect -674 153 -662 187
rect -628 153 -616 187
rect -674 119 -616 153
rect -674 85 -662 119
rect -628 85 -616 119
rect -674 51 -616 85
rect -674 17 -662 51
rect -628 17 -616 51
rect -674 -17 -616 17
rect -674 -51 -662 -17
rect -628 -51 -616 -17
rect -674 -85 -616 -51
rect -674 -119 -662 -85
rect -628 -119 -616 -85
rect -674 -153 -616 -119
rect -674 -187 -662 -153
rect -628 -187 -616 -153
rect -674 -200 -616 -187
rect -416 187 -358 200
rect -416 153 -404 187
rect -370 153 -358 187
rect -416 119 -358 153
rect -416 85 -404 119
rect -370 85 -358 119
rect -416 51 -358 85
rect -416 17 -404 51
rect -370 17 -358 51
rect -416 -17 -358 17
rect -416 -51 -404 -17
rect -370 -51 -358 -17
rect -416 -85 -358 -51
rect -416 -119 -404 -85
rect -370 -119 -358 -85
rect -416 -153 -358 -119
rect -416 -187 -404 -153
rect -370 -187 -358 -153
rect -416 -200 -358 -187
rect -158 187 -100 200
rect -158 153 -146 187
rect -112 153 -100 187
rect -158 119 -100 153
rect -158 85 -146 119
rect -112 85 -100 119
rect -158 51 -100 85
rect -158 17 -146 51
rect -112 17 -100 51
rect -158 -17 -100 17
rect -158 -51 -146 -17
rect -112 -51 -100 -17
rect -158 -85 -100 -51
rect -158 -119 -146 -85
rect -112 -119 -100 -85
rect -158 -153 -100 -119
rect -158 -187 -146 -153
rect -112 -187 -100 -153
rect -158 -200 -100 -187
rect 100 187 158 200
rect 100 153 112 187
rect 146 153 158 187
rect 100 119 158 153
rect 100 85 112 119
rect 146 85 158 119
rect 100 51 158 85
rect 100 17 112 51
rect 146 17 158 51
rect 100 -17 158 17
rect 100 -51 112 -17
rect 146 -51 158 -17
rect 100 -85 158 -51
rect 100 -119 112 -85
rect 146 -119 158 -85
rect 100 -153 158 -119
rect 100 -187 112 -153
rect 146 -187 158 -153
rect 100 -200 158 -187
rect 358 187 416 200
rect 358 153 370 187
rect 404 153 416 187
rect 358 119 416 153
rect 358 85 370 119
rect 404 85 416 119
rect 358 51 416 85
rect 358 17 370 51
rect 404 17 416 51
rect 358 -17 416 17
rect 358 -51 370 -17
rect 404 -51 416 -17
rect 358 -85 416 -51
rect 358 -119 370 -85
rect 404 -119 416 -85
rect 358 -153 416 -119
rect 358 -187 370 -153
rect 404 -187 416 -153
rect 358 -200 416 -187
rect 616 187 674 200
rect 616 153 628 187
rect 662 153 674 187
rect 616 119 674 153
rect 616 85 628 119
rect 662 85 674 119
rect 616 51 674 85
rect 616 17 628 51
rect 662 17 674 51
rect 616 -17 674 17
rect 616 -51 628 -17
rect 662 -51 674 -17
rect 616 -85 674 -51
rect 616 -119 628 -85
rect 662 -119 674 -85
rect 616 -153 674 -119
rect 616 -187 628 -153
rect 662 -187 674 -153
rect 616 -200 674 -187
rect 874 187 932 200
rect 874 153 886 187
rect 920 153 932 187
rect 874 119 932 153
rect 874 85 886 119
rect 920 85 932 119
rect 874 51 932 85
rect 874 17 886 51
rect 920 17 932 51
rect 874 -17 932 17
rect 874 -51 886 -17
rect 920 -51 932 -17
rect 874 -85 932 -51
rect 874 -119 886 -85
rect 920 -119 932 -85
rect 874 -153 932 -119
rect 874 -187 886 -153
rect 920 -187 932 -153
rect 874 -200 932 -187
<< pdiffc >>
rect -920 153 -886 187
rect -920 85 -886 119
rect -920 17 -886 51
rect -920 -51 -886 -17
rect -920 -119 -886 -85
rect -920 -187 -886 -153
rect -662 153 -628 187
rect -662 85 -628 119
rect -662 17 -628 51
rect -662 -51 -628 -17
rect -662 -119 -628 -85
rect -662 -187 -628 -153
rect -404 153 -370 187
rect -404 85 -370 119
rect -404 17 -370 51
rect -404 -51 -370 -17
rect -404 -119 -370 -85
rect -404 -187 -370 -153
rect -146 153 -112 187
rect -146 85 -112 119
rect -146 17 -112 51
rect -146 -51 -112 -17
rect -146 -119 -112 -85
rect -146 -187 -112 -153
rect 112 153 146 187
rect 112 85 146 119
rect 112 17 146 51
rect 112 -51 146 -17
rect 112 -119 146 -85
rect 112 -187 146 -153
rect 370 153 404 187
rect 370 85 404 119
rect 370 17 404 51
rect 370 -51 404 -17
rect 370 -119 404 -85
rect 370 -187 404 -153
rect 628 153 662 187
rect 628 85 662 119
rect 628 17 662 51
rect 628 -51 662 -17
rect 628 -119 662 -85
rect 628 -187 662 -153
rect 886 153 920 187
rect 886 85 920 119
rect 886 17 920 51
rect 886 -51 920 -17
rect 886 -119 920 -85
rect 886 -187 920 -153
<< poly >>
rect -840 281 -708 297
rect -840 264 -791 281
rect -874 247 -791 264
rect -757 264 -708 281
rect -582 281 -450 297
rect -582 264 -533 281
rect -757 247 -674 264
rect -874 200 -674 247
rect -616 247 -533 264
rect -499 264 -450 281
rect -324 281 -192 297
rect -324 264 -275 281
rect -499 247 -416 264
rect -616 200 -416 247
rect -358 247 -275 264
rect -241 264 -192 281
rect -66 281 66 297
rect -66 264 -17 281
rect -241 247 -158 264
rect -358 200 -158 247
rect -100 247 -17 264
rect 17 264 66 281
rect 192 281 324 297
rect 192 264 241 281
rect 17 247 100 264
rect -100 200 100 247
rect 158 247 241 264
rect 275 264 324 281
rect 450 281 582 297
rect 450 264 499 281
rect 275 247 358 264
rect 158 200 358 247
rect 416 247 499 264
rect 533 264 582 281
rect 708 281 840 297
rect 708 264 757 281
rect 533 247 616 264
rect 416 200 616 247
rect 674 247 757 264
rect 791 264 840 281
rect 791 247 874 264
rect 674 200 874 247
rect -874 -247 -674 -200
rect -874 -264 -791 -247
rect -840 -281 -791 -264
rect -757 -264 -674 -247
rect -616 -247 -416 -200
rect -616 -264 -533 -247
rect -757 -281 -708 -264
rect -840 -297 -708 -281
rect -582 -281 -533 -264
rect -499 -264 -416 -247
rect -358 -247 -158 -200
rect -358 -264 -275 -247
rect -499 -281 -450 -264
rect -582 -297 -450 -281
rect -324 -281 -275 -264
rect -241 -264 -158 -247
rect -100 -247 100 -200
rect -100 -264 -17 -247
rect -241 -281 -192 -264
rect -324 -297 -192 -281
rect -66 -281 -17 -264
rect 17 -264 100 -247
rect 158 -247 358 -200
rect 158 -264 241 -247
rect 17 -281 66 -264
rect -66 -297 66 -281
rect 192 -281 241 -264
rect 275 -264 358 -247
rect 416 -247 616 -200
rect 416 -264 499 -247
rect 275 -281 324 -264
rect 192 -297 324 -281
rect 450 -281 499 -264
rect 533 -264 616 -247
rect 674 -247 874 -200
rect 674 -264 757 -247
rect 533 -281 582 -264
rect 450 -297 582 -281
rect 708 -281 757 -264
rect 791 -264 874 -247
rect 791 -281 840 -264
rect 708 -297 840 -281
<< polycont >>
rect -791 247 -757 281
rect -533 247 -499 281
rect -275 247 -241 281
rect -17 247 17 281
rect 241 247 275 281
rect 499 247 533 281
rect 757 247 791 281
rect -791 -281 -757 -247
rect -533 -281 -499 -247
rect -275 -281 -241 -247
rect -17 -281 17 -247
rect 241 -281 275 -247
rect 499 -281 533 -247
rect 757 -281 791 -247
<< locali >>
rect -840 247 -791 281
rect -757 247 -708 281
rect -582 247 -533 281
rect -499 247 -450 281
rect -324 247 -275 281
rect -241 247 -192 281
rect -66 247 -17 281
rect 17 247 66 281
rect 192 247 241 281
rect 275 247 324 281
rect 450 247 499 281
rect 533 247 582 281
rect 708 247 757 281
rect 791 247 840 281
rect -920 187 -886 204
rect -920 119 -886 127
rect -920 51 -886 55
rect -920 -55 -886 -51
rect -920 -127 -886 -119
rect -920 -204 -886 -187
rect -662 187 -628 204
rect -662 119 -628 127
rect -662 51 -628 55
rect -662 -55 -628 -51
rect -662 -127 -628 -119
rect -662 -204 -628 -187
rect -404 187 -370 204
rect -404 119 -370 127
rect -404 51 -370 55
rect -404 -55 -370 -51
rect -404 -127 -370 -119
rect -404 -204 -370 -187
rect -146 187 -112 204
rect -146 119 -112 127
rect -146 51 -112 55
rect -146 -55 -112 -51
rect -146 -127 -112 -119
rect -146 -204 -112 -187
rect 112 187 146 204
rect 112 119 146 127
rect 112 51 146 55
rect 112 -55 146 -51
rect 112 -127 146 -119
rect 112 -204 146 -187
rect 370 187 404 204
rect 370 119 404 127
rect 370 51 404 55
rect 370 -55 404 -51
rect 370 -127 404 -119
rect 370 -204 404 -187
rect 628 187 662 204
rect 628 119 662 127
rect 628 51 662 55
rect 628 -55 662 -51
rect 628 -127 662 -119
rect 628 -204 662 -187
rect 886 187 920 204
rect 886 119 920 127
rect 886 51 920 55
rect 886 -55 920 -51
rect 886 -127 920 -119
rect 886 -204 920 -187
rect -840 -281 -791 -247
rect -757 -281 -708 -247
rect -582 -281 -533 -247
rect -499 -281 -450 -247
rect -324 -281 -275 -247
rect -241 -281 -192 -247
rect -66 -281 -17 -247
rect 17 -281 66 -247
rect 192 -281 241 -247
rect 275 -281 324 -247
rect 450 -281 499 -247
rect 533 -281 582 -247
rect 708 -281 757 -247
rect 791 -281 840 -247
<< viali >>
rect -791 247 -757 281
rect -533 247 -499 281
rect -275 247 -241 281
rect -17 247 17 281
rect 241 247 275 281
rect 499 247 533 281
rect 757 247 791 281
rect -920 153 -886 161
rect -920 127 -886 153
rect -920 85 -886 89
rect -920 55 -886 85
rect -920 -17 -886 17
rect -920 -85 -886 -55
rect -920 -89 -886 -85
rect -920 -153 -886 -127
rect -920 -161 -886 -153
rect -662 153 -628 161
rect -662 127 -628 153
rect -662 85 -628 89
rect -662 55 -628 85
rect -662 -17 -628 17
rect -662 -85 -628 -55
rect -662 -89 -628 -85
rect -662 -153 -628 -127
rect -662 -161 -628 -153
rect -404 153 -370 161
rect -404 127 -370 153
rect -404 85 -370 89
rect -404 55 -370 85
rect -404 -17 -370 17
rect -404 -85 -370 -55
rect -404 -89 -370 -85
rect -404 -153 -370 -127
rect -404 -161 -370 -153
rect -146 153 -112 161
rect -146 127 -112 153
rect -146 85 -112 89
rect -146 55 -112 85
rect -146 -17 -112 17
rect -146 -85 -112 -55
rect -146 -89 -112 -85
rect -146 -153 -112 -127
rect -146 -161 -112 -153
rect 112 153 146 161
rect 112 127 146 153
rect 112 85 146 89
rect 112 55 146 85
rect 112 -17 146 17
rect 112 -85 146 -55
rect 112 -89 146 -85
rect 112 -153 146 -127
rect 112 -161 146 -153
rect 370 153 404 161
rect 370 127 404 153
rect 370 85 404 89
rect 370 55 404 85
rect 370 -17 404 17
rect 370 -85 404 -55
rect 370 -89 404 -85
rect 370 -153 404 -127
rect 370 -161 404 -153
rect 628 153 662 161
rect 628 127 662 153
rect 628 85 662 89
rect 628 55 662 85
rect 628 -17 662 17
rect 628 -85 662 -55
rect 628 -89 662 -85
rect 628 -153 662 -127
rect 628 -161 662 -153
rect 886 153 920 161
rect 886 127 920 153
rect 886 85 920 89
rect 886 55 920 85
rect 886 -17 920 17
rect 886 -85 920 -55
rect 886 -89 920 -85
rect 886 -153 920 -127
rect 886 -161 920 -153
rect -791 -281 -757 -247
rect -533 -281 -499 -247
rect -275 -281 -241 -247
rect -17 -281 17 -247
rect 241 -281 275 -247
rect 499 -281 533 -247
rect 757 -281 791 -247
<< metal1 >>
rect -828 281 -720 287
rect -828 247 -791 281
rect -757 247 -720 281
rect -828 241 -720 247
rect -570 281 -462 287
rect -570 247 -533 281
rect -499 247 -462 281
rect -570 241 -462 247
rect -312 281 -204 287
rect -312 247 -275 281
rect -241 247 -204 281
rect -312 241 -204 247
rect -54 281 54 287
rect -54 247 -17 281
rect 17 247 54 281
rect -54 241 54 247
rect 204 281 312 287
rect 204 247 241 281
rect 275 247 312 281
rect 204 241 312 247
rect 462 281 570 287
rect 462 247 499 281
rect 533 247 570 281
rect 462 241 570 247
rect 720 281 828 287
rect 720 247 757 281
rect 791 247 828 281
rect 720 241 828 247
rect -926 161 -880 200
rect -926 127 -920 161
rect -886 127 -880 161
rect -926 89 -880 127
rect -926 55 -920 89
rect -886 55 -880 89
rect -926 17 -880 55
rect -926 -17 -920 17
rect -886 -17 -880 17
rect -926 -55 -880 -17
rect -926 -89 -920 -55
rect -886 -89 -880 -55
rect -926 -127 -880 -89
rect -926 -161 -920 -127
rect -886 -161 -880 -127
rect -926 -200 -880 -161
rect -668 161 -622 200
rect -668 127 -662 161
rect -628 127 -622 161
rect -668 89 -622 127
rect -668 55 -662 89
rect -628 55 -622 89
rect -668 17 -622 55
rect -668 -17 -662 17
rect -628 -17 -622 17
rect -668 -55 -622 -17
rect -668 -89 -662 -55
rect -628 -89 -622 -55
rect -668 -127 -622 -89
rect -668 -161 -662 -127
rect -628 -161 -622 -127
rect -668 -200 -622 -161
rect -410 161 -364 200
rect -410 127 -404 161
rect -370 127 -364 161
rect -410 89 -364 127
rect -410 55 -404 89
rect -370 55 -364 89
rect -410 17 -364 55
rect -410 -17 -404 17
rect -370 -17 -364 17
rect -410 -55 -364 -17
rect -410 -89 -404 -55
rect -370 -89 -364 -55
rect -410 -127 -364 -89
rect -410 -161 -404 -127
rect -370 -161 -364 -127
rect -410 -200 -364 -161
rect -152 161 -106 200
rect -152 127 -146 161
rect -112 127 -106 161
rect -152 89 -106 127
rect -152 55 -146 89
rect -112 55 -106 89
rect -152 17 -106 55
rect -152 -17 -146 17
rect -112 -17 -106 17
rect -152 -55 -106 -17
rect -152 -89 -146 -55
rect -112 -89 -106 -55
rect -152 -127 -106 -89
rect -152 -161 -146 -127
rect -112 -161 -106 -127
rect -152 -200 -106 -161
rect 106 161 152 200
rect 106 127 112 161
rect 146 127 152 161
rect 106 89 152 127
rect 106 55 112 89
rect 146 55 152 89
rect 106 17 152 55
rect 106 -17 112 17
rect 146 -17 152 17
rect 106 -55 152 -17
rect 106 -89 112 -55
rect 146 -89 152 -55
rect 106 -127 152 -89
rect 106 -161 112 -127
rect 146 -161 152 -127
rect 106 -200 152 -161
rect 364 161 410 200
rect 364 127 370 161
rect 404 127 410 161
rect 364 89 410 127
rect 364 55 370 89
rect 404 55 410 89
rect 364 17 410 55
rect 364 -17 370 17
rect 404 -17 410 17
rect 364 -55 410 -17
rect 364 -89 370 -55
rect 404 -89 410 -55
rect 364 -127 410 -89
rect 364 -161 370 -127
rect 404 -161 410 -127
rect 364 -200 410 -161
rect 622 161 668 200
rect 622 127 628 161
rect 662 127 668 161
rect 622 89 668 127
rect 622 55 628 89
rect 662 55 668 89
rect 622 17 668 55
rect 622 -17 628 17
rect 662 -17 668 17
rect 622 -55 668 -17
rect 622 -89 628 -55
rect 662 -89 668 -55
rect 622 -127 668 -89
rect 622 -161 628 -127
rect 662 -161 668 -127
rect 622 -200 668 -161
rect 880 161 926 200
rect 880 127 886 161
rect 920 127 926 161
rect 880 89 926 127
rect 880 55 886 89
rect 920 55 926 89
rect 880 17 926 55
rect 880 -17 886 17
rect 920 -17 926 17
rect 880 -55 926 -17
rect 880 -89 886 -55
rect 920 -89 926 -55
rect 880 -127 926 -89
rect 880 -161 886 -127
rect 920 -161 926 -127
rect 880 -200 926 -161
rect -828 -247 -720 -241
rect -828 -281 -791 -247
rect -757 -281 -720 -247
rect -828 -287 -720 -281
rect -570 -247 -462 -241
rect -570 -281 -533 -247
rect -499 -281 -462 -247
rect -570 -287 -462 -281
rect -312 -247 -204 -241
rect -312 -281 -275 -247
rect -241 -281 -204 -247
rect -312 -287 -204 -281
rect -54 -247 54 -241
rect -54 -281 -17 -247
rect 17 -281 54 -247
rect -54 -287 54 -281
rect 204 -247 312 -241
rect 204 -281 241 -247
rect 275 -281 312 -247
rect 204 -287 312 -281
rect 462 -247 570 -241
rect 462 -281 499 -247
rect 533 -281 570 -247
rect 462 -287 570 -281
rect 720 -247 828 -241
rect 720 -281 757 -247
rect 791 -281 828 -247
rect 720 -287 828 -281
<< end >>
