magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -11495 -2057 11495 2057
<< pwell >>
rect -10235 -735 10235 735
<< nmos >>
rect -10151 109 -9191 709
rect -9133 109 -8173 709
rect -8115 109 -7155 709
rect -7097 109 -6137 709
rect -6079 109 -5119 709
rect -5061 109 -4101 709
rect -4043 109 -3083 709
rect -3025 109 -2065 709
rect -2007 109 -1047 709
rect -989 109 -29 709
rect 29 109 989 709
rect 1047 109 2007 709
rect 2065 109 3025 709
rect 3083 109 4043 709
rect 4101 109 5061 709
rect 5119 109 6079 709
rect 6137 109 7097 709
rect 7155 109 8115 709
rect 8173 109 9133 709
rect 9191 109 10151 709
rect -10151 -709 -9191 -109
rect -9133 -709 -8173 -109
rect -8115 -709 -7155 -109
rect -7097 -709 -6137 -109
rect -6079 -709 -5119 -109
rect -5061 -709 -4101 -109
rect -4043 -709 -3083 -109
rect -3025 -709 -2065 -109
rect -2007 -709 -1047 -109
rect -989 -709 -29 -109
rect 29 -709 989 -109
rect 1047 -709 2007 -109
rect 2065 -709 3025 -109
rect 3083 -709 4043 -109
rect 4101 -709 5061 -109
rect 5119 -709 6079 -109
rect 6137 -709 7097 -109
rect 7155 -709 8115 -109
rect 8173 -709 9133 -109
rect 9191 -709 10151 -109
<< ndiff >>
rect -10209 664 -10151 709
rect -10209 630 -10197 664
rect -10163 630 -10151 664
rect -10209 596 -10151 630
rect -10209 562 -10197 596
rect -10163 562 -10151 596
rect -10209 528 -10151 562
rect -10209 494 -10197 528
rect -10163 494 -10151 528
rect -10209 460 -10151 494
rect -10209 426 -10197 460
rect -10163 426 -10151 460
rect -10209 392 -10151 426
rect -10209 358 -10197 392
rect -10163 358 -10151 392
rect -10209 324 -10151 358
rect -10209 290 -10197 324
rect -10163 290 -10151 324
rect -10209 256 -10151 290
rect -10209 222 -10197 256
rect -10163 222 -10151 256
rect -10209 188 -10151 222
rect -10209 154 -10197 188
rect -10163 154 -10151 188
rect -10209 109 -10151 154
rect -9191 664 -9133 709
rect -9191 630 -9179 664
rect -9145 630 -9133 664
rect -9191 596 -9133 630
rect -9191 562 -9179 596
rect -9145 562 -9133 596
rect -9191 528 -9133 562
rect -9191 494 -9179 528
rect -9145 494 -9133 528
rect -9191 460 -9133 494
rect -9191 426 -9179 460
rect -9145 426 -9133 460
rect -9191 392 -9133 426
rect -9191 358 -9179 392
rect -9145 358 -9133 392
rect -9191 324 -9133 358
rect -9191 290 -9179 324
rect -9145 290 -9133 324
rect -9191 256 -9133 290
rect -9191 222 -9179 256
rect -9145 222 -9133 256
rect -9191 188 -9133 222
rect -9191 154 -9179 188
rect -9145 154 -9133 188
rect -9191 109 -9133 154
rect -8173 664 -8115 709
rect -8173 630 -8161 664
rect -8127 630 -8115 664
rect -8173 596 -8115 630
rect -8173 562 -8161 596
rect -8127 562 -8115 596
rect -8173 528 -8115 562
rect -8173 494 -8161 528
rect -8127 494 -8115 528
rect -8173 460 -8115 494
rect -8173 426 -8161 460
rect -8127 426 -8115 460
rect -8173 392 -8115 426
rect -8173 358 -8161 392
rect -8127 358 -8115 392
rect -8173 324 -8115 358
rect -8173 290 -8161 324
rect -8127 290 -8115 324
rect -8173 256 -8115 290
rect -8173 222 -8161 256
rect -8127 222 -8115 256
rect -8173 188 -8115 222
rect -8173 154 -8161 188
rect -8127 154 -8115 188
rect -8173 109 -8115 154
rect -7155 664 -7097 709
rect -7155 630 -7143 664
rect -7109 630 -7097 664
rect -7155 596 -7097 630
rect -7155 562 -7143 596
rect -7109 562 -7097 596
rect -7155 528 -7097 562
rect -7155 494 -7143 528
rect -7109 494 -7097 528
rect -7155 460 -7097 494
rect -7155 426 -7143 460
rect -7109 426 -7097 460
rect -7155 392 -7097 426
rect -7155 358 -7143 392
rect -7109 358 -7097 392
rect -7155 324 -7097 358
rect -7155 290 -7143 324
rect -7109 290 -7097 324
rect -7155 256 -7097 290
rect -7155 222 -7143 256
rect -7109 222 -7097 256
rect -7155 188 -7097 222
rect -7155 154 -7143 188
rect -7109 154 -7097 188
rect -7155 109 -7097 154
rect -6137 664 -6079 709
rect -6137 630 -6125 664
rect -6091 630 -6079 664
rect -6137 596 -6079 630
rect -6137 562 -6125 596
rect -6091 562 -6079 596
rect -6137 528 -6079 562
rect -6137 494 -6125 528
rect -6091 494 -6079 528
rect -6137 460 -6079 494
rect -6137 426 -6125 460
rect -6091 426 -6079 460
rect -6137 392 -6079 426
rect -6137 358 -6125 392
rect -6091 358 -6079 392
rect -6137 324 -6079 358
rect -6137 290 -6125 324
rect -6091 290 -6079 324
rect -6137 256 -6079 290
rect -6137 222 -6125 256
rect -6091 222 -6079 256
rect -6137 188 -6079 222
rect -6137 154 -6125 188
rect -6091 154 -6079 188
rect -6137 109 -6079 154
rect -5119 664 -5061 709
rect -5119 630 -5107 664
rect -5073 630 -5061 664
rect -5119 596 -5061 630
rect -5119 562 -5107 596
rect -5073 562 -5061 596
rect -5119 528 -5061 562
rect -5119 494 -5107 528
rect -5073 494 -5061 528
rect -5119 460 -5061 494
rect -5119 426 -5107 460
rect -5073 426 -5061 460
rect -5119 392 -5061 426
rect -5119 358 -5107 392
rect -5073 358 -5061 392
rect -5119 324 -5061 358
rect -5119 290 -5107 324
rect -5073 290 -5061 324
rect -5119 256 -5061 290
rect -5119 222 -5107 256
rect -5073 222 -5061 256
rect -5119 188 -5061 222
rect -5119 154 -5107 188
rect -5073 154 -5061 188
rect -5119 109 -5061 154
rect -4101 664 -4043 709
rect -4101 630 -4089 664
rect -4055 630 -4043 664
rect -4101 596 -4043 630
rect -4101 562 -4089 596
rect -4055 562 -4043 596
rect -4101 528 -4043 562
rect -4101 494 -4089 528
rect -4055 494 -4043 528
rect -4101 460 -4043 494
rect -4101 426 -4089 460
rect -4055 426 -4043 460
rect -4101 392 -4043 426
rect -4101 358 -4089 392
rect -4055 358 -4043 392
rect -4101 324 -4043 358
rect -4101 290 -4089 324
rect -4055 290 -4043 324
rect -4101 256 -4043 290
rect -4101 222 -4089 256
rect -4055 222 -4043 256
rect -4101 188 -4043 222
rect -4101 154 -4089 188
rect -4055 154 -4043 188
rect -4101 109 -4043 154
rect -3083 664 -3025 709
rect -3083 630 -3071 664
rect -3037 630 -3025 664
rect -3083 596 -3025 630
rect -3083 562 -3071 596
rect -3037 562 -3025 596
rect -3083 528 -3025 562
rect -3083 494 -3071 528
rect -3037 494 -3025 528
rect -3083 460 -3025 494
rect -3083 426 -3071 460
rect -3037 426 -3025 460
rect -3083 392 -3025 426
rect -3083 358 -3071 392
rect -3037 358 -3025 392
rect -3083 324 -3025 358
rect -3083 290 -3071 324
rect -3037 290 -3025 324
rect -3083 256 -3025 290
rect -3083 222 -3071 256
rect -3037 222 -3025 256
rect -3083 188 -3025 222
rect -3083 154 -3071 188
rect -3037 154 -3025 188
rect -3083 109 -3025 154
rect -2065 664 -2007 709
rect -2065 630 -2053 664
rect -2019 630 -2007 664
rect -2065 596 -2007 630
rect -2065 562 -2053 596
rect -2019 562 -2007 596
rect -2065 528 -2007 562
rect -2065 494 -2053 528
rect -2019 494 -2007 528
rect -2065 460 -2007 494
rect -2065 426 -2053 460
rect -2019 426 -2007 460
rect -2065 392 -2007 426
rect -2065 358 -2053 392
rect -2019 358 -2007 392
rect -2065 324 -2007 358
rect -2065 290 -2053 324
rect -2019 290 -2007 324
rect -2065 256 -2007 290
rect -2065 222 -2053 256
rect -2019 222 -2007 256
rect -2065 188 -2007 222
rect -2065 154 -2053 188
rect -2019 154 -2007 188
rect -2065 109 -2007 154
rect -1047 664 -989 709
rect -1047 630 -1035 664
rect -1001 630 -989 664
rect -1047 596 -989 630
rect -1047 562 -1035 596
rect -1001 562 -989 596
rect -1047 528 -989 562
rect -1047 494 -1035 528
rect -1001 494 -989 528
rect -1047 460 -989 494
rect -1047 426 -1035 460
rect -1001 426 -989 460
rect -1047 392 -989 426
rect -1047 358 -1035 392
rect -1001 358 -989 392
rect -1047 324 -989 358
rect -1047 290 -1035 324
rect -1001 290 -989 324
rect -1047 256 -989 290
rect -1047 222 -1035 256
rect -1001 222 -989 256
rect -1047 188 -989 222
rect -1047 154 -1035 188
rect -1001 154 -989 188
rect -1047 109 -989 154
rect -29 664 29 709
rect -29 630 -17 664
rect 17 630 29 664
rect -29 596 29 630
rect -29 562 -17 596
rect 17 562 29 596
rect -29 528 29 562
rect -29 494 -17 528
rect 17 494 29 528
rect -29 460 29 494
rect -29 426 -17 460
rect 17 426 29 460
rect -29 392 29 426
rect -29 358 -17 392
rect 17 358 29 392
rect -29 324 29 358
rect -29 290 -17 324
rect 17 290 29 324
rect -29 256 29 290
rect -29 222 -17 256
rect 17 222 29 256
rect -29 188 29 222
rect -29 154 -17 188
rect 17 154 29 188
rect -29 109 29 154
rect 989 664 1047 709
rect 989 630 1001 664
rect 1035 630 1047 664
rect 989 596 1047 630
rect 989 562 1001 596
rect 1035 562 1047 596
rect 989 528 1047 562
rect 989 494 1001 528
rect 1035 494 1047 528
rect 989 460 1047 494
rect 989 426 1001 460
rect 1035 426 1047 460
rect 989 392 1047 426
rect 989 358 1001 392
rect 1035 358 1047 392
rect 989 324 1047 358
rect 989 290 1001 324
rect 1035 290 1047 324
rect 989 256 1047 290
rect 989 222 1001 256
rect 1035 222 1047 256
rect 989 188 1047 222
rect 989 154 1001 188
rect 1035 154 1047 188
rect 989 109 1047 154
rect 2007 664 2065 709
rect 2007 630 2019 664
rect 2053 630 2065 664
rect 2007 596 2065 630
rect 2007 562 2019 596
rect 2053 562 2065 596
rect 2007 528 2065 562
rect 2007 494 2019 528
rect 2053 494 2065 528
rect 2007 460 2065 494
rect 2007 426 2019 460
rect 2053 426 2065 460
rect 2007 392 2065 426
rect 2007 358 2019 392
rect 2053 358 2065 392
rect 2007 324 2065 358
rect 2007 290 2019 324
rect 2053 290 2065 324
rect 2007 256 2065 290
rect 2007 222 2019 256
rect 2053 222 2065 256
rect 2007 188 2065 222
rect 2007 154 2019 188
rect 2053 154 2065 188
rect 2007 109 2065 154
rect 3025 664 3083 709
rect 3025 630 3037 664
rect 3071 630 3083 664
rect 3025 596 3083 630
rect 3025 562 3037 596
rect 3071 562 3083 596
rect 3025 528 3083 562
rect 3025 494 3037 528
rect 3071 494 3083 528
rect 3025 460 3083 494
rect 3025 426 3037 460
rect 3071 426 3083 460
rect 3025 392 3083 426
rect 3025 358 3037 392
rect 3071 358 3083 392
rect 3025 324 3083 358
rect 3025 290 3037 324
rect 3071 290 3083 324
rect 3025 256 3083 290
rect 3025 222 3037 256
rect 3071 222 3083 256
rect 3025 188 3083 222
rect 3025 154 3037 188
rect 3071 154 3083 188
rect 3025 109 3083 154
rect 4043 664 4101 709
rect 4043 630 4055 664
rect 4089 630 4101 664
rect 4043 596 4101 630
rect 4043 562 4055 596
rect 4089 562 4101 596
rect 4043 528 4101 562
rect 4043 494 4055 528
rect 4089 494 4101 528
rect 4043 460 4101 494
rect 4043 426 4055 460
rect 4089 426 4101 460
rect 4043 392 4101 426
rect 4043 358 4055 392
rect 4089 358 4101 392
rect 4043 324 4101 358
rect 4043 290 4055 324
rect 4089 290 4101 324
rect 4043 256 4101 290
rect 4043 222 4055 256
rect 4089 222 4101 256
rect 4043 188 4101 222
rect 4043 154 4055 188
rect 4089 154 4101 188
rect 4043 109 4101 154
rect 5061 664 5119 709
rect 5061 630 5073 664
rect 5107 630 5119 664
rect 5061 596 5119 630
rect 5061 562 5073 596
rect 5107 562 5119 596
rect 5061 528 5119 562
rect 5061 494 5073 528
rect 5107 494 5119 528
rect 5061 460 5119 494
rect 5061 426 5073 460
rect 5107 426 5119 460
rect 5061 392 5119 426
rect 5061 358 5073 392
rect 5107 358 5119 392
rect 5061 324 5119 358
rect 5061 290 5073 324
rect 5107 290 5119 324
rect 5061 256 5119 290
rect 5061 222 5073 256
rect 5107 222 5119 256
rect 5061 188 5119 222
rect 5061 154 5073 188
rect 5107 154 5119 188
rect 5061 109 5119 154
rect 6079 664 6137 709
rect 6079 630 6091 664
rect 6125 630 6137 664
rect 6079 596 6137 630
rect 6079 562 6091 596
rect 6125 562 6137 596
rect 6079 528 6137 562
rect 6079 494 6091 528
rect 6125 494 6137 528
rect 6079 460 6137 494
rect 6079 426 6091 460
rect 6125 426 6137 460
rect 6079 392 6137 426
rect 6079 358 6091 392
rect 6125 358 6137 392
rect 6079 324 6137 358
rect 6079 290 6091 324
rect 6125 290 6137 324
rect 6079 256 6137 290
rect 6079 222 6091 256
rect 6125 222 6137 256
rect 6079 188 6137 222
rect 6079 154 6091 188
rect 6125 154 6137 188
rect 6079 109 6137 154
rect 7097 664 7155 709
rect 7097 630 7109 664
rect 7143 630 7155 664
rect 7097 596 7155 630
rect 7097 562 7109 596
rect 7143 562 7155 596
rect 7097 528 7155 562
rect 7097 494 7109 528
rect 7143 494 7155 528
rect 7097 460 7155 494
rect 7097 426 7109 460
rect 7143 426 7155 460
rect 7097 392 7155 426
rect 7097 358 7109 392
rect 7143 358 7155 392
rect 7097 324 7155 358
rect 7097 290 7109 324
rect 7143 290 7155 324
rect 7097 256 7155 290
rect 7097 222 7109 256
rect 7143 222 7155 256
rect 7097 188 7155 222
rect 7097 154 7109 188
rect 7143 154 7155 188
rect 7097 109 7155 154
rect 8115 664 8173 709
rect 8115 630 8127 664
rect 8161 630 8173 664
rect 8115 596 8173 630
rect 8115 562 8127 596
rect 8161 562 8173 596
rect 8115 528 8173 562
rect 8115 494 8127 528
rect 8161 494 8173 528
rect 8115 460 8173 494
rect 8115 426 8127 460
rect 8161 426 8173 460
rect 8115 392 8173 426
rect 8115 358 8127 392
rect 8161 358 8173 392
rect 8115 324 8173 358
rect 8115 290 8127 324
rect 8161 290 8173 324
rect 8115 256 8173 290
rect 8115 222 8127 256
rect 8161 222 8173 256
rect 8115 188 8173 222
rect 8115 154 8127 188
rect 8161 154 8173 188
rect 8115 109 8173 154
rect 9133 664 9191 709
rect 9133 630 9145 664
rect 9179 630 9191 664
rect 9133 596 9191 630
rect 9133 562 9145 596
rect 9179 562 9191 596
rect 9133 528 9191 562
rect 9133 494 9145 528
rect 9179 494 9191 528
rect 9133 460 9191 494
rect 9133 426 9145 460
rect 9179 426 9191 460
rect 9133 392 9191 426
rect 9133 358 9145 392
rect 9179 358 9191 392
rect 9133 324 9191 358
rect 9133 290 9145 324
rect 9179 290 9191 324
rect 9133 256 9191 290
rect 9133 222 9145 256
rect 9179 222 9191 256
rect 9133 188 9191 222
rect 9133 154 9145 188
rect 9179 154 9191 188
rect 9133 109 9191 154
rect 10151 664 10209 709
rect 10151 630 10163 664
rect 10197 630 10209 664
rect 10151 596 10209 630
rect 10151 562 10163 596
rect 10197 562 10209 596
rect 10151 528 10209 562
rect 10151 494 10163 528
rect 10197 494 10209 528
rect 10151 460 10209 494
rect 10151 426 10163 460
rect 10197 426 10209 460
rect 10151 392 10209 426
rect 10151 358 10163 392
rect 10197 358 10209 392
rect 10151 324 10209 358
rect 10151 290 10163 324
rect 10197 290 10209 324
rect 10151 256 10209 290
rect 10151 222 10163 256
rect 10197 222 10209 256
rect 10151 188 10209 222
rect 10151 154 10163 188
rect 10197 154 10209 188
rect 10151 109 10209 154
rect -10209 -154 -10151 -109
rect -10209 -188 -10197 -154
rect -10163 -188 -10151 -154
rect -10209 -222 -10151 -188
rect -10209 -256 -10197 -222
rect -10163 -256 -10151 -222
rect -10209 -290 -10151 -256
rect -10209 -324 -10197 -290
rect -10163 -324 -10151 -290
rect -10209 -358 -10151 -324
rect -10209 -392 -10197 -358
rect -10163 -392 -10151 -358
rect -10209 -426 -10151 -392
rect -10209 -460 -10197 -426
rect -10163 -460 -10151 -426
rect -10209 -494 -10151 -460
rect -10209 -528 -10197 -494
rect -10163 -528 -10151 -494
rect -10209 -562 -10151 -528
rect -10209 -596 -10197 -562
rect -10163 -596 -10151 -562
rect -10209 -630 -10151 -596
rect -10209 -664 -10197 -630
rect -10163 -664 -10151 -630
rect -10209 -709 -10151 -664
rect -9191 -154 -9133 -109
rect -9191 -188 -9179 -154
rect -9145 -188 -9133 -154
rect -9191 -222 -9133 -188
rect -9191 -256 -9179 -222
rect -9145 -256 -9133 -222
rect -9191 -290 -9133 -256
rect -9191 -324 -9179 -290
rect -9145 -324 -9133 -290
rect -9191 -358 -9133 -324
rect -9191 -392 -9179 -358
rect -9145 -392 -9133 -358
rect -9191 -426 -9133 -392
rect -9191 -460 -9179 -426
rect -9145 -460 -9133 -426
rect -9191 -494 -9133 -460
rect -9191 -528 -9179 -494
rect -9145 -528 -9133 -494
rect -9191 -562 -9133 -528
rect -9191 -596 -9179 -562
rect -9145 -596 -9133 -562
rect -9191 -630 -9133 -596
rect -9191 -664 -9179 -630
rect -9145 -664 -9133 -630
rect -9191 -709 -9133 -664
rect -8173 -154 -8115 -109
rect -8173 -188 -8161 -154
rect -8127 -188 -8115 -154
rect -8173 -222 -8115 -188
rect -8173 -256 -8161 -222
rect -8127 -256 -8115 -222
rect -8173 -290 -8115 -256
rect -8173 -324 -8161 -290
rect -8127 -324 -8115 -290
rect -8173 -358 -8115 -324
rect -8173 -392 -8161 -358
rect -8127 -392 -8115 -358
rect -8173 -426 -8115 -392
rect -8173 -460 -8161 -426
rect -8127 -460 -8115 -426
rect -8173 -494 -8115 -460
rect -8173 -528 -8161 -494
rect -8127 -528 -8115 -494
rect -8173 -562 -8115 -528
rect -8173 -596 -8161 -562
rect -8127 -596 -8115 -562
rect -8173 -630 -8115 -596
rect -8173 -664 -8161 -630
rect -8127 -664 -8115 -630
rect -8173 -709 -8115 -664
rect -7155 -154 -7097 -109
rect -7155 -188 -7143 -154
rect -7109 -188 -7097 -154
rect -7155 -222 -7097 -188
rect -7155 -256 -7143 -222
rect -7109 -256 -7097 -222
rect -7155 -290 -7097 -256
rect -7155 -324 -7143 -290
rect -7109 -324 -7097 -290
rect -7155 -358 -7097 -324
rect -7155 -392 -7143 -358
rect -7109 -392 -7097 -358
rect -7155 -426 -7097 -392
rect -7155 -460 -7143 -426
rect -7109 -460 -7097 -426
rect -7155 -494 -7097 -460
rect -7155 -528 -7143 -494
rect -7109 -528 -7097 -494
rect -7155 -562 -7097 -528
rect -7155 -596 -7143 -562
rect -7109 -596 -7097 -562
rect -7155 -630 -7097 -596
rect -7155 -664 -7143 -630
rect -7109 -664 -7097 -630
rect -7155 -709 -7097 -664
rect -6137 -154 -6079 -109
rect -6137 -188 -6125 -154
rect -6091 -188 -6079 -154
rect -6137 -222 -6079 -188
rect -6137 -256 -6125 -222
rect -6091 -256 -6079 -222
rect -6137 -290 -6079 -256
rect -6137 -324 -6125 -290
rect -6091 -324 -6079 -290
rect -6137 -358 -6079 -324
rect -6137 -392 -6125 -358
rect -6091 -392 -6079 -358
rect -6137 -426 -6079 -392
rect -6137 -460 -6125 -426
rect -6091 -460 -6079 -426
rect -6137 -494 -6079 -460
rect -6137 -528 -6125 -494
rect -6091 -528 -6079 -494
rect -6137 -562 -6079 -528
rect -6137 -596 -6125 -562
rect -6091 -596 -6079 -562
rect -6137 -630 -6079 -596
rect -6137 -664 -6125 -630
rect -6091 -664 -6079 -630
rect -6137 -709 -6079 -664
rect -5119 -154 -5061 -109
rect -5119 -188 -5107 -154
rect -5073 -188 -5061 -154
rect -5119 -222 -5061 -188
rect -5119 -256 -5107 -222
rect -5073 -256 -5061 -222
rect -5119 -290 -5061 -256
rect -5119 -324 -5107 -290
rect -5073 -324 -5061 -290
rect -5119 -358 -5061 -324
rect -5119 -392 -5107 -358
rect -5073 -392 -5061 -358
rect -5119 -426 -5061 -392
rect -5119 -460 -5107 -426
rect -5073 -460 -5061 -426
rect -5119 -494 -5061 -460
rect -5119 -528 -5107 -494
rect -5073 -528 -5061 -494
rect -5119 -562 -5061 -528
rect -5119 -596 -5107 -562
rect -5073 -596 -5061 -562
rect -5119 -630 -5061 -596
rect -5119 -664 -5107 -630
rect -5073 -664 -5061 -630
rect -5119 -709 -5061 -664
rect -4101 -154 -4043 -109
rect -4101 -188 -4089 -154
rect -4055 -188 -4043 -154
rect -4101 -222 -4043 -188
rect -4101 -256 -4089 -222
rect -4055 -256 -4043 -222
rect -4101 -290 -4043 -256
rect -4101 -324 -4089 -290
rect -4055 -324 -4043 -290
rect -4101 -358 -4043 -324
rect -4101 -392 -4089 -358
rect -4055 -392 -4043 -358
rect -4101 -426 -4043 -392
rect -4101 -460 -4089 -426
rect -4055 -460 -4043 -426
rect -4101 -494 -4043 -460
rect -4101 -528 -4089 -494
rect -4055 -528 -4043 -494
rect -4101 -562 -4043 -528
rect -4101 -596 -4089 -562
rect -4055 -596 -4043 -562
rect -4101 -630 -4043 -596
rect -4101 -664 -4089 -630
rect -4055 -664 -4043 -630
rect -4101 -709 -4043 -664
rect -3083 -154 -3025 -109
rect -3083 -188 -3071 -154
rect -3037 -188 -3025 -154
rect -3083 -222 -3025 -188
rect -3083 -256 -3071 -222
rect -3037 -256 -3025 -222
rect -3083 -290 -3025 -256
rect -3083 -324 -3071 -290
rect -3037 -324 -3025 -290
rect -3083 -358 -3025 -324
rect -3083 -392 -3071 -358
rect -3037 -392 -3025 -358
rect -3083 -426 -3025 -392
rect -3083 -460 -3071 -426
rect -3037 -460 -3025 -426
rect -3083 -494 -3025 -460
rect -3083 -528 -3071 -494
rect -3037 -528 -3025 -494
rect -3083 -562 -3025 -528
rect -3083 -596 -3071 -562
rect -3037 -596 -3025 -562
rect -3083 -630 -3025 -596
rect -3083 -664 -3071 -630
rect -3037 -664 -3025 -630
rect -3083 -709 -3025 -664
rect -2065 -154 -2007 -109
rect -2065 -188 -2053 -154
rect -2019 -188 -2007 -154
rect -2065 -222 -2007 -188
rect -2065 -256 -2053 -222
rect -2019 -256 -2007 -222
rect -2065 -290 -2007 -256
rect -2065 -324 -2053 -290
rect -2019 -324 -2007 -290
rect -2065 -358 -2007 -324
rect -2065 -392 -2053 -358
rect -2019 -392 -2007 -358
rect -2065 -426 -2007 -392
rect -2065 -460 -2053 -426
rect -2019 -460 -2007 -426
rect -2065 -494 -2007 -460
rect -2065 -528 -2053 -494
rect -2019 -528 -2007 -494
rect -2065 -562 -2007 -528
rect -2065 -596 -2053 -562
rect -2019 -596 -2007 -562
rect -2065 -630 -2007 -596
rect -2065 -664 -2053 -630
rect -2019 -664 -2007 -630
rect -2065 -709 -2007 -664
rect -1047 -154 -989 -109
rect -1047 -188 -1035 -154
rect -1001 -188 -989 -154
rect -1047 -222 -989 -188
rect -1047 -256 -1035 -222
rect -1001 -256 -989 -222
rect -1047 -290 -989 -256
rect -1047 -324 -1035 -290
rect -1001 -324 -989 -290
rect -1047 -358 -989 -324
rect -1047 -392 -1035 -358
rect -1001 -392 -989 -358
rect -1047 -426 -989 -392
rect -1047 -460 -1035 -426
rect -1001 -460 -989 -426
rect -1047 -494 -989 -460
rect -1047 -528 -1035 -494
rect -1001 -528 -989 -494
rect -1047 -562 -989 -528
rect -1047 -596 -1035 -562
rect -1001 -596 -989 -562
rect -1047 -630 -989 -596
rect -1047 -664 -1035 -630
rect -1001 -664 -989 -630
rect -1047 -709 -989 -664
rect -29 -154 29 -109
rect -29 -188 -17 -154
rect 17 -188 29 -154
rect -29 -222 29 -188
rect -29 -256 -17 -222
rect 17 -256 29 -222
rect -29 -290 29 -256
rect -29 -324 -17 -290
rect 17 -324 29 -290
rect -29 -358 29 -324
rect -29 -392 -17 -358
rect 17 -392 29 -358
rect -29 -426 29 -392
rect -29 -460 -17 -426
rect 17 -460 29 -426
rect -29 -494 29 -460
rect -29 -528 -17 -494
rect 17 -528 29 -494
rect -29 -562 29 -528
rect -29 -596 -17 -562
rect 17 -596 29 -562
rect -29 -630 29 -596
rect -29 -664 -17 -630
rect 17 -664 29 -630
rect -29 -709 29 -664
rect 989 -154 1047 -109
rect 989 -188 1001 -154
rect 1035 -188 1047 -154
rect 989 -222 1047 -188
rect 989 -256 1001 -222
rect 1035 -256 1047 -222
rect 989 -290 1047 -256
rect 989 -324 1001 -290
rect 1035 -324 1047 -290
rect 989 -358 1047 -324
rect 989 -392 1001 -358
rect 1035 -392 1047 -358
rect 989 -426 1047 -392
rect 989 -460 1001 -426
rect 1035 -460 1047 -426
rect 989 -494 1047 -460
rect 989 -528 1001 -494
rect 1035 -528 1047 -494
rect 989 -562 1047 -528
rect 989 -596 1001 -562
rect 1035 -596 1047 -562
rect 989 -630 1047 -596
rect 989 -664 1001 -630
rect 1035 -664 1047 -630
rect 989 -709 1047 -664
rect 2007 -154 2065 -109
rect 2007 -188 2019 -154
rect 2053 -188 2065 -154
rect 2007 -222 2065 -188
rect 2007 -256 2019 -222
rect 2053 -256 2065 -222
rect 2007 -290 2065 -256
rect 2007 -324 2019 -290
rect 2053 -324 2065 -290
rect 2007 -358 2065 -324
rect 2007 -392 2019 -358
rect 2053 -392 2065 -358
rect 2007 -426 2065 -392
rect 2007 -460 2019 -426
rect 2053 -460 2065 -426
rect 2007 -494 2065 -460
rect 2007 -528 2019 -494
rect 2053 -528 2065 -494
rect 2007 -562 2065 -528
rect 2007 -596 2019 -562
rect 2053 -596 2065 -562
rect 2007 -630 2065 -596
rect 2007 -664 2019 -630
rect 2053 -664 2065 -630
rect 2007 -709 2065 -664
rect 3025 -154 3083 -109
rect 3025 -188 3037 -154
rect 3071 -188 3083 -154
rect 3025 -222 3083 -188
rect 3025 -256 3037 -222
rect 3071 -256 3083 -222
rect 3025 -290 3083 -256
rect 3025 -324 3037 -290
rect 3071 -324 3083 -290
rect 3025 -358 3083 -324
rect 3025 -392 3037 -358
rect 3071 -392 3083 -358
rect 3025 -426 3083 -392
rect 3025 -460 3037 -426
rect 3071 -460 3083 -426
rect 3025 -494 3083 -460
rect 3025 -528 3037 -494
rect 3071 -528 3083 -494
rect 3025 -562 3083 -528
rect 3025 -596 3037 -562
rect 3071 -596 3083 -562
rect 3025 -630 3083 -596
rect 3025 -664 3037 -630
rect 3071 -664 3083 -630
rect 3025 -709 3083 -664
rect 4043 -154 4101 -109
rect 4043 -188 4055 -154
rect 4089 -188 4101 -154
rect 4043 -222 4101 -188
rect 4043 -256 4055 -222
rect 4089 -256 4101 -222
rect 4043 -290 4101 -256
rect 4043 -324 4055 -290
rect 4089 -324 4101 -290
rect 4043 -358 4101 -324
rect 4043 -392 4055 -358
rect 4089 -392 4101 -358
rect 4043 -426 4101 -392
rect 4043 -460 4055 -426
rect 4089 -460 4101 -426
rect 4043 -494 4101 -460
rect 4043 -528 4055 -494
rect 4089 -528 4101 -494
rect 4043 -562 4101 -528
rect 4043 -596 4055 -562
rect 4089 -596 4101 -562
rect 4043 -630 4101 -596
rect 4043 -664 4055 -630
rect 4089 -664 4101 -630
rect 4043 -709 4101 -664
rect 5061 -154 5119 -109
rect 5061 -188 5073 -154
rect 5107 -188 5119 -154
rect 5061 -222 5119 -188
rect 5061 -256 5073 -222
rect 5107 -256 5119 -222
rect 5061 -290 5119 -256
rect 5061 -324 5073 -290
rect 5107 -324 5119 -290
rect 5061 -358 5119 -324
rect 5061 -392 5073 -358
rect 5107 -392 5119 -358
rect 5061 -426 5119 -392
rect 5061 -460 5073 -426
rect 5107 -460 5119 -426
rect 5061 -494 5119 -460
rect 5061 -528 5073 -494
rect 5107 -528 5119 -494
rect 5061 -562 5119 -528
rect 5061 -596 5073 -562
rect 5107 -596 5119 -562
rect 5061 -630 5119 -596
rect 5061 -664 5073 -630
rect 5107 -664 5119 -630
rect 5061 -709 5119 -664
rect 6079 -154 6137 -109
rect 6079 -188 6091 -154
rect 6125 -188 6137 -154
rect 6079 -222 6137 -188
rect 6079 -256 6091 -222
rect 6125 -256 6137 -222
rect 6079 -290 6137 -256
rect 6079 -324 6091 -290
rect 6125 -324 6137 -290
rect 6079 -358 6137 -324
rect 6079 -392 6091 -358
rect 6125 -392 6137 -358
rect 6079 -426 6137 -392
rect 6079 -460 6091 -426
rect 6125 -460 6137 -426
rect 6079 -494 6137 -460
rect 6079 -528 6091 -494
rect 6125 -528 6137 -494
rect 6079 -562 6137 -528
rect 6079 -596 6091 -562
rect 6125 -596 6137 -562
rect 6079 -630 6137 -596
rect 6079 -664 6091 -630
rect 6125 -664 6137 -630
rect 6079 -709 6137 -664
rect 7097 -154 7155 -109
rect 7097 -188 7109 -154
rect 7143 -188 7155 -154
rect 7097 -222 7155 -188
rect 7097 -256 7109 -222
rect 7143 -256 7155 -222
rect 7097 -290 7155 -256
rect 7097 -324 7109 -290
rect 7143 -324 7155 -290
rect 7097 -358 7155 -324
rect 7097 -392 7109 -358
rect 7143 -392 7155 -358
rect 7097 -426 7155 -392
rect 7097 -460 7109 -426
rect 7143 -460 7155 -426
rect 7097 -494 7155 -460
rect 7097 -528 7109 -494
rect 7143 -528 7155 -494
rect 7097 -562 7155 -528
rect 7097 -596 7109 -562
rect 7143 -596 7155 -562
rect 7097 -630 7155 -596
rect 7097 -664 7109 -630
rect 7143 -664 7155 -630
rect 7097 -709 7155 -664
rect 8115 -154 8173 -109
rect 8115 -188 8127 -154
rect 8161 -188 8173 -154
rect 8115 -222 8173 -188
rect 8115 -256 8127 -222
rect 8161 -256 8173 -222
rect 8115 -290 8173 -256
rect 8115 -324 8127 -290
rect 8161 -324 8173 -290
rect 8115 -358 8173 -324
rect 8115 -392 8127 -358
rect 8161 -392 8173 -358
rect 8115 -426 8173 -392
rect 8115 -460 8127 -426
rect 8161 -460 8173 -426
rect 8115 -494 8173 -460
rect 8115 -528 8127 -494
rect 8161 -528 8173 -494
rect 8115 -562 8173 -528
rect 8115 -596 8127 -562
rect 8161 -596 8173 -562
rect 8115 -630 8173 -596
rect 8115 -664 8127 -630
rect 8161 -664 8173 -630
rect 8115 -709 8173 -664
rect 9133 -154 9191 -109
rect 9133 -188 9145 -154
rect 9179 -188 9191 -154
rect 9133 -222 9191 -188
rect 9133 -256 9145 -222
rect 9179 -256 9191 -222
rect 9133 -290 9191 -256
rect 9133 -324 9145 -290
rect 9179 -324 9191 -290
rect 9133 -358 9191 -324
rect 9133 -392 9145 -358
rect 9179 -392 9191 -358
rect 9133 -426 9191 -392
rect 9133 -460 9145 -426
rect 9179 -460 9191 -426
rect 9133 -494 9191 -460
rect 9133 -528 9145 -494
rect 9179 -528 9191 -494
rect 9133 -562 9191 -528
rect 9133 -596 9145 -562
rect 9179 -596 9191 -562
rect 9133 -630 9191 -596
rect 9133 -664 9145 -630
rect 9179 -664 9191 -630
rect 9133 -709 9191 -664
rect 10151 -154 10209 -109
rect 10151 -188 10163 -154
rect 10197 -188 10209 -154
rect 10151 -222 10209 -188
rect 10151 -256 10163 -222
rect 10197 -256 10209 -222
rect 10151 -290 10209 -256
rect 10151 -324 10163 -290
rect 10197 -324 10209 -290
rect 10151 -358 10209 -324
rect 10151 -392 10163 -358
rect 10197 -392 10209 -358
rect 10151 -426 10209 -392
rect 10151 -460 10163 -426
rect 10197 -460 10209 -426
rect 10151 -494 10209 -460
rect 10151 -528 10163 -494
rect 10197 -528 10209 -494
rect 10151 -562 10209 -528
rect 10151 -596 10163 -562
rect 10197 -596 10209 -562
rect 10151 -630 10209 -596
rect 10151 -664 10163 -630
rect 10197 -664 10209 -630
rect 10151 -709 10209 -664
<< ndiffc >>
rect -10197 630 -10163 664
rect -10197 562 -10163 596
rect -10197 494 -10163 528
rect -10197 426 -10163 460
rect -10197 358 -10163 392
rect -10197 290 -10163 324
rect -10197 222 -10163 256
rect -10197 154 -10163 188
rect -9179 630 -9145 664
rect -9179 562 -9145 596
rect -9179 494 -9145 528
rect -9179 426 -9145 460
rect -9179 358 -9145 392
rect -9179 290 -9145 324
rect -9179 222 -9145 256
rect -9179 154 -9145 188
rect -8161 630 -8127 664
rect -8161 562 -8127 596
rect -8161 494 -8127 528
rect -8161 426 -8127 460
rect -8161 358 -8127 392
rect -8161 290 -8127 324
rect -8161 222 -8127 256
rect -8161 154 -8127 188
rect -7143 630 -7109 664
rect -7143 562 -7109 596
rect -7143 494 -7109 528
rect -7143 426 -7109 460
rect -7143 358 -7109 392
rect -7143 290 -7109 324
rect -7143 222 -7109 256
rect -7143 154 -7109 188
rect -6125 630 -6091 664
rect -6125 562 -6091 596
rect -6125 494 -6091 528
rect -6125 426 -6091 460
rect -6125 358 -6091 392
rect -6125 290 -6091 324
rect -6125 222 -6091 256
rect -6125 154 -6091 188
rect -5107 630 -5073 664
rect -5107 562 -5073 596
rect -5107 494 -5073 528
rect -5107 426 -5073 460
rect -5107 358 -5073 392
rect -5107 290 -5073 324
rect -5107 222 -5073 256
rect -5107 154 -5073 188
rect -4089 630 -4055 664
rect -4089 562 -4055 596
rect -4089 494 -4055 528
rect -4089 426 -4055 460
rect -4089 358 -4055 392
rect -4089 290 -4055 324
rect -4089 222 -4055 256
rect -4089 154 -4055 188
rect -3071 630 -3037 664
rect -3071 562 -3037 596
rect -3071 494 -3037 528
rect -3071 426 -3037 460
rect -3071 358 -3037 392
rect -3071 290 -3037 324
rect -3071 222 -3037 256
rect -3071 154 -3037 188
rect -2053 630 -2019 664
rect -2053 562 -2019 596
rect -2053 494 -2019 528
rect -2053 426 -2019 460
rect -2053 358 -2019 392
rect -2053 290 -2019 324
rect -2053 222 -2019 256
rect -2053 154 -2019 188
rect -1035 630 -1001 664
rect -1035 562 -1001 596
rect -1035 494 -1001 528
rect -1035 426 -1001 460
rect -1035 358 -1001 392
rect -1035 290 -1001 324
rect -1035 222 -1001 256
rect -1035 154 -1001 188
rect -17 630 17 664
rect -17 562 17 596
rect -17 494 17 528
rect -17 426 17 460
rect -17 358 17 392
rect -17 290 17 324
rect -17 222 17 256
rect -17 154 17 188
rect 1001 630 1035 664
rect 1001 562 1035 596
rect 1001 494 1035 528
rect 1001 426 1035 460
rect 1001 358 1035 392
rect 1001 290 1035 324
rect 1001 222 1035 256
rect 1001 154 1035 188
rect 2019 630 2053 664
rect 2019 562 2053 596
rect 2019 494 2053 528
rect 2019 426 2053 460
rect 2019 358 2053 392
rect 2019 290 2053 324
rect 2019 222 2053 256
rect 2019 154 2053 188
rect 3037 630 3071 664
rect 3037 562 3071 596
rect 3037 494 3071 528
rect 3037 426 3071 460
rect 3037 358 3071 392
rect 3037 290 3071 324
rect 3037 222 3071 256
rect 3037 154 3071 188
rect 4055 630 4089 664
rect 4055 562 4089 596
rect 4055 494 4089 528
rect 4055 426 4089 460
rect 4055 358 4089 392
rect 4055 290 4089 324
rect 4055 222 4089 256
rect 4055 154 4089 188
rect 5073 630 5107 664
rect 5073 562 5107 596
rect 5073 494 5107 528
rect 5073 426 5107 460
rect 5073 358 5107 392
rect 5073 290 5107 324
rect 5073 222 5107 256
rect 5073 154 5107 188
rect 6091 630 6125 664
rect 6091 562 6125 596
rect 6091 494 6125 528
rect 6091 426 6125 460
rect 6091 358 6125 392
rect 6091 290 6125 324
rect 6091 222 6125 256
rect 6091 154 6125 188
rect 7109 630 7143 664
rect 7109 562 7143 596
rect 7109 494 7143 528
rect 7109 426 7143 460
rect 7109 358 7143 392
rect 7109 290 7143 324
rect 7109 222 7143 256
rect 7109 154 7143 188
rect 8127 630 8161 664
rect 8127 562 8161 596
rect 8127 494 8161 528
rect 8127 426 8161 460
rect 8127 358 8161 392
rect 8127 290 8161 324
rect 8127 222 8161 256
rect 8127 154 8161 188
rect 9145 630 9179 664
rect 9145 562 9179 596
rect 9145 494 9179 528
rect 9145 426 9179 460
rect 9145 358 9179 392
rect 9145 290 9179 324
rect 9145 222 9179 256
rect 9145 154 9179 188
rect 10163 630 10197 664
rect 10163 562 10197 596
rect 10163 494 10197 528
rect 10163 426 10197 460
rect 10163 358 10197 392
rect 10163 290 10197 324
rect 10163 222 10197 256
rect 10163 154 10197 188
rect -10197 -188 -10163 -154
rect -10197 -256 -10163 -222
rect -10197 -324 -10163 -290
rect -10197 -392 -10163 -358
rect -10197 -460 -10163 -426
rect -10197 -528 -10163 -494
rect -10197 -596 -10163 -562
rect -10197 -664 -10163 -630
rect -9179 -188 -9145 -154
rect -9179 -256 -9145 -222
rect -9179 -324 -9145 -290
rect -9179 -392 -9145 -358
rect -9179 -460 -9145 -426
rect -9179 -528 -9145 -494
rect -9179 -596 -9145 -562
rect -9179 -664 -9145 -630
rect -8161 -188 -8127 -154
rect -8161 -256 -8127 -222
rect -8161 -324 -8127 -290
rect -8161 -392 -8127 -358
rect -8161 -460 -8127 -426
rect -8161 -528 -8127 -494
rect -8161 -596 -8127 -562
rect -8161 -664 -8127 -630
rect -7143 -188 -7109 -154
rect -7143 -256 -7109 -222
rect -7143 -324 -7109 -290
rect -7143 -392 -7109 -358
rect -7143 -460 -7109 -426
rect -7143 -528 -7109 -494
rect -7143 -596 -7109 -562
rect -7143 -664 -7109 -630
rect -6125 -188 -6091 -154
rect -6125 -256 -6091 -222
rect -6125 -324 -6091 -290
rect -6125 -392 -6091 -358
rect -6125 -460 -6091 -426
rect -6125 -528 -6091 -494
rect -6125 -596 -6091 -562
rect -6125 -664 -6091 -630
rect -5107 -188 -5073 -154
rect -5107 -256 -5073 -222
rect -5107 -324 -5073 -290
rect -5107 -392 -5073 -358
rect -5107 -460 -5073 -426
rect -5107 -528 -5073 -494
rect -5107 -596 -5073 -562
rect -5107 -664 -5073 -630
rect -4089 -188 -4055 -154
rect -4089 -256 -4055 -222
rect -4089 -324 -4055 -290
rect -4089 -392 -4055 -358
rect -4089 -460 -4055 -426
rect -4089 -528 -4055 -494
rect -4089 -596 -4055 -562
rect -4089 -664 -4055 -630
rect -3071 -188 -3037 -154
rect -3071 -256 -3037 -222
rect -3071 -324 -3037 -290
rect -3071 -392 -3037 -358
rect -3071 -460 -3037 -426
rect -3071 -528 -3037 -494
rect -3071 -596 -3037 -562
rect -3071 -664 -3037 -630
rect -2053 -188 -2019 -154
rect -2053 -256 -2019 -222
rect -2053 -324 -2019 -290
rect -2053 -392 -2019 -358
rect -2053 -460 -2019 -426
rect -2053 -528 -2019 -494
rect -2053 -596 -2019 -562
rect -2053 -664 -2019 -630
rect -1035 -188 -1001 -154
rect -1035 -256 -1001 -222
rect -1035 -324 -1001 -290
rect -1035 -392 -1001 -358
rect -1035 -460 -1001 -426
rect -1035 -528 -1001 -494
rect -1035 -596 -1001 -562
rect -1035 -664 -1001 -630
rect -17 -188 17 -154
rect -17 -256 17 -222
rect -17 -324 17 -290
rect -17 -392 17 -358
rect -17 -460 17 -426
rect -17 -528 17 -494
rect -17 -596 17 -562
rect -17 -664 17 -630
rect 1001 -188 1035 -154
rect 1001 -256 1035 -222
rect 1001 -324 1035 -290
rect 1001 -392 1035 -358
rect 1001 -460 1035 -426
rect 1001 -528 1035 -494
rect 1001 -596 1035 -562
rect 1001 -664 1035 -630
rect 2019 -188 2053 -154
rect 2019 -256 2053 -222
rect 2019 -324 2053 -290
rect 2019 -392 2053 -358
rect 2019 -460 2053 -426
rect 2019 -528 2053 -494
rect 2019 -596 2053 -562
rect 2019 -664 2053 -630
rect 3037 -188 3071 -154
rect 3037 -256 3071 -222
rect 3037 -324 3071 -290
rect 3037 -392 3071 -358
rect 3037 -460 3071 -426
rect 3037 -528 3071 -494
rect 3037 -596 3071 -562
rect 3037 -664 3071 -630
rect 4055 -188 4089 -154
rect 4055 -256 4089 -222
rect 4055 -324 4089 -290
rect 4055 -392 4089 -358
rect 4055 -460 4089 -426
rect 4055 -528 4089 -494
rect 4055 -596 4089 -562
rect 4055 -664 4089 -630
rect 5073 -188 5107 -154
rect 5073 -256 5107 -222
rect 5073 -324 5107 -290
rect 5073 -392 5107 -358
rect 5073 -460 5107 -426
rect 5073 -528 5107 -494
rect 5073 -596 5107 -562
rect 5073 -664 5107 -630
rect 6091 -188 6125 -154
rect 6091 -256 6125 -222
rect 6091 -324 6125 -290
rect 6091 -392 6125 -358
rect 6091 -460 6125 -426
rect 6091 -528 6125 -494
rect 6091 -596 6125 -562
rect 6091 -664 6125 -630
rect 7109 -188 7143 -154
rect 7109 -256 7143 -222
rect 7109 -324 7143 -290
rect 7109 -392 7143 -358
rect 7109 -460 7143 -426
rect 7109 -528 7143 -494
rect 7109 -596 7143 -562
rect 7109 -664 7143 -630
rect 8127 -188 8161 -154
rect 8127 -256 8161 -222
rect 8127 -324 8161 -290
rect 8127 -392 8161 -358
rect 8127 -460 8161 -426
rect 8127 -528 8161 -494
rect 8127 -596 8161 -562
rect 8127 -664 8161 -630
rect 9145 -188 9179 -154
rect 9145 -256 9179 -222
rect 9145 -324 9179 -290
rect 9145 -392 9179 -358
rect 9145 -460 9179 -426
rect 9145 -528 9179 -494
rect 9145 -596 9179 -562
rect 9145 -664 9179 -630
rect 10163 -188 10197 -154
rect 10163 -256 10197 -222
rect 10163 -324 10197 -290
rect 10163 -392 10197 -358
rect 10163 -460 10197 -426
rect 10163 -528 10197 -494
rect 10163 -596 10197 -562
rect 10163 -664 10197 -630
<< poly >>
rect -9965 781 -9377 797
rect -9965 764 -9926 781
rect -10151 747 -9926 764
rect -9892 747 -9858 781
rect -9824 747 -9790 781
rect -9756 747 -9722 781
rect -9688 747 -9654 781
rect -9620 747 -9586 781
rect -9552 747 -9518 781
rect -9484 747 -9450 781
rect -9416 764 -9377 781
rect -8947 781 -8359 797
rect -8947 764 -8908 781
rect -9416 747 -9191 764
rect -10151 709 -9191 747
rect -9133 747 -8908 764
rect -8874 747 -8840 781
rect -8806 747 -8772 781
rect -8738 747 -8704 781
rect -8670 747 -8636 781
rect -8602 747 -8568 781
rect -8534 747 -8500 781
rect -8466 747 -8432 781
rect -8398 764 -8359 781
rect -7929 781 -7341 797
rect -7929 764 -7890 781
rect -8398 747 -8173 764
rect -9133 709 -8173 747
rect -8115 747 -7890 764
rect -7856 747 -7822 781
rect -7788 747 -7754 781
rect -7720 747 -7686 781
rect -7652 747 -7618 781
rect -7584 747 -7550 781
rect -7516 747 -7482 781
rect -7448 747 -7414 781
rect -7380 764 -7341 781
rect -6911 781 -6323 797
rect -6911 764 -6872 781
rect -7380 747 -7155 764
rect -8115 709 -7155 747
rect -7097 747 -6872 764
rect -6838 747 -6804 781
rect -6770 747 -6736 781
rect -6702 747 -6668 781
rect -6634 747 -6600 781
rect -6566 747 -6532 781
rect -6498 747 -6464 781
rect -6430 747 -6396 781
rect -6362 764 -6323 781
rect -5893 781 -5305 797
rect -5893 764 -5854 781
rect -6362 747 -6137 764
rect -7097 709 -6137 747
rect -6079 747 -5854 764
rect -5820 747 -5786 781
rect -5752 747 -5718 781
rect -5684 747 -5650 781
rect -5616 747 -5582 781
rect -5548 747 -5514 781
rect -5480 747 -5446 781
rect -5412 747 -5378 781
rect -5344 764 -5305 781
rect -4875 781 -4287 797
rect -4875 764 -4836 781
rect -5344 747 -5119 764
rect -6079 709 -5119 747
rect -5061 747 -4836 764
rect -4802 747 -4768 781
rect -4734 747 -4700 781
rect -4666 747 -4632 781
rect -4598 747 -4564 781
rect -4530 747 -4496 781
rect -4462 747 -4428 781
rect -4394 747 -4360 781
rect -4326 764 -4287 781
rect -3857 781 -3269 797
rect -3857 764 -3818 781
rect -4326 747 -4101 764
rect -5061 709 -4101 747
rect -4043 747 -3818 764
rect -3784 747 -3750 781
rect -3716 747 -3682 781
rect -3648 747 -3614 781
rect -3580 747 -3546 781
rect -3512 747 -3478 781
rect -3444 747 -3410 781
rect -3376 747 -3342 781
rect -3308 764 -3269 781
rect -2839 781 -2251 797
rect -2839 764 -2800 781
rect -3308 747 -3083 764
rect -4043 709 -3083 747
rect -3025 747 -2800 764
rect -2766 747 -2732 781
rect -2698 747 -2664 781
rect -2630 747 -2596 781
rect -2562 747 -2528 781
rect -2494 747 -2460 781
rect -2426 747 -2392 781
rect -2358 747 -2324 781
rect -2290 764 -2251 781
rect -1821 781 -1233 797
rect -1821 764 -1782 781
rect -2290 747 -2065 764
rect -3025 709 -2065 747
rect -2007 747 -1782 764
rect -1748 747 -1714 781
rect -1680 747 -1646 781
rect -1612 747 -1578 781
rect -1544 747 -1510 781
rect -1476 747 -1442 781
rect -1408 747 -1374 781
rect -1340 747 -1306 781
rect -1272 764 -1233 781
rect -803 781 -215 797
rect -803 764 -764 781
rect -1272 747 -1047 764
rect -2007 709 -1047 747
rect -989 747 -764 764
rect -730 747 -696 781
rect -662 747 -628 781
rect -594 747 -560 781
rect -526 747 -492 781
rect -458 747 -424 781
rect -390 747 -356 781
rect -322 747 -288 781
rect -254 764 -215 781
rect 215 781 803 797
rect 215 764 254 781
rect -254 747 -29 764
rect -989 709 -29 747
rect 29 747 254 764
rect 288 747 322 781
rect 356 747 390 781
rect 424 747 458 781
rect 492 747 526 781
rect 560 747 594 781
rect 628 747 662 781
rect 696 747 730 781
rect 764 764 803 781
rect 1233 781 1821 797
rect 1233 764 1272 781
rect 764 747 989 764
rect 29 709 989 747
rect 1047 747 1272 764
rect 1306 747 1340 781
rect 1374 747 1408 781
rect 1442 747 1476 781
rect 1510 747 1544 781
rect 1578 747 1612 781
rect 1646 747 1680 781
rect 1714 747 1748 781
rect 1782 764 1821 781
rect 2251 781 2839 797
rect 2251 764 2290 781
rect 1782 747 2007 764
rect 1047 709 2007 747
rect 2065 747 2290 764
rect 2324 747 2358 781
rect 2392 747 2426 781
rect 2460 747 2494 781
rect 2528 747 2562 781
rect 2596 747 2630 781
rect 2664 747 2698 781
rect 2732 747 2766 781
rect 2800 764 2839 781
rect 3269 781 3857 797
rect 3269 764 3308 781
rect 2800 747 3025 764
rect 2065 709 3025 747
rect 3083 747 3308 764
rect 3342 747 3376 781
rect 3410 747 3444 781
rect 3478 747 3512 781
rect 3546 747 3580 781
rect 3614 747 3648 781
rect 3682 747 3716 781
rect 3750 747 3784 781
rect 3818 764 3857 781
rect 4287 781 4875 797
rect 4287 764 4326 781
rect 3818 747 4043 764
rect 3083 709 4043 747
rect 4101 747 4326 764
rect 4360 747 4394 781
rect 4428 747 4462 781
rect 4496 747 4530 781
rect 4564 747 4598 781
rect 4632 747 4666 781
rect 4700 747 4734 781
rect 4768 747 4802 781
rect 4836 764 4875 781
rect 5305 781 5893 797
rect 5305 764 5344 781
rect 4836 747 5061 764
rect 4101 709 5061 747
rect 5119 747 5344 764
rect 5378 747 5412 781
rect 5446 747 5480 781
rect 5514 747 5548 781
rect 5582 747 5616 781
rect 5650 747 5684 781
rect 5718 747 5752 781
rect 5786 747 5820 781
rect 5854 764 5893 781
rect 6323 781 6911 797
rect 6323 764 6362 781
rect 5854 747 6079 764
rect 5119 709 6079 747
rect 6137 747 6362 764
rect 6396 747 6430 781
rect 6464 747 6498 781
rect 6532 747 6566 781
rect 6600 747 6634 781
rect 6668 747 6702 781
rect 6736 747 6770 781
rect 6804 747 6838 781
rect 6872 764 6911 781
rect 7341 781 7929 797
rect 7341 764 7380 781
rect 6872 747 7097 764
rect 6137 709 7097 747
rect 7155 747 7380 764
rect 7414 747 7448 781
rect 7482 747 7516 781
rect 7550 747 7584 781
rect 7618 747 7652 781
rect 7686 747 7720 781
rect 7754 747 7788 781
rect 7822 747 7856 781
rect 7890 764 7929 781
rect 8359 781 8947 797
rect 8359 764 8398 781
rect 7890 747 8115 764
rect 7155 709 8115 747
rect 8173 747 8398 764
rect 8432 747 8466 781
rect 8500 747 8534 781
rect 8568 747 8602 781
rect 8636 747 8670 781
rect 8704 747 8738 781
rect 8772 747 8806 781
rect 8840 747 8874 781
rect 8908 764 8947 781
rect 9377 781 9965 797
rect 9377 764 9416 781
rect 8908 747 9133 764
rect 8173 709 9133 747
rect 9191 747 9416 764
rect 9450 747 9484 781
rect 9518 747 9552 781
rect 9586 747 9620 781
rect 9654 747 9688 781
rect 9722 747 9756 781
rect 9790 747 9824 781
rect 9858 747 9892 781
rect 9926 764 9965 781
rect 9926 747 10151 764
rect 9191 709 10151 747
rect -10151 71 -9191 109
rect -10151 54 -9926 71
rect -9965 37 -9926 54
rect -9892 37 -9858 71
rect -9824 37 -9790 71
rect -9756 37 -9722 71
rect -9688 37 -9654 71
rect -9620 37 -9586 71
rect -9552 37 -9518 71
rect -9484 37 -9450 71
rect -9416 54 -9191 71
rect -9133 71 -8173 109
rect -9133 54 -8908 71
rect -9416 37 -9377 54
rect -9965 21 -9377 37
rect -8947 37 -8908 54
rect -8874 37 -8840 71
rect -8806 37 -8772 71
rect -8738 37 -8704 71
rect -8670 37 -8636 71
rect -8602 37 -8568 71
rect -8534 37 -8500 71
rect -8466 37 -8432 71
rect -8398 54 -8173 71
rect -8115 71 -7155 109
rect -8115 54 -7890 71
rect -8398 37 -8359 54
rect -8947 21 -8359 37
rect -7929 37 -7890 54
rect -7856 37 -7822 71
rect -7788 37 -7754 71
rect -7720 37 -7686 71
rect -7652 37 -7618 71
rect -7584 37 -7550 71
rect -7516 37 -7482 71
rect -7448 37 -7414 71
rect -7380 54 -7155 71
rect -7097 71 -6137 109
rect -7097 54 -6872 71
rect -7380 37 -7341 54
rect -7929 21 -7341 37
rect -6911 37 -6872 54
rect -6838 37 -6804 71
rect -6770 37 -6736 71
rect -6702 37 -6668 71
rect -6634 37 -6600 71
rect -6566 37 -6532 71
rect -6498 37 -6464 71
rect -6430 37 -6396 71
rect -6362 54 -6137 71
rect -6079 71 -5119 109
rect -6079 54 -5854 71
rect -6362 37 -6323 54
rect -6911 21 -6323 37
rect -5893 37 -5854 54
rect -5820 37 -5786 71
rect -5752 37 -5718 71
rect -5684 37 -5650 71
rect -5616 37 -5582 71
rect -5548 37 -5514 71
rect -5480 37 -5446 71
rect -5412 37 -5378 71
rect -5344 54 -5119 71
rect -5061 71 -4101 109
rect -5061 54 -4836 71
rect -5344 37 -5305 54
rect -5893 21 -5305 37
rect -4875 37 -4836 54
rect -4802 37 -4768 71
rect -4734 37 -4700 71
rect -4666 37 -4632 71
rect -4598 37 -4564 71
rect -4530 37 -4496 71
rect -4462 37 -4428 71
rect -4394 37 -4360 71
rect -4326 54 -4101 71
rect -4043 71 -3083 109
rect -4043 54 -3818 71
rect -4326 37 -4287 54
rect -4875 21 -4287 37
rect -3857 37 -3818 54
rect -3784 37 -3750 71
rect -3716 37 -3682 71
rect -3648 37 -3614 71
rect -3580 37 -3546 71
rect -3512 37 -3478 71
rect -3444 37 -3410 71
rect -3376 37 -3342 71
rect -3308 54 -3083 71
rect -3025 71 -2065 109
rect -3025 54 -2800 71
rect -3308 37 -3269 54
rect -3857 21 -3269 37
rect -2839 37 -2800 54
rect -2766 37 -2732 71
rect -2698 37 -2664 71
rect -2630 37 -2596 71
rect -2562 37 -2528 71
rect -2494 37 -2460 71
rect -2426 37 -2392 71
rect -2358 37 -2324 71
rect -2290 54 -2065 71
rect -2007 71 -1047 109
rect -2007 54 -1782 71
rect -2290 37 -2251 54
rect -2839 21 -2251 37
rect -1821 37 -1782 54
rect -1748 37 -1714 71
rect -1680 37 -1646 71
rect -1612 37 -1578 71
rect -1544 37 -1510 71
rect -1476 37 -1442 71
rect -1408 37 -1374 71
rect -1340 37 -1306 71
rect -1272 54 -1047 71
rect -989 71 -29 109
rect -989 54 -764 71
rect -1272 37 -1233 54
rect -1821 21 -1233 37
rect -803 37 -764 54
rect -730 37 -696 71
rect -662 37 -628 71
rect -594 37 -560 71
rect -526 37 -492 71
rect -458 37 -424 71
rect -390 37 -356 71
rect -322 37 -288 71
rect -254 54 -29 71
rect 29 71 989 109
rect 29 54 254 71
rect -254 37 -215 54
rect -803 21 -215 37
rect 215 37 254 54
rect 288 37 322 71
rect 356 37 390 71
rect 424 37 458 71
rect 492 37 526 71
rect 560 37 594 71
rect 628 37 662 71
rect 696 37 730 71
rect 764 54 989 71
rect 1047 71 2007 109
rect 1047 54 1272 71
rect 764 37 803 54
rect 215 21 803 37
rect 1233 37 1272 54
rect 1306 37 1340 71
rect 1374 37 1408 71
rect 1442 37 1476 71
rect 1510 37 1544 71
rect 1578 37 1612 71
rect 1646 37 1680 71
rect 1714 37 1748 71
rect 1782 54 2007 71
rect 2065 71 3025 109
rect 2065 54 2290 71
rect 1782 37 1821 54
rect 1233 21 1821 37
rect 2251 37 2290 54
rect 2324 37 2358 71
rect 2392 37 2426 71
rect 2460 37 2494 71
rect 2528 37 2562 71
rect 2596 37 2630 71
rect 2664 37 2698 71
rect 2732 37 2766 71
rect 2800 54 3025 71
rect 3083 71 4043 109
rect 3083 54 3308 71
rect 2800 37 2839 54
rect 2251 21 2839 37
rect 3269 37 3308 54
rect 3342 37 3376 71
rect 3410 37 3444 71
rect 3478 37 3512 71
rect 3546 37 3580 71
rect 3614 37 3648 71
rect 3682 37 3716 71
rect 3750 37 3784 71
rect 3818 54 4043 71
rect 4101 71 5061 109
rect 4101 54 4326 71
rect 3818 37 3857 54
rect 3269 21 3857 37
rect 4287 37 4326 54
rect 4360 37 4394 71
rect 4428 37 4462 71
rect 4496 37 4530 71
rect 4564 37 4598 71
rect 4632 37 4666 71
rect 4700 37 4734 71
rect 4768 37 4802 71
rect 4836 54 5061 71
rect 5119 71 6079 109
rect 5119 54 5344 71
rect 4836 37 4875 54
rect 4287 21 4875 37
rect 5305 37 5344 54
rect 5378 37 5412 71
rect 5446 37 5480 71
rect 5514 37 5548 71
rect 5582 37 5616 71
rect 5650 37 5684 71
rect 5718 37 5752 71
rect 5786 37 5820 71
rect 5854 54 6079 71
rect 6137 71 7097 109
rect 6137 54 6362 71
rect 5854 37 5893 54
rect 5305 21 5893 37
rect 6323 37 6362 54
rect 6396 37 6430 71
rect 6464 37 6498 71
rect 6532 37 6566 71
rect 6600 37 6634 71
rect 6668 37 6702 71
rect 6736 37 6770 71
rect 6804 37 6838 71
rect 6872 54 7097 71
rect 7155 71 8115 109
rect 7155 54 7380 71
rect 6872 37 6911 54
rect 6323 21 6911 37
rect 7341 37 7380 54
rect 7414 37 7448 71
rect 7482 37 7516 71
rect 7550 37 7584 71
rect 7618 37 7652 71
rect 7686 37 7720 71
rect 7754 37 7788 71
rect 7822 37 7856 71
rect 7890 54 8115 71
rect 8173 71 9133 109
rect 8173 54 8398 71
rect 7890 37 7929 54
rect 7341 21 7929 37
rect 8359 37 8398 54
rect 8432 37 8466 71
rect 8500 37 8534 71
rect 8568 37 8602 71
rect 8636 37 8670 71
rect 8704 37 8738 71
rect 8772 37 8806 71
rect 8840 37 8874 71
rect 8908 54 9133 71
rect 9191 71 10151 109
rect 9191 54 9416 71
rect 8908 37 8947 54
rect 8359 21 8947 37
rect 9377 37 9416 54
rect 9450 37 9484 71
rect 9518 37 9552 71
rect 9586 37 9620 71
rect 9654 37 9688 71
rect 9722 37 9756 71
rect 9790 37 9824 71
rect 9858 37 9892 71
rect 9926 54 10151 71
rect 9926 37 9965 54
rect 9377 21 9965 37
rect -9965 -37 -9377 -21
rect -9965 -54 -9926 -37
rect -10151 -71 -9926 -54
rect -9892 -71 -9858 -37
rect -9824 -71 -9790 -37
rect -9756 -71 -9722 -37
rect -9688 -71 -9654 -37
rect -9620 -71 -9586 -37
rect -9552 -71 -9518 -37
rect -9484 -71 -9450 -37
rect -9416 -54 -9377 -37
rect -8947 -37 -8359 -21
rect -8947 -54 -8908 -37
rect -9416 -71 -9191 -54
rect -10151 -109 -9191 -71
rect -9133 -71 -8908 -54
rect -8874 -71 -8840 -37
rect -8806 -71 -8772 -37
rect -8738 -71 -8704 -37
rect -8670 -71 -8636 -37
rect -8602 -71 -8568 -37
rect -8534 -71 -8500 -37
rect -8466 -71 -8432 -37
rect -8398 -54 -8359 -37
rect -7929 -37 -7341 -21
rect -7929 -54 -7890 -37
rect -8398 -71 -8173 -54
rect -9133 -109 -8173 -71
rect -8115 -71 -7890 -54
rect -7856 -71 -7822 -37
rect -7788 -71 -7754 -37
rect -7720 -71 -7686 -37
rect -7652 -71 -7618 -37
rect -7584 -71 -7550 -37
rect -7516 -71 -7482 -37
rect -7448 -71 -7414 -37
rect -7380 -54 -7341 -37
rect -6911 -37 -6323 -21
rect -6911 -54 -6872 -37
rect -7380 -71 -7155 -54
rect -8115 -109 -7155 -71
rect -7097 -71 -6872 -54
rect -6838 -71 -6804 -37
rect -6770 -71 -6736 -37
rect -6702 -71 -6668 -37
rect -6634 -71 -6600 -37
rect -6566 -71 -6532 -37
rect -6498 -71 -6464 -37
rect -6430 -71 -6396 -37
rect -6362 -54 -6323 -37
rect -5893 -37 -5305 -21
rect -5893 -54 -5854 -37
rect -6362 -71 -6137 -54
rect -7097 -109 -6137 -71
rect -6079 -71 -5854 -54
rect -5820 -71 -5786 -37
rect -5752 -71 -5718 -37
rect -5684 -71 -5650 -37
rect -5616 -71 -5582 -37
rect -5548 -71 -5514 -37
rect -5480 -71 -5446 -37
rect -5412 -71 -5378 -37
rect -5344 -54 -5305 -37
rect -4875 -37 -4287 -21
rect -4875 -54 -4836 -37
rect -5344 -71 -5119 -54
rect -6079 -109 -5119 -71
rect -5061 -71 -4836 -54
rect -4802 -71 -4768 -37
rect -4734 -71 -4700 -37
rect -4666 -71 -4632 -37
rect -4598 -71 -4564 -37
rect -4530 -71 -4496 -37
rect -4462 -71 -4428 -37
rect -4394 -71 -4360 -37
rect -4326 -54 -4287 -37
rect -3857 -37 -3269 -21
rect -3857 -54 -3818 -37
rect -4326 -71 -4101 -54
rect -5061 -109 -4101 -71
rect -4043 -71 -3818 -54
rect -3784 -71 -3750 -37
rect -3716 -71 -3682 -37
rect -3648 -71 -3614 -37
rect -3580 -71 -3546 -37
rect -3512 -71 -3478 -37
rect -3444 -71 -3410 -37
rect -3376 -71 -3342 -37
rect -3308 -54 -3269 -37
rect -2839 -37 -2251 -21
rect -2839 -54 -2800 -37
rect -3308 -71 -3083 -54
rect -4043 -109 -3083 -71
rect -3025 -71 -2800 -54
rect -2766 -71 -2732 -37
rect -2698 -71 -2664 -37
rect -2630 -71 -2596 -37
rect -2562 -71 -2528 -37
rect -2494 -71 -2460 -37
rect -2426 -71 -2392 -37
rect -2358 -71 -2324 -37
rect -2290 -54 -2251 -37
rect -1821 -37 -1233 -21
rect -1821 -54 -1782 -37
rect -2290 -71 -2065 -54
rect -3025 -109 -2065 -71
rect -2007 -71 -1782 -54
rect -1748 -71 -1714 -37
rect -1680 -71 -1646 -37
rect -1612 -71 -1578 -37
rect -1544 -71 -1510 -37
rect -1476 -71 -1442 -37
rect -1408 -71 -1374 -37
rect -1340 -71 -1306 -37
rect -1272 -54 -1233 -37
rect -803 -37 -215 -21
rect -803 -54 -764 -37
rect -1272 -71 -1047 -54
rect -2007 -109 -1047 -71
rect -989 -71 -764 -54
rect -730 -71 -696 -37
rect -662 -71 -628 -37
rect -594 -71 -560 -37
rect -526 -71 -492 -37
rect -458 -71 -424 -37
rect -390 -71 -356 -37
rect -322 -71 -288 -37
rect -254 -54 -215 -37
rect 215 -37 803 -21
rect 215 -54 254 -37
rect -254 -71 -29 -54
rect -989 -109 -29 -71
rect 29 -71 254 -54
rect 288 -71 322 -37
rect 356 -71 390 -37
rect 424 -71 458 -37
rect 492 -71 526 -37
rect 560 -71 594 -37
rect 628 -71 662 -37
rect 696 -71 730 -37
rect 764 -54 803 -37
rect 1233 -37 1821 -21
rect 1233 -54 1272 -37
rect 764 -71 989 -54
rect 29 -109 989 -71
rect 1047 -71 1272 -54
rect 1306 -71 1340 -37
rect 1374 -71 1408 -37
rect 1442 -71 1476 -37
rect 1510 -71 1544 -37
rect 1578 -71 1612 -37
rect 1646 -71 1680 -37
rect 1714 -71 1748 -37
rect 1782 -54 1821 -37
rect 2251 -37 2839 -21
rect 2251 -54 2290 -37
rect 1782 -71 2007 -54
rect 1047 -109 2007 -71
rect 2065 -71 2290 -54
rect 2324 -71 2358 -37
rect 2392 -71 2426 -37
rect 2460 -71 2494 -37
rect 2528 -71 2562 -37
rect 2596 -71 2630 -37
rect 2664 -71 2698 -37
rect 2732 -71 2766 -37
rect 2800 -54 2839 -37
rect 3269 -37 3857 -21
rect 3269 -54 3308 -37
rect 2800 -71 3025 -54
rect 2065 -109 3025 -71
rect 3083 -71 3308 -54
rect 3342 -71 3376 -37
rect 3410 -71 3444 -37
rect 3478 -71 3512 -37
rect 3546 -71 3580 -37
rect 3614 -71 3648 -37
rect 3682 -71 3716 -37
rect 3750 -71 3784 -37
rect 3818 -54 3857 -37
rect 4287 -37 4875 -21
rect 4287 -54 4326 -37
rect 3818 -71 4043 -54
rect 3083 -109 4043 -71
rect 4101 -71 4326 -54
rect 4360 -71 4394 -37
rect 4428 -71 4462 -37
rect 4496 -71 4530 -37
rect 4564 -71 4598 -37
rect 4632 -71 4666 -37
rect 4700 -71 4734 -37
rect 4768 -71 4802 -37
rect 4836 -54 4875 -37
rect 5305 -37 5893 -21
rect 5305 -54 5344 -37
rect 4836 -71 5061 -54
rect 4101 -109 5061 -71
rect 5119 -71 5344 -54
rect 5378 -71 5412 -37
rect 5446 -71 5480 -37
rect 5514 -71 5548 -37
rect 5582 -71 5616 -37
rect 5650 -71 5684 -37
rect 5718 -71 5752 -37
rect 5786 -71 5820 -37
rect 5854 -54 5893 -37
rect 6323 -37 6911 -21
rect 6323 -54 6362 -37
rect 5854 -71 6079 -54
rect 5119 -109 6079 -71
rect 6137 -71 6362 -54
rect 6396 -71 6430 -37
rect 6464 -71 6498 -37
rect 6532 -71 6566 -37
rect 6600 -71 6634 -37
rect 6668 -71 6702 -37
rect 6736 -71 6770 -37
rect 6804 -71 6838 -37
rect 6872 -54 6911 -37
rect 7341 -37 7929 -21
rect 7341 -54 7380 -37
rect 6872 -71 7097 -54
rect 6137 -109 7097 -71
rect 7155 -71 7380 -54
rect 7414 -71 7448 -37
rect 7482 -71 7516 -37
rect 7550 -71 7584 -37
rect 7618 -71 7652 -37
rect 7686 -71 7720 -37
rect 7754 -71 7788 -37
rect 7822 -71 7856 -37
rect 7890 -54 7929 -37
rect 8359 -37 8947 -21
rect 8359 -54 8398 -37
rect 7890 -71 8115 -54
rect 7155 -109 8115 -71
rect 8173 -71 8398 -54
rect 8432 -71 8466 -37
rect 8500 -71 8534 -37
rect 8568 -71 8602 -37
rect 8636 -71 8670 -37
rect 8704 -71 8738 -37
rect 8772 -71 8806 -37
rect 8840 -71 8874 -37
rect 8908 -54 8947 -37
rect 9377 -37 9965 -21
rect 9377 -54 9416 -37
rect 8908 -71 9133 -54
rect 8173 -109 9133 -71
rect 9191 -71 9416 -54
rect 9450 -71 9484 -37
rect 9518 -71 9552 -37
rect 9586 -71 9620 -37
rect 9654 -71 9688 -37
rect 9722 -71 9756 -37
rect 9790 -71 9824 -37
rect 9858 -71 9892 -37
rect 9926 -54 9965 -37
rect 9926 -71 10151 -54
rect 9191 -109 10151 -71
rect -10151 -747 -9191 -709
rect -10151 -764 -9926 -747
rect -9965 -781 -9926 -764
rect -9892 -781 -9858 -747
rect -9824 -781 -9790 -747
rect -9756 -781 -9722 -747
rect -9688 -781 -9654 -747
rect -9620 -781 -9586 -747
rect -9552 -781 -9518 -747
rect -9484 -781 -9450 -747
rect -9416 -764 -9191 -747
rect -9133 -747 -8173 -709
rect -9133 -764 -8908 -747
rect -9416 -781 -9377 -764
rect -9965 -797 -9377 -781
rect -8947 -781 -8908 -764
rect -8874 -781 -8840 -747
rect -8806 -781 -8772 -747
rect -8738 -781 -8704 -747
rect -8670 -781 -8636 -747
rect -8602 -781 -8568 -747
rect -8534 -781 -8500 -747
rect -8466 -781 -8432 -747
rect -8398 -764 -8173 -747
rect -8115 -747 -7155 -709
rect -8115 -764 -7890 -747
rect -8398 -781 -8359 -764
rect -8947 -797 -8359 -781
rect -7929 -781 -7890 -764
rect -7856 -781 -7822 -747
rect -7788 -781 -7754 -747
rect -7720 -781 -7686 -747
rect -7652 -781 -7618 -747
rect -7584 -781 -7550 -747
rect -7516 -781 -7482 -747
rect -7448 -781 -7414 -747
rect -7380 -764 -7155 -747
rect -7097 -747 -6137 -709
rect -7097 -764 -6872 -747
rect -7380 -781 -7341 -764
rect -7929 -797 -7341 -781
rect -6911 -781 -6872 -764
rect -6838 -781 -6804 -747
rect -6770 -781 -6736 -747
rect -6702 -781 -6668 -747
rect -6634 -781 -6600 -747
rect -6566 -781 -6532 -747
rect -6498 -781 -6464 -747
rect -6430 -781 -6396 -747
rect -6362 -764 -6137 -747
rect -6079 -747 -5119 -709
rect -6079 -764 -5854 -747
rect -6362 -781 -6323 -764
rect -6911 -797 -6323 -781
rect -5893 -781 -5854 -764
rect -5820 -781 -5786 -747
rect -5752 -781 -5718 -747
rect -5684 -781 -5650 -747
rect -5616 -781 -5582 -747
rect -5548 -781 -5514 -747
rect -5480 -781 -5446 -747
rect -5412 -781 -5378 -747
rect -5344 -764 -5119 -747
rect -5061 -747 -4101 -709
rect -5061 -764 -4836 -747
rect -5344 -781 -5305 -764
rect -5893 -797 -5305 -781
rect -4875 -781 -4836 -764
rect -4802 -781 -4768 -747
rect -4734 -781 -4700 -747
rect -4666 -781 -4632 -747
rect -4598 -781 -4564 -747
rect -4530 -781 -4496 -747
rect -4462 -781 -4428 -747
rect -4394 -781 -4360 -747
rect -4326 -764 -4101 -747
rect -4043 -747 -3083 -709
rect -4043 -764 -3818 -747
rect -4326 -781 -4287 -764
rect -4875 -797 -4287 -781
rect -3857 -781 -3818 -764
rect -3784 -781 -3750 -747
rect -3716 -781 -3682 -747
rect -3648 -781 -3614 -747
rect -3580 -781 -3546 -747
rect -3512 -781 -3478 -747
rect -3444 -781 -3410 -747
rect -3376 -781 -3342 -747
rect -3308 -764 -3083 -747
rect -3025 -747 -2065 -709
rect -3025 -764 -2800 -747
rect -3308 -781 -3269 -764
rect -3857 -797 -3269 -781
rect -2839 -781 -2800 -764
rect -2766 -781 -2732 -747
rect -2698 -781 -2664 -747
rect -2630 -781 -2596 -747
rect -2562 -781 -2528 -747
rect -2494 -781 -2460 -747
rect -2426 -781 -2392 -747
rect -2358 -781 -2324 -747
rect -2290 -764 -2065 -747
rect -2007 -747 -1047 -709
rect -2007 -764 -1782 -747
rect -2290 -781 -2251 -764
rect -2839 -797 -2251 -781
rect -1821 -781 -1782 -764
rect -1748 -781 -1714 -747
rect -1680 -781 -1646 -747
rect -1612 -781 -1578 -747
rect -1544 -781 -1510 -747
rect -1476 -781 -1442 -747
rect -1408 -781 -1374 -747
rect -1340 -781 -1306 -747
rect -1272 -764 -1047 -747
rect -989 -747 -29 -709
rect -989 -764 -764 -747
rect -1272 -781 -1233 -764
rect -1821 -797 -1233 -781
rect -803 -781 -764 -764
rect -730 -781 -696 -747
rect -662 -781 -628 -747
rect -594 -781 -560 -747
rect -526 -781 -492 -747
rect -458 -781 -424 -747
rect -390 -781 -356 -747
rect -322 -781 -288 -747
rect -254 -764 -29 -747
rect 29 -747 989 -709
rect 29 -764 254 -747
rect -254 -781 -215 -764
rect -803 -797 -215 -781
rect 215 -781 254 -764
rect 288 -781 322 -747
rect 356 -781 390 -747
rect 424 -781 458 -747
rect 492 -781 526 -747
rect 560 -781 594 -747
rect 628 -781 662 -747
rect 696 -781 730 -747
rect 764 -764 989 -747
rect 1047 -747 2007 -709
rect 1047 -764 1272 -747
rect 764 -781 803 -764
rect 215 -797 803 -781
rect 1233 -781 1272 -764
rect 1306 -781 1340 -747
rect 1374 -781 1408 -747
rect 1442 -781 1476 -747
rect 1510 -781 1544 -747
rect 1578 -781 1612 -747
rect 1646 -781 1680 -747
rect 1714 -781 1748 -747
rect 1782 -764 2007 -747
rect 2065 -747 3025 -709
rect 2065 -764 2290 -747
rect 1782 -781 1821 -764
rect 1233 -797 1821 -781
rect 2251 -781 2290 -764
rect 2324 -781 2358 -747
rect 2392 -781 2426 -747
rect 2460 -781 2494 -747
rect 2528 -781 2562 -747
rect 2596 -781 2630 -747
rect 2664 -781 2698 -747
rect 2732 -781 2766 -747
rect 2800 -764 3025 -747
rect 3083 -747 4043 -709
rect 3083 -764 3308 -747
rect 2800 -781 2839 -764
rect 2251 -797 2839 -781
rect 3269 -781 3308 -764
rect 3342 -781 3376 -747
rect 3410 -781 3444 -747
rect 3478 -781 3512 -747
rect 3546 -781 3580 -747
rect 3614 -781 3648 -747
rect 3682 -781 3716 -747
rect 3750 -781 3784 -747
rect 3818 -764 4043 -747
rect 4101 -747 5061 -709
rect 4101 -764 4326 -747
rect 3818 -781 3857 -764
rect 3269 -797 3857 -781
rect 4287 -781 4326 -764
rect 4360 -781 4394 -747
rect 4428 -781 4462 -747
rect 4496 -781 4530 -747
rect 4564 -781 4598 -747
rect 4632 -781 4666 -747
rect 4700 -781 4734 -747
rect 4768 -781 4802 -747
rect 4836 -764 5061 -747
rect 5119 -747 6079 -709
rect 5119 -764 5344 -747
rect 4836 -781 4875 -764
rect 4287 -797 4875 -781
rect 5305 -781 5344 -764
rect 5378 -781 5412 -747
rect 5446 -781 5480 -747
rect 5514 -781 5548 -747
rect 5582 -781 5616 -747
rect 5650 -781 5684 -747
rect 5718 -781 5752 -747
rect 5786 -781 5820 -747
rect 5854 -764 6079 -747
rect 6137 -747 7097 -709
rect 6137 -764 6362 -747
rect 5854 -781 5893 -764
rect 5305 -797 5893 -781
rect 6323 -781 6362 -764
rect 6396 -781 6430 -747
rect 6464 -781 6498 -747
rect 6532 -781 6566 -747
rect 6600 -781 6634 -747
rect 6668 -781 6702 -747
rect 6736 -781 6770 -747
rect 6804 -781 6838 -747
rect 6872 -764 7097 -747
rect 7155 -747 8115 -709
rect 7155 -764 7380 -747
rect 6872 -781 6911 -764
rect 6323 -797 6911 -781
rect 7341 -781 7380 -764
rect 7414 -781 7448 -747
rect 7482 -781 7516 -747
rect 7550 -781 7584 -747
rect 7618 -781 7652 -747
rect 7686 -781 7720 -747
rect 7754 -781 7788 -747
rect 7822 -781 7856 -747
rect 7890 -764 8115 -747
rect 8173 -747 9133 -709
rect 8173 -764 8398 -747
rect 7890 -781 7929 -764
rect 7341 -797 7929 -781
rect 8359 -781 8398 -764
rect 8432 -781 8466 -747
rect 8500 -781 8534 -747
rect 8568 -781 8602 -747
rect 8636 -781 8670 -747
rect 8704 -781 8738 -747
rect 8772 -781 8806 -747
rect 8840 -781 8874 -747
rect 8908 -764 9133 -747
rect 9191 -747 10151 -709
rect 9191 -764 9416 -747
rect 8908 -781 8947 -764
rect 8359 -797 8947 -781
rect 9377 -781 9416 -764
rect 9450 -781 9484 -747
rect 9518 -781 9552 -747
rect 9586 -781 9620 -747
rect 9654 -781 9688 -747
rect 9722 -781 9756 -747
rect 9790 -781 9824 -747
rect 9858 -781 9892 -747
rect 9926 -764 10151 -747
rect 9926 -781 9965 -764
rect 9377 -797 9965 -781
<< polycont >>
rect -9926 747 -9892 781
rect -9858 747 -9824 781
rect -9790 747 -9756 781
rect -9722 747 -9688 781
rect -9654 747 -9620 781
rect -9586 747 -9552 781
rect -9518 747 -9484 781
rect -9450 747 -9416 781
rect -8908 747 -8874 781
rect -8840 747 -8806 781
rect -8772 747 -8738 781
rect -8704 747 -8670 781
rect -8636 747 -8602 781
rect -8568 747 -8534 781
rect -8500 747 -8466 781
rect -8432 747 -8398 781
rect -7890 747 -7856 781
rect -7822 747 -7788 781
rect -7754 747 -7720 781
rect -7686 747 -7652 781
rect -7618 747 -7584 781
rect -7550 747 -7516 781
rect -7482 747 -7448 781
rect -7414 747 -7380 781
rect -6872 747 -6838 781
rect -6804 747 -6770 781
rect -6736 747 -6702 781
rect -6668 747 -6634 781
rect -6600 747 -6566 781
rect -6532 747 -6498 781
rect -6464 747 -6430 781
rect -6396 747 -6362 781
rect -5854 747 -5820 781
rect -5786 747 -5752 781
rect -5718 747 -5684 781
rect -5650 747 -5616 781
rect -5582 747 -5548 781
rect -5514 747 -5480 781
rect -5446 747 -5412 781
rect -5378 747 -5344 781
rect -4836 747 -4802 781
rect -4768 747 -4734 781
rect -4700 747 -4666 781
rect -4632 747 -4598 781
rect -4564 747 -4530 781
rect -4496 747 -4462 781
rect -4428 747 -4394 781
rect -4360 747 -4326 781
rect -3818 747 -3784 781
rect -3750 747 -3716 781
rect -3682 747 -3648 781
rect -3614 747 -3580 781
rect -3546 747 -3512 781
rect -3478 747 -3444 781
rect -3410 747 -3376 781
rect -3342 747 -3308 781
rect -2800 747 -2766 781
rect -2732 747 -2698 781
rect -2664 747 -2630 781
rect -2596 747 -2562 781
rect -2528 747 -2494 781
rect -2460 747 -2426 781
rect -2392 747 -2358 781
rect -2324 747 -2290 781
rect -1782 747 -1748 781
rect -1714 747 -1680 781
rect -1646 747 -1612 781
rect -1578 747 -1544 781
rect -1510 747 -1476 781
rect -1442 747 -1408 781
rect -1374 747 -1340 781
rect -1306 747 -1272 781
rect -764 747 -730 781
rect -696 747 -662 781
rect -628 747 -594 781
rect -560 747 -526 781
rect -492 747 -458 781
rect -424 747 -390 781
rect -356 747 -322 781
rect -288 747 -254 781
rect 254 747 288 781
rect 322 747 356 781
rect 390 747 424 781
rect 458 747 492 781
rect 526 747 560 781
rect 594 747 628 781
rect 662 747 696 781
rect 730 747 764 781
rect 1272 747 1306 781
rect 1340 747 1374 781
rect 1408 747 1442 781
rect 1476 747 1510 781
rect 1544 747 1578 781
rect 1612 747 1646 781
rect 1680 747 1714 781
rect 1748 747 1782 781
rect 2290 747 2324 781
rect 2358 747 2392 781
rect 2426 747 2460 781
rect 2494 747 2528 781
rect 2562 747 2596 781
rect 2630 747 2664 781
rect 2698 747 2732 781
rect 2766 747 2800 781
rect 3308 747 3342 781
rect 3376 747 3410 781
rect 3444 747 3478 781
rect 3512 747 3546 781
rect 3580 747 3614 781
rect 3648 747 3682 781
rect 3716 747 3750 781
rect 3784 747 3818 781
rect 4326 747 4360 781
rect 4394 747 4428 781
rect 4462 747 4496 781
rect 4530 747 4564 781
rect 4598 747 4632 781
rect 4666 747 4700 781
rect 4734 747 4768 781
rect 4802 747 4836 781
rect 5344 747 5378 781
rect 5412 747 5446 781
rect 5480 747 5514 781
rect 5548 747 5582 781
rect 5616 747 5650 781
rect 5684 747 5718 781
rect 5752 747 5786 781
rect 5820 747 5854 781
rect 6362 747 6396 781
rect 6430 747 6464 781
rect 6498 747 6532 781
rect 6566 747 6600 781
rect 6634 747 6668 781
rect 6702 747 6736 781
rect 6770 747 6804 781
rect 6838 747 6872 781
rect 7380 747 7414 781
rect 7448 747 7482 781
rect 7516 747 7550 781
rect 7584 747 7618 781
rect 7652 747 7686 781
rect 7720 747 7754 781
rect 7788 747 7822 781
rect 7856 747 7890 781
rect 8398 747 8432 781
rect 8466 747 8500 781
rect 8534 747 8568 781
rect 8602 747 8636 781
rect 8670 747 8704 781
rect 8738 747 8772 781
rect 8806 747 8840 781
rect 8874 747 8908 781
rect 9416 747 9450 781
rect 9484 747 9518 781
rect 9552 747 9586 781
rect 9620 747 9654 781
rect 9688 747 9722 781
rect 9756 747 9790 781
rect 9824 747 9858 781
rect 9892 747 9926 781
rect -9926 37 -9892 71
rect -9858 37 -9824 71
rect -9790 37 -9756 71
rect -9722 37 -9688 71
rect -9654 37 -9620 71
rect -9586 37 -9552 71
rect -9518 37 -9484 71
rect -9450 37 -9416 71
rect -8908 37 -8874 71
rect -8840 37 -8806 71
rect -8772 37 -8738 71
rect -8704 37 -8670 71
rect -8636 37 -8602 71
rect -8568 37 -8534 71
rect -8500 37 -8466 71
rect -8432 37 -8398 71
rect -7890 37 -7856 71
rect -7822 37 -7788 71
rect -7754 37 -7720 71
rect -7686 37 -7652 71
rect -7618 37 -7584 71
rect -7550 37 -7516 71
rect -7482 37 -7448 71
rect -7414 37 -7380 71
rect -6872 37 -6838 71
rect -6804 37 -6770 71
rect -6736 37 -6702 71
rect -6668 37 -6634 71
rect -6600 37 -6566 71
rect -6532 37 -6498 71
rect -6464 37 -6430 71
rect -6396 37 -6362 71
rect -5854 37 -5820 71
rect -5786 37 -5752 71
rect -5718 37 -5684 71
rect -5650 37 -5616 71
rect -5582 37 -5548 71
rect -5514 37 -5480 71
rect -5446 37 -5412 71
rect -5378 37 -5344 71
rect -4836 37 -4802 71
rect -4768 37 -4734 71
rect -4700 37 -4666 71
rect -4632 37 -4598 71
rect -4564 37 -4530 71
rect -4496 37 -4462 71
rect -4428 37 -4394 71
rect -4360 37 -4326 71
rect -3818 37 -3784 71
rect -3750 37 -3716 71
rect -3682 37 -3648 71
rect -3614 37 -3580 71
rect -3546 37 -3512 71
rect -3478 37 -3444 71
rect -3410 37 -3376 71
rect -3342 37 -3308 71
rect -2800 37 -2766 71
rect -2732 37 -2698 71
rect -2664 37 -2630 71
rect -2596 37 -2562 71
rect -2528 37 -2494 71
rect -2460 37 -2426 71
rect -2392 37 -2358 71
rect -2324 37 -2290 71
rect -1782 37 -1748 71
rect -1714 37 -1680 71
rect -1646 37 -1612 71
rect -1578 37 -1544 71
rect -1510 37 -1476 71
rect -1442 37 -1408 71
rect -1374 37 -1340 71
rect -1306 37 -1272 71
rect -764 37 -730 71
rect -696 37 -662 71
rect -628 37 -594 71
rect -560 37 -526 71
rect -492 37 -458 71
rect -424 37 -390 71
rect -356 37 -322 71
rect -288 37 -254 71
rect 254 37 288 71
rect 322 37 356 71
rect 390 37 424 71
rect 458 37 492 71
rect 526 37 560 71
rect 594 37 628 71
rect 662 37 696 71
rect 730 37 764 71
rect 1272 37 1306 71
rect 1340 37 1374 71
rect 1408 37 1442 71
rect 1476 37 1510 71
rect 1544 37 1578 71
rect 1612 37 1646 71
rect 1680 37 1714 71
rect 1748 37 1782 71
rect 2290 37 2324 71
rect 2358 37 2392 71
rect 2426 37 2460 71
rect 2494 37 2528 71
rect 2562 37 2596 71
rect 2630 37 2664 71
rect 2698 37 2732 71
rect 2766 37 2800 71
rect 3308 37 3342 71
rect 3376 37 3410 71
rect 3444 37 3478 71
rect 3512 37 3546 71
rect 3580 37 3614 71
rect 3648 37 3682 71
rect 3716 37 3750 71
rect 3784 37 3818 71
rect 4326 37 4360 71
rect 4394 37 4428 71
rect 4462 37 4496 71
rect 4530 37 4564 71
rect 4598 37 4632 71
rect 4666 37 4700 71
rect 4734 37 4768 71
rect 4802 37 4836 71
rect 5344 37 5378 71
rect 5412 37 5446 71
rect 5480 37 5514 71
rect 5548 37 5582 71
rect 5616 37 5650 71
rect 5684 37 5718 71
rect 5752 37 5786 71
rect 5820 37 5854 71
rect 6362 37 6396 71
rect 6430 37 6464 71
rect 6498 37 6532 71
rect 6566 37 6600 71
rect 6634 37 6668 71
rect 6702 37 6736 71
rect 6770 37 6804 71
rect 6838 37 6872 71
rect 7380 37 7414 71
rect 7448 37 7482 71
rect 7516 37 7550 71
rect 7584 37 7618 71
rect 7652 37 7686 71
rect 7720 37 7754 71
rect 7788 37 7822 71
rect 7856 37 7890 71
rect 8398 37 8432 71
rect 8466 37 8500 71
rect 8534 37 8568 71
rect 8602 37 8636 71
rect 8670 37 8704 71
rect 8738 37 8772 71
rect 8806 37 8840 71
rect 8874 37 8908 71
rect 9416 37 9450 71
rect 9484 37 9518 71
rect 9552 37 9586 71
rect 9620 37 9654 71
rect 9688 37 9722 71
rect 9756 37 9790 71
rect 9824 37 9858 71
rect 9892 37 9926 71
rect -9926 -71 -9892 -37
rect -9858 -71 -9824 -37
rect -9790 -71 -9756 -37
rect -9722 -71 -9688 -37
rect -9654 -71 -9620 -37
rect -9586 -71 -9552 -37
rect -9518 -71 -9484 -37
rect -9450 -71 -9416 -37
rect -8908 -71 -8874 -37
rect -8840 -71 -8806 -37
rect -8772 -71 -8738 -37
rect -8704 -71 -8670 -37
rect -8636 -71 -8602 -37
rect -8568 -71 -8534 -37
rect -8500 -71 -8466 -37
rect -8432 -71 -8398 -37
rect -7890 -71 -7856 -37
rect -7822 -71 -7788 -37
rect -7754 -71 -7720 -37
rect -7686 -71 -7652 -37
rect -7618 -71 -7584 -37
rect -7550 -71 -7516 -37
rect -7482 -71 -7448 -37
rect -7414 -71 -7380 -37
rect -6872 -71 -6838 -37
rect -6804 -71 -6770 -37
rect -6736 -71 -6702 -37
rect -6668 -71 -6634 -37
rect -6600 -71 -6566 -37
rect -6532 -71 -6498 -37
rect -6464 -71 -6430 -37
rect -6396 -71 -6362 -37
rect -5854 -71 -5820 -37
rect -5786 -71 -5752 -37
rect -5718 -71 -5684 -37
rect -5650 -71 -5616 -37
rect -5582 -71 -5548 -37
rect -5514 -71 -5480 -37
rect -5446 -71 -5412 -37
rect -5378 -71 -5344 -37
rect -4836 -71 -4802 -37
rect -4768 -71 -4734 -37
rect -4700 -71 -4666 -37
rect -4632 -71 -4598 -37
rect -4564 -71 -4530 -37
rect -4496 -71 -4462 -37
rect -4428 -71 -4394 -37
rect -4360 -71 -4326 -37
rect -3818 -71 -3784 -37
rect -3750 -71 -3716 -37
rect -3682 -71 -3648 -37
rect -3614 -71 -3580 -37
rect -3546 -71 -3512 -37
rect -3478 -71 -3444 -37
rect -3410 -71 -3376 -37
rect -3342 -71 -3308 -37
rect -2800 -71 -2766 -37
rect -2732 -71 -2698 -37
rect -2664 -71 -2630 -37
rect -2596 -71 -2562 -37
rect -2528 -71 -2494 -37
rect -2460 -71 -2426 -37
rect -2392 -71 -2358 -37
rect -2324 -71 -2290 -37
rect -1782 -71 -1748 -37
rect -1714 -71 -1680 -37
rect -1646 -71 -1612 -37
rect -1578 -71 -1544 -37
rect -1510 -71 -1476 -37
rect -1442 -71 -1408 -37
rect -1374 -71 -1340 -37
rect -1306 -71 -1272 -37
rect -764 -71 -730 -37
rect -696 -71 -662 -37
rect -628 -71 -594 -37
rect -560 -71 -526 -37
rect -492 -71 -458 -37
rect -424 -71 -390 -37
rect -356 -71 -322 -37
rect -288 -71 -254 -37
rect 254 -71 288 -37
rect 322 -71 356 -37
rect 390 -71 424 -37
rect 458 -71 492 -37
rect 526 -71 560 -37
rect 594 -71 628 -37
rect 662 -71 696 -37
rect 730 -71 764 -37
rect 1272 -71 1306 -37
rect 1340 -71 1374 -37
rect 1408 -71 1442 -37
rect 1476 -71 1510 -37
rect 1544 -71 1578 -37
rect 1612 -71 1646 -37
rect 1680 -71 1714 -37
rect 1748 -71 1782 -37
rect 2290 -71 2324 -37
rect 2358 -71 2392 -37
rect 2426 -71 2460 -37
rect 2494 -71 2528 -37
rect 2562 -71 2596 -37
rect 2630 -71 2664 -37
rect 2698 -71 2732 -37
rect 2766 -71 2800 -37
rect 3308 -71 3342 -37
rect 3376 -71 3410 -37
rect 3444 -71 3478 -37
rect 3512 -71 3546 -37
rect 3580 -71 3614 -37
rect 3648 -71 3682 -37
rect 3716 -71 3750 -37
rect 3784 -71 3818 -37
rect 4326 -71 4360 -37
rect 4394 -71 4428 -37
rect 4462 -71 4496 -37
rect 4530 -71 4564 -37
rect 4598 -71 4632 -37
rect 4666 -71 4700 -37
rect 4734 -71 4768 -37
rect 4802 -71 4836 -37
rect 5344 -71 5378 -37
rect 5412 -71 5446 -37
rect 5480 -71 5514 -37
rect 5548 -71 5582 -37
rect 5616 -71 5650 -37
rect 5684 -71 5718 -37
rect 5752 -71 5786 -37
rect 5820 -71 5854 -37
rect 6362 -71 6396 -37
rect 6430 -71 6464 -37
rect 6498 -71 6532 -37
rect 6566 -71 6600 -37
rect 6634 -71 6668 -37
rect 6702 -71 6736 -37
rect 6770 -71 6804 -37
rect 6838 -71 6872 -37
rect 7380 -71 7414 -37
rect 7448 -71 7482 -37
rect 7516 -71 7550 -37
rect 7584 -71 7618 -37
rect 7652 -71 7686 -37
rect 7720 -71 7754 -37
rect 7788 -71 7822 -37
rect 7856 -71 7890 -37
rect 8398 -71 8432 -37
rect 8466 -71 8500 -37
rect 8534 -71 8568 -37
rect 8602 -71 8636 -37
rect 8670 -71 8704 -37
rect 8738 -71 8772 -37
rect 8806 -71 8840 -37
rect 8874 -71 8908 -37
rect 9416 -71 9450 -37
rect 9484 -71 9518 -37
rect 9552 -71 9586 -37
rect 9620 -71 9654 -37
rect 9688 -71 9722 -37
rect 9756 -71 9790 -37
rect 9824 -71 9858 -37
rect 9892 -71 9926 -37
rect -9926 -781 -9892 -747
rect -9858 -781 -9824 -747
rect -9790 -781 -9756 -747
rect -9722 -781 -9688 -747
rect -9654 -781 -9620 -747
rect -9586 -781 -9552 -747
rect -9518 -781 -9484 -747
rect -9450 -781 -9416 -747
rect -8908 -781 -8874 -747
rect -8840 -781 -8806 -747
rect -8772 -781 -8738 -747
rect -8704 -781 -8670 -747
rect -8636 -781 -8602 -747
rect -8568 -781 -8534 -747
rect -8500 -781 -8466 -747
rect -8432 -781 -8398 -747
rect -7890 -781 -7856 -747
rect -7822 -781 -7788 -747
rect -7754 -781 -7720 -747
rect -7686 -781 -7652 -747
rect -7618 -781 -7584 -747
rect -7550 -781 -7516 -747
rect -7482 -781 -7448 -747
rect -7414 -781 -7380 -747
rect -6872 -781 -6838 -747
rect -6804 -781 -6770 -747
rect -6736 -781 -6702 -747
rect -6668 -781 -6634 -747
rect -6600 -781 -6566 -747
rect -6532 -781 -6498 -747
rect -6464 -781 -6430 -747
rect -6396 -781 -6362 -747
rect -5854 -781 -5820 -747
rect -5786 -781 -5752 -747
rect -5718 -781 -5684 -747
rect -5650 -781 -5616 -747
rect -5582 -781 -5548 -747
rect -5514 -781 -5480 -747
rect -5446 -781 -5412 -747
rect -5378 -781 -5344 -747
rect -4836 -781 -4802 -747
rect -4768 -781 -4734 -747
rect -4700 -781 -4666 -747
rect -4632 -781 -4598 -747
rect -4564 -781 -4530 -747
rect -4496 -781 -4462 -747
rect -4428 -781 -4394 -747
rect -4360 -781 -4326 -747
rect -3818 -781 -3784 -747
rect -3750 -781 -3716 -747
rect -3682 -781 -3648 -747
rect -3614 -781 -3580 -747
rect -3546 -781 -3512 -747
rect -3478 -781 -3444 -747
rect -3410 -781 -3376 -747
rect -3342 -781 -3308 -747
rect -2800 -781 -2766 -747
rect -2732 -781 -2698 -747
rect -2664 -781 -2630 -747
rect -2596 -781 -2562 -747
rect -2528 -781 -2494 -747
rect -2460 -781 -2426 -747
rect -2392 -781 -2358 -747
rect -2324 -781 -2290 -747
rect -1782 -781 -1748 -747
rect -1714 -781 -1680 -747
rect -1646 -781 -1612 -747
rect -1578 -781 -1544 -747
rect -1510 -781 -1476 -747
rect -1442 -781 -1408 -747
rect -1374 -781 -1340 -747
rect -1306 -781 -1272 -747
rect -764 -781 -730 -747
rect -696 -781 -662 -747
rect -628 -781 -594 -747
rect -560 -781 -526 -747
rect -492 -781 -458 -747
rect -424 -781 -390 -747
rect -356 -781 -322 -747
rect -288 -781 -254 -747
rect 254 -781 288 -747
rect 322 -781 356 -747
rect 390 -781 424 -747
rect 458 -781 492 -747
rect 526 -781 560 -747
rect 594 -781 628 -747
rect 662 -781 696 -747
rect 730 -781 764 -747
rect 1272 -781 1306 -747
rect 1340 -781 1374 -747
rect 1408 -781 1442 -747
rect 1476 -781 1510 -747
rect 1544 -781 1578 -747
rect 1612 -781 1646 -747
rect 1680 -781 1714 -747
rect 1748 -781 1782 -747
rect 2290 -781 2324 -747
rect 2358 -781 2392 -747
rect 2426 -781 2460 -747
rect 2494 -781 2528 -747
rect 2562 -781 2596 -747
rect 2630 -781 2664 -747
rect 2698 -781 2732 -747
rect 2766 -781 2800 -747
rect 3308 -781 3342 -747
rect 3376 -781 3410 -747
rect 3444 -781 3478 -747
rect 3512 -781 3546 -747
rect 3580 -781 3614 -747
rect 3648 -781 3682 -747
rect 3716 -781 3750 -747
rect 3784 -781 3818 -747
rect 4326 -781 4360 -747
rect 4394 -781 4428 -747
rect 4462 -781 4496 -747
rect 4530 -781 4564 -747
rect 4598 -781 4632 -747
rect 4666 -781 4700 -747
rect 4734 -781 4768 -747
rect 4802 -781 4836 -747
rect 5344 -781 5378 -747
rect 5412 -781 5446 -747
rect 5480 -781 5514 -747
rect 5548 -781 5582 -747
rect 5616 -781 5650 -747
rect 5684 -781 5718 -747
rect 5752 -781 5786 -747
rect 5820 -781 5854 -747
rect 6362 -781 6396 -747
rect 6430 -781 6464 -747
rect 6498 -781 6532 -747
rect 6566 -781 6600 -747
rect 6634 -781 6668 -747
rect 6702 -781 6736 -747
rect 6770 -781 6804 -747
rect 6838 -781 6872 -747
rect 7380 -781 7414 -747
rect 7448 -781 7482 -747
rect 7516 -781 7550 -747
rect 7584 -781 7618 -747
rect 7652 -781 7686 -747
rect 7720 -781 7754 -747
rect 7788 -781 7822 -747
rect 7856 -781 7890 -747
rect 8398 -781 8432 -747
rect 8466 -781 8500 -747
rect 8534 -781 8568 -747
rect 8602 -781 8636 -747
rect 8670 -781 8704 -747
rect 8738 -781 8772 -747
rect 8806 -781 8840 -747
rect 8874 -781 8908 -747
rect 9416 -781 9450 -747
rect 9484 -781 9518 -747
rect 9552 -781 9586 -747
rect 9620 -781 9654 -747
rect 9688 -781 9722 -747
rect 9756 -781 9790 -747
rect 9824 -781 9858 -747
rect 9892 -781 9926 -747
<< locali >>
rect -9965 747 -9926 781
rect -9892 747 -9868 781
rect -9824 747 -9796 781
rect -9756 747 -9724 781
rect -9688 747 -9654 781
rect -9618 747 -9586 781
rect -9546 747 -9518 781
rect -9474 747 -9450 781
rect -9416 747 -9377 781
rect -8947 747 -8908 781
rect -8874 747 -8850 781
rect -8806 747 -8778 781
rect -8738 747 -8706 781
rect -8670 747 -8636 781
rect -8600 747 -8568 781
rect -8528 747 -8500 781
rect -8456 747 -8432 781
rect -8398 747 -8359 781
rect -7929 747 -7890 781
rect -7856 747 -7832 781
rect -7788 747 -7760 781
rect -7720 747 -7688 781
rect -7652 747 -7618 781
rect -7582 747 -7550 781
rect -7510 747 -7482 781
rect -7438 747 -7414 781
rect -7380 747 -7341 781
rect -6911 747 -6872 781
rect -6838 747 -6814 781
rect -6770 747 -6742 781
rect -6702 747 -6670 781
rect -6634 747 -6600 781
rect -6564 747 -6532 781
rect -6492 747 -6464 781
rect -6420 747 -6396 781
rect -6362 747 -6323 781
rect -5893 747 -5854 781
rect -5820 747 -5796 781
rect -5752 747 -5724 781
rect -5684 747 -5652 781
rect -5616 747 -5582 781
rect -5546 747 -5514 781
rect -5474 747 -5446 781
rect -5402 747 -5378 781
rect -5344 747 -5305 781
rect -4875 747 -4836 781
rect -4802 747 -4778 781
rect -4734 747 -4706 781
rect -4666 747 -4634 781
rect -4598 747 -4564 781
rect -4528 747 -4496 781
rect -4456 747 -4428 781
rect -4384 747 -4360 781
rect -4326 747 -4287 781
rect -3857 747 -3818 781
rect -3784 747 -3760 781
rect -3716 747 -3688 781
rect -3648 747 -3616 781
rect -3580 747 -3546 781
rect -3510 747 -3478 781
rect -3438 747 -3410 781
rect -3366 747 -3342 781
rect -3308 747 -3269 781
rect -2839 747 -2800 781
rect -2766 747 -2742 781
rect -2698 747 -2670 781
rect -2630 747 -2598 781
rect -2562 747 -2528 781
rect -2492 747 -2460 781
rect -2420 747 -2392 781
rect -2348 747 -2324 781
rect -2290 747 -2251 781
rect -1821 747 -1782 781
rect -1748 747 -1724 781
rect -1680 747 -1652 781
rect -1612 747 -1580 781
rect -1544 747 -1510 781
rect -1474 747 -1442 781
rect -1402 747 -1374 781
rect -1330 747 -1306 781
rect -1272 747 -1233 781
rect -803 747 -764 781
rect -730 747 -706 781
rect -662 747 -634 781
rect -594 747 -562 781
rect -526 747 -492 781
rect -456 747 -424 781
rect -384 747 -356 781
rect -312 747 -288 781
rect -254 747 -215 781
rect 215 747 254 781
rect 288 747 312 781
rect 356 747 384 781
rect 424 747 456 781
rect 492 747 526 781
rect 562 747 594 781
rect 634 747 662 781
rect 706 747 730 781
rect 764 747 803 781
rect 1233 747 1272 781
rect 1306 747 1330 781
rect 1374 747 1402 781
rect 1442 747 1474 781
rect 1510 747 1544 781
rect 1580 747 1612 781
rect 1652 747 1680 781
rect 1724 747 1748 781
rect 1782 747 1821 781
rect 2251 747 2290 781
rect 2324 747 2348 781
rect 2392 747 2420 781
rect 2460 747 2492 781
rect 2528 747 2562 781
rect 2598 747 2630 781
rect 2670 747 2698 781
rect 2742 747 2766 781
rect 2800 747 2839 781
rect 3269 747 3308 781
rect 3342 747 3366 781
rect 3410 747 3438 781
rect 3478 747 3510 781
rect 3546 747 3580 781
rect 3616 747 3648 781
rect 3688 747 3716 781
rect 3760 747 3784 781
rect 3818 747 3857 781
rect 4287 747 4326 781
rect 4360 747 4384 781
rect 4428 747 4456 781
rect 4496 747 4528 781
rect 4564 747 4598 781
rect 4634 747 4666 781
rect 4706 747 4734 781
rect 4778 747 4802 781
rect 4836 747 4875 781
rect 5305 747 5344 781
rect 5378 747 5402 781
rect 5446 747 5474 781
rect 5514 747 5546 781
rect 5582 747 5616 781
rect 5652 747 5684 781
rect 5724 747 5752 781
rect 5796 747 5820 781
rect 5854 747 5893 781
rect 6323 747 6362 781
rect 6396 747 6420 781
rect 6464 747 6492 781
rect 6532 747 6564 781
rect 6600 747 6634 781
rect 6670 747 6702 781
rect 6742 747 6770 781
rect 6814 747 6838 781
rect 6872 747 6911 781
rect 7341 747 7380 781
rect 7414 747 7438 781
rect 7482 747 7510 781
rect 7550 747 7582 781
rect 7618 747 7652 781
rect 7688 747 7720 781
rect 7760 747 7788 781
rect 7832 747 7856 781
rect 7890 747 7929 781
rect 8359 747 8398 781
rect 8432 747 8456 781
rect 8500 747 8528 781
rect 8568 747 8600 781
rect 8636 747 8670 781
rect 8706 747 8738 781
rect 8778 747 8806 781
rect 8850 747 8874 781
rect 8908 747 8947 781
rect 9377 747 9416 781
rect 9450 747 9474 781
rect 9518 747 9546 781
rect 9586 747 9618 781
rect 9654 747 9688 781
rect 9724 747 9756 781
rect 9796 747 9824 781
rect 9868 747 9892 781
rect 9926 747 9965 781
rect -10197 678 -10163 713
rect -10197 606 -10163 630
rect -10197 534 -10163 562
rect -10197 462 -10163 494
rect -10197 392 -10163 426
rect -10197 324 -10163 356
rect -10197 256 -10163 284
rect -10197 188 -10163 212
rect -10197 105 -10163 140
rect -9179 678 -9145 713
rect -9179 606 -9145 630
rect -9179 534 -9145 562
rect -9179 462 -9145 494
rect -9179 392 -9145 426
rect -9179 324 -9145 356
rect -9179 256 -9145 284
rect -9179 188 -9145 212
rect -9179 105 -9145 140
rect -8161 678 -8127 713
rect -8161 606 -8127 630
rect -8161 534 -8127 562
rect -8161 462 -8127 494
rect -8161 392 -8127 426
rect -8161 324 -8127 356
rect -8161 256 -8127 284
rect -8161 188 -8127 212
rect -8161 105 -8127 140
rect -7143 678 -7109 713
rect -7143 606 -7109 630
rect -7143 534 -7109 562
rect -7143 462 -7109 494
rect -7143 392 -7109 426
rect -7143 324 -7109 356
rect -7143 256 -7109 284
rect -7143 188 -7109 212
rect -7143 105 -7109 140
rect -6125 678 -6091 713
rect -6125 606 -6091 630
rect -6125 534 -6091 562
rect -6125 462 -6091 494
rect -6125 392 -6091 426
rect -6125 324 -6091 356
rect -6125 256 -6091 284
rect -6125 188 -6091 212
rect -6125 105 -6091 140
rect -5107 678 -5073 713
rect -5107 606 -5073 630
rect -5107 534 -5073 562
rect -5107 462 -5073 494
rect -5107 392 -5073 426
rect -5107 324 -5073 356
rect -5107 256 -5073 284
rect -5107 188 -5073 212
rect -5107 105 -5073 140
rect -4089 678 -4055 713
rect -4089 606 -4055 630
rect -4089 534 -4055 562
rect -4089 462 -4055 494
rect -4089 392 -4055 426
rect -4089 324 -4055 356
rect -4089 256 -4055 284
rect -4089 188 -4055 212
rect -4089 105 -4055 140
rect -3071 678 -3037 713
rect -3071 606 -3037 630
rect -3071 534 -3037 562
rect -3071 462 -3037 494
rect -3071 392 -3037 426
rect -3071 324 -3037 356
rect -3071 256 -3037 284
rect -3071 188 -3037 212
rect -3071 105 -3037 140
rect -2053 678 -2019 713
rect -2053 606 -2019 630
rect -2053 534 -2019 562
rect -2053 462 -2019 494
rect -2053 392 -2019 426
rect -2053 324 -2019 356
rect -2053 256 -2019 284
rect -2053 188 -2019 212
rect -2053 105 -2019 140
rect -1035 678 -1001 713
rect -1035 606 -1001 630
rect -1035 534 -1001 562
rect -1035 462 -1001 494
rect -1035 392 -1001 426
rect -1035 324 -1001 356
rect -1035 256 -1001 284
rect -1035 188 -1001 212
rect -1035 105 -1001 140
rect -17 678 17 713
rect -17 606 17 630
rect -17 534 17 562
rect -17 462 17 494
rect -17 392 17 426
rect -17 324 17 356
rect -17 256 17 284
rect -17 188 17 212
rect -17 105 17 140
rect 1001 678 1035 713
rect 1001 606 1035 630
rect 1001 534 1035 562
rect 1001 462 1035 494
rect 1001 392 1035 426
rect 1001 324 1035 356
rect 1001 256 1035 284
rect 1001 188 1035 212
rect 1001 105 1035 140
rect 2019 678 2053 713
rect 2019 606 2053 630
rect 2019 534 2053 562
rect 2019 462 2053 494
rect 2019 392 2053 426
rect 2019 324 2053 356
rect 2019 256 2053 284
rect 2019 188 2053 212
rect 2019 105 2053 140
rect 3037 678 3071 713
rect 3037 606 3071 630
rect 3037 534 3071 562
rect 3037 462 3071 494
rect 3037 392 3071 426
rect 3037 324 3071 356
rect 3037 256 3071 284
rect 3037 188 3071 212
rect 3037 105 3071 140
rect 4055 678 4089 713
rect 4055 606 4089 630
rect 4055 534 4089 562
rect 4055 462 4089 494
rect 4055 392 4089 426
rect 4055 324 4089 356
rect 4055 256 4089 284
rect 4055 188 4089 212
rect 4055 105 4089 140
rect 5073 678 5107 713
rect 5073 606 5107 630
rect 5073 534 5107 562
rect 5073 462 5107 494
rect 5073 392 5107 426
rect 5073 324 5107 356
rect 5073 256 5107 284
rect 5073 188 5107 212
rect 5073 105 5107 140
rect 6091 678 6125 713
rect 6091 606 6125 630
rect 6091 534 6125 562
rect 6091 462 6125 494
rect 6091 392 6125 426
rect 6091 324 6125 356
rect 6091 256 6125 284
rect 6091 188 6125 212
rect 6091 105 6125 140
rect 7109 678 7143 713
rect 7109 606 7143 630
rect 7109 534 7143 562
rect 7109 462 7143 494
rect 7109 392 7143 426
rect 7109 324 7143 356
rect 7109 256 7143 284
rect 7109 188 7143 212
rect 7109 105 7143 140
rect 8127 678 8161 713
rect 8127 606 8161 630
rect 8127 534 8161 562
rect 8127 462 8161 494
rect 8127 392 8161 426
rect 8127 324 8161 356
rect 8127 256 8161 284
rect 8127 188 8161 212
rect 8127 105 8161 140
rect 9145 678 9179 713
rect 9145 606 9179 630
rect 9145 534 9179 562
rect 9145 462 9179 494
rect 9145 392 9179 426
rect 9145 324 9179 356
rect 9145 256 9179 284
rect 9145 188 9179 212
rect 9145 105 9179 140
rect 10163 678 10197 713
rect 10163 606 10197 630
rect 10163 534 10197 562
rect 10163 462 10197 494
rect 10163 392 10197 426
rect 10163 324 10197 356
rect 10163 256 10197 284
rect 10163 188 10197 212
rect 10163 105 10197 140
rect -9965 37 -9926 71
rect -9892 37 -9868 71
rect -9824 37 -9796 71
rect -9756 37 -9724 71
rect -9688 37 -9654 71
rect -9618 37 -9586 71
rect -9546 37 -9518 71
rect -9474 37 -9450 71
rect -9416 37 -9377 71
rect -8947 37 -8908 71
rect -8874 37 -8850 71
rect -8806 37 -8778 71
rect -8738 37 -8706 71
rect -8670 37 -8636 71
rect -8600 37 -8568 71
rect -8528 37 -8500 71
rect -8456 37 -8432 71
rect -8398 37 -8359 71
rect -7929 37 -7890 71
rect -7856 37 -7832 71
rect -7788 37 -7760 71
rect -7720 37 -7688 71
rect -7652 37 -7618 71
rect -7582 37 -7550 71
rect -7510 37 -7482 71
rect -7438 37 -7414 71
rect -7380 37 -7341 71
rect -6911 37 -6872 71
rect -6838 37 -6814 71
rect -6770 37 -6742 71
rect -6702 37 -6670 71
rect -6634 37 -6600 71
rect -6564 37 -6532 71
rect -6492 37 -6464 71
rect -6420 37 -6396 71
rect -6362 37 -6323 71
rect -5893 37 -5854 71
rect -5820 37 -5796 71
rect -5752 37 -5724 71
rect -5684 37 -5652 71
rect -5616 37 -5582 71
rect -5546 37 -5514 71
rect -5474 37 -5446 71
rect -5402 37 -5378 71
rect -5344 37 -5305 71
rect -4875 37 -4836 71
rect -4802 37 -4778 71
rect -4734 37 -4706 71
rect -4666 37 -4634 71
rect -4598 37 -4564 71
rect -4528 37 -4496 71
rect -4456 37 -4428 71
rect -4384 37 -4360 71
rect -4326 37 -4287 71
rect -3857 37 -3818 71
rect -3784 37 -3760 71
rect -3716 37 -3688 71
rect -3648 37 -3616 71
rect -3580 37 -3546 71
rect -3510 37 -3478 71
rect -3438 37 -3410 71
rect -3366 37 -3342 71
rect -3308 37 -3269 71
rect -2839 37 -2800 71
rect -2766 37 -2742 71
rect -2698 37 -2670 71
rect -2630 37 -2598 71
rect -2562 37 -2528 71
rect -2492 37 -2460 71
rect -2420 37 -2392 71
rect -2348 37 -2324 71
rect -2290 37 -2251 71
rect -1821 37 -1782 71
rect -1748 37 -1724 71
rect -1680 37 -1652 71
rect -1612 37 -1580 71
rect -1544 37 -1510 71
rect -1474 37 -1442 71
rect -1402 37 -1374 71
rect -1330 37 -1306 71
rect -1272 37 -1233 71
rect -803 37 -764 71
rect -730 37 -706 71
rect -662 37 -634 71
rect -594 37 -562 71
rect -526 37 -492 71
rect -456 37 -424 71
rect -384 37 -356 71
rect -312 37 -288 71
rect -254 37 -215 71
rect 215 37 254 71
rect 288 37 312 71
rect 356 37 384 71
rect 424 37 456 71
rect 492 37 526 71
rect 562 37 594 71
rect 634 37 662 71
rect 706 37 730 71
rect 764 37 803 71
rect 1233 37 1272 71
rect 1306 37 1330 71
rect 1374 37 1402 71
rect 1442 37 1474 71
rect 1510 37 1544 71
rect 1580 37 1612 71
rect 1652 37 1680 71
rect 1724 37 1748 71
rect 1782 37 1821 71
rect 2251 37 2290 71
rect 2324 37 2348 71
rect 2392 37 2420 71
rect 2460 37 2492 71
rect 2528 37 2562 71
rect 2598 37 2630 71
rect 2670 37 2698 71
rect 2742 37 2766 71
rect 2800 37 2839 71
rect 3269 37 3308 71
rect 3342 37 3366 71
rect 3410 37 3438 71
rect 3478 37 3510 71
rect 3546 37 3580 71
rect 3616 37 3648 71
rect 3688 37 3716 71
rect 3760 37 3784 71
rect 3818 37 3857 71
rect 4287 37 4326 71
rect 4360 37 4384 71
rect 4428 37 4456 71
rect 4496 37 4528 71
rect 4564 37 4598 71
rect 4634 37 4666 71
rect 4706 37 4734 71
rect 4778 37 4802 71
rect 4836 37 4875 71
rect 5305 37 5344 71
rect 5378 37 5402 71
rect 5446 37 5474 71
rect 5514 37 5546 71
rect 5582 37 5616 71
rect 5652 37 5684 71
rect 5724 37 5752 71
rect 5796 37 5820 71
rect 5854 37 5893 71
rect 6323 37 6362 71
rect 6396 37 6420 71
rect 6464 37 6492 71
rect 6532 37 6564 71
rect 6600 37 6634 71
rect 6670 37 6702 71
rect 6742 37 6770 71
rect 6814 37 6838 71
rect 6872 37 6911 71
rect 7341 37 7380 71
rect 7414 37 7438 71
rect 7482 37 7510 71
rect 7550 37 7582 71
rect 7618 37 7652 71
rect 7688 37 7720 71
rect 7760 37 7788 71
rect 7832 37 7856 71
rect 7890 37 7929 71
rect 8359 37 8398 71
rect 8432 37 8456 71
rect 8500 37 8528 71
rect 8568 37 8600 71
rect 8636 37 8670 71
rect 8706 37 8738 71
rect 8778 37 8806 71
rect 8850 37 8874 71
rect 8908 37 8947 71
rect 9377 37 9416 71
rect 9450 37 9474 71
rect 9518 37 9546 71
rect 9586 37 9618 71
rect 9654 37 9688 71
rect 9724 37 9756 71
rect 9796 37 9824 71
rect 9868 37 9892 71
rect 9926 37 9965 71
rect -9965 -71 -9926 -37
rect -9892 -71 -9868 -37
rect -9824 -71 -9796 -37
rect -9756 -71 -9724 -37
rect -9688 -71 -9654 -37
rect -9618 -71 -9586 -37
rect -9546 -71 -9518 -37
rect -9474 -71 -9450 -37
rect -9416 -71 -9377 -37
rect -8947 -71 -8908 -37
rect -8874 -71 -8850 -37
rect -8806 -71 -8778 -37
rect -8738 -71 -8706 -37
rect -8670 -71 -8636 -37
rect -8600 -71 -8568 -37
rect -8528 -71 -8500 -37
rect -8456 -71 -8432 -37
rect -8398 -71 -8359 -37
rect -7929 -71 -7890 -37
rect -7856 -71 -7832 -37
rect -7788 -71 -7760 -37
rect -7720 -71 -7688 -37
rect -7652 -71 -7618 -37
rect -7582 -71 -7550 -37
rect -7510 -71 -7482 -37
rect -7438 -71 -7414 -37
rect -7380 -71 -7341 -37
rect -6911 -71 -6872 -37
rect -6838 -71 -6814 -37
rect -6770 -71 -6742 -37
rect -6702 -71 -6670 -37
rect -6634 -71 -6600 -37
rect -6564 -71 -6532 -37
rect -6492 -71 -6464 -37
rect -6420 -71 -6396 -37
rect -6362 -71 -6323 -37
rect -5893 -71 -5854 -37
rect -5820 -71 -5796 -37
rect -5752 -71 -5724 -37
rect -5684 -71 -5652 -37
rect -5616 -71 -5582 -37
rect -5546 -71 -5514 -37
rect -5474 -71 -5446 -37
rect -5402 -71 -5378 -37
rect -5344 -71 -5305 -37
rect -4875 -71 -4836 -37
rect -4802 -71 -4778 -37
rect -4734 -71 -4706 -37
rect -4666 -71 -4634 -37
rect -4598 -71 -4564 -37
rect -4528 -71 -4496 -37
rect -4456 -71 -4428 -37
rect -4384 -71 -4360 -37
rect -4326 -71 -4287 -37
rect -3857 -71 -3818 -37
rect -3784 -71 -3760 -37
rect -3716 -71 -3688 -37
rect -3648 -71 -3616 -37
rect -3580 -71 -3546 -37
rect -3510 -71 -3478 -37
rect -3438 -71 -3410 -37
rect -3366 -71 -3342 -37
rect -3308 -71 -3269 -37
rect -2839 -71 -2800 -37
rect -2766 -71 -2742 -37
rect -2698 -71 -2670 -37
rect -2630 -71 -2598 -37
rect -2562 -71 -2528 -37
rect -2492 -71 -2460 -37
rect -2420 -71 -2392 -37
rect -2348 -71 -2324 -37
rect -2290 -71 -2251 -37
rect -1821 -71 -1782 -37
rect -1748 -71 -1724 -37
rect -1680 -71 -1652 -37
rect -1612 -71 -1580 -37
rect -1544 -71 -1510 -37
rect -1474 -71 -1442 -37
rect -1402 -71 -1374 -37
rect -1330 -71 -1306 -37
rect -1272 -71 -1233 -37
rect -803 -71 -764 -37
rect -730 -71 -706 -37
rect -662 -71 -634 -37
rect -594 -71 -562 -37
rect -526 -71 -492 -37
rect -456 -71 -424 -37
rect -384 -71 -356 -37
rect -312 -71 -288 -37
rect -254 -71 -215 -37
rect 215 -71 254 -37
rect 288 -71 312 -37
rect 356 -71 384 -37
rect 424 -71 456 -37
rect 492 -71 526 -37
rect 562 -71 594 -37
rect 634 -71 662 -37
rect 706 -71 730 -37
rect 764 -71 803 -37
rect 1233 -71 1272 -37
rect 1306 -71 1330 -37
rect 1374 -71 1402 -37
rect 1442 -71 1474 -37
rect 1510 -71 1544 -37
rect 1580 -71 1612 -37
rect 1652 -71 1680 -37
rect 1724 -71 1748 -37
rect 1782 -71 1821 -37
rect 2251 -71 2290 -37
rect 2324 -71 2348 -37
rect 2392 -71 2420 -37
rect 2460 -71 2492 -37
rect 2528 -71 2562 -37
rect 2598 -71 2630 -37
rect 2670 -71 2698 -37
rect 2742 -71 2766 -37
rect 2800 -71 2839 -37
rect 3269 -71 3308 -37
rect 3342 -71 3366 -37
rect 3410 -71 3438 -37
rect 3478 -71 3510 -37
rect 3546 -71 3580 -37
rect 3616 -71 3648 -37
rect 3688 -71 3716 -37
rect 3760 -71 3784 -37
rect 3818 -71 3857 -37
rect 4287 -71 4326 -37
rect 4360 -71 4384 -37
rect 4428 -71 4456 -37
rect 4496 -71 4528 -37
rect 4564 -71 4598 -37
rect 4634 -71 4666 -37
rect 4706 -71 4734 -37
rect 4778 -71 4802 -37
rect 4836 -71 4875 -37
rect 5305 -71 5344 -37
rect 5378 -71 5402 -37
rect 5446 -71 5474 -37
rect 5514 -71 5546 -37
rect 5582 -71 5616 -37
rect 5652 -71 5684 -37
rect 5724 -71 5752 -37
rect 5796 -71 5820 -37
rect 5854 -71 5893 -37
rect 6323 -71 6362 -37
rect 6396 -71 6420 -37
rect 6464 -71 6492 -37
rect 6532 -71 6564 -37
rect 6600 -71 6634 -37
rect 6670 -71 6702 -37
rect 6742 -71 6770 -37
rect 6814 -71 6838 -37
rect 6872 -71 6911 -37
rect 7341 -71 7380 -37
rect 7414 -71 7438 -37
rect 7482 -71 7510 -37
rect 7550 -71 7582 -37
rect 7618 -71 7652 -37
rect 7688 -71 7720 -37
rect 7760 -71 7788 -37
rect 7832 -71 7856 -37
rect 7890 -71 7929 -37
rect 8359 -71 8398 -37
rect 8432 -71 8456 -37
rect 8500 -71 8528 -37
rect 8568 -71 8600 -37
rect 8636 -71 8670 -37
rect 8706 -71 8738 -37
rect 8778 -71 8806 -37
rect 8850 -71 8874 -37
rect 8908 -71 8947 -37
rect 9377 -71 9416 -37
rect 9450 -71 9474 -37
rect 9518 -71 9546 -37
rect 9586 -71 9618 -37
rect 9654 -71 9688 -37
rect 9724 -71 9756 -37
rect 9796 -71 9824 -37
rect 9868 -71 9892 -37
rect 9926 -71 9965 -37
rect -10197 -140 -10163 -105
rect -10197 -212 -10163 -188
rect -10197 -284 -10163 -256
rect -10197 -356 -10163 -324
rect -10197 -426 -10163 -392
rect -10197 -494 -10163 -462
rect -10197 -562 -10163 -534
rect -10197 -630 -10163 -606
rect -10197 -713 -10163 -678
rect -9179 -140 -9145 -105
rect -9179 -212 -9145 -188
rect -9179 -284 -9145 -256
rect -9179 -356 -9145 -324
rect -9179 -426 -9145 -392
rect -9179 -494 -9145 -462
rect -9179 -562 -9145 -534
rect -9179 -630 -9145 -606
rect -9179 -713 -9145 -678
rect -8161 -140 -8127 -105
rect -8161 -212 -8127 -188
rect -8161 -284 -8127 -256
rect -8161 -356 -8127 -324
rect -8161 -426 -8127 -392
rect -8161 -494 -8127 -462
rect -8161 -562 -8127 -534
rect -8161 -630 -8127 -606
rect -8161 -713 -8127 -678
rect -7143 -140 -7109 -105
rect -7143 -212 -7109 -188
rect -7143 -284 -7109 -256
rect -7143 -356 -7109 -324
rect -7143 -426 -7109 -392
rect -7143 -494 -7109 -462
rect -7143 -562 -7109 -534
rect -7143 -630 -7109 -606
rect -7143 -713 -7109 -678
rect -6125 -140 -6091 -105
rect -6125 -212 -6091 -188
rect -6125 -284 -6091 -256
rect -6125 -356 -6091 -324
rect -6125 -426 -6091 -392
rect -6125 -494 -6091 -462
rect -6125 -562 -6091 -534
rect -6125 -630 -6091 -606
rect -6125 -713 -6091 -678
rect -5107 -140 -5073 -105
rect -5107 -212 -5073 -188
rect -5107 -284 -5073 -256
rect -5107 -356 -5073 -324
rect -5107 -426 -5073 -392
rect -5107 -494 -5073 -462
rect -5107 -562 -5073 -534
rect -5107 -630 -5073 -606
rect -5107 -713 -5073 -678
rect -4089 -140 -4055 -105
rect -4089 -212 -4055 -188
rect -4089 -284 -4055 -256
rect -4089 -356 -4055 -324
rect -4089 -426 -4055 -392
rect -4089 -494 -4055 -462
rect -4089 -562 -4055 -534
rect -4089 -630 -4055 -606
rect -4089 -713 -4055 -678
rect -3071 -140 -3037 -105
rect -3071 -212 -3037 -188
rect -3071 -284 -3037 -256
rect -3071 -356 -3037 -324
rect -3071 -426 -3037 -392
rect -3071 -494 -3037 -462
rect -3071 -562 -3037 -534
rect -3071 -630 -3037 -606
rect -3071 -713 -3037 -678
rect -2053 -140 -2019 -105
rect -2053 -212 -2019 -188
rect -2053 -284 -2019 -256
rect -2053 -356 -2019 -324
rect -2053 -426 -2019 -392
rect -2053 -494 -2019 -462
rect -2053 -562 -2019 -534
rect -2053 -630 -2019 -606
rect -2053 -713 -2019 -678
rect -1035 -140 -1001 -105
rect -1035 -212 -1001 -188
rect -1035 -284 -1001 -256
rect -1035 -356 -1001 -324
rect -1035 -426 -1001 -392
rect -1035 -494 -1001 -462
rect -1035 -562 -1001 -534
rect -1035 -630 -1001 -606
rect -1035 -713 -1001 -678
rect -17 -140 17 -105
rect -17 -212 17 -188
rect -17 -284 17 -256
rect -17 -356 17 -324
rect -17 -426 17 -392
rect -17 -494 17 -462
rect -17 -562 17 -534
rect -17 -630 17 -606
rect -17 -713 17 -678
rect 1001 -140 1035 -105
rect 1001 -212 1035 -188
rect 1001 -284 1035 -256
rect 1001 -356 1035 -324
rect 1001 -426 1035 -392
rect 1001 -494 1035 -462
rect 1001 -562 1035 -534
rect 1001 -630 1035 -606
rect 1001 -713 1035 -678
rect 2019 -140 2053 -105
rect 2019 -212 2053 -188
rect 2019 -284 2053 -256
rect 2019 -356 2053 -324
rect 2019 -426 2053 -392
rect 2019 -494 2053 -462
rect 2019 -562 2053 -534
rect 2019 -630 2053 -606
rect 2019 -713 2053 -678
rect 3037 -140 3071 -105
rect 3037 -212 3071 -188
rect 3037 -284 3071 -256
rect 3037 -356 3071 -324
rect 3037 -426 3071 -392
rect 3037 -494 3071 -462
rect 3037 -562 3071 -534
rect 3037 -630 3071 -606
rect 3037 -713 3071 -678
rect 4055 -140 4089 -105
rect 4055 -212 4089 -188
rect 4055 -284 4089 -256
rect 4055 -356 4089 -324
rect 4055 -426 4089 -392
rect 4055 -494 4089 -462
rect 4055 -562 4089 -534
rect 4055 -630 4089 -606
rect 4055 -713 4089 -678
rect 5073 -140 5107 -105
rect 5073 -212 5107 -188
rect 5073 -284 5107 -256
rect 5073 -356 5107 -324
rect 5073 -426 5107 -392
rect 5073 -494 5107 -462
rect 5073 -562 5107 -534
rect 5073 -630 5107 -606
rect 5073 -713 5107 -678
rect 6091 -140 6125 -105
rect 6091 -212 6125 -188
rect 6091 -284 6125 -256
rect 6091 -356 6125 -324
rect 6091 -426 6125 -392
rect 6091 -494 6125 -462
rect 6091 -562 6125 -534
rect 6091 -630 6125 -606
rect 6091 -713 6125 -678
rect 7109 -140 7143 -105
rect 7109 -212 7143 -188
rect 7109 -284 7143 -256
rect 7109 -356 7143 -324
rect 7109 -426 7143 -392
rect 7109 -494 7143 -462
rect 7109 -562 7143 -534
rect 7109 -630 7143 -606
rect 7109 -713 7143 -678
rect 8127 -140 8161 -105
rect 8127 -212 8161 -188
rect 8127 -284 8161 -256
rect 8127 -356 8161 -324
rect 8127 -426 8161 -392
rect 8127 -494 8161 -462
rect 8127 -562 8161 -534
rect 8127 -630 8161 -606
rect 8127 -713 8161 -678
rect 9145 -140 9179 -105
rect 9145 -212 9179 -188
rect 9145 -284 9179 -256
rect 9145 -356 9179 -324
rect 9145 -426 9179 -392
rect 9145 -494 9179 -462
rect 9145 -562 9179 -534
rect 9145 -630 9179 -606
rect 9145 -713 9179 -678
rect 10163 -140 10197 -105
rect 10163 -212 10197 -188
rect 10163 -284 10197 -256
rect 10163 -356 10197 -324
rect 10163 -426 10197 -392
rect 10163 -494 10197 -462
rect 10163 -562 10197 -534
rect 10163 -630 10197 -606
rect 10163 -713 10197 -678
rect -9965 -781 -9926 -747
rect -9892 -781 -9868 -747
rect -9824 -781 -9796 -747
rect -9756 -781 -9724 -747
rect -9688 -781 -9654 -747
rect -9618 -781 -9586 -747
rect -9546 -781 -9518 -747
rect -9474 -781 -9450 -747
rect -9416 -781 -9377 -747
rect -8947 -781 -8908 -747
rect -8874 -781 -8850 -747
rect -8806 -781 -8778 -747
rect -8738 -781 -8706 -747
rect -8670 -781 -8636 -747
rect -8600 -781 -8568 -747
rect -8528 -781 -8500 -747
rect -8456 -781 -8432 -747
rect -8398 -781 -8359 -747
rect -7929 -781 -7890 -747
rect -7856 -781 -7832 -747
rect -7788 -781 -7760 -747
rect -7720 -781 -7688 -747
rect -7652 -781 -7618 -747
rect -7582 -781 -7550 -747
rect -7510 -781 -7482 -747
rect -7438 -781 -7414 -747
rect -7380 -781 -7341 -747
rect -6911 -781 -6872 -747
rect -6838 -781 -6814 -747
rect -6770 -781 -6742 -747
rect -6702 -781 -6670 -747
rect -6634 -781 -6600 -747
rect -6564 -781 -6532 -747
rect -6492 -781 -6464 -747
rect -6420 -781 -6396 -747
rect -6362 -781 -6323 -747
rect -5893 -781 -5854 -747
rect -5820 -781 -5796 -747
rect -5752 -781 -5724 -747
rect -5684 -781 -5652 -747
rect -5616 -781 -5582 -747
rect -5546 -781 -5514 -747
rect -5474 -781 -5446 -747
rect -5402 -781 -5378 -747
rect -5344 -781 -5305 -747
rect -4875 -781 -4836 -747
rect -4802 -781 -4778 -747
rect -4734 -781 -4706 -747
rect -4666 -781 -4634 -747
rect -4598 -781 -4564 -747
rect -4528 -781 -4496 -747
rect -4456 -781 -4428 -747
rect -4384 -781 -4360 -747
rect -4326 -781 -4287 -747
rect -3857 -781 -3818 -747
rect -3784 -781 -3760 -747
rect -3716 -781 -3688 -747
rect -3648 -781 -3616 -747
rect -3580 -781 -3546 -747
rect -3510 -781 -3478 -747
rect -3438 -781 -3410 -747
rect -3366 -781 -3342 -747
rect -3308 -781 -3269 -747
rect -2839 -781 -2800 -747
rect -2766 -781 -2742 -747
rect -2698 -781 -2670 -747
rect -2630 -781 -2598 -747
rect -2562 -781 -2528 -747
rect -2492 -781 -2460 -747
rect -2420 -781 -2392 -747
rect -2348 -781 -2324 -747
rect -2290 -781 -2251 -747
rect -1821 -781 -1782 -747
rect -1748 -781 -1724 -747
rect -1680 -781 -1652 -747
rect -1612 -781 -1580 -747
rect -1544 -781 -1510 -747
rect -1474 -781 -1442 -747
rect -1402 -781 -1374 -747
rect -1330 -781 -1306 -747
rect -1272 -781 -1233 -747
rect -803 -781 -764 -747
rect -730 -781 -706 -747
rect -662 -781 -634 -747
rect -594 -781 -562 -747
rect -526 -781 -492 -747
rect -456 -781 -424 -747
rect -384 -781 -356 -747
rect -312 -781 -288 -747
rect -254 -781 -215 -747
rect 215 -781 254 -747
rect 288 -781 312 -747
rect 356 -781 384 -747
rect 424 -781 456 -747
rect 492 -781 526 -747
rect 562 -781 594 -747
rect 634 -781 662 -747
rect 706 -781 730 -747
rect 764 -781 803 -747
rect 1233 -781 1272 -747
rect 1306 -781 1330 -747
rect 1374 -781 1402 -747
rect 1442 -781 1474 -747
rect 1510 -781 1544 -747
rect 1580 -781 1612 -747
rect 1652 -781 1680 -747
rect 1724 -781 1748 -747
rect 1782 -781 1821 -747
rect 2251 -781 2290 -747
rect 2324 -781 2348 -747
rect 2392 -781 2420 -747
rect 2460 -781 2492 -747
rect 2528 -781 2562 -747
rect 2598 -781 2630 -747
rect 2670 -781 2698 -747
rect 2742 -781 2766 -747
rect 2800 -781 2839 -747
rect 3269 -781 3308 -747
rect 3342 -781 3366 -747
rect 3410 -781 3438 -747
rect 3478 -781 3510 -747
rect 3546 -781 3580 -747
rect 3616 -781 3648 -747
rect 3688 -781 3716 -747
rect 3760 -781 3784 -747
rect 3818 -781 3857 -747
rect 4287 -781 4326 -747
rect 4360 -781 4384 -747
rect 4428 -781 4456 -747
rect 4496 -781 4528 -747
rect 4564 -781 4598 -747
rect 4634 -781 4666 -747
rect 4706 -781 4734 -747
rect 4778 -781 4802 -747
rect 4836 -781 4875 -747
rect 5305 -781 5344 -747
rect 5378 -781 5402 -747
rect 5446 -781 5474 -747
rect 5514 -781 5546 -747
rect 5582 -781 5616 -747
rect 5652 -781 5684 -747
rect 5724 -781 5752 -747
rect 5796 -781 5820 -747
rect 5854 -781 5893 -747
rect 6323 -781 6362 -747
rect 6396 -781 6420 -747
rect 6464 -781 6492 -747
rect 6532 -781 6564 -747
rect 6600 -781 6634 -747
rect 6670 -781 6702 -747
rect 6742 -781 6770 -747
rect 6814 -781 6838 -747
rect 6872 -781 6911 -747
rect 7341 -781 7380 -747
rect 7414 -781 7438 -747
rect 7482 -781 7510 -747
rect 7550 -781 7582 -747
rect 7618 -781 7652 -747
rect 7688 -781 7720 -747
rect 7760 -781 7788 -747
rect 7832 -781 7856 -747
rect 7890 -781 7929 -747
rect 8359 -781 8398 -747
rect 8432 -781 8456 -747
rect 8500 -781 8528 -747
rect 8568 -781 8600 -747
rect 8636 -781 8670 -747
rect 8706 -781 8738 -747
rect 8778 -781 8806 -747
rect 8850 -781 8874 -747
rect 8908 -781 8947 -747
rect 9377 -781 9416 -747
rect 9450 -781 9474 -747
rect 9518 -781 9546 -747
rect 9586 -781 9618 -747
rect 9654 -781 9688 -747
rect 9724 -781 9756 -747
rect 9796 -781 9824 -747
rect 9868 -781 9892 -747
rect 9926 -781 9965 -747
<< viali >>
rect -9868 747 -9858 781
rect -9858 747 -9834 781
rect -9796 747 -9790 781
rect -9790 747 -9762 781
rect -9724 747 -9722 781
rect -9722 747 -9690 781
rect -9652 747 -9620 781
rect -9620 747 -9618 781
rect -9580 747 -9552 781
rect -9552 747 -9546 781
rect -9508 747 -9484 781
rect -9484 747 -9474 781
rect -8850 747 -8840 781
rect -8840 747 -8816 781
rect -8778 747 -8772 781
rect -8772 747 -8744 781
rect -8706 747 -8704 781
rect -8704 747 -8672 781
rect -8634 747 -8602 781
rect -8602 747 -8600 781
rect -8562 747 -8534 781
rect -8534 747 -8528 781
rect -8490 747 -8466 781
rect -8466 747 -8456 781
rect -7832 747 -7822 781
rect -7822 747 -7798 781
rect -7760 747 -7754 781
rect -7754 747 -7726 781
rect -7688 747 -7686 781
rect -7686 747 -7654 781
rect -7616 747 -7584 781
rect -7584 747 -7582 781
rect -7544 747 -7516 781
rect -7516 747 -7510 781
rect -7472 747 -7448 781
rect -7448 747 -7438 781
rect -6814 747 -6804 781
rect -6804 747 -6780 781
rect -6742 747 -6736 781
rect -6736 747 -6708 781
rect -6670 747 -6668 781
rect -6668 747 -6636 781
rect -6598 747 -6566 781
rect -6566 747 -6564 781
rect -6526 747 -6498 781
rect -6498 747 -6492 781
rect -6454 747 -6430 781
rect -6430 747 -6420 781
rect -5796 747 -5786 781
rect -5786 747 -5762 781
rect -5724 747 -5718 781
rect -5718 747 -5690 781
rect -5652 747 -5650 781
rect -5650 747 -5618 781
rect -5580 747 -5548 781
rect -5548 747 -5546 781
rect -5508 747 -5480 781
rect -5480 747 -5474 781
rect -5436 747 -5412 781
rect -5412 747 -5402 781
rect -4778 747 -4768 781
rect -4768 747 -4744 781
rect -4706 747 -4700 781
rect -4700 747 -4672 781
rect -4634 747 -4632 781
rect -4632 747 -4600 781
rect -4562 747 -4530 781
rect -4530 747 -4528 781
rect -4490 747 -4462 781
rect -4462 747 -4456 781
rect -4418 747 -4394 781
rect -4394 747 -4384 781
rect -3760 747 -3750 781
rect -3750 747 -3726 781
rect -3688 747 -3682 781
rect -3682 747 -3654 781
rect -3616 747 -3614 781
rect -3614 747 -3582 781
rect -3544 747 -3512 781
rect -3512 747 -3510 781
rect -3472 747 -3444 781
rect -3444 747 -3438 781
rect -3400 747 -3376 781
rect -3376 747 -3366 781
rect -2742 747 -2732 781
rect -2732 747 -2708 781
rect -2670 747 -2664 781
rect -2664 747 -2636 781
rect -2598 747 -2596 781
rect -2596 747 -2564 781
rect -2526 747 -2494 781
rect -2494 747 -2492 781
rect -2454 747 -2426 781
rect -2426 747 -2420 781
rect -2382 747 -2358 781
rect -2358 747 -2348 781
rect -1724 747 -1714 781
rect -1714 747 -1690 781
rect -1652 747 -1646 781
rect -1646 747 -1618 781
rect -1580 747 -1578 781
rect -1578 747 -1546 781
rect -1508 747 -1476 781
rect -1476 747 -1474 781
rect -1436 747 -1408 781
rect -1408 747 -1402 781
rect -1364 747 -1340 781
rect -1340 747 -1330 781
rect -706 747 -696 781
rect -696 747 -672 781
rect -634 747 -628 781
rect -628 747 -600 781
rect -562 747 -560 781
rect -560 747 -528 781
rect -490 747 -458 781
rect -458 747 -456 781
rect -418 747 -390 781
rect -390 747 -384 781
rect -346 747 -322 781
rect -322 747 -312 781
rect 312 747 322 781
rect 322 747 346 781
rect 384 747 390 781
rect 390 747 418 781
rect 456 747 458 781
rect 458 747 490 781
rect 528 747 560 781
rect 560 747 562 781
rect 600 747 628 781
rect 628 747 634 781
rect 672 747 696 781
rect 696 747 706 781
rect 1330 747 1340 781
rect 1340 747 1364 781
rect 1402 747 1408 781
rect 1408 747 1436 781
rect 1474 747 1476 781
rect 1476 747 1508 781
rect 1546 747 1578 781
rect 1578 747 1580 781
rect 1618 747 1646 781
rect 1646 747 1652 781
rect 1690 747 1714 781
rect 1714 747 1724 781
rect 2348 747 2358 781
rect 2358 747 2382 781
rect 2420 747 2426 781
rect 2426 747 2454 781
rect 2492 747 2494 781
rect 2494 747 2526 781
rect 2564 747 2596 781
rect 2596 747 2598 781
rect 2636 747 2664 781
rect 2664 747 2670 781
rect 2708 747 2732 781
rect 2732 747 2742 781
rect 3366 747 3376 781
rect 3376 747 3400 781
rect 3438 747 3444 781
rect 3444 747 3472 781
rect 3510 747 3512 781
rect 3512 747 3544 781
rect 3582 747 3614 781
rect 3614 747 3616 781
rect 3654 747 3682 781
rect 3682 747 3688 781
rect 3726 747 3750 781
rect 3750 747 3760 781
rect 4384 747 4394 781
rect 4394 747 4418 781
rect 4456 747 4462 781
rect 4462 747 4490 781
rect 4528 747 4530 781
rect 4530 747 4562 781
rect 4600 747 4632 781
rect 4632 747 4634 781
rect 4672 747 4700 781
rect 4700 747 4706 781
rect 4744 747 4768 781
rect 4768 747 4778 781
rect 5402 747 5412 781
rect 5412 747 5436 781
rect 5474 747 5480 781
rect 5480 747 5508 781
rect 5546 747 5548 781
rect 5548 747 5580 781
rect 5618 747 5650 781
rect 5650 747 5652 781
rect 5690 747 5718 781
rect 5718 747 5724 781
rect 5762 747 5786 781
rect 5786 747 5796 781
rect 6420 747 6430 781
rect 6430 747 6454 781
rect 6492 747 6498 781
rect 6498 747 6526 781
rect 6564 747 6566 781
rect 6566 747 6598 781
rect 6636 747 6668 781
rect 6668 747 6670 781
rect 6708 747 6736 781
rect 6736 747 6742 781
rect 6780 747 6804 781
rect 6804 747 6814 781
rect 7438 747 7448 781
rect 7448 747 7472 781
rect 7510 747 7516 781
rect 7516 747 7544 781
rect 7582 747 7584 781
rect 7584 747 7616 781
rect 7654 747 7686 781
rect 7686 747 7688 781
rect 7726 747 7754 781
rect 7754 747 7760 781
rect 7798 747 7822 781
rect 7822 747 7832 781
rect 8456 747 8466 781
rect 8466 747 8490 781
rect 8528 747 8534 781
rect 8534 747 8562 781
rect 8600 747 8602 781
rect 8602 747 8634 781
rect 8672 747 8704 781
rect 8704 747 8706 781
rect 8744 747 8772 781
rect 8772 747 8778 781
rect 8816 747 8840 781
rect 8840 747 8850 781
rect 9474 747 9484 781
rect 9484 747 9508 781
rect 9546 747 9552 781
rect 9552 747 9580 781
rect 9618 747 9620 781
rect 9620 747 9652 781
rect 9690 747 9722 781
rect 9722 747 9724 781
rect 9762 747 9790 781
rect 9790 747 9796 781
rect 9834 747 9858 781
rect 9858 747 9868 781
rect -10197 664 -10163 678
rect -10197 644 -10163 664
rect -10197 596 -10163 606
rect -10197 572 -10163 596
rect -10197 528 -10163 534
rect -10197 500 -10163 528
rect -10197 460 -10163 462
rect -10197 428 -10163 460
rect -10197 358 -10163 390
rect -10197 356 -10163 358
rect -10197 290 -10163 318
rect -10197 284 -10163 290
rect -10197 222 -10163 246
rect -10197 212 -10163 222
rect -10197 154 -10163 174
rect -10197 140 -10163 154
rect -9179 664 -9145 678
rect -9179 644 -9145 664
rect -9179 596 -9145 606
rect -9179 572 -9145 596
rect -9179 528 -9145 534
rect -9179 500 -9145 528
rect -9179 460 -9145 462
rect -9179 428 -9145 460
rect -9179 358 -9145 390
rect -9179 356 -9145 358
rect -9179 290 -9145 318
rect -9179 284 -9145 290
rect -9179 222 -9145 246
rect -9179 212 -9145 222
rect -9179 154 -9145 174
rect -9179 140 -9145 154
rect -8161 664 -8127 678
rect -8161 644 -8127 664
rect -8161 596 -8127 606
rect -8161 572 -8127 596
rect -8161 528 -8127 534
rect -8161 500 -8127 528
rect -8161 460 -8127 462
rect -8161 428 -8127 460
rect -8161 358 -8127 390
rect -8161 356 -8127 358
rect -8161 290 -8127 318
rect -8161 284 -8127 290
rect -8161 222 -8127 246
rect -8161 212 -8127 222
rect -8161 154 -8127 174
rect -8161 140 -8127 154
rect -7143 664 -7109 678
rect -7143 644 -7109 664
rect -7143 596 -7109 606
rect -7143 572 -7109 596
rect -7143 528 -7109 534
rect -7143 500 -7109 528
rect -7143 460 -7109 462
rect -7143 428 -7109 460
rect -7143 358 -7109 390
rect -7143 356 -7109 358
rect -7143 290 -7109 318
rect -7143 284 -7109 290
rect -7143 222 -7109 246
rect -7143 212 -7109 222
rect -7143 154 -7109 174
rect -7143 140 -7109 154
rect -6125 664 -6091 678
rect -6125 644 -6091 664
rect -6125 596 -6091 606
rect -6125 572 -6091 596
rect -6125 528 -6091 534
rect -6125 500 -6091 528
rect -6125 460 -6091 462
rect -6125 428 -6091 460
rect -6125 358 -6091 390
rect -6125 356 -6091 358
rect -6125 290 -6091 318
rect -6125 284 -6091 290
rect -6125 222 -6091 246
rect -6125 212 -6091 222
rect -6125 154 -6091 174
rect -6125 140 -6091 154
rect -5107 664 -5073 678
rect -5107 644 -5073 664
rect -5107 596 -5073 606
rect -5107 572 -5073 596
rect -5107 528 -5073 534
rect -5107 500 -5073 528
rect -5107 460 -5073 462
rect -5107 428 -5073 460
rect -5107 358 -5073 390
rect -5107 356 -5073 358
rect -5107 290 -5073 318
rect -5107 284 -5073 290
rect -5107 222 -5073 246
rect -5107 212 -5073 222
rect -5107 154 -5073 174
rect -5107 140 -5073 154
rect -4089 664 -4055 678
rect -4089 644 -4055 664
rect -4089 596 -4055 606
rect -4089 572 -4055 596
rect -4089 528 -4055 534
rect -4089 500 -4055 528
rect -4089 460 -4055 462
rect -4089 428 -4055 460
rect -4089 358 -4055 390
rect -4089 356 -4055 358
rect -4089 290 -4055 318
rect -4089 284 -4055 290
rect -4089 222 -4055 246
rect -4089 212 -4055 222
rect -4089 154 -4055 174
rect -4089 140 -4055 154
rect -3071 664 -3037 678
rect -3071 644 -3037 664
rect -3071 596 -3037 606
rect -3071 572 -3037 596
rect -3071 528 -3037 534
rect -3071 500 -3037 528
rect -3071 460 -3037 462
rect -3071 428 -3037 460
rect -3071 358 -3037 390
rect -3071 356 -3037 358
rect -3071 290 -3037 318
rect -3071 284 -3037 290
rect -3071 222 -3037 246
rect -3071 212 -3037 222
rect -3071 154 -3037 174
rect -3071 140 -3037 154
rect -2053 664 -2019 678
rect -2053 644 -2019 664
rect -2053 596 -2019 606
rect -2053 572 -2019 596
rect -2053 528 -2019 534
rect -2053 500 -2019 528
rect -2053 460 -2019 462
rect -2053 428 -2019 460
rect -2053 358 -2019 390
rect -2053 356 -2019 358
rect -2053 290 -2019 318
rect -2053 284 -2019 290
rect -2053 222 -2019 246
rect -2053 212 -2019 222
rect -2053 154 -2019 174
rect -2053 140 -2019 154
rect -1035 664 -1001 678
rect -1035 644 -1001 664
rect -1035 596 -1001 606
rect -1035 572 -1001 596
rect -1035 528 -1001 534
rect -1035 500 -1001 528
rect -1035 460 -1001 462
rect -1035 428 -1001 460
rect -1035 358 -1001 390
rect -1035 356 -1001 358
rect -1035 290 -1001 318
rect -1035 284 -1001 290
rect -1035 222 -1001 246
rect -1035 212 -1001 222
rect -1035 154 -1001 174
rect -1035 140 -1001 154
rect -17 664 17 678
rect -17 644 17 664
rect -17 596 17 606
rect -17 572 17 596
rect -17 528 17 534
rect -17 500 17 528
rect -17 460 17 462
rect -17 428 17 460
rect -17 358 17 390
rect -17 356 17 358
rect -17 290 17 318
rect -17 284 17 290
rect -17 222 17 246
rect -17 212 17 222
rect -17 154 17 174
rect -17 140 17 154
rect 1001 664 1035 678
rect 1001 644 1035 664
rect 1001 596 1035 606
rect 1001 572 1035 596
rect 1001 528 1035 534
rect 1001 500 1035 528
rect 1001 460 1035 462
rect 1001 428 1035 460
rect 1001 358 1035 390
rect 1001 356 1035 358
rect 1001 290 1035 318
rect 1001 284 1035 290
rect 1001 222 1035 246
rect 1001 212 1035 222
rect 1001 154 1035 174
rect 1001 140 1035 154
rect 2019 664 2053 678
rect 2019 644 2053 664
rect 2019 596 2053 606
rect 2019 572 2053 596
rect 2019 528 2053 534
rect 2019 500 2053 528
rect 2019 460 2053 462
rect 2019 428 2053 460
rect 2019 358 2053 390
rect 2019 356 2053 358
rect 2019 290 2053 318
rect 2019 284 2053 290
rect 2019 222 2053 246
rect 2019 212 2053 222
rect 2019 154 2053 174
rect 2019 140 2053 154
rect 3037 664 3071 678
rect 3037 644 3071 664
rect 3037 596 3071 606
rect 3037 572 3071 596
rect 3037 528 3071 534
rect 3037 500 3071 528
rect 3037 460 3071 462
rect 3037 428 3071 460
rect 3037 358 3071 390
rect 3037 356 3071 358
rect 3037 290 3071 318
rect 3037 284 3071 290
rect 3037 222 3071 246
rect 3037 212 3071 222
rect 3037 154 3071 174
rect 3037 140 3071 154
rect 4055 664 4089 678
rect 4055 644 4089 664
rect 4055 596 4089 606
rect 4055 572 4089 596
rect 4055 528 4089 534
rect 4055 500 4089 528
rect 4055 460 4089 462
rect 4055 428 4089 460
rect 4055 358 4089 390
rect 4055 356 4089 358
rect 4055 290 4089 318
rect 4055 284 4089 290
rect 4055 222 4089 246
rect 4055 212 4089 222
rect 4055 154 4089 174
rect 4055 140 4089 154
rect 5073 664 5107 678
rect 5073 644 5107 664
rect 5073 596 5107 606
rect 5073 572 5107 596
rect 5073 528 5107 534
rect 5073 500 5107 528
rect 5073 460 5107 462
rect 5073 428 5107 460
rect 5073 358 5107 390
rect 5073 356 5107 358
rect 5073 290 5107 318
rect 5073 284 5107 290
rect 5073 222 5107 246
rect 5073 212 5107 222
rect 5073 154 5107 174
rect 5073 140 5107 154
rect 6091 664 6125 678
rect 6091 644 6125 664
rect 6091 596 6125 606
rect 6091 572 6125 596
rect 6091 528 6125 534
rect 6091 500 6125 528
rect 6091 460 6125 462
rect 6091 428 6125 460
rect 6091 358 6125 390
rect 6091 356 6125 358
rect 6091 290 6125 318
rect 6091 284 6125 290
rect 6091 222 6125 246
rect 6091 212 6125 222
rect 6091 154 6125 174
rect 6091 140 6125 154
rect 7109 664 7143 678
rect 7109 644 7143 664
rect 7109 596 7143 606
rect 7109 572 7143 596
rect 7109 528 7143 534
rect 7109 500 7143 528
rect 7109 460 7143 462
rect 7109 428 7143 460
rect 7109 358 7143 390
rect 7109 356 7143 358
rect 7109 290 7143 318
rect 7109 284 7143 290
rect 7109 222 7143 246
rect 7109 212 7143 222
rect 7109 154 7143 174
rect 7109 140 7143 154
rect 8127 664 8161 678
rect 8127 644 8161 664
rect 8127 596 8161 606
rect 8127 572 8161 596
rect 8127 528 8161 534
rect 8127 500 8161 528
rect 8127 460 8161 462
rect 8127 428 8161 460
rect 8127 358 8161 390
rect 8127 356 8161 358
rect 8127 290 8161 318
rect 8127 284 8161 290
rect 8127 222 8161 246
rect 8127 212 8161 222
rect 8127 154 8161 174
rect 8127 140 8161 154
rect 9145 664 9179 678
rect 9145 644 9179 664
rect 9145 596 9179 606
rect 9145 572 9179 596
rect 9145 528 9179 534
rect 9145 500 9179 528
rect 9145 460 9179 462
rect 9145 428 9179 460
rect 9145 358 9179 390
rect 9145 356 9179 358
rect 9145 290 9179 318
rect 9145 284 9179 290
rect 9145 222 9179 246
rect 9145 212 9179 222
rect 9145 154 9179 174
rect 9145 140 9179 154
rect 10163 664 10197 678
rect 10163 644 10197 664
rect 10163 596 10197 606
rect 10163 572 10197 596
rect 10163 528 10197 534
rect 10163 500 10197 528
rect 10163 460 10197 462
rect 10163 428 10197 460
rect 10163 358 10197 390
rect 10163 356 10197 358
rect 10163 290 10197 318
rect 10163 284 10197 290
rect 10163 222 10197 246
rect 10163 212 10197 222
rect 10163 154 10197 174
rect 10163 140 10197 154
rect -9868 37 -9858 71
rect -9858 37 -9834 71
rect -9796 37 -9790 71
rect -9790 37 -9762 71
rect -9724 37 -9722 71
rect -9722 37 -9690 71
rect -9652 37 -9620 71
rect -9620 37 -9618 71
rect -9580 37 -9552 71
rect -9552 37 -9546 71
rect -9508 37 -9484 71
rect -9484 37 -9474 71
rect -8850 37 -8840 71
rect -8840 37 -8816 71
rect -8778 37 -8772 71
rect -8772 37 -8744 71
rect -8706 37 -8704 71
rect -8704 37 -8672 71
rect -8634 37 -8602 71
rect -8602 37 -8600 71
rect -8562 37 -8534 71
rect -8534 37 -8528 71
rect -8490 37 -8466 71
rect -8466 37 -8456 71
rect -7832 37 -7822 71
rect -7822 37 -7798 71
rect -7760 37 -7754 71
rect -7754 37 -7726 71
rect -7688 37 -7686 71
rect -7686 37 -7654 71
rect -7616 37 -7584 71
rect -7584 37 -7582 71
rect -7544 37 -7516 71
rect -7516 37 -7510 71
rect -7472 37 -7448 71
rect -7448 37 -7438 71
rect -6814 37 -6804 71
rect -6804 37 -6780 71
rect -6742 37 -6736 71
rect -6736 37 -6708 71
rect -6670 37 -6668 71
rect -6668 37 -6636 71
rect -6598 37 -6566 71
rect -6566 37 -6564 71
rect -6526 37 -6498 71
rect -6498 37 -6492 71
rect -6454 37 -6430 71
rect -6430 37 -6420 71
rect -5796 37 -5786 71
rect -5786 37 -5762 71
rect -5724 37 -5718 71
rect -5718 37 -5690 71
rect -5652 37 -5650 71
rect -5650 37 -5618 71
rect -5580 37 -5548 71
rect -5548 37 -5546 71
rect -5508 37 -5480 71
rect -5480 37 -5474 71
rect -5436 37 -5412 71
rect -5412 37 -5402 71
rect -4778 37 -4768 71
rect -4768 37 -4744 71
rect -4706 37 -4700 71
rect -4700 37 -4672 71
rect -4634 37 -4632 71
rect -4632 37 -4600 71
rect -4562 37 -4530 71
rect -4530 37 -4528 71
rect -4490 37 -4462 71
rect -4462 37 -4456 71
rect -4418 37 -4394 71
rect -4394 37 -4384 71
rect -3760 37 -3750 71
rect -3750 37 -3726 71
rect -3688 37 -3682 71
rect -3682 37 -3654 71
rect -3616 37 -3614 71
rect -3614 37 -3582 71
rect -3544 37 -3512 71
rect -3512 37 -3510 71
rect -3472 37 -3444 71
rect -3444 37 -3438 71
rect -3400 37 -3376 71
rect -3376 37 -3366 71
rect -2742 37 -2732 71
rect -2732 37 -2708 71
rect -2670 37 -2664 71
rect -2664 37 -2636 71
rect -2598 37 -2596 71
rect -2596 37 -2564 71
rect -2526 37 -2494 71
rect -2494 37 -2492 71
rect -2454 37 -2426 71
rect -2426 37 -2420 71
rect -2382 37 -2358 71
rect -2358 37 -2348 71
rect -1724 37 -1714 71
rect -1714 37 -1690 71
rect -1652 37 -1646 71
rect -1646 37 -1618 71
rect -1580 37 -1578 71
rect -1578 37 -1546 71
rect -1508 37 -1476 71
rect -1476 37 -1474 71
rect -1436 37 -1408 71
rect -1408 37 -1402 71
rect -1364 37 -1340 71
rect -1340 37 -1330 71
rect -706 37 -696 71
rect -696 37 -672 71
rect -634 37 -628 71
rect -628 37 -600 71
rect -562 37 -560 71
rect -560 37 -528 71
rect -490 37 -458 71
rect -458 37 -456 71
rect -418 37 -390 71
rect -390 37 -384 71
rect -346 37 -322 71
rect -322 37 -312 71
rect 312 37 322 71
rect 322 37 346 71
rect 384 37 390 71
rect 390 37 418 71
rect 456 37 458 71
rect 458 37 490 71
rect 528 37 560 71
rect 560 37 562 71
rect 600 37 628 71
rect 628 37 634 71
rect 672 37 696 71
rect 696 37 706 71
rect 1330 37 1340 71
rect 1340 37 1364 71
rect 1402 37 1408 71
rect 1408 37 1436 71
rect 1474 37 1476 71
rect 1476 37 1508 71
rect 1546 37 1578 71
rect 1578 37 1580 71
rect 1618 37 1646 71
rect 1646 37 1652 71
rect 1690 37 1714 71
rect 1714 37 1724 71
rect 2348 37 2358 71
rect 2358 37 2382 71
rect 2420 37 2426 71
rect 2426 37 2454 71
rect 2492 37 2494 71
rect 2494 37 2526 71
rect 2564 37 2596 71
rect 2596 37 2598 71
rect 2636 37 2664 71
rect 2664 37 2670 71
rect 2708 37 2732 71
rect 2732 37 2742 71
rect 3366 37 3376 71
rect 3376 37 3400 71
rect 3438 37 3444 71
rect 3444 37 3472 71
rect 3510 37 3512 71
rect 3512 37 3544 71
rect 3582 37 3614 71
rect 3614 37 3616 71
rect 3654 37 3682 71
rect 3682 37 3688 71
rect 3726 37 3750 71
rect 3750 37 3760 71
rect 4384 37 4394 71
rect 4394 37 4418 71
rect 4456 37 4462 71
rect 4462 37 4490 71
rect 4528 37 4530 71
rect 4530 37 4562 71
rect 4600 37 4632 71
rect 4632 37 4634 71
rect 4672 37 4700 71
rect 4700 37 4706 71
rect 4744 37 4768 71
rect 4768 37 4778 71
rect 5402 37 5412 71
rect 5412 37 5436 71
rect 5474 37 5480 71
rect 5480 37 5508 71
rect 5546 37 5548 71
rect 5548 37 5580 71
rect 5618 37 5650 71
rect 5650 37 5652 71
rect 5690 37 5718 71
rect 5718 37 5724 71
rect 5762 37 5786 71
rect 5786 37 5796 71
rect 6420 37 6430 71
rect 6430 37 6454 71
rect 6492 37 6498 71
rect 6498 37 6526 71
rect 6564 37 6566 71
rect 6566 37 6598 71
rect 6636 37 6668 71
rect 6668 37 6670 71
rect 6708 37 6736 71
rect 6736 37 6742 71
rect 6780 37 6804 71
rect 6804 37 6814 71
rect 7438 37 7448 71
rect 7448 37 7472 71
rect 7510 37 7516 71
rect 7516 37 7544 71
rect 7582 37 7584 71
rect 7584 37 7616 71
rect 7654 37 7686 71
rect 7686 37 7688 71
rect 7726 37 7754 71
rect 7754 37 7760 71
rect 7798 37 7822 71
rect 7822 37 7832 71
rect 8456 37 8466 71
rect 8466 37 8490 71
rect 8528 37 8534 71
rect 8534 37 8562 71
rect 8600 37 8602 71
rect 8602 37 8634 71
rect 8672 37 8704 71
rect 8704 37 8706 71
rect 8744 37 8772 71
rect 8772 37 8778 71
rect 8816 37 8840 71
rect 8840 37 8850 71
rect 9474 37 9484 71
rect 9484 37 9508 71
rect 9546 37 9552 71
rect 9552 37 9580 71
rect 9618 37 9620 71
rect 9620 37 9652 71
rect 9690 37 9722 71
rect 9722 37 9724 71
rect 9762 37 9790 71
rect 9790 37 9796 71
rect 9834 37 9858 71
rect 9858 37 9868 71
rect -9868 -71 -9858 -37
rect -9858 -71 -9834 -37
rect -9796 -71 -9790 -37
rect -9790 -71 -9762 -37
rect -9724 -71 -9722 -37
rect -9722 -71 -9690 -37
rect -9652 -71 -9620 -37
rect -9620 -71 -9618 -37
rect -9580 -71 -9552 -37
rect -9552 -71 -9546 -37
rect -9508 -71 -9484 -37
rect -9484 -71 -9474 -37
rect -8850 -71 -8840 -37
rect -8840 -71 -8816 -37
rect -8778 -71 -8772 -37
rect -8772 -71 -8744 -37
rect -8706 -71 -8704 -37
rect -8704 -71 -8672 -37
rect -8634 -71 -8602 -37
rect -8602 -71 -8600 -37
rect -8562 -71 -8534 -37
rect -8534 -71 -8528 -37
rect -8490 -71 -8466 -37
rect -8466 -71 -8456 -37
rect -7832 -71 -7822 -37
rect -7822 -71 -7798 -37
rect -7760 -71 -7754 -37
rect -7754 -71 -7726 -37
rect -7688 -71 -7686 -37
rect -7686 -71 -7654 -37
rect -7616 -71 -7584 -37
rect -7584 -71 -7582 -37
rect -7544 -71 -7516 -37
rect -7516 -71 -7510 -37
rect -7472 -71 -7448 -37
rect -7448 -71 -7438 -37
rect -6814 -71 -6804 -37
rect -6804 -71 -6780 -37
rect -6742 -71 -6736 -37
rect -6736 -71 -6708 -37
rect -6670 -71 -6668 -37
rect -6668 -71 -6636 -37
rect -6598 -71 -6566 -37
rect -6566 -71 -6564 -37
rect -6526 -71 -6498 -37
rect -6498 -71 -6492 -37
rect -6454 -71 -6430 -37
rect -6430 -71 -6420 -37
rect -5796 -71 -5786 -37
rect -5786 -71 -5762 -37
rect -5724 -71 -5718 -37
rect -5718 -71 -5690 -37
rect -5652 -71 -5650 -37
rect -5650 -71 -5618 -37
rect -5580 -71 -5548 -37
rect -5548 -71 -5546 -37
rect -5508 -71 -5480 -37
rect -5480 -71 -5474 -37
rect -5436 -71 -5412 -37
rect -5412 -71 -5402 -37
rect -4778 -71 -4768 -37
rect -4768 -71 -4744 -37
rect -4706 -71 -4700 -37
rect -4700 -71 -4672 -37
rect -4634 -71 -4632 -37
rect -4632 -71 -4600 -37
rect -4562 -71 -4530 -37
rect -4530 -71 -4528 -37
rect -4490 -71 -4462 -37
rect -4462 -71 -4456 -37
rect -4418 -71 -4394 -37
rect -4394 -71 -4384 -37
rect -3760 -71 -3750 -37
rect -3750 -71 -3726 -37
rect -3688 -71 -3682 -37
rect -3682 -71 -3654 -37
rect -3616 -71 -3614 -37
rect -3614 -71 -3582 -37
rect -3544 -71 -3512 -37
rect -3512 -71 -3510 -37
rect -3472 -71 -3444 -37
rect -3444 -71 -3438 -37
rect -3400 -71 -3376 -37
rect -3376 -71 -3366 -37
rect -2742 -71 -2732 -37
rect -2732 -71 -2708 -37
rect -2670 -71 -2664 -37
rect -2664 -71 -2636 -37
rect -2598 -71 -2596 -37
rect -2596 -71 -2564 -37
rect -2526 -71 -2494 -37
rect -2494 -71 -2492 -37
rect -2454 -71 -2426 -37
rect -2426 -71 -2420 -37
rect -2382 -71 -2358 -37
rect -2358 -71 -2348 -37
rect -1724 -71 -1714 -37
rect -1714 -71 -1690 -37
rect -1652 -71 -1646 -37
rect -1646 -71 -1618 -37
rect -1580 -71 -1578 -37
rect -1578 -71 -1546 -37
rect -1508 -71 -1476 -37
rect -1476 -71 -1474 -37
rect -1436 -71 -1408 -37
rect -1408 -71 -1402 -37
rect -1364 -71 -1340 -37
rect -1340 -71 -1330 -37
rect -706 -71 -696 -37
rect -696 -71 -672 -37
rect -634 -71 -628 -37
rect -628 -71 -600 -37
rect -562 -71 -560 -37
rect -560 -71 -528 -37
rect -490 -71 -458 -37
rect -458 -71 -456 -37
rect -418 -71 -390 -37
rect -390 -71 -384 -37
rect -346 -71 -322 -37
rect -322 -71 -312 -37
rect 312 -71 322 -37
rect 322 -71 346 -37
rect 384 -71 390 -37
rect 390 -71 418 -37
rect 456 -71 458 -37
rect 458 -71 490 -37
rect 528 -71 560 -37
rect 560 -71 562 -37
rect 600 -71 628 -37
rect 628 -71 634 -37
rect 672 -71 696 -37
rect 696 -71 706 -37
rect 1330 -71 1340 -37
rect 1340 -71 1364 -37
rect 1402 -71 1408 -37
rect 1408 -71 1436 -37
rect 1474 -71 1476 -37
rect 1476 -71 1508 -37
rect 1546 -71 1578 -37
rect 1578 -71 1580 -37
rect 1618 -71 1646 -37
rect 1646 -71 1652 -37
rect 1690 -71 1714 -37
rect 1714 -71 1724 -37
rect 2348 -71 2358 -37
rect 2358 -71 2382 -37
rect 2420 -71 2426 -37
rect 2426 -71 2454 -37
rect 2492 -71 2494 -37
rect 2494 -71 2526 -37
rect 2564 -71 2596 -37
rect 2596 -71 2598 -37
rect 2636 -71 2664 -37
rect 2664 -71 2670 -37
rect 2708 -71 2732 -37
rect 2732 -71 2742 -37
rect 3366 -71 3376 -37
rect 3376 -71 3400 -37
rect 3438 -71 3444 -37
rect 3444 -71 3472 -37
rect 3510 -71 3512 -37
rect 3512 -71 3544 -37
rect 3582 -71 3614 -37
rect 3614 -71 3616 -37
rect 3654 -71 3682 -37
rect 3682 -71 3688 -37
rect 3726 -71 3750 -37
rect 3750 -71 3760 -37
rect 4384 -71 4394 -37
rect 4394 -71 4418 -37
rect 4456 -71 4462 -37
rect 4462 -71 4490 -37
rect 4528 -71 4530 -37
rect 4530 -71 4562 -37
rect 4600 -71 4632 -37
rect 4632 -71 4634 -37
rect 4672 -71 4700 -37
rect 4700 -71 4706 -37
rect 4744 -71 4768 -37
rect 4768 -71 4778 -37
rect 5402 -71 5412 -37
rect 5412 -71 5436 -37
rect 5474 -71 5480 -37
rect 5480 -71 5508 -37
rect 5546 -71 5548 -37
rect 5548 -71 5580 -37
rect 5618 -71 5650 -37
rect 5650 -71 5652 -37
rect 5690 -71 5718 -37
rect 5718 -71 5724 -37
rect 5762 -71 5786 -37
rect 5786 -71 5796 -37
rect 6420 -71 6430 -37
rect 6430 -71 6454 -37
rect 6492 -71 6498 -37
rect 6498 -71 6526 -37
rect 6564 -71 6566 -37
rect 6566 -71 6598 -37
rect 6636 -71 6668 -37
rect 6668 -71 6670 -37
rect 6708 -71 6736 -37
rect 6736 -71 6742 -37
rect 6780 -71 6804 -37
rect 6804 -71 6814 -37
rect 7438 -71 7448 -37
rect 7448 -71 7472 -37
rect 7510 -71 7516 -37
rect 7516 -71 7544 -37
rect 7582 -71 7584 -37
rect 7584 -71 7616 -37
rect 7654 -71 7686 -37
rect 7686 -71 7688 -37
rect 7726 -71 7754 -37
rect 7754 -71 7760 -37
rect 7798 -71 7822 -37
rect 7822 -71 7832 -37
rect 8456 -71 8466 -37
rect 8466 -71 8490 -37
rect 8528 -71 8534 -37
rect 8534 -71 8562 -37
rect 8600 -71 8602 -37
rect 8602 -71 8634 -37
rect 8672 -71 8704 -37
rect 8704 -71 8706 -37
rect 8744 -71 8772 -37
rect 8772 -71 8778 -37
rect 8816 -71 8840 -37
rect 8840 -71 8850 -37
rect 9474 -71 9484 -37
rect 9484 -71 9508 -37
rect 9546 -71 9552 -37
rect 9552 -71 9580 -37
rect 9618 -71 9620 -37
rect 9620 -71 9652 -37
rect 9690 -71 9722 -37
rect 9722 -71 9724 -37
rect 9762 -71 9790 -37
rect 9790 -71 9796 -37
rect 9834 -71 9858 -37
rect 9858 -71 9868 -37
rect -10197 -154 -10163 -140
rect -10197 -174 -10163 -154
rect -10197 -222 -10163 -212
rect -10197 -246 -10163 -222
rect -10197 -290 -10163 -284
rect -10197 -318 -10163 -290
rect -10197 -358 -10163 -356
rect -10197 -390 -10163 -358
rect -10197 -460 -10163 -428
rect -10197 -462 -10163 -460
rect -10197 -528 -10163 -500
rect -10197 -534 -10163 -528
rect -10197 -596 -10163 -572
rect -10197 -606 -10163 -596
rect -10197 -664 -10163 -644
rect -10197 -678 -10163 -664
rect -9179 -154 -9145 -140
rect -9179 -174 -9145 -154
rect -9179 -222 -9145 -212
rect -9179 -246 -9145 -222
rect -9179 -290 -9145 -284
rect -9179 -318 -9145 -290
rect -9179 -358 -9145 -356
rect -9179 -390 -9145 -358
rect -9179 -460 -9145 -428
rect -9179 -462 -9145 -460
rect -9179 -528 -9145 -500
rect -9179 -534 -9145 -528
rect -9179 -596 -9145 -572
rect -9179 -606 -9145 -596
rect -9179 -664 -9145 -644
rect -9179 -678 -9145 -664
rect -8161 -154 -8127 -140
rect -8161 -174 -8127 -154
rect -8161 -222 -8127 -212
rect -8161 -246 -8127 -222
rect -8161 -290 -8127 -284
rect -8161 -318 -8127 -290
rect -8161 -358 -8127 -356
rect -8161 -390 -8127 -358
rect -8161 -460 -8127 -428
rect -8161 -462 -8127 -460
rect -8161 -528 -8127 -500
rect -8161 -534 -8127 -528
rect -8161 -596 -8127 -572
rect -8161 -606 -8127 -596
rect -8161 -664 -8127 -644
rect -8161 -678 -8127 -664
rect -7143 -154 -7109 -140
rect -7143 -174 -7109 -154
rect -7143 -222 -7109 -212
rect -7143 -246 -7109 -222
rect -7143 -290 -7109 -284
rect -7143 -318 -7109 -290
rect -7143 -358 -7109 -356
rect -7143 -390 -7109 -358
rect -7143 -460 -7109 -428
rect -7143 -462 -7109 -460
rect -7143 -528 -7109 -500
rect -7143 -534 -7109 -528
rect -7143 -596 -7109 -572
rect -7143 -606 -7109 -596
rect -7143 -664 -7109 -644
rect -7143 -678 -7109 -664
rect -6125 -154 -6091 -140
rect -6125 -174 -6091 -154
rect -6125 -222 -6091 -212
rect -6125 -246 -6091 -222
rect -6125 -290 -6091 -284
rect -6125 -318 -6091 -290
rect -6125 -358 -6091 -356
rect -6125 -390 -6091 -358
rect -6125 -460 -6091 -428
rect -6125 -462 -6091 -460
rect -6125 -528 -6091 -500
rect -6125 -534 -6091 -528
rect -6125 -596 -6091 -572
rect -6125 -606 -6091 -596
rect -6125 -664 -6091 -644
rect -6125 -678 -6091 -664
rect -5107 -154 -5073 -140
rect -5107 -174 -5073 -154
rect -5107 -222 -5073 -212
rect -5107 -246 -5073 -222
rect -5107 -290 -5073 -284
rect -5107 -318 -5073 -290
rect -5107 -358 -5073 -356
rect -5107 -390 -5073 -358
rect -5107 -460 -5073 -428
rect -5107 -462 -5073 -460
rect -5107 -528 -5073 -500
rect -5107 -534 -5073 -528
rect -5107 -596 -5073 -572
rect -5107 -606 -5073 -596
rect -5107 -664 -5073 -644
rect -5107 -678 -5073 -664
rect -4089 -154 -4055 -140
rect -4089 -174 -4055 -154
rect -4089 -222 -4055 -212
rect -4089 -246 -4055 -222
rect -4089 -290 -4055 -284
rect -4089 -318 -4055 -290
rect -4089 -358 -4055 -356
rect -4089 -390 -4055 -358
rect -4089 -460 -4055 -428
rect -4089 -462 -4055 -460
rect -4089 -528 -4055 -500
rect -4089 -534 -4055 -528
rect -4089 -596 -4055 -572
rect -4089 -606 -4055 -596
rect -4089 -664 -4055 -644
rect -4089 -678 -4055 -664
rect -3071 -154 -3037 -140
rect -3071 -174 -3037 -154
rect -3071 -222 -3037 -212
rect -3071 -246 -3037 -222
rect -3071 -290 -3037 -284
rect -3071 -318 -3037 -290
rect -3071 -358 -3037 -356
rect -3071 -390 -3037 -358
rect -3071 -460 -3037 -428
rect -3071 -462 -3037 -460
rect -3071 -528 -3037 -500
rect -3071 -534 -3037 -528
rect -3071 -596 -3037 -572
rect -3071 -606 -3037 -596
rect -3071 -664 -3037 -644
rect -3071 -678 -3037 -664
rect -2053 -154 -2019 -140
rect -2053 -174 -2019 -154
rect -2053 -222 -2019 -212
rect -2053 -246 -2019 -222
rect -2053 -290 -2019 -284
rect -2053 -318 -2019 -290
rect -2053 -358 -2019 -356
rect -2053 -390 -2019 -358
rect -2053 -460 -2019 -428
rect -2053 -462 -2019 -460
rect -2053 -528 -2019 -500
rect -2053 -534 -2019 -528
rect -2053 -596 -2019 -572
rect -2053 -606 -2019 -596
rect -2053 -664 -2019 -644
rect -2053 -678 -2019 -664
rect -1035 -154 -1001 -140
rect -1035 -174 -1001 -154
rect -1035 -222 -1001 -212
rect -1035 -246 -1001 -222
rect -1035 -290 -1001 -284
rect -1035 -318 -1001 -290
rect -1035 -358 -1001 -356
rect -1035 -390 -1001 -358
rect -1035 -460 -1001 -428
rect -1035 -462 -1001 -460
rect -1035 -528 -1001 -500
rect -1035 -534 -1001 -528
rect -1035 -596 -1001 -572
rect -1035 -606 -1001 -596
rect -1035 -664 -1001 -644
rect -1035 -678 -1001 -664
rect -17 -154 17 -140
rect -17 -174 17 -154
rect -17 -222 17 -212
rect -17 -246 17 -222
rect -17 -290 17 -284
rect -17 -318 17 -290
rect -17 -358 17 -356
rect -17 -390 17 -358
rect -17 -460 17 -428
rect -17 -462 17 -460
rect -17 -528 17 -500
rect -17 -534 17 -528
rect -17 -596 17 -572
rect -17 -606 17 -596
rect -17 -664 17 -644
rect -17 -678 17 -664
rect 1001 -154 1035 -140
rect 1001 -174 1035 -154
rect 1001 -222 1035 -212
rect 1001 -246 1035 -222
rect 1001 -290 1035 -284
rect 1001 -318 1035 -290
rect 1001 -358 1035 -356
rect 1001 -390 1035 -358
rect 1001 -460 1035 -428
rect 1001 -462 1035 -460
rect 1001 -528 1035 -500
rect 1001 -534 1035 -528
rect 1001 -596 1035 -572
rect 1001 -606 1035 -596
rect 1001 -664 1035 -644
rect 1001 -678 1035 -664
rect 2019 -154 2053 -140
rect 2019 -174 2053 -154
rect 2019 -222 2053 -212
rect 2019 -246 2053 -222
rect 2019 -290 2053 -284
rect 2019 -318 2053 -290
rect 2019 -358 2053 -356
rect 2019 -390 2053 -358
rect 2019 -460 2053 -428
rect 2019 -462 2053 -460
rect 2019 -528 2053 -500
rect 2019 -534 2053 -528
rect 2019 -596 2053 -572
rect 2019 -606 2053 -596
rect 2019 -664 2053 -644
rect 2019 -678 2053 -664
rect 3037 -154 3071 -140
rect 3037 -174 3071 -154
rect 3037 -222 3071 -212
rect 3037 -246 3071 -222
rect 3037 -290 3071 -284
rect 3037 -318 3071 -290
rect 3037 -358 3071 -356
rect 3037 -390 3071 -358
rect 3037 -460 3071 -428
rect 3037 -462 3071 -460
rect 3037 -528 3071 -500
rect 3037 -534 3071 -528
rect 3037 -596 3071 -572
rect 3037 -606 3071 -596
rect 3037 -664 3071 -644
rect 3037 -678 3071 -664
rect 4055 -154 4089 -140
rect 4055 -174 4089 -154
rect 4055 -222 4089 -212
rect 4055 -246 4089 -222
rect 4055 -290 4089 -284
rect 4055 -318 4089 -290
rect 4055 -358 4089 -356
rect 4055 -390 4089 -358
rect 4055 -460 4089 -428
rect 4055 -462 4089 -460
rect 4055 -528 4089 -500
rect 4055 -534 4089 -528
rect 4055 -596 4089 -572
rect 4055 -606 4089 -596
rect 4055 -664 4089 -644
rect 4055 -678 4089 -664
rect 5073 -154 5107 -140
rect 5073 -174 5107 -154
rect 5073 -222 5107 -212
rect 5073 -246 5107 -222
rect 5073 -290 5107 -284
rect 5073 -318 5107 -290
rect 5073 -358 5107 -356
rect 5073 -390 5107 -358
rect 5073 -460 5107 -428
rect 5073 -462 5107 -460
rect 5073 -528 5107 -500
rect 5073 -534 5107 -528
rect 5073 -596 5107 -572
rect 5073 -606 5107 -596
rect 5073 -664 5107 -644
rect 5073 -678 5107 -664
rect 6091 -154 6125 -140
rect 6091 -174 6125 -154
rect 6091 -222 6125 -212
rect 6091 -246 6125 -222
rect 6091 -290 6125 -284
rect 6091 -318 6125 -290
rect 6091 -358 6125 -356
rect 6091 -390 6125 -358
rect 6091 -460 6125 -428
rect 6091 -462 6125 -460
rect 6091 -528 6125 -500
rect 6091 -534 6125 -528
rect 6091 -596 6125 -572
rect 6091 -606 6125 -596
rect 6091 -664 6125 -644
rect 6091 -678 6125 -664
rect 7109 -154 7143 -140
rect 7109 -174 7143 -154
rect 7109 -222 7143 -212
rect 7109 -246 7143 -222
rect 7109 -290 7143 -284
rect 7109 -318 7143 -290
rect 7109 -358 7143 -356
rect 7109 -390 7143 -358
rect 7109 -460 7143 -428
rect 7109 -462 7143 -460
rect 7109 -528 7143 -500
rect 7109 -534 7143 -528
rect 7109 -596 7143 -572
rect 7109 -606 7143 -596
rect 7109 -664 7143 -644
rect 7109 -678 7143 -664
rect 8127 -154 8161 -140
rect 8127 -174 8161 -154
rect 8127 -222 8161 -212
rect 8127 -246 8161 -222
rect 8127 -290 8161 -284
rect 8127 -318 8161 -290
rect 8127 -358 8161 -356
rect 8127 -390 8161 -358
rect 8127 -460 8161 -428
rect 8127 -462 8161 -460
rect 8127 -528 8161 -500
rect 8127 -534 8161 -528
rect 8127 -596 8161 -572
rect 8127 -606 8161 -596
rect 8127 -664 8161 -644
rect 8127 -678 8161 -664
rect 9145 -154 9179 -140
rect 9145 -174 9179 -154
rect 9145 -222 9179 -212
rect 9145 -246 9179 -222
rect 9145 -290 9179 -284
rect 9145 -318 9179 -290
rect 9145 -358 9179 -356
rect 9145 -390 9179 -358
rect 9145 -460 9179 -428
rect 9145 -462 9179 -460
rect 9145 -528 9179 -500
rect 9145 -534 9179 -528
rect 9145 -596 9179 -572
rect 9145 -606 9179 -596
rect 9145 -664 9179 -644
rect 9145 -678 9179 -664
rect 10163 -154 10197 -140
rect 10163 -174 10197 -154
rect 10163 -222 10197 -212
rect 10163 -246 10197 -222
rect 10163 -290 10197 -284
rect 10163 -318 10197 -290
rect 10163 -358 10197 -356
rect 10163 -390 10197 -358
rect 10163 -460 10197 -428
rect 10163 -462 10197 -460
rect 10163 -528 10197 -500
rect 10163 -534 10197 -528
rect 10163 -596 10197 -572
rect 10163 -606 10197 -596
rect 10163 -664 10197 -644
rect 10163 -678 10197 -664
rect -9868 -781 -9858 -747
rect -9858 -781 -9834 -747
rect -9796 -781 -9790 -747
rect -9790 -781 -9762 -747
rect -9724 -781 -9722 -747
rect -9722 -781 -9690 -747
rect -9652 -781 -9620 -747
rect -9620 -781 -9618 -747
rect -9580 -781 -9552 -747
rect -9552 -781 -9546 -747
rect -9508 -781 -9484 -747
rect -9484 -781 -9474 -747
rect -8850 -781 -8840 -747
rect -8840 -781 -8816 -747
rect -8778 -781 -8772 -747
rect -8772 -781 -8744 -747
rect -8706 -781 -8704 -747
rect -8704 -781 -8672 -747
rect -8634 -781 -8602 -747
rect -8602 -781 -8600 -747
rect -8562 -781 -8534 -747
rect -8534 -781 -8528 -747
rect -8490 -781 -8466 -747
rect -8466 -781 -8456 -747
rect -7832 -781 -7822 -747
rect -7822 -781 -7798 -747
rect -7760 -781 -7754 -747
rect -7754 -781 -7726 -747
rect -7688 -781 -7686 -747
rect -7686 -781 -7654 -747
rect -7616 -781 -7584 -747
rect -7584 -781 -7582 -747
rect -7544 -781 -7516 -747
rect -7516 -781 -7510 -747
rect -7472 -781 -7448 -747
rect -7448 -781 -7438 -747
rect -6814 -781 -6804 -747
rect -6804 -781 -6780 -747
rect -6742 -781 -6736 -747
rect -6736 -781 -6708 -747
rect -6670 -781 -6668 -747
rect -6668 -781 -6636 -747
rect -6598 -781 -6566 -747
rect -6566 -781 -6564 -747
rect -6526 -781 -6498 -747
rect -6498 -781 -6492 -747
rect -6454 -781 -6430 -747
rect -6430 -781 -6420 -747
rect -5796 -781 -5786 -747
rect -5786 -781 -5762 -747
rect -5724 -781 -5718 -747
rect -5718 -781 -5690 -747
rect -5652 -781 -5650 -747
rect -5650 -781 -5618 -747
rect -5580 -781 -5548 -747
rect -5548 -781 -5546 -747
rect -5508 -781 -5480 -747
rect -5480 -781 -5474 -747
rect -5436 -781 -5412 -747
rect -5412 -781 -5402 -747
rect -4778 -781 -4768 -747
rect -4768 -781 -4744 -747
rect -4706 -781 -4700 -747
rect -4700 -781 -4672 -747
rect -4634 -781 -4632 -747
rect -4632 -781 -4600 -747
rect -4562 -781 -4530 -747
rect -4530 -781 -4528 -747
rect -4490 -781 -4462 -747
rect -4462 -781 -4456 -747
rect -4418 -781 -4394 -747
rect -4394 -781 -4384 -747
rect -3760 -781 -3750 -747
rect -3750 -781 -3726 -747
rect -3688 -781 -3682 -747
rect -3682 -781 -3654 -747
rect -3616 -781 -3614 -747
rect -3614 -781 -3582 -747
rect -3544 -781 -3512 -747
rect -3512 -781 -3510 -747
rect -3472 -781 -3444 -747
rect -3444 -781 -3438 -747
rect -3400 -781 -3376 -747
rect -3376 -781 -3366 -747
rect -2742 -781 -2732 -747
rect -2732 -781 -2708 -747
rect -2670 -781 -2664 -747
rect -2664 -781 -2636 -747
rect -2598 -781 -2596 -747
rect -2596 -781 -2564 -747
rect -2526 -781 -2494 -747
rect -2494 -781 -2492 -747
rect -2454 -781 -2426 -747
rect -2426 -781 -2420 -747
rect -2382 -781 -2358 -747
rect -2358 -781 -2348 -747
rect -1724 -781 -1714 -747
rect -1714 -781 -1690 -747
rect -1652 -781 -1646 -747
rect -1646 -781 -1618 -747
rect -1580 -781 -1578 -747
rect -1578 -781 -1546 -747
rect -1508 -781 -1476 -747
rect -1476 -781 -1474 -747
rect -1436 -781 -1408 -747
rect -1408 -781 -1402 -747
rect -1364 -781 -1340 -747
rect -1340 -781 -1330 -747
rect -706 -781 -696 -747
rect -696 -781 -672 -747
rect -634 -781 -628 -747
rect -628 -781 -600 -747
rect -562 -781 -560 -747
rect -560 -781 -528 -747
rect -490 -781 -458 -747
rect -458 -781 -456 -747
rect -418 -781 -390 -747
rect -390 -781 -384 -747
rect -346 -781 -322 -747
rect -322 -781 -312 -747
rect 312 -781 322 -747
rect 322 -781 346 -747
rect 384 -781 390 -747
rect 390 -781 418 -747
rect 456 -781 458 -747
rect 458 -781 490 -747
rect 528 -781 560 -747
rect 560 -781 562 -747
rect 600 -781 628 -747
rect 628 -781 634 -747
rect 672 -781 696 -747
rect 696 -781 706 -747
rect 1330 -781 1340 -747
rect 1340 -781 1364 -747
rect 1402 -781 1408 -747
rect 1408 -781 1436 -747
rect 1474 -781 1476 -747
rect 1476 -781 1508 -747
rect 1546 -781 1578 -747
rect 1578 -781 1580 -747
rect 1618 -781 1646 -747
rect 1646 -781 1652 -747
rect 1690 -781 1714 -747
rect 1714 -781 1724 -747
rect 2348 -781 2358 -747
rect 2358 -781 2382 -747
rect 2420 -781 2426 -747
rect 2426 -781 2454 -747
rect 2492 -781 2494 -747
rect 2494 -781 2526 -747
rect 2564 -781 2596 -747
rect 2596 -781 2598 -747
rect 2636 -781 2664 -747
rect 2664 -781 2670 -747
rect 2708 -781 2732 -747
rect 2732 -781 2742 -747
rect 3366 -781 3376 -747
rect 3376 -781 3400 -747
rect 3438 -781 3444 -747
rect 3444 -781 3472 -747
rect 3510 -781 3512 -747
rect 3512 -781 3544 -747
rect 3582 -781 3614 -747
rect 3614 -781 3616 -747
rect 3654 -781 3682 -747
rect 3682 -781 3688 -747
rect 3726 -781 3750 -747
rect 3750 -781 3760 -747
rect 4384 -781 4394 -747
rect 4394 -781 4418 -747
rect 4456 -781 4462 -747
rect 4462 -781 4490 -747
rect 4528 -781 4530 -747
rect 4530 -781 4562 -747
rect 4600 -781 4632 -747
rect 4632 -781 4634 -747
rect 4672 -781 4700 -747
rect 4700 -781 4706 -747
rect 4744 -781 4768 -747
rect 4768 -781 4778 -747
rect 5402 -781 5412 -747
rect 5412 -781 5436 -747
rect 5474 -781 5480 -747
rect 5480 -781 5508 -747
rect 5546 -781 5548 -747
rect 5548 -781 5580 -747
rect 5618 -781 5650 -747
rect 5650 -781 5652 -747
rect 5690 -781 5718 -747
rect 5718 -781 5724 -747
rect 5762 -781 5786 -747
rect 5786 -781 5796 -747
rect 6420 -781 6430 -747
rect 6430 -781 6454 -747
rect 6492 -781 6498 -747
rect 6498 -781 6526 -747
rect 6564 -781 6566 -747
rect 6566 -781 6598 -747
rect 6636 -781 6668 -747
rect 6668 -781 6670 -747
rect 6708 -781 6736 -747
rect 6736 -781 6742 -747
rect 6780 -781 6804 -747
rect 6804 -781 6814 -747
rect 7438 -781 7448 -747
rect 7448 -781 7472 -747
rect 7510 -781 7516 -747
rect 7516 -781 7544 -747
rect 7582 -781 7584 -747
rect 7584 -781 7616 -747
rect 7654 -781 7686 -747
rect 7686 -781 7688 -747
rect 7726 -781 7754 -747
rect 7754 -781 7760 -747
rect 7798 -781 7822 -747
rect 7822 -781 7832 -747
rect 8456 -781 8466 -747
rect 8466 -781 8490 -747
rect 8528 -781 8534 -747
rect 8534 -781 8562 -747
rect 8600 -781 8602 -747
rect 8602 -781 8634 -747
rect 8672 -781 8704 -747
rect 8704 -781 8706 -747
rect 8744 -781 8772 -747
rect 8772 -781 8778 -747
rect 8816 -781 8840 -747
rect 8840 -781 8850 -747
rect 9474 -781 9484 -747
rect 9484 -781 9508 -747
rect 9546 -781 9552 -747
rect 9552 -781 9580 -747
rect 9618 -781 9620 -747
rect 9620 -781 9652 -747
rect 9690 -781 9722 -747
rect 9722 -781 9724 -747
rect 9762 -781 9790 -747
rect 9790 -781 9796 -747
rect 9834 -781 9858 -747
rect 9858 -781 9868 -747
<< metal1 >>
rect -9915 781 -9427 787
rect -9915 747 -9868 781
rect -9834 747 -9796 781
rect -9762 747 -9724 781
rect -9690 747 -9652 781
rect -9618 747 -9580 781
rect -9546 747 -9508 781
rect -9474 747 -9427 781
rect -9915 741 -9427 747
rect -8897 781 -8409 787
rect -8897 747 -8850 781
rect -8816 747 -8778 781
rect -8744 747 -8706 781
rect -8672 747 -8634 781
rect -8600 747 -8562 781
rect -8528 747 -8490 781
rect -8456 747 -8409 781
rect -8897 741 -8409 747
rect -7879 781 -7391 787
rect -7879 747 -7832 781
rect -7798 747 -7760 781
rect -7726 747 -7688 781
rect -7654 747 -7616 781
rect -7582 747 -7544 781
rect -7510 747 -7472 781
rect -7438 747 -7391 781
rect -7879 741 -7391 747
rect -6861 781 -6373 787
rect -6861 747 -6814 781
rect -6780 747 -6742 781
rect -6708 747 -6670 781
rect -6636 747 -6598 781
rect -6564 747 -6526 781
rect -6492 747 -6454 781
rect -6420 747 -6373 781
rect -6861 741 -6373 747
rect -5843 781 -5355 787
rect -5843 747 -5796 781
rect -5762 747 -5724 781
rect -5690 747 -5652 781
rect -5618 747 -5580 781
rect -5546 747 -5508 781
rect -5474 747 -5436 781
rect -5402 747 -5355 781
rect -5843 741 -5355 747
rect -4825 781 -4337 787
rect -4825 747 -4778 781
rect -4744 747 -4706 781
rect -4672 747 -4634 781
rect -4600 747 -4562 781
rect -4528 747 -4490 781
rect -4456 747 -4418 781
rect -4384 747 -4337 781
rect -4825 741 -4337 747
rect -3807 781 -3319 787
rect -3807 747 -3760 781
rect -3726 747 -3688 781
rect -3654 747 -3616 781
rect -3582 747 -3544 781
rect -3510 747 -3472 781
rect -3438 747 -3400 781
rect -3366 747 -3319 781
rect -3807 741 -3319 747
rect -2789 781 -2301 787
rect -2789 747 -2742 781
rect -2708 747 -2670 781
rect -2636 747 -2598 781
rect -2564 747 -2526 781
rect -2492 747 -2454 781
rect -2420 747 -2382 781
rect -2348 747 -2301 781
rect -2789 741 -2301 747
rect -1771 781 -1283 787
rect -1771 747 -1724 781
rect -1690 747 -1652 781
rect -1618 747 -1580 781
rect -1546 747 -1508 781
rect -1474 747 -1436 781
rect -1402 747 -1364 781
rect -1330 747 -1283 781
rect -1771 741 -1283 747
rect -753 781 -265 787
rect -753 747 -706 781
rect -672 747 -634 781
rect -600 747 -562 781
rect -528 747 -490 781
rect -456 747 -418 781
rect -384 747 -346 781
rect -312 747 -265 781
rect -753 741 -265 747
rect 265 781 753 787
rect 265 747 312 781
rect 346 747 384 781
rect 418 747 456 781
rect 490 747 528 781
rect 562 747 600 781
rect 634 747 672 781
rect 706 747 753 781
rect 265 741 753 747
rect 1283 781 1771 787
rect 1283 747 1330 781
rect 1364 747 1402 781
rect 1436 747 1474 781
rect 1508 747 1546 781
rect 1580 747 1618 781
rect 1652 747 1690 781
rect 1724 747 1771 781
rect 1283 741 1771 747
rect 2301 781 2789 787
rect 2301 747 2348 781
rect 2382 747 2420 781
rect 2454 747 2492 781
rect 2526 747 2564 781
rect 2598 747 2636 781
rect 2670 747 2708 781
rect 2742 747 2789 781
rect 2301 741 2789 747
rect 3319 781 3807 787
rect 3319 747 3366 781
rect 3400 747 3438 781
rect 3472 747 3510 781
rect 3544 747 3582 781
rect 3616 747 3654 781
rect 3688 747 3726 781
rect 3760 747 3807 781
rect 3319 741 3807 747
rect 4337 781 4825 787
rect 4337 747 4384 781
rect 4418 747 4456 781
rect 4490 747 4528 781
rect 4562 747 4600 781
rect 4634 747 4672 781
rect 4706 747 4744 781
rect 4778 747 4825 781
rect 4337 741 4825 747
rect 5355 781 5843 787
rect 5355 747 5402 781
rect 5436 747 5474 781
rect 5508 747 5546 781
rect 5580 747 5618 781
rect 5652 747 5690 781
rect 5724 747 5762 781
rect 5796 747 5843 781
rect 5355 741 5843 747
rect 6373 781 6861 787
rect 6373 747 6420 781
rect 6454 747 6492 781
rect 6526 747 6564 781
rect 6598 747 6636 781
rect 6670 747 6708 781
rect 6742 747 6780 781
rect 6814 747 6861 781
rect 6373 741 6861 747
rect 7391 781 7879 787
rect 7391 747 7438 781
rect 7472 747 7510 781
rect 7544 747 7582 781
rect 7616 747 7654 781
rect 7688 747 7726 781
rect 7760 747 7798 781
rect 7832 747 7879 781
rect 7391 741 7879 747
rect 8409 781 8897 787
rect 8409 747 8456 781
rect 8490 747 8528 781
rect 8562 747 8600 781
rect 8634 747 8672 781
rect 8706 747 8744 781
rect 8778 747 8816 781
rect 8850 747 8897 781
rect 8409 741 8897 747
rect 9427 781 9915 787
rect 9427 747 9474 781
rect 9508 747 9546 781
rect 9580 747 9618 781
rect 9652 747 9690 781
rect 9724 747 9762 781
rect 9796 747 9834 781
rect 9868 747 9915 781
rect 9427 741 9915 747
rect -10203 678 -10157 709
rect -10203 644 -10197 678
rect -10163 644 -10157 678
rect -10203 606 -10157 644
rect -10203 572 -10197 606
rect -10163 572 -10157 606
rect -10203 534 -10157 572
rect -10203 500 -10197 534
rect -10163 500 -10157 534
rect -10203 462 -10157 500
rect -10203 428 -10197 462
rect -10163 428 -10157 462
rect -10203 390 -10157 428
rect -10203 356 -10197 390
rect -10163 356 -10157 390
rect -10203 318 -10157 356
rect -10203 284 -10197 318
rect -10163 284 -10157 318
rect -10203 246 -10157 284
rect -10203 212 -10197 246
rect -10163 212 -10157 246
rect -10203 174 -10157 212
rect -10203 140 -10197 174
rect -10163 140 -10157 174
rect -10203 109 -10157 140
rect -9185 678 -9139 709
rect -9185 644 -9179 678
rect -9145 644 -9139 678
rect -9185 606 -9139 644
rect -9185 572 -9179 606
rect -9145 572 -9139 606
rect -9185 534 -9139 572
rect -9185 500 -9179 534
rect -9145 500 -9139 534
rect -9185 462 -9139 500
rect -9185 428 -9179 462
rect -9145 428 -9139 462
rect -9185 390 -9139 428
rect -9185 356 -9179 390
rect -9145 356 -9139 390
rect -9185 318 -9139 356
rect -9185 284 -9179 318
rect -9145 284 -9139 318
rect -9185 246 -9139 284
rect -9185 212 -9179 246
rect -9145 212 -9139 246
rect -9185 174 -9139 212
rect -9185 140 -9179 174
rect -9145 140 -9139 174
rect -9185 109 -9139 140
rect -8167 678 -8121 709
rect -8167 644 -8161 678
rect -8127 644 -8121 678
rect -8167 606 -8121 644
rect -8167 572 -8161 606
rect -8127 572 -8121 606
rect -8167 534 -8121 572
rect -8167 500 -8161 534
rect -8127 500 -8121 534
rect -8167 462 -8121 500
rect -8167 428 -8161 462
rect -8127 428 -8121 462
rect -8167 390 -8121 428
rect -8167 356 -8161 390
rect -8127 356 -8121 390
rect -8167 318 -8121 356
rect -8167 284 -8161 318
rect -8127 284 -8121 318
rect -8167 246 -8121 284
rect -8167 212 -8161 246
rect -8127 212 -8121 246
rect -8167 174 -8121 212
rect -8167 140 -8161 174
rect -8127 140 -8121 174
rect -8167 109 -8121 140
rect -7149 678 -7103 709
rect -7149 644 -7143 678
rect -7109 644 -7103 678
rect -7149 606 -7103 644
rect -7149 572 -7143 606
rect -7109 572 -7103 606
rect -7149 534 -7103 572
rect -7149 500 -7143 534
rect -7109 500 -7103 534
rect -7149 462 -7103 500
rect -7149 428 -7143 462
rect -7109 428 -7103 462
rect -7149 390 -7103 428
rect -7149 356 -7143 390
rect -7109 356 -7103 390
rect -7149 318 -7103 356
rect -7149 284 -7143 318
rect -7109 284 -7103 318
rect -7149 246 -7103 284
rect -7149 212 -7143 246
rect -7109 212 -7103 246
rect -7149 174 -7103 212
rect -7149 140 -7143 174
rect -7109 140 -7103 174
rect -7149 109 -7103 140
rect -6131 678 -6085 709
rect -6131 644 -6125 678
rect -6091 644 -6085 678
rect -6131 606 -6085 644
rect -6131 572 -6125 606
rect -6091 572 -6085 606
rect -6131 534 -6085 572
rect -6131 500 -6125 534
rect -6091 500 -6085 534
rect -6131 462 -6085 500
rect -6131 428 -6125 462
rect -6091 428 -6085 462
rect -6131 390 -6085 428
rect -6131 356 -6125 390
rect -6091 356 -6085 390
rect -6131 318 -6085 356
rect -6131 284 -6125 318
rect -6091 284 -6085 318
rect -6131 246 -6085 284
rect -6131 212 -6125 246
rect -6091 212 -6085 246
rect -6131 174 -6085 212
rect -6131 140 -6125 174
rect -6091 140 -6085 174
rect -6131 109 -6085 140
rect -5113 678 -5067 709
rect -5113 644 -5107 678
rect -5073 644 -5067 678
rect -5113 606 -5067 644
rect -5113 572 -5107 606
rect -5073 572 -5067 606
rect -5113 534 -5067 572
rect -5113 500 -5107 534
rect -5073 500 -5067 534
rect -5113 462 -5067 500
rect -5113 428 -5107 462
rect -5073 428 -5067 462
rect -5113 390 -5067 428
rect -5113 356 -5107 390
rect -5073 356 -5067 390
rect -5113 318 -5067 356
rect -5113 284 -5107 318
rect -5073 284 -5067 318
rect -5113 246 -5067 284
rect -5113 212 -5107 246
rect -5073 212 -5067 246
rect -5113 174 -5067 212
rect -5113 140 -5107 174
rect -5073 140 -5067 174
rect -5113 109 -5067 140
rect -4095 678 -4049 709
rect -4095 644 -4089 678
rect -4055 644 -4049 678
rect -4095 606 -4049 644
rect -4095 572 -4089 606
rect -4055 572 -4049 606
rect -4095 534 -4049 572
rect -4095 500 -4089 534
rect -4055 500 -4049 534
rect -4095 462 -4049 500
rect -4095 428 -4089 462
rect -4055 428 -4049 462
rect -4095 390 -4049 428
rect -4095 356 -4089 390
rect -4055 356 -4049 390
rect -4095 318 -4049 356
rect -4095 284 -4089 318
rect -4055 284 -4049 318
rect -4095 246 -4049 284
rect -4095 212 -4089 246
rect -4055 212 -4049 246
rect -4095 174 -4049 212
rect -4095 140 -4089 174
rect -4055 140 -4049 174
rect -4095 109 -4049 140
rect -3077 678 -3031 709
rect -3077 644 -3071 678
rect -3037 644 -3031 678
rect -3077 606 -3031 644
rect -3077 572 -3071 606
rect -3037 572 -3031 606
rect -3077 534 -3031 572
rect -3077 500 -3071 534
rect -3037 500 -3031 534
rect -3077 462 -3031 500
rect -3077 428 -3071 462
rect -3037 428 -3031 462
rect -3077 390 -3031 428
rect -3077 356 -3071 390
rect -3037 356 -3031 390
rect -3077 318 -3031 356
rect -3077 284 -3071 318
rect -3037 284 -3031 318
rect -3077 246 -3031 284
rect -3077 212 -3071 246
rect -3037 212 -3031 246
rect -3077 174 -3031 212
rect -3077 140 -3071 174
rect -3037 140 -3031 174
rect -3077 109 -3031 140
rect -2059 678 -2013 709
rect -2059 644 -2053 678
rect -2019 644 -2013 678
rect -2059 606 -2013 644
rect -2059 572 -2053 606
rect -2019 572 -2013 606
rect -2059 534 -2013 572
rect -2059 500 -2053 534
rect -2019 500 -2013 534
rect -2059 462 -2013 500
rect -2059 428 -2053 462
rect -2019 428 -2013 462
rect -2059 390 -2013 428
rect -2059 356 -2053 390
rect -2019 356 -2013 390
rect -2059 318 -2013 356
rect -2059 284 -2053 318
rect -2019 284 -2013 318
rect -2059 246 -2013 284
rect -2059 212 -2053 246
rect -2019 212 -2013 246
rect -2059 174 -2013 212
rect -2059 140 -2053 174
rect -2019 140 -2013 174
rect -2059 109 -2013 140
rect -1041 678 -995 709
rect -1041 644 -1035 678
rect -1001 644 -995 678
rect -1041 606 -995 644
rect -1041 572 -1035 606
rect -1001 572 -995 606
rect -1041 534 -995 572
rect -1041 500 -1035 534
rect -1001 500 -995 534
rect -1041 462 -995 500
rect -1041 428 -1035 462
rect -1001 428 -995 462
rect -1041 390 -995 428
rect -1041 356 -1035 390
rect -1001 356 -995 390
rect -1041 318 -995 356
rect -1041 284 -1035 318
rect -1001 284 -995 318
rect -1041 246 -995 284
rect -1041 212 -1035 246
rect -1001 212 -995 246
rect -1041 174 -995 212
rect -1041 140 -1035 174
rect -1001 140 -995 174
rect -1041 109 -995 140
rect -23 678 23 709
rect -23 644 -17 678
rect 17 644 23 678
rect -23 606 23 644
rect -23 572 -17 606
rect 17 572 23 606
rect -23 534 23 572
rect -23 500 -17 534
rect 17 500 23 534
rect -23 462 23 500
rect -23 428 -17 462
rect 17 428 23 462
rect -23 390 23 428
rect -23 356 -17 390
rect 17 356 23 390
rect -23 318 23 356
rect -23 284 -17 318
rect 17 284 23 318
rect -23 246 23 284
rect -23 212 -17 246
rect 17 212 23 246
rect -23 174 23 212
rect -23 140 -17 174
rect 17 140 23 174
rect -23 109 23 140
rect 995 678 1041 709
rect 995 644 1001 678
rect 1035 644 1041 678
rect 995 606 1041 644
rect 995 572 1001 606
rect 1035 572 1041 606
rect 995 534 1041 572
rect 995 500 1001 534
rect 1035 500 1041 534
rect 995 462 1041 500
rect 995 428 1001 462
rect 1035 428 1041 462
rect 995 390 1041 428
rect 995 356 1001 390
rect 1035 356 1041 390
rect 995 318 1041 356
rect 995 284 1001 318
rect 1035 284 1041 318
rect 995 246 1041 284
rect 995 212 1001 246
rect 1035 212 1041 246
rect 995 174 1041 212
rect 995 140 1001 174
rect 1035 140 1041 174
rect 995 109 1041 140
rect 2013 678 2059 709
rect 2013 644 2019 678
rect 2053 644 2059 678
rect 2013 606 2059 644
rect 2013 572 2019 606
rect 2053 572 2059 606
rect 2013 534 2059 572
rect 2013 500 2019 534
rect 2053 500 2059 534
rect 2013 462 2059 500
rect 2013 428 2019 462
rect 2053 428 2059 462
rect 2013 390 2059 428
rect 2013 356 2019 390
rect 2053 356 2059 390
rect 2013 318 2059 356
rect 2013 284 2019 318
rect 2053 284 2059 318
rect 2013 246 2059 284
rect 2013 212 2019 246
rect 2053 212 2059 246
rect 2013 174 2059 212
rect 2013 140 2019 174
rect 2053 140 2059 174
rect 2013 109 2059 140
rect 3031 678 3077 709
rect 3031 644 3037 678
rect 3071 644 3077 678
rect 3031 606 3077 644
rect 3031 572 3037 606
rect 3071 572 3077 606
rect 3031 534 3077 572
rect 3031 500 3037 534
rect 3071 500 3077 534
rect 3031 462 3077 500
rect 3031 428 3037 462
rect 3071 428 3077 462
rect 3031 390 3077 428
rect 3031 356 3037 390
rect 3071 356 3077 390
rect 3031 318 3077 356
rect 3031 284 3037 318
rect 3071 284 3077 318
rect 3031 246 3077 284
rect 3031 212 3037 246
rect 3071 212 3077 246
rect 3031 174 3077 212
rect 3031 140 3037 174
rect 3071 140 3077 174
rect 3031 109 3077 140
rect 4049 678 4095 709
rect 4049 644 4055 678
rect 4089 644 4095 678
rect 4049 606 4095 644
rect 4049 572 4055 606
rect 4089 572 4095 606
rect 4049 534 4095 572
rect 4049 500 4055 534
rect 4089 500 4095 534
rect 4049 462 4095 500
rect 4049 428 4055 462
rect 4089 428 4095 462
rect 4049 390 4095 428
rect 4049 356 4055 390
rect 4089 356 4095 390
rect 4049 318 4095 356
rect 4049 284 4055 318
rect 4089 284 4095 318
rect 4049 246 4095 284
rect 4049 212 4055 246
rect 4089 212 4095 246
rect 4049 174 4095 212
rect 4049 140 4055 174
rect 4089 140 4095 174
rect 4049 109 4095 140
rect 5067 678 5113 709
rect 5067 644 5073 678
rect 5107 644 5113 678
rect 5067 606 5113 644
rect 5067 572 5073 606
rect 5107 572 5113 606
rect 5067 534 5113 572
rect 5067 500 5073 534
rect 5107 500 5113 534
rect 5067 462 5113 500
rect 5067 428 5073 462
rect 5107 428 5113 462
rect 5067 390 5113 428
rect 5067 356 5073 390
rect 5107 356 5113 390
rect 5067 318 5113 356
rect 5067 284 5073 318
rect 5107 284 5113 318
rect 5067 246 5113 284
rect 5067 212 5073 246
rect 5107 212 5113 246
rect 5067 174 5113 212
rect 5067 140 5073 174
rect 5107 140 5113 174
rect 5067 109 5113 140
rect 6085 678 6131 709
rect 6085 644 6091 678
rect 6125 644 6131 678
rect 6085 606 6131 644
rect 6085 572 6091 606
rect 6125 572 6131 606
rect 6085 534 6131 572
rect 6085 500 6091 534
rect 6125 500 6131 534
rect 6085 462 6131 500
rect 6085 428 6091 462
rect 6125 428 6131 462
rect 6085 390 6131 428
rect 6085 356 6091 390
rect 6125 356 6131 390
rect 6085 318 6131 356
rect 6085 284 6091 318
rect 6125 284 6131 318
rect 6085 246 6131 284
rect 6085 212 6091 246
rect 6125 212 6131 246
rect 6085 174 6131 212
rect 6085 140 6091 174
rect 6125 140 6131 174
rect 6085 109 6131 140
rect 7103 678 7149 709
rect 7103 644 7109 678
rect 7143 644 7149 678
rect 7103 606 7149 644
rect 7103 572 7109 606
rect 7143 572 7149 606
rect 7103 534 7149 572
rect 7103 500 7109 534
rect 7143 500 7149 534
rect 7103 462 7149 500
rect 7103 428 7109 462
rect 7143 428 7149 462
rect 7103 390 7149 428
rect 7103 356 7109 390
rect 7143 356 7149 390
rect 7103 318 7149 356
rect 7103 284 7109 318
rect 7143 284 7149 318
rect 7103 246 7149 284
rect 7103 212 7109 246
rect 7143 212 7149 246
rect 7103 174 7149 212
rect 7103 140 7109 174
rect 7143 140 7149 174
rect 7103 109 7149 140
rect 8121 678 8167 709
rect 8121 644 8127 678
rect 8161 644 8167 678
rect 8121 606 8167 644
rect 8121 572 8127 606
rect 8161 572 8167 606
rect 8121 534 8167 572
rect 8121 500 8127 534
rect 8161 500 8167 534
rect 8121 462 8167 500
rect 8121 428 8127 462
rect 8161 428 8167 462
rect 8121 390 8167 428
rect 8121 356 8127 390
rect 8161 356 8167 390
rect 8121 318 8167 356
rect 8121 284 8127 318
rect 8161 284 8167 318
rect 8121 246 8167 284
rect 8121 212 8127 246
rect 8161 212 8167 246
rect 8121 174 8167 212
rect 8121 140 8127 174
rect 8161 140 8167 174
rect 8121 109 8167 140
rect 9139 678 9185 709
rect 9139 644 9145 678
rect 9179 644 9185 678
rect 9139 606 9185 644
rect 9139 572 9145 606
rect 9179 572 9185 606
rect 9139 534 9185 572
rect 9139 500 9145 534
rect 9179 500 9185 534
rect 9139 462 9185 500
rect 9139 428 9145 462
rect 9179 428 9185 462
rect 9139 390 9185 428
rect 9139 356 9145 390
rect 9179 356 9185 390
rect 9139 318 9185 356
rect 9139 284 9145 318
rect 9179 284 9185 318
rect 9139 246 9185 284
rect 9139 212 9145 246
rect 9179 212 9185 246
rect 9139 174 9185 212
rect 9139 140 9145 174
rect 9179 140 9185 174
rect 9139 109 9185 140
rect 10157 678 10203 709
rect 10157 644 10163 678
rect 10197 644 10203 678
rect 10157 606 10203 644
rect 10157 572 10163 606
rect 10197 572 10203 606
rect 10157 534 10203 572
rect 10157 500 10163 534
rect 10197 500 10203 534
rect 10157 462 10203 500
rect 10157 428 10163 462
rect 10197 428 10203 462
rect 10157 390 10203 428
rect 10157 356 10163 390
rect 10197 356 10203 390
rect 10157 318 10203 356
rect 10157 284 10163 318
rect 10197 284 10203 318
rect 10157 246 10203 284
rect 10157 212 10163 246
rect 10197 212 10203 246
rect 10157 174 10203 212
rect 10157 140 10163 174
rect 10197 140 10203 174
rect 10157 109 10203 140
rect -9915 71 -9427 77
rect -9915 37 -9868 71
rect -9834 37 -9796 71
rect -9762 37 -9724 71
rect -9690 37 -9652 71
rect -9618 37 -9580 71
rect -9546 37 -9508 71
rect -9474 37 -9427 71
rect -9915 31 -9427 37
rect -8897 71 -8409 77
rect -8897 37 -8850 71
rect -8816 37 -8778 71
rect -8744 37 -8706 71
rect -8672 37 -8634 71
rect -8600 37 -8562 71
rect -8528 37 -8490 71
rect -8456 37 -8409 71
rect -8897 31 -8409 37
rect -7879 71 -7391 77
rect -7879 37 -7832 71
rect -7798 37 -7760 71
rect -7726 37 -7688 71
rect -7654 37 -7616 71
rect -7582 37 -7544 71
rect -7510 37 -7472 71
rect -7438 37 -7391 71
rect -7879 31 -7391 37
rect -6861 71 -6373 77
rect -6861 37 -6814 71
rect -6780 37 -6742 71
rect -6708 37 -6670 71
rect -6636 37 -6598 71
rect -6564 37 -6526 71
rect -6492 37 -6454 71
rect -6420 37 -6373 71
rect -6861 31 -6373 37
rect -5843 71 -5355 77
rect -5843 37 -5796 71
rect -5762 37 -5724 71
rect -5690 37 -5652 71
rect -5618 37 -5580 71
rect -5546 37 -5508 71
rect -5474 37 -5436 71
rect -5402 37 -5355 71
rect -5843 31 -5355 37
rect -4825 71 -4337 77
rect -4825 37 -4778 71
rect -4744 37 -4706 71
rect -4672 37 -4634 71
rect -4600 37 -4562 71
rect -4528 37 -4490 71
rect -4456 37 -4418 71
rect -4384 37 -4337 71
rect -4825 31 -4337 37
rect -3807 71 -3319 77
rect -3807 37 -3760 71
rect -3726 37 -3688 71
rect -3654 37 -3616 71
rect -3582 37 -3544 71
rect -3510 37 -3472 71
rect -3438 37 -3400 71
rect -3366 37 -3319 71
rect -3807 31 -3319 37
rect -2789 71 -2301 77
rect -2789 37 -2742 71
rect -2708 37 -2670 71
rect -2636 37 -2598 71
rect -2564 37 -2526 71
rect -2492 37 -2454 71
rect -2420 37 -2382 71
rect -2348 37 -2301 71
rect -2789 31 -2301 37
rect -1771 71 -1283 77
rect -1771 37 -1724 71
rect -1690 37 -1652 71
rect -1618 37 -1580 71
rect -1546 37 -1508 71
rect -1474 37 -1436 71
rect -1402 37 -1364 71
rect -1330 37 -1283 71
rect -1771 31 -1283 37
rect -753 71 -265 77
rect -753 37 -706 71
rect -672 37 -634 71
rect -600 37 -562 71
rect -528 37 -490 71
rect -456 37 -418 71
rect -384 37 -346 71
rect -312 37 -265 71
rect -753 31 -265 37
rect 265 71 753 77
rect 265 37 312 71
rect 346 37 384 71
rect 418 37 456 71
rect 490 37 528 71
rect 562 37 600 71
rect 634 37 672 71
rect 706 37 753 71
rect 265 31 753 37
rect 1283 71 1771 77
rect 1283 37 1330 71
rect 1364 37 1402 71
rect 1436 37 1474 71
rect 1508 37 1546 71
rect 1580 37 1618 71
rect 1652 37 1690 71
rect 1724 37 1771 71
rect 1283 31 1771 37
rect 2301 71 2789 77
rect 2301 37 2348 71
rect 2382 37 2420 71
rect 2454 37 2492 71
rect 2526 37 2564 71
rect 2598 37 2636 71
rect 2670 37 2708 71
rect 2742 37 2789 71
rect 2301 31 2789 37
rect 3319 71 3807 77
rect 3319 37 3366 71
rect 3400 37 3438 71
rect 3472 37 3510 71
rect 3544 37 3582 71
rect 3616 37 3654 71
rect 3688 37 3726 71
rect 3760 37 3807 71
rect 3319 31 3807 37
rect 4337 71 4825 77
rect 4337 37 4384 71
rect 4418 37 4456 71
rect 4490 37 4528 71
rect 4562 37 4600 71
rect 4634 37 4672 71
rect 4706 37 4744 71
rect 4778 37 4825 71
rect 4337 31 4825 37
rect 5355 71 5843 77
rect 5355 37 5402 71
rect 5436 37 5474 71
rect 5508 37 5546 71
rect 5580 37 5618 71
rect 5652 37 5690 71
rect 5724 37 5762 71
rect 5796 37 5843 71
rect 5355 31 5843 37
rect 6373 71 6861 77
rect 6373 37 6420 71
rect 6454 37 6492 71
rect 6526 37 6564 71
rect 6598 37 6636 71
rect 6670 37 6708 71
rect 6742 37 6780 71
rect 6814 37 6861 71
rect 6373 31 6861 37
rect 7391 71 7879 77
rect 7391 37 7438 71
rect 7472 37 7510 71
rect 7544 37 7582 71
rect 7616 37 7654 71
rect 7688 37 7726 71
rect 7760 37 7798 71
rect 7832 37 7879 71
rect 7391 31 7879 37
rect 8409 71 8897 77
rect 8409 37 8456 71
rect 8490 37 8528 71
rect 8562 37 8600 71
rect 8634 37 8672 71
rect 8706 37 8744 71
rect 8778 37 8816 71
rect 8850 37 8897 71
rect 8409 31 8897 37
rect 9427 71 9915 77
rect 9427 37 9474 71
rect 9508 37 9546 71
rect 9580 37 9618 71
rect 9652 37 9690 71
rect 9724 37 9762 71
rect 9796 37 9834 71
rect 9868 37 9915 71
rect 9427 31 9915 37
rect -9915 -37 -9427 -31
rect -9915 -71 -9868 -37
rect -9834 -71 -9796 -37
rect -9762 -71 -9724 -37
rect -9690 -71 -9652 -37
rect -9618 -71 -9580 -37
rect -9546 -71 -9508 -37
rect -9474 -71 -9427 -37
rect -9915 -77 -9427 -71
rect -8897 -37 -8409 -31
rect -8897 -71 -8850 -37
rect -8816 -71 -8778 -37
rect -8744 -71 -8706 -37
rect -8672 -71 -8634 -37
rect -8600 -71 -8562 -37
rect -8528 -71 -8490 -37
rect -8456 -71 -8409 -37
rect -8897 -77 -8409 -71
rect -7879 -37 -7391 -31
rect -7879 -71 -7832 -37
rect -7798 -71 -7760 -37
rect -7726 -71 -7688 -37
rect -7654 -71 -7616 -37
rect -7582 -71 -7544 -37
rect -7510 -71 -7472 -37
rect -7438 -71 -7391 -37
rect -7879 -77 -7391 -71
rect -6861 -37 -6373 -31
rect -6861 -71 -6814 -37
rect -6780 -71 -6742 -37
rect -6708 -71 -6670 -37
rect -6636 -71 -6598 -37
rect -6564 -71 -6526 -37
rect -6492 -71 -6454 -37
rect -6420 -71 -6373 -37
rect -6861 -77 -6373 -71
rect -5843 -37 -5355 -31
rect -5843 -71 -5796 -37
rect -5762 -71 -5724 -37
rect -5690 -71 -5652 -37
rect -5618 -71 -5580 -37
rect -5546 -71 -5508 -37
rect -5474 -71 -5436 -37
rect -5402 -71 -5355 -37
rect -5843 -77 -5355 -71
rect -4825 -37 -4337 -31
rect -4825 -71 -4778 -37
rect -4744 -71 -4706 -37
rect -4672 -71 -4634 -37
rect -4600 -71 -4562 -37
rect -4528 -71 -4490 -37
rect -4456 -71 -4418 -37
rect -4384 -71 -4337 -37
rect -4825 -77 -4337 -71
rect -3807 -37 -3319 -31
rect -3807 -71 -3760 -37
rect -3726 -71 -3688 -37
rect -3654 -71 -3616 -37
rect -3582 -71 -3544 -37
rect -3510 -71 -3472 -37
rect -3438 -71 -3400 -37
rect -3366 -71 -3319 -37
rect -3807 -77 -3319 -71
rect -2789 -37 -2301 -31
rect -2789 -71 -2742 -37
rect -2708 -71 -2670 -37
rect -2636 -71 -2598 -37
rect -2564 -71 -2526 -37
rect -2492 -71 -2454 -37
rect -2420 -71 -2382 -37
rect -2348 -71 -2301 -37
rect -2789 -77 -2301 -71
rect -1771 -37 -1283 -31
rect -1771 -71 -1724 -37
rect -1690 -71 -1652 -37
rect -1618 -71 -1580 -37
rect -1546 -71 -1508 -37
rect -1474 -71 -1436 -37
rect -1402 -71 -1364 -37
rect -1330 -71 -1283 -37
rect -1771 -77 -1283 -71
rect -753 -37 -265 -31
rect -753 -71 -706 -37
rect -672 -71 -634 -37
rect -600 -71 -562 -37
rect -528 -71 -490 -37
rect -456 -71 -418 -37
rect -384 -71 -346 -37
rect -312 -71 -265 -37
rect -753 -77 -265 -71
rect 265 -37 753 -31
rect 265 -71 312 -37
rect 346 -71 384 -37
rect 418 -71 456 -37
rect 490 -71 528 -37
rect 562 -71 600 -37
rect 634 -71 672 -37
rect 706 -71 753 -37
rect 265 -77 753 -71
rect 1283 -37 1771 -31
rect 1283 -71 1330 -37
rect 1364 -71 1402 -37
rect 1436 -71 1474 -37
rect 1508 -71 1546 -37
rect 1580 -71 1618 -37
rect 1652 -71 1690 -37
rect 1724 -71 1771 -37
rect 1283 -77 1771 -71
rect 2301 -37 2789 -31
rect 2301 -71 2348 -37
rect 2382 -71 2420 -37
rect 2454 -71 2492 -37
rect 2526 -71 2564 -37
rect 2598 -71 2636 -37
rect 2670 -71 2708 -37
rect 2742 -71 2789 -37
rect 2301 -77 2789 -71
rect 3319 -37 3807 -31
rect 3319 -71 3366 -37
rect 3400 -71 3438 -37
rect 3472 -71 3510 -37
rect 3544 -71 3582 -37
rect 3616 -71 3654 -37
rect 3688 -71 3726 -37
rect 3760 -71 3807 -37
rect 3319 -77 3807 -71
rect 4337 -37 4825 -31
rect 4337 -71 4384 -37
rect 4418 -71 4456 -37
rect 4490 -71 4528 -37
rect 4562 -71 4600 -37
rect 4634 -71 4672 -37
rect 4706 -71 4744 -37
rect 4778 -71 4825 -37
rect 4337 -77 4825 -71
rect 5355 -37 5843 -31
rect 5355 -71 5402 -37
rect 5436 -71 5474 -37
rect 5508 -71 5546 -37
rect 5580 -71 5618 -37
rect 5652 -71 5690 -37
rect 5724 -71 5762 -37
rect 5796 -71 5843 -37
rect 5355 -77 5843 -71
rect 6373 -37 6861 -31
rect 6373 -71 6420 -37
rect 6454 -71 6492 -37
rect 6526 -71 6564 -37
rect 6598 -71 6636 -37
rect 6670 -71 6708 -37
rect 6742 -71 6780 -37
rect 6814 -71 6861 -37
rect 6373 -77 6861 -71
rect 7391 -37 7879 -31
rect 7391 -71 7438 -37
rect 7472 -71 7510 -37
rect 7544 -71 7582 -37
rect 7616 -71 7654 -37
rect 7688 -71 7726 -37
rect 7760 -71 7798 -37
rect 7832 -71 7879 -37
rect 7391 -77 7879 -71
rect 8409 -37 8897 -31
rect 8409 -71 8456 -37
rect 8490 -71 8528 -37
rect 8562 -71 8600 -37
rect 8634 -71 8672 -37
rect 8706 -71 8744 -37
rect 8778 -71 8816 -37
rect 8850 -71 8897 -37
rect 8409 -77 8897 -71
rect 9427 -37 9915 -31
rect 9427 -71 9474 -37
rect 9508 -71 9546 -37
rect 9580 -71 9618 -37
rect 9652 -71 9690 -37
rect 9724 -71 9762 -37
rect 9796 -71 9834 -37
rect 9868 -71 9915 -37
rect 9427 -77 9915 -71
rect -10203 -140 -10157 -109
rect -10203 -174 -10197 -140
rect -10163 -174 -10157 -140
rect -10203 -212 -10157 -174
rect -10203 -246 -10197 -212
rect -10163 -246 -10157 -212
rect -10203 -284 -10157 -246
rect -10203 -318 -10197 -284
rect -10163 -318 -10157 -284
rect -10203 -356 -10157 -318
rect -10203 -390 -10197 -356
rect -10163 -390 -10157 -356
rect -10203 -428 -10157 -390
rect -10203 -462 -10197 -428
rect -10163 -462 -10157 -428
rect -10203 -500 -10157 -462
rect -10203 -534 -10197 -500
rect -10163 -534 -10157 -500
rect -10203 -572 -10157 -534
rect -10203 -606 -10197 -572
rect -10163 -606 -10157 -572
rect -10203 -644 -10157 -606
rect -10203 -678 -10197 -644
rect -10163 -678 -10157 -644
rect -10203 -709 -10157 -678
rect -9185 -140 -9139 -109
rect -9185 -174 -9179 -140
rect -9145 -174 -9139 -140
rect -9185 -212 -9139 -174
rect -9185 -246 -9179 -212
rect -9145 -246 -9139 -212
rect -9185 -284 -9139 -246
rect -9185 -318 -9179 -284
rect -9145 -318 -9139 -284
rect -9185 -356 -9139 -318
rect -9185 -390 -9179 -356
rect -9145 -390 -9139 -356
rect -9185 -428 -9139 -390
rect -9185 -462 -9179 -428
rect -9145 -462 -9139 -428
rect -9185 -500 -9139 -462
rect -9185 -534 -9179 -500
rect -9145 -534 -9139 -500
rect -9185 -572 -9139 -534
rect -9185 -606 -9179 -572
rect -9145 -606 -9139 -572
rect -9185 -644 -9139 -606
rect -9185 -678 -9179 -644
rect -9145 -678 -9139 -644
rect -9185 -709 -9139 -678
rect -8167 -140 -8121 -109
rect -8167 -174 -8161 -140
rect -8127 -174 -8121 -140
rect -8167 -212 -8121 -174
rect -8167 -246 -8161 -212
rect -8127 -246 -8121 -212
rect -8167 -284 -8121 -246
rect -8167 -318 -8161 -284
rect -8127 -318 -8121 -284
rect -8167 -356 -8121 -318
rect -8167 -390 -8161 -356
rect -8127 -390 -8121 -356
rect -8167 -428 -8121 -390
rect -8167 -462 -8161 -428
rect -8127 -462 -8121 -428
rect -8167 -500 -8121 -462
rect -8167 -534 -8161 -500
rect -8127 -534 -8121 -500
rect -8167 -572 -8121 -534
rect -8167 -606 -8161 -572
rect -8127 -606 -8121 -572
rect -8167 -644 -8121 -606
rect -8167 -678 -8161 -644
rect -8127 -678 -8121 -644
rect -8167 -709 -8121 -678
rect -7149 -140 -7103 -109
rect -7149 -174 -7143 -140
rect -7109 -174 -7103 -140
rect -7149 -212 -7103 -174
rect -7149 -246 -7143 -212
rect -7109 -246 -7103 -212
rect -7149 -284 -7103 -246
rect -7149 -318 -7143 -284
rect -7109 -318 -7103 -284
rect -7149 -356 -7103 -318
rect -7149 -390 -7143 -356
rect -7109 -390 -7103 -356
rect -7149 -428 -7103 -390
rect -7149 -462 -7143 -428
rect -7109 -462 -7103 -428
rect -7149 -500 -7103 -462
rect -7149 -534 -7143 -500
rect -7109 -534 -7103 -500
rect -7149 -572 -7103 -534
rect -7149 -606 -7143 -572
rect -7109 -606 -7103 -572
rect -7149 -644 -7103 -606
rect -7149 -678 -7143 -644
rect -7109 -678 -7103 -644
rect -7149 -709 -7103 -678
rect -6131 -140 -6085 -109
rect -6131 -174 -6125 -140
rect -6091 -174 -6085 -140
rect -6131 -212 -6085 -174
rect -6131 -246 -6125 -212
rect -6091 -246 -6085 -212
rect -6131 -284 -6085 -246
rect -6131 -318 -6125 -284
rect -6091 -318 -6085 -284
rect -6131 -356 -6085 -318
rect -6131 -390 -6125 -356
rect -6091 -390 -6085 -356
rect -6131 -428 -6085 -390
rect -6131 -462 -6125 -428
rect -6091 -462 -6085 -428
rect -6131 -500 -6085 -462
rect -6131 -534 -6125 -500
rect -6091 -534 -6085 -500
rect -6131 -572 -6085 -534
rect -6131 -606 -6125 -572
rect -6091 -606 -6085 -572
rect -6131 -644 -6085 -606
rect -6131 -678 -6125 -644
rect -6091 -678 -6085 -644
rect -6131 -709 -6085 -678
rect -5113 -140 -5067 -109
rect -5113 -174 -5107 -140
rect -5073 -174 -5067 -140
rect -5113 -212 -5067 -174
rect -5113 -246 -5107 -212
rect -5073 -246 -5067 -212
rect -5113 -284 -5067 -246
rect -5113 -318 -5107 -284
rect -5073 -318 -5067 -284
rect -5113 -356 -5067 -318
rect -5113 -390 -5107 -356
rect -5073 -390 -5067 -356
rect -5113 -428 -5067 -390
rect -5113 -462 -5107 -428
rect -5073 -462 -5067 -428
rect -5113 -500 -5067 -462
rect -5113 -534 -5107 -500
rect -5073 -534 -5067 -500
rect -5113 -572 -5067 -534
rect -5113 -606 -5107 -572
rect -5073 -606 -5067 -572
rect -5113 -644 -5067 -606
rect -5113 -678 -5107 -644
rect -5073 -678 -5067 -644
rect -5113 -709 -5067 -678
rect -4095 -140 -4049 -109
rect -4095 -174 -4089 -140
rect -4055 -174 -4049 -140
rect -4095 -212 -4049 -174
rect -4095 -246 -4089 -212
rect -4055 -246 -4049 -212
rect -4095 -284 -4049 -246
rect -4095 -318 -4089 -284
rect -4055 -318 -4049 -284
rect -4095 -356 -4049 -318
rect -4095 -390 -4089 -356
rect -4055 -390 -4049 -356
rect -4095 -428 -4049 -390
rect -4095 -462 -4089 -428
rect -4055 -462 -4049 -428
rect -4095 -500 -4049 -462
rect -4095 -534 -4089 -500
rect -4055 -534 -4049 -500
rect -4095 -572 -4049 -534
rect -4095 -606 -4089 -572
rect -4055 -606 -4049 -572
rect -4095 -644 -4049 -606
rect -4095 -678 -4089 -644
rect -4055 -678 -4049 -644
rect -4095 -709 -4049 -678
rect -3077 -140 -3031 -109
rect -3077 -174 -3071 -140
rect -3037 -174 -3031 -140
rect -3077 -212 -3031 -174
rect -3077 -246 -3071 -212
rect -3037 -246 -3031 -212
rect -3077 -284 -3031 -246
rect -3077 -318 -3071 -284
rect -3037 -318 -3031 -284
rect -3077 -356 -3031 -318
rect -3077 -390 -3071 -356
rect -3037 -390 -3031 -356
rect -3077 -428 -3031 -390
rect -3077 -462 -3071 -428
rect -3037 -462 -3031 -428
rect -3077 -500 -3031 -462
rect -3077 -534 -3071 -500
rect -3037 -534 -3031 -500
rect -3077 -572 -3031 -534
rect -3077 -606 -3071 -572
rect -3037 -606 -3031 -572
rect -3077 -644 -3031 -606
rect -3077 -678 -3071 -644
rect -3037 -678 -3031 -644
rect -3077 -709 -3031 -678
rect -2059 -140 -2013 -109
rect -2059 -174 -2053 -140
rect -2019 -174 -2013 -140
rect -2059 -212 -2013 -174
rect -2059 -246 -2053 -212
rect -2019 -246 -2013 -212
rect -2059 -284 -2013 -246
rect -2059 -318 -2053 -284
rect -2019 -318 -2013 -284
rect -2059 -356 -2013 -318
rect -2059 -390 -2053 -356
rect -2019 -390 -2013 -356
rect -2059 -428 -2013 -390
rect -2059 -462 -2053 -428
rect -2019 -462 -2013 -428
rect -2059 -500 -2013 -462
rect -2059 -534 -2053 -500
rect -2019 -534 -2013 -500
rect -2059 -572 -2013 -534
rect -2059 -606 -2053 -572
rect -2019 -606 -2013 -572
rect -2059 -644 -2013 -606
rect -2059 -678 -2053 -644
rect -2019 -678 -2013 -644
rect -2059 -709 -2013 -678
rect -1041 -140 -995 -109
rect -1041 -174 -1035 -140
rect -1001 -174 -995 -140
rect -1041 -212 -995 -174
rect -1041 -246 -1035 -212
rect -1001 -246 -995 -212
rect -1041 -284 -995 -246
rect -1041 -318 -1035 -284
rect -1001 -318 -995 -284
rect -1041 -356 -995 -318
rect -1041 -390 -1035 -356
rect -1001 -390 -995 -356
rect -1041 -428 -995 -390
rect -1041 -462 -1035 -428
rect -1001 -462 -995 -428
rect -1041 -500 -995 -462
rect -1041 -534 -1035 -500
rect -1001 -534 -995 -500
rect -1041 -572 -995 -534
rect -1041 -606 -1035 -572
rect -1001 -606 -995 -572
rect -1041 -644 -995 -606
rect -1041 -678 -1035 -644
rect -1001 -678 -995 -644
rect -1041 -709 -995 -678
rect -23 -140 23 -109
rect -23 -174 -17 -140
rect 17 -174 23 -140
rect -23 -212 23 -174
rect -23 -246 -17 -212
rect 17 -246 23 -212
rect -23 -284 23 -246
rect -23 -318 -17 -284
rect 17 -318 23 -284
rect -23 -356 23 -318
rect -23 -390 -17 -356
rect 17 -390 23 -356
rect -23 -428 23 -390
rect -23 -462 -17 -428
rect 17 -462 23 -428
rect -23 -500 23 -462
rect -23 -534 -17 -500
rect 17 -534 23 -500
rect -23 -572 23 -534
rect -23 -606 -17 -572
rect 17 -606 23 -572
rect -23 -644 23 -606
rect -23 -678 -17 -644
rect 17 -678 23 -644
rect -23 -709 23 -678
rect 995 -140 1041 -109
rect 995 -174 1001 -140
rect 1035 -174 1041 -140
rect 995 -212 1041 -174
rect 995 -246 1001 -212
rect 1035 -246 1041 -212
rect 995 -284 1041 -246
rect 995 -318 1001 -284
rect 1035 -318 1041 -284
rect 995 -356 1041 -318
rect 995 -390 1001 -356
rect 1035 -390 1041 -356
rect 995 -428 1041 -390
rect 995 -462 1001 -428
rect 1035 -462 1041 -428
rect 995 -500 1041 -462
rect 995 -534 1001 -500
rect 1035 -534 1041 -500
rect 995 -572 1041 -534
rect 995 -606 1001 -572
rect 1035 -606 1041 -572
rect 995 -644 1041 -606
rect 995 -678 1001 -644
rect 1035 -678 1041 -644
rect 995 -709 1041 -678
rect 2013 -140 2059 -109
rect 2013 -174 2019 -140
rect 2053 -174 2059 -140
rect 2013 -212 2059 -174
rect 2013 -246 2019 -212
rect 2053 -246 2059 -212
rect 2013 -284 2059 -246
rect 2013 -318 2019 -284
rect 2053 -318 2059 -284
rect 2013 -356 2059 -318
rect 2013 -390 2019 -356
rect 2053 -390 2059 -356
rect 2013 -428 2059 -390
rect 2013 -462 2019 -428
rect 2053 -462 2059 -428
rect 2013 -500 2059 -462
rect 2013 -534 2019 -500
rect 2053 -534 2059 -500
rect 2013 -572 2059 -534
rect 2013 -606 2019 -572
rect 2053 -606 2059 -572
rect 2013 -644 2059 -606
rect 2013 -678 2019 -644
rect 2053 -678 2059 -644
rect 2013 -709 2059 -678
rect 3031 -140 3077 -109
rect 3031 -174 3037 -140
rect 3071 -174 3077 -140
rect 3031 -212 3077 -174
rect 3031 -246 3037 -212
rect 3071 -246 3077 -212
rect 3031 -284 3077 -246
rect 3031 -318 3037 -284
rect 3071 -318 3077 -284
rect 3031 -356 3077 -318
rect 3031 -390 3037 -356
rect 3071 -390 3077 -356
rect 3031 -428 3077 -390
rect 3031 -462 3037 -428
rect 3071 -462 3077 -428
rect 3031 -500 3077 -462
rect 3031 -534 3037 -500
rect 3071 -534 3077 -500
rect 3031 -572 3077 -534
rect 3031 -606 3037 -572
rect 3071 -606 3077 -572
rect 3031 -644 3077 -606
rect 3031 -678 3037 -644
rect 3071 -678 3077 -644
rect 3031 -709 3077 -678
rect 4049 -140 4095 -109
rect 4049 -174 4055 -140
rect 4089 -174 4095 -140
rect 4049 -212 4095 -174
rect 4049 -246 4055 -212
rect 4089 -246 4095 -212
rect 4049 -284 4095 -246
rect 4049 -318 4055 -284
rect 4089 -318 4095 -284
rect 4049 -356 4095 -318
rect 4049 -390 4055 -356
rect 4089 -390 4095 -356
rect 4049 -428 4095 -390
rect 4049 -462 4055 -428
rect 4089 -462 4095 -428
rect 4049 -500 4095 -462
rect 4049 -534 4055 -500
rect 4089 -534 4095 -500
rect 4049 -572 4095 -534
rect 4049 -606 4055 -572
rect 4089 -606 4095 -572
rect 4049 -644 4095 -606
rect 4049 -678 4055 -644
rect 4089 -678 4095 -644
rect 4049 -709 4095 -678
rect 5067 -140 5113 -109
rect 5067 -174 5073 -140
rect 5107 -174 5113 -140
rect 5067 -212 5113 -174
rect 5067 -246 5073 -212
rect 5107 -246 5113 -212
rect 5067 -284 5113 -246
rect 5067 -318 5073 -284
rect 5107 -318 5113 -284
rect 5067 -356 5113 -318
rect 5067 -390 5073 -356
rect 5107 -390 5113 -356
rect 5067 -428 5113 -390
rect 5067 -462 5073 -428
rect 5107 -462 5113 -428
rect 5067 -500 5113 -462
rect 5067 -534 5073 -500
rect 5107 -534 5113 -500
rect 5067 -572 5113 -534
rect 5067 -606 5073 -572
rect 5107 -606 5113 -572
rect 5067 -644 5113 -606
rect 5067 -678 5073 -644
rect 5107 -678 5113 -644
rect 5067 -709 5113 -678
rect 6085 -140 6131 -109
rect 6085 -174 6091 -140
rect 6125 -174 6131 -140
rect 6085 -212 6131 -174
rect 6085 -246 6091 -212
rect 6125 -246 6131 -212
rect 6085 -284 6131 -246
rect 6085 -318 6091 -284
rect 6125 -318 6131 -284
rect 6085 -356 6131 -318
rect 6085 -390 6091 -356
rect 6125 -390 6131 -356
rect 6085 -428 6131 -390
rect 6085 -462 6091 -428
rect 6125 -462 6131 -428
rect 6085 -500 6131 -462
rect 6085 -534 6091 -500
rect 6125 -534 6131 -500
rect 6085 -572 6131 -534
rect 6085 -606 6091 -572
rect 6125 -606 6131 -572
rect 6085 -644 6131 -606
rect 6085 -678 6091 -644
rect 6125 -678 6131 -644
rect 6085 -709 6131 -678
rect 7103 -140 7149 -109
rect 7103 -174 7109 -140
rect 7143 -174 7149 -140
rect 7103 -212 7149 -174
rect 7103 -246 7109 -212
rect 7143 -246 7149 -212
rect 7103 -284 7149 -246
rect 7103 -318 7109 -284
rect 7143 -318 7149 -284
rect 7103 -356 7149 -318
rect 7103 -390 7109 -356
rect 7143 -390 7149 -356
rect 7103 -428 7149 -390
rect 7103 -462 7109 -428
rect 7143 -462 7149 -428
rect 7103 -500 7149 -462
rect 7103 -534 7109 -500
rect 7143 -534 7149 -500
rect 7103 -572 7149 -534
rect 7103 -606 7109 -572
rect 7143 -606 7149 -572
rect 7103 -644 7149 -606
rect 7103 -678 7109 -644
rect 7143 -678 7149 -644
rect 7103 -709 7149 -678
rect 8121 -140 8167 -109
rect 8121 -174 8127 -140
rect 8161 -174 8167 -140
rect 8121 -212 8167 -174
rect 8121 -246 8127 -212
rect 8161 -246 8167 -212
rect 8121 -284 8167 -246
rect 8121 -318 8127 -284
rect 8161 -318 8167 -284
rect 8121 -356 8167 -318
rect 8121 -390 8127 -356
rect 8161 -390 8167 -356
rect 8121 -428 8167 -390
rect 8121 -462 8127 -428
rect 8161 -462 8167 -428
rect 8121 -500 8167 -462
rect 8121 -534 8127 -500
rect 8161 -534 8167 -500
rect 8121 -572 8167 -534
rect 8121 -606 8127 -572
rect 8161 -606 8167 -572
rect 8121 -644 8167 -606
rect 8121 -678 8127 -644
rect 8161 -678 8167 -644
rect 8121 -709 8167 -678
rect 9139 -140 9185 -109
rect 9139 -174 9145 -140
rect 9179 -174 9185 -140
rect 9139 -212 9185 -174
rect 9139 -246 9145 -212
rect 9179 -246 9185 -212
rect 9139 -284 9185 -246
rect 9139 -318 9145 -284
rect 9179 -318 9185 -284
rect 9139 -356 9185 -318
rect 9139 -390 9145 -356
rect 9179 -390 9185 -356
rect 9139 -428 9185 -390
rect 9139 -462 9145 -428
rect 9179 -462 9185 -428
rect 9139 -500 9185 -462
rect 9139 -534 9145 -500
rect 9179 -534 9185 -500
rect 9139 -572 9185 -534
rect 9139 -606 9145 -572
rect 9179 -606 9185 -572
rect 9139 -644 9185 -606
rect 9139 -678 9145 -644
rect 9179 -678 9185 -644
rect 9139 -709 9185 -678
rect 10157 -140 10203 -109
rect 10157 -174 10163 -140
rect 10197 -174 10203 -140
rect 10157 -212 10203 -174
rect 10157 -246 10163 -212
rect 10197 -246 10203 -212
rect 10157 -284 10203 -246
rect 10157 -318 10163 -284
rect 10197 -318 10203 -284
rect 10157 -356 10203 -318
rect 10157 -390 10163 -356
rect 10197 -390 10203 -356
rect 10157 -428 10203 -390
rect 10157 -462 10163 -428
rect 10197 -462 10203 -428
rect 10157 -500 10203 -462
rect 10157 -534 10163 -500
rect 10197 -534 10203 -500
rect 10157 -572 10203 -534
rect 10157 -606 10163 -572
rect 10197 -606 10203 -572
rect 10157 -644 10203 -606
rect 10157 -678 10163 -644
rect 10197 -678 10203 -644
rect 10157 -709 10203 -678
rect -9915 -747 -9427 -741
rect -9915 -781 -9868 -747
rect -9834 -781 -9796 -747
rect -9762 -781 -9724 -747
rect -9690 -781 -9652 -747
rect -9618 -781 -9580 -747
rect -9546 -781 -9508 -747
rect -9474 -781 -9427 -747
rect -9915 -787 -9427 -781
rect -8897 -747 -8409 -741
rect -8897 -781 -8850 -747
rect -8816 -781 -8778 -747
rect -8744 -781 -8706 -747
rect -8672 -781 -8634 -747
rect -8600 -781 -8562 -747
rect -8528 -781 -8490 -747
rect -8456 -781 -8409 -747
rect -8897 -787 -8409 -781
rect -7879 -747 -7391 -741
rect -7879 -781 -7832 -747
rect -7798 -781 -7760 -747
rect -7726 -781 -7688 -747
rect -7654 -781 -7616 -747
rect -7582 -781 -7544 -747
rect -7510 -781 -7472 -747
rect -7438 -781 -7391 -747
rect -7879 -787 -7391 -781
rect -6861 -747 -6373 -741
rect -6861 -781 -6814 -747
rect -6780 -781 -6742 -747
rect -6708 -781 -6670 -747
rect -6636 -781 -6598 -747
rect -6564 -781 -6526 -747
rect -6492 -781 -6454 -747
rect -6420 -781 -6373 -747
rect -6861 -787 -6373 -781
rect -5843 -747 -5355 -741
rect -5843 -781 -5796 -747
rect -5762 -781 -5724 -747
rect -5690 -781 -5652 -747
rect -5618 -781 -5580 -747
rect -5546 -781 -5508 -747
rect -5474 -781 -5436 -747
rect -5402 -781 -5355 -747
rect -5843 -787 -5355 -781
rect -4825 -747 -4337 -741
rect -4825 -781 -4778 -747
rect -4744 -781 -4706 -747
rect -4672 -781 -4634 -747
rect -4600 -781 -4562 -747
rect -4528 -781 -4490 -747
rect -4456 -781 -4418 -747
rect -4384 -781 -4337 -747
rect -4825 -787 -4337 -781
rect -3807 -747 -3319 -741
rect -3807 -781 -3760 -747
rect -3726 -781 -3688 -747
rect -3654 -781 -3616 -747
rect -3582 -781 -3544 -747
rect -3510 -781 -3472 -747
rect -3438 -781 -3400 -747
rect -3366 -781 -3319 -747
rect -3807 -787 -3319 -781
rect -2789 -747 -2301 -741
rect -2789 -781 -2742 -747
rect -2708 -781 -2670 -747
rect -2636 -781 -2598 -747
rect -2564 -781 -2526 -747
rect -2492 -781 -2454 -747
rect -2420 -781 -2382 -747
rect -2348 -781 -2301 -747
rect -2789 -787 -2301 -781
rect -1771 -747 -1283 -741
rect -1771 -781 -1724 -747
rect -1690 -781 -1652 -747
rect -1618 -781 -1580 -747
rect -1546 -781 -1508 -747
rect -1474 -781 -1436 -747
rect -1402 -781 -1364 -747
rect -1330 -781 -1283 -747
rect -1771 -787 -1283 -781
rect -753 -747 -265 -741
rect -753 -781 -706 -747
rect -672 -781 -634 -747
rect -600 -781 -562 -747
rect -528 -781 -490 -747
rect -456 -781 -418 -747
rect -384 -781 -346 -747
rect -312 -781 -265 -747
rect -753 -787 -265 -781
rect 265 -747 753 -741
rect 265 -781 312 -747
rect 346 -781 384 -747
rect 418 -781 456 -747
rect 490 -781 528 -747
rect 562 -781 600 -747
rect 634 -781 672 -747
rect 706 -781 753 -747
rect 265 -787 753 -781
rect 1283 -747 1771 -741
rect 1283 -781 1330 -747
rect 1364 -781 1402 -747
rect 1436 -781 1474 -747
rect 1508 -781 1546 -747
rect 1580 -781 1618 -747
rect 1652 -781 1690 -747
rect 1724 -781 1771 -747
rect 1283 -787 1771 -781
rect 2301 -747 2789 -741
rect 2301 -781 2348 -747
rect 2382 -781 2420 -747
rect 2454 -781 2492 -747
rect 2526 -781 2564 -747
rect 2598 -781 2636 -747
rect 2670 -781 2708 -747
rect 2742 -781 2789 -747
rect 2301 -787 2789 -781
rect 3319 -747 3807 -741
rect 3319 -781 3366 -747
rect 3400 -781 3438 -747
rect 3472 -781 3510 -747
rect 3544 -781 3582 -747
rect 3616 -781 3654 -747
rect 3688 -781 3726 -747
rect 3760 -781 3807 -747
rect 3319 -787 3807 -781
rect 4337 -747 4825 -741
rect 4337 -781 4384 -747
rect 4418 -781 4456 -747
rect 4490 -781 4528 -747
rect 4562 -781 4600 -747
rect 4634 -781 4672 -747
rect 4706 -781 4744 -747
rect 4778 -781 4825 -747
rect 4337 -787 4825 -781
rect 5355 -747 5843 -741
rect 5355 -781 5402 -747
rect 5436 -781 5474 -747
rect 5508 -781 5546 -747
rect 5580 -781 5618 -747
rect 5652 -781 5690 -747
rect 5724 -781 5762 -747
rect 5796 -781 5843 -747
rect 5355 -787 5843 -781
rect 6373 -747 6861 -741
rect 6373 -781 6420 -747
rect 6454 -781 6492 -747
rect 6526 -781 6564 -747
rect 6598 -781 6636 -747
rect 6670 -781 6708 -747
rect 6742 -781 6780 -747
rect 6814 -781 6861 -747
rect 6373 -787 6861 -781
rect 7391 -747 7879 -741
rect 7391 -781 7438 -747
rect 7472 -781 7510 -747
rect 7544 -781 7582 -747
rect 7616 -781 7654 -747
rect 7688 -781 7726 -747
rect 7760 -781 7798 -747
rect 7832 -781 7879 -747
rect 7391 -787 7879 -781
rect 8409 -747 8897 -741
rect 8409 -781 8456 -747
rect 8490 -781 8528 -747
rect 8562 -781 8600 -747
rect 8634 -781 8672 -747
rect 8706 -781 8744 -747
rect 8778 -781 8816 -747
rect 8850 -781 8897 -747
rect 8409 -787 8897 -781
rect 9427 -747 9915 -741
rect 9427 -781 9474 -747
rect 9508 -781 9546 -747
rect 9580 -781 9618 -747
rect 9652 -781 9690 -747
rect 9724 -781 9762 -747
rect 9796 -781 9834 -747
rect 9868 -781 9915 -747
rect 9427 -787 9915 -781
<< end >>
