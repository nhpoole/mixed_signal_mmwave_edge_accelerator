magic
tech sky130A
timestamp 1626065694
<< checkpaint >>
rect -717 -717 717 717
<< metal4 >>
rect -87 59 87 87
rect -87 -59 -59 59
rect 59 -59 87 59
rect -87 -87 87 -59
<< via4 >>
rect -59 -59 59 59
<< metal5 >>
rect -87 59 87 87
rect -87 -59 -59 59
rect 59 -59 87 59
rect -87 -87 87 -59
<< end >>
