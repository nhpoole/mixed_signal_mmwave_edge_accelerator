* Stimulus file.

.param Itail=1u Ibias=1u vcmdes=1 vincm=1 vsig=0 vdd=1.8 Wp=16 Wn=2 Wpcm=64 Wncm=4 Wbias=1
+ Lbias=3.2 nfactorL=1 nfactorW=6 K=1 K2=0.5

vdd VDD GND 'vdd'
vip vip GND dc 'vincm+vsig' ac 0.5 0
vim vim GND dc 'vincm-vsig' ac 0.5 180
vocm vocm GND 'vcmdes'

.control
options savecurrents
save all
+ @m.xm5.msky130_fd_pr__nfet_01v8[id]
+ @m.xm5.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm7.msky130_fd_pr__nfet_01v8[id]
+ @m.xm7.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm10.msky130_fd_pr__nfet_01v8[id]
+ @m.xm10.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm12.msky130_fd_pr__pfet_01v8[id]
+ @m.xm12.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm12.msky130_fd_pr__pfet_01v8[cgd]
+ @m.xm15.msky130_fd_pr__pfet_01v8_lvt[id]
+ @m.xm15.msky130_fd_pr__pfet_01v8_lvt[vth]
+ @m.xm15.msky130_fd_pr__pfet_01v8_lvt[cgd]
+ @m.xm27.msky130_fd_pr__nfet_01v8[id]
+ @m.xm27.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm31.msky130_fd_pr__pfet_01v8[id]
+ @m.xm31.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm31.msky130_fd_pr__pfet_01v8[cgd]
+ @m.xm32.msky130_fd_pr__pfet_01v8_lvt[id]
+ @m.xm32.msky130_fd_pr__pfet_01v8_lvt[vth]
+ @m.xm32.msky130_fd_pr__pfet_01v8_lvt[cgd]
+ @m.xm33.msky130_fd_pr__pfet_01v8_lvt[id]
+ @m.xm33.msky130_fd_pr__pfet_01v8_lvt[vth]
+ @m.xm34.msky130_fd_pr__pfet_01v8_lvt[id]
+ @m.xm34.msky130_fd_pr__pfet_01v8_lvt[vth]
+ @m.xm35.msky130_fd_pr__pfet_01v8_lvt[id]
+ @m.xm35.msky130_fd_pr__pfet_01v8_lvt[vth]
+ @m.xm36.msky130_fd_pr__pfet_01v8[id]
+ @m.xm36.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm37.msky130_fd_pr__pfet_01v8[id]
+ @m.xm37.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm38.msky130_fd_pr__pfet_01v8[id]
+ @m.xm38.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm39.msky130_fd_pr__pfet_01v8[id]
+ @m.xm39.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm40.msky130_fd_pr__pfet_01v8[id]
+ @m.xm40.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm41.msky130_fd_pr__nfet_01v8[id]
+ @m.xm41.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm42.msky130_fd_pr__nfet_01v8[id]
+ @m.xm42.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm43.msky130_fd_pr__nfet_01v8[id]
+ @m.xm43.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm44.msky130_fd_pr__nfet_01v8[id]
+ @m.xm44.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm45.msky130_fd_pr__nfet_01v8[id]
+ @m.xm45.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm51.msky130_fd_pr__nfet_01v8_lvt[id]
+ @m.xm51.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @m.xm51.msky130_fd_pr__nfet_01v8_lvt[cgd]
+ @m.xm53.msky130_fd_pr__nfet_01v8_lvt[id]
+ @m.xm53.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @m.xm53.msky130_fd_pr__nfet_01v8_lvt[cgd]

+ @m.xm1.msky130_fd_pr__pfet_01v8_lvt[id]
+ @m.xm1.msky130_fd_pr__pfet_01v8_lvt[vth]
+ @m.xm1.msky130_fd_pr__pfet_01v8_lvt[cgd]
+ @m.xm2.msky130_fd_pr__nfet_01v8[id]
+ @m.xm2.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm3.msky130_fd_pr__pfet_01v8_lvt[id]
+ @m.xm3.msky130_fd_pr__pfet_01v8_lvt[vth]
+ @m.xm3.msky130_fd_pr__pfet_01v8_lvt[cgd]
+ @m.xm4.msky130_fd_pr__nfet_01v8[id]
+ @m.xm4.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm6.msky130_fd_pr__pfet_01v8[id]
+ @m.xm6.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm8.msky130_fd_pr__nfet_01v8[id]
+ @m.xm8.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm8.msky130_fd_pr__nfet_01v8[cgd]
+ @m.xm9.msky130_fd_pr__nfet_01v8[id]
+ @m.xm9.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm9.msky130_fd_pr__nfet_01v8[cgd]
+ @m.xm11.msky130_fd_pr__nfet_01v8[id]
+ @m.xm11.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm11.msky130_fd_pr__nfet_01v8[cgd]
+ @m.xm13.msky130_fd_pr__pfet_01v8_lvt[id]
+ @m.xm13.msky130_fd_pr__pfet_01v8_lvt[vth]
+ @m.xm14.msky130_fd_pr__pfet_01v8_lvt[id]
+ @m.xm14.msky130_fd_pr__pfet_01v8_lvt[vth]
+ @m.xm16.msky130_fd_pr__pfet_01v8[id]
+ @m.xm16.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm17.msky130_fd_pr__nfet_01v8_lvt[id]
+ @m.xm17.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @m.xm18.msky130_fd_pr__nfet_01v8_lvt[id]
+ @m.xm18.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @m.xm19.msky130_fd_pr__nfet_01v8_lvt[id]
+ @m.xm19.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @m.xm20.msky130_fd_pr__nfet_01v8_lvt[id]
+ @m.xm20.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @m.xm21.msky130_fd_pr__nfet_01v8[id]
+ @m.xm21.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm22.msky130_fd_pr__nfet_01v8[id]
+ @m.xm22.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm23.msky130_fd_pr__pfet_01v8[id]
+ @m.xm23.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm24.msky130_fd_pr__pfet_01v8[id]
+ @m.xm24.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm25.msky130_fd_pr__pfet_01v8[id]
+ @m.xm25.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm26.msky130_fd_pr__nfet_01v8[id]
+ @m.xm26.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm28.msky130_fd_pr__nfet_01v8[id]
+ @m.xm28.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm28.msky130_fd_pr__nfet_01v8[cgd]
+ @m.xm29.msky130_fd_pr__nfet_01v8[id]
+ @m.xm29.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm30.msky130_fd_pr__pfet_01v8[id]
+ @m.xm30.msky130_fd_pr__pfet_01v8[vth]

op
run
print all
write diff_fold_casc_ota_twostage_op.raw

*dc vip 0.5 1.5 0.01
*run
*write diff_fold_casc_ota_dc.raw

ac dec 100 0.1 1g
*save v(vop_casc) v(vom_casc)
*plot v(vop) v(vom) vm(vop) vm(vom) vp(vop) vp(vom) vdb(vop) vdb(vom)
run
write diff_fold_casc_ota_twostage_ac.raw
quit
.endc