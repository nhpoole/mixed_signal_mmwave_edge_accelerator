magic
tech sky130A
magscale 1 2
timestamp 1624185512
<< nwell >>
rect 17382 14696 41898 29438
<< pwell >>
rect -238 -2078 4438 978
rect 4682 -2178 41998 13938
<< nmos >>
rect 332 42 532 442
rect 590 42 790 442
rect 848 42 1048 442
rect 1106 42 1306 442
rect 1364 42 1564 442
rect 1622 42 1822 442
rect 1880 42 2080 442
rect 2138 42 2338 442
rect 2396 42 2596 442
rect 2654 42 2854 442
rect 2912 42 3112 442
rect 3170 42 3370 442
rect 3428 42 3628 442
rect 3686 42 3886 442
rect 332 -958 532 -558
rect 590 -958 790 -558
rect 848 -958 1048 -558
rect 1106 -958 1306 -558
rect 1364 -958 1564 -558
rect 1622 -958 1822 -558
rect 1880 -958 2080 -558
rect 2138 -958 2338 -558
rect 2396 -958 2596 -558
rect 2654 -958 2854 -558
rect 2912 -958 3112 -558
rect 3170 -958 3370 -558
rect 3428 -958 3628 -558
rect 3686 -958 3886 -558
rect 19668 12444 20628 13044
rect 20686 12444 21646 13044
rect 21704 12444 22664 13044
rect 22722 12444 23682 13044
rect 23740 12444 24700 13044
rect 24758 12444 25718 13044
rect 25776 12444 26736 13044
rect 26794 12444 27754 13044
rect 27812 12444 28772 13044
rect 28830 12444 29790 13044
rect 29848 12444 30808 13044
rect 30866 12444 31826 13044
rect 31884 12444 32844 13044
rect 32902 12444 33862 13044
rect 33920 12444 34880 13044
rect 34938 12444 35898 13044
rect 35956 12444 36916 13044
rect 36974 12444 37934 13044
rect 37992 12444 38952 13044
rect 39010 12444 39970 13044
rect 19668 11626 20628 12226
rect 20686 11626 21646 12226
rect 21704 11626 22664 12226
rect 22722 11626 23682 12226
rect 23740 11626 24700 12226
rect 24758 11626 25718 12226
rect 25776 11626 26736 12226
rect 26794 11626 27754 12226
rect 27812 11626 28772 12226
rect 28830 11626 29790 12226
rect 29848 11626 30808 12226
rect 30866 11626 31826 12226
rect 31884 11626 32844 12226
rect 32902 11626 33862 12226
rect 33920 11626 34880 12226
rect 34938 11626 35898 12226
rect 35956 11626 36916 12226
rect 36974 11626 37934 12226
rect 37992 11626 38952 12226
rect 39010 11626 39970 12226
rect 19668 10248 20628 10848
rect 20686 10248 21646 10848
rect 21704 10248 22664 10848
rect 22722 10248 23682 10848
rect 23740 10248 24700 10848
rect 24758 10248 25718 10848
rect 25776 10248 26736 10848
rect 26794 10248 27754 10848
rect 27812 10248 28772 10848
rect 28830 10248 29790 10848
rect 29848 10248 30808 10848
rect 30866 10248 31826 10848
rect 31884 10248 32844 10848
rect 32902 10248 33862 10848
rect 33920 10248 34880 10848
rect 34938 10248 35898 10848
rect 35956 10248 36916 10848
rect 36974 10248 37934 10848
rect 37992 10248 38952 10848
rect 39010 10248 39970 10848
rect 19668 9016 20628 9616
rect 20686 9016 21646 9616
rect 21704 9016 22664 9616
rect 22722 9016 23682 9616
rect 23740 9016 24700 9616
rect 24758 9016 25718 9616
rect 25776 9016 26736 9616
rect 26794 9016 27754 9616
rect 27812 9016 28772 9616
rect 28830 9016 29790 9616
rect 29848 9016 30808 9616
rect 30866 9016 31826 9616
rect 31884 9016 32844 9616
rect 32902 9016 33862 9616
rect 33920 9016 34880 9616
rect 34938 9016 35898 9616
rect 35956 9016 36916 9616
rect 36974 9016 37934 9616
rect 37992 9016 38952 9616
rect 39010 9016 39970 9616
rect 19666 7782 20626 8382
rect 20684 7782 21644 8382
rect 21702 7782 22662 8382
rect 22720 7782 23680 8382
rect 23738 7782 24698 8382
rect 24756 7782 25716 8382
rect 25774 7782 26734 8382
rect 26792 7782 27752 8382
rect 27810 7782 28770 8382
rect 28828 7782 29788 8382
rect 29846 7782 30806 8382
rect 30864 7782 31824 8382
rect 31882 7782 32842 8382
rect 32900 7782 33860 8382
rect 33918 7782 34878 8382
rect 34936 7782 35896 8382
rect 35954 7782 36914 8382
rect 36972 7782 37932 8382
rect 37990 7782 38950 8382
rect 39008 7782 39968 8382
rect 19666 6548 20626 7148
rect 20684 6548 21644 7148
rect 21702 6548 22662 7148
rect 22720 6548 23680 7148
rect 23738 6548 24698 7148
rect 24756 6548 25716 7148
rect 25774 6548 26734 7148
rect 26792 6548 27752 7148
rect 27810 6548 28770 7148
rect 28828 6548 29788 7148
rect 29846 6548 30806 7148
rect 30864 6548 31824 7148
rect 31882 6548 32842 7148
rect 32900 6548 33860 7148
rect 33918 6548 34878 7148
rect 34936 6548 35896 7148
rect 35954 6548 36914 7148
rect 36972 6548 37932 7148
rect 37990 6548 38950 7148
rect 39008 6548 39968 7148
rect 19666 5316 20626 5916
rect 20684 5316 21644 5916
rect 21702 5316 22662 5916
rect 22720 5316 23680 5916
rect 23738 5316 24698 5916
rect 24756 5316 25716 5916
rect 25774 5316 26734 5916
rect 26792 5316 27752 5916
rect 27810 5316 28770 5916
rect 28828 5316 29788 5916
rect 29846 5316 30806 5916
rect 30864 5316 31824 5916
rect 31882 5316 32842 5916
rect 32900 5316 33860 5916
rect 33918 5316 34878 5916
rect 34936 5316 35896 5916
rect 35954 5316 36914 5916
rect 36972 5316 37932 5916
rect 37990 5316 38950 5916
rect 39008 5316 39968 5916
rect 19666 4082 20626 4682
rect 20684 4082 21644 4682
rect 21702 4082 22662 4682
rect 22720 4082 23680 4682
rect 23738 4082 24698 4682
rect 24756 4082 25716 4682
rect 25774 4082 26734 4682
rect 26792 4082 27752 4682
rect 27810 4082 28770 4682
rect 28828 4082 29788 4682
rect 29846 4082 30806 4682
rect 30864 4082 31824 4682
rect 31882 4082 32842 4682
rect 32900 4082 33860 4682
rect 33918 4082 34878 4682
rect 34936 4082 35896 4682
rect 35954 4082 36914 4682
rect 36972 4082 37932 4682
rect 37990 4082 38950 4682
rect 39008 4082 39968 4682
rect 19666 2848 20626 3448
rect 20684 2848 21644 3448
rect 21702 2848 22662 3448
rect 22720 2848 23680 3448
rect 23738 2848 24698 3448
rect 24756 2848 25716 3448
rect 25774 2848 26734 3448
rect 26792 2848 27752 3448
rect 27810 2848 28770 3448
rect 28828 2848 29788 3448
rect 29846 2848 30806 3448
rect 30864 2848 31824 3448
rect 31882 2848 32842 3448
rect 32900 2848 33860 3448
rect 33918 2848 34878 3448
rect 34936 2848 35896 3448
rect 35954 2848 36914 3448
rect 36972 2848 37932 3448
rect 37990 2848 38950 3448
rect 39008 2848 39968 3448
rect 19666 1616 20626 2216
rect 20684 1616 21644 2216
rect 21702 1616 22662 2216
rect 22720 1616 23680 2216
rect 23738 1616 24698 2216
rect 24756 1616 25716 2216
rect 25774 1616 26734 2216
rect 26792 1616 27752 2216
rect 27810 1616 28770 2216
rect 28828 1616 29788 2216
rect 29846 1616 30806 2216
rect 30864 1616 31824 2216
rect 31882 1616 32842 2216
rect 32900 1616 33860 2216
rect 33918 1616 34878 2216
rect 34936 1616 35896 2216
rect 35954 1616 36914 2216
rect 36972 1616 37932 2216
rect 37990 1616 38950 2216
rect 39008 1616 39968 2216
rect 19666 382 20626 982
rect 20684 382 21644 982
rect 21702 382 22662 982
rect 22720 382 23680 982
rect 23738 382 24698 982
rect 24756 382 25716 982
rect 25774 382 26734 982
rect 26792 382 27752 982
rect 27810 382 28770 982
rect 28828 382 29788 982
rect 29846 382 30806 982
rect 30864 382 31824 982
rect 31882 382 32842 982
rect 32900 382 33860 982
rect 33918 382 34878 982
rect 34936 382 35896 982
rect 35954 382 36914 982
rect 36972 382 37932 982
rect 37990 382 38950 982
rect 39008 382 39968 982
rect 7036 -660 7996 -60
rect 8054 -660 9014 -60
rect 9072 -660 10032 -60
rect 10090 -660 11050 -60
rect 11108 -660 12068 -60
rect 12126 -660 13086 -60
rect 13144 -660 14104 -60
rect 14162 -660 15122 -60
rect 15180 -660 16140 -60
rect 16198 -660 17158 -60
rect 19666 -850 20626 -250
rect 20684 -850 21644 -250
rect 21702 -850 22662 -250
rect 22720 -850 23680 -250
rect 23738 -850 24698 -250
rect 24756 -850 25716 -250
rect 25774 -850 26734 -250
rect 26792 -850 27752 -250
rect 27810 -850 28770 -250
rect 28828 -850 29788 -250
rect 29846 -850 30806 -250
rect 30864 -850 31824 -250
rect 31882 -850 32842 -250
rect 32900 -850 33860 -250
rect 33918 -850 34878 -250
rect 34936 -850 35896 -250
rect 35954 -850 36914 -250
rect 36972 -850 37932 -250
rect 37990 -850 38950 -250
rect 39008 -850 39968 -250
<< pmos >>
rect 24560 19408 25520 20008
rect 25578 19408 26538 20008
rect 26596 19408 27556 20008
rect 27614 19408 28574 20008
rect 28632 19408 29592 20008
rect 29650 19408 30610 20008
rect 30668 19408 31628 20008
rect 31686 19408 32646 20008
rect 32704 19408 33664 20008
rect 33722 19408 34682 20008
rect 34740 19408 35700 20008
rect 35758 19408 36718 20008
rect 36776 19408 37736 20008
rect 37794 19408 38754 20008
rect 38812 19408 39772 20008
rect 24560 18152 25520 18752
rect 25578 18152 26538 18752
rect 26596 18152 27556 18752
rect 27614 18152 28574 18752
rect 28632 18152 29592 18752
rect 29650 18152 30610 18752
rect 30668 18152 31628 18752
rect 31686 18152 32646 18752
rect 32704 18152 33664 18752
rect 33722 18152 34682 18752
rect 34740 18152 35700 18752
rect 35758 18152 36718 18752
rect 36776 18152 37736 18752
rect 37794 18152 38754 18752
rect 38812 18152 39772 18752
rect 24560 16896 25520 17496
rect 25578 16896 26538 17496
rect 26596 16896 27556 17496
rect 27614 16896 28574 17496
rect 28632 16896 29592 17496
rect 29650 16896 30610 17496
rect 30668 16896 31628 17496
rect 31686 16896 32646 17496
rect 32704 16896 33664 17496
rect 33722 16896 34682 17496
rect 34740 16896 35700 17496
rect 35758 16896 36718 17496
rect 36776 16896 37736 17496
rect 37794 16896 38754 17496
rect 38812 16896 39772 17496
rect 24560 15640 25520 16240
rect 25578 15640 26538 16240
rect 26596 15640 27556 16240
rect 27614 15640 28574 16240
rect 28632 15640 29592 16240
rect 29650 15640 30610 16240
rect 30668 15640 31628 16240
rect 31686 15640 32646 16240
rect 32704 15640 33664 16240
rect 33722 15640 34682 16240
rect 34740 15640 35700 16240
rect 35758 15640 36718 16240
rect 36776 15640 37736 16240
rect 37794 15640 38754 16240
rect 38812 15640 39772 16240
<< pmoslvt >>
rect 23574 25954 24534 26554
rect 24592 25954 25552 26554
rect 25610 25954 26570 26554
rect 26628 25954 27588 26554
rect 27646 25954 28606 26554
rect 28664 25954 29624 26554
rect 29682 25954 30642 26554
rect 30700 25954 31660 26554
rect 31718 25954 32678 26554
rect 32736 25954 33696 26554
rect 33754 25954 34714 26554
rect 34772 25954 35732 26554
rect 35790 25954 36750 26554
rect 36808 25954 37768 26554
rect 37826 25954 38786 26554
rect 38844 25954 39804 26554
rect 23574 24818 24534 25418
rect 24592 24818 25552 25418
rect 25610 24818 26570 25418
rect 26628 24818 27588 25418
rect 27646 24818 28606 25418
rect 28664 24818 29624 25418
rect 29682 24818 30642 25418
rect 30700 24818 31660 25418
rect 31718 24818 32678 25418
rect 32736 24818 33696 25418
rect 33754 24818 34714 25418
rect 34772 24818 35732 25418
rect 35790 24818 36750 25418
rect 36808 24818 37768 25418
rect 37826 24818 38786 25418
rect 38844 24818 39804 25418
rect 23574 23682 24534 24282
rect 24592 23682 25552 24282
rect 25610 23682 26570 24282
rect 26628 23682 27588 24282
rect 27646 23682 28606 24282
rect 28664 23682 29624 24282
rect 29682 23682 30642 24282
rect 30700 23682 31660 24282
rect 31718 23682 32678 24282
rect 32736 23682 33696 24282
rect 33754 23682 34714 24282
rect 34772 23682 35732 24282
rect 35790 23682 36750 24282
rect 36808 23682 37768 24282
rect 37826 23682 38786 24282
rect 38844 23682 39804 24282
rect 24768 22044 25728 22644
rect 25786 22044 26746 22644
rect 26804 22044 27764 22644
rect 27822 22044 28782 22644
rect 28840 22044 29800 22644
rect 29858 22044 30818 22644
rect 30876 22044 31836 22644
rect 31894 22044 32854 22644
rect 32912 22044 33872 22644
rect 33930 22044 34890 22644
rect 34948 22044 35908 22644
rect 35966 22044 36926 22644
rect 36984 22044 37944 22644
rect 38002 22044 38962 22644
rect 24768 21012 25728 21612
rect 25786 21012 26746 21612
rect 26804 21012 27764 21612
rect 27822 21012 28782 21612
rect 28840 21012 29800 21612
rect 29858 21012 30818 21612
rect 30876 21012 31836 21612
rect 31894 21012 32854 21612
rect 32912 21012 33872 21612
rect 33930 21012 34890 21612
rect 34948 21012 35908 21612
rect 35966 21012 36926 21612
rect 36984 21012 37944 21612
rect 38002 21012 38962 21612
rect 19256 19304 20216 19904
rect 20274 19304 21234 19904
rect 21292 19304 22252 19904
rect 22310 19304 23270 19904
rect 19256 18272 20216 18872
rect 20274 18272 21234 18872
rect 21292 18272 22252 18872
rect 22310 18272 23270 18872
rect 19256 17240 20216 17840
rect 20274 17240 21234 17840
rect 21292 17240 22252 17840
rect 22310 17240 23270 17840
rect 19256 16208 20216 16808
rect 20274 16208 21234 16808
rect 21292 16208 22252 16808
rect 22310 16208 23270 16808
<< nmoslvt >>
rect 7902 11968 8862 12568
rect 8920 11968 9880 12568
rect 9938 11968 10898 12568
rect 10956 11968 11916 12568
rect 11974 11968 12934 12568
rect 12992 11968 13952 12568
rect 14010 11968 14970 12568
rect 15028 11968 15988 12568
rect 16046 11968 17006 12568
rect 7902 11150 8862 11750
rect 8920 11150 9880 11750
rect 9938 11150 10898 11750
rect 10956 11150 11916 11750
rect 11974 11150 12934 11750
rect 12992 11150 13952 11750
rect 14010 11150 14970 11750
rect 15028 11150 15988 11750
rect 16046 11150 17006 11750
rect 7902 10332 8862 10932
rect 8920 10332 9880 10932
rect 9938 10332 10898 10932
rect 10956 10332 11916 10932
rect 11974 10332 12934 10932
rect 12992 10332 13952 10932
rect 14010 10332 14970 10932
rect 15028 10332 15988 10932
rect 16046 10332 17006 10932
rect 7902 9514 8862 10114
rect 8920 9514 9880 10114
rect 9938 9514 10898 10114
rect 10956 9514 11916 10114
rect 11974 9514 12934 10114
rect 12992 9514 13952 10114
rect 14010 9514 14970 10114
rect 15028 9514 15988 10114
rect 16046 9514 17006 10114
rect 7902 8696 8862 9296
rect 8920 8696 9880 9296
rect 9938 8696 10898 9296
rect 10956 8696 11916 9296
rect 11974 8696 12934 9296
rect 12992 8696 13952 9296
rect 14010 8696 14970 9296
rect 15028 8696 15988 9296
rect 16046 8696 17006 9296
rect 7902 7878 8862 8478
rect 8920 7878 9880 8478
rect 9938 7878 10898 8478
rect 10956 7878 11916 8478
rect 11974 7878 12934 8478
rect 12992 7878 13952 8478
rect 14010 7878 14970 8478
rect 15028 7878 15988 8478
rect 16046 7878 17006 8478
rect 7902 7060 8862 7660
rect 8920 7060 9880 7660
rect 9938 7060 10898 7660
rect 10956 7060 11916 7660
rect 11974 7060 12934 7660
rect 12992 7060 13952 7660
rect 14010 7060 14970 7660
rect 15028 7060 15988 7660
rect 16046 7060 17006 7660
rect 7902 6242 8862 6842
rect 8920 6242 9880 6842
rect 9938 6242 10898 6842
rect 10956 6242 11916 6842
rect 11974 6242 12934 6842
rect 12992 6242 13952 6842
rect 14010 6242 14970 6842
rect 15028 6242 15988 6842
rect 16046 6242 17006 6842
rect 6578 4218 7538 4818
rect 7596 4218 8556 4818
rect 8614 4218 9574 4818
rect 9632 4218 10592 4818
rect 10650 4218 11610 4818
rect 11668 4218 12628 4818
rect 12686 4218 13646 4818
rect 13704 4218 14664 4818
rect 14722 4218 15682 4818
rect 15740 4218 16700 4818
rect 16758 4218 17718 4818
rect 6578 3106 7538 3706
rect 7596 3106 8556 3706
rect 8614 3106 9574 3706
rect 9632 3106 10592 3706
rect 10650 3106 11610 3706
rect 11668 3106 12628 3706
rect 12686 3106 13646 3706
rect 13704 3106 14664 3706
rect 14722 3106 15682 3706
rect 15740 3106 16700 3706
rect 16758 3106 17718 3706
rect 6578 1994 7538 2594
rect 7596 1994 8556 2594
rect 8614 1994 9574 2594
rect 9632 1994 10592 2594
rect 10650 1994 11610 2594
rect 11668 1994 12628 2594
rect 12686 1994 13646 2594
rect 13704 1994 14664 2594
rect 14722 1994 15682 2594
rect 15740 1994 16700 2594
rect 16758 1994 17718 2594
rect 6578 882 7538 1482
rect 7596 882 8556 1482
rect 8614 882 9574 1482
rect 9632 882 10592 1482
rect 10650 882 11610 1482
rect 11668 882 12628 1482
rect 12686 882 13646 1482
rect 13704 882 14664 1482
rect 14722 882 15682 1482
rect 15740 882 16700 1482
rect 16758 882 17718 1482
<< ndiff >>
rect 274 430 332 442
rect 274 54 286 430
rect 320 54 332 430
rect 274 42 332 54
rect 532 430 590 442
rect 532 54 544 430
rect 578 54 590 430
rect 532 42 590 54
rect 790 430 848 442
rect 790 54 802 430
rect 836 54 848 430
rect 790 42 848 54
rect 1048 430 1106 442
rect 1048 54 1060 430
rect 1094 54 1106 430
rect 1048 42 1106 54
rect 1306 430 1364 442
rect 1306 54 1318 430
rect 1352 54 1364 430
rect 1306 42 1364 54
rect 1564 430 1622 442
rect 1564 54 1576 430
rect 1610 54 1622 430
rect 1564 42 1622 54
rect 1822 430 1880 442
rect 1822 54 1834 430
rect 1868 54 1880 430
rect 1822 42 1880 54
rect 2080 430 2138 442
rect 2080 54 2092 430
rect 2126 54 2138 430
rect 2080 42 2138 54
rect 2338 430 2396 442
rect 2338 54 2350 430
rect 2384 54 2396 430
rect 2338 42 2396 54
rect 2596 430 2654 442
rect 2596 54 2608 430
rect 2642 54 2654 430
rect 2596 42 2654 54
rect 2854 430 2912 442
rect 2854 54 2866 430
rect 2900 54 2912 430
rect 2854 42 2912 54
rect 3112 430 3170 442
rect 3112 54 3124 430
rect 3158 54 3170 430
rect 3112 42 3170 54
rect 3370 430 3428 442
rect 3370 54 3382 430
rect 3416 54 3428 430
rect 3370 42 3428 54
rect 3628 430 3686 442
rect 3628 54 3640 430
rect 3674 54 3686 430
rect 3628 42 3686 54
rect 3886 430 3944 442
rect 3886 54 3898 430
rect 3932 54 3944 430
rect 3886 42 3944 54
rect 274 -570 332 -558
rect 274 -946 286 -570
rect 320 -946 332 -570
rect 274 -958 332 -946
rect 532 -570 590 -558
rect 532 -946 544 -570
rect 578 -946 590 -570
rect 532 -958 590 -946
rect 790 -570 848 -558
rect 790 -946 802 -570
rect 836 -946 848 -570
rect 790 -958 848 -946
rect 1048 -570 1106 -558
rect 1048 -946 1060 -570
rect 1094 -946 1106 -570
rect 1048 -958 1106 -946
rect 1306 -570 1364 -558
rect 1306 -946 1318 -570
rect 1352 -946 1364 -570
rect 1306 -958 1364 -946
rect 1564 -570 1622 -558
rect 1564 -946 1576 -570
rect 1610 -946 1622 -570
rect 1564 -958 1622 -946
rect 1822 -570 1880 -558
rect 1822 -946 1834 -570
rect 1868 -946 1880 -570
rect 1822 -958 1880 -946
rect 2080 -570 2138 -558
rect 2080 -946 2092 -570
rect 2126 -946 2138 -570
rect 2080 -958 2138 -946
rect 2338 -570 2396 -558
rect 2338 -946 2350 -570
rect 2384 -946 2396 -570
rect 2338 -958 2396 -946
rect 2596 -570 2654 -558
rect 2596 -946 2608 -570
rect 2642 -946 2654 -570
rect 2596 -958 2654 -946
rect 2854 -570 2912 -558
rect 2854 -946 2866 -570
rect 2900 -946 2912 -570
rect 2854 -958 2912 -946
rect 3112 -570 3170 -558
rect 3112 -946 3124 -570
rect 3158 -946 3170 -570
rect 3112 -958 3170 -946
rect 3370 -570 3428 -558
rect 3370 -946 3382 -570
rect 3416 -946 3428 -570
rect 3370 -958 3428 -946
rect 3628 -570 3686 -558
rect 3628 -946 3640 -570
rect 3674 -946 3686 -570
rect 3628 -958 3686 -946
rect 3886 -570 3944 -558
rect 3886 -946 3898 -570
rect 3932 -946 3944 -570
rect 3886 -958 3944 -946
rect 19610 13032 19668 13044
rect 7844 12556 7902 12568
rect 7844 11980 7856 12556
rect 7890 11980 7902 12556
rect 7844 11968 7902 11980
rect 8862 12556 8920 12568
rect 8862 11980 8874 12556
rect 8908 11980 8920 12556
rect 8862 11968 8920 11980
rect 9880 12556 9938 12568
rect 9880 11980 9892 12556
rect 9926 11980 9938 12556
rect 9880 11968 9938 11980
rect 10898 12556 10956 12568
rect 10898 11980 10910 12556
rect 10944 11980 10956 12556
rect 10898 11968 10956 11980
rect 11916 12556 11974 12568
rect 11916 11980 11928 12556
rect 11962 11980 11974 12556
rect 11916 11968 11974 11980
rect 12934 12556 12992 12568
rect 12934 11980 12946 12556
rect 12980 11980 12992 12556
rect 12934 11968 12992 11980
rect 13952 12556 14010 12568
rect 13952 11980 13964 12556
rect 13998 11980 14010 12556
rect 13952 11968 14010 11980
rect 14970 12556 15028 12568
rect 14970 11980 14982 12556
rect 15016 11980 15028 12556
rect 14970 11968 15028 11980
rect 15988 12556 16046 12568
rect 15988 11980 16000 12556
rect 16034 11980 16046 12556
rect 15988 11968 16046 11980
rect 17006 12556 17064 12568
rect 17006 11980 17018 12556
rect 17052 11980 17064 12556
rect 19610 12456 19622 13032
rect 19656 12456 19668 13032
rect 19610 12444 19668 12456
rect 20628 13032 20686 13044
rect 20628 12456 20640 13032
rect 20674 12456 20686 13032
rect 20628 12444 20686 12456
rect 21646 13032 21704 13044
rect 21646 12456 21658 13032
rect 21692 12456 21704 13032
rect 21646 12444 21704 12456
rect 22664 13032 22722 13044
rect 22664 12456 22676 13032
rect 22710 12456 22722 13032
rect 22664 12444 22722 12456
rect 23682 13032 23740 13044
rect 23682 12456 23694 13032
rect 23728 12456 23740 13032
rect 23682 12444 23740 12456
rect 24700 13032 24758 13044
rect 24700 12456 24712 13032
rect 24746 12456 24758 13032
rect 24700 12444 24758 12456
rect 25718 13032 25776 13044
rect 25718 12456 25730 13032
rect 25764 12456 25776 13032
rect 25718 12444 25776 12456
rect 26736 13032 26794 13044
rect 26736 12456 26748 13032
rect 26782 12456 26794 13032
rect 26736 12444 26794 12456
rect 27754 13032 27812 13044
rect 27754 12456 27766 13032
rect 27800 12456 27812 13032
rect 27754 12444 27812 12456
rect 28772 13032 28830 13044
rect 28772 12456 28784 13032
rect 28818 12456 28830 13032
rect 28772 12444 28830 12456
rect 29790 13032 29848 13044
rect 29790 12456 29802 13032
rect 29836 12456 29848 13032
rect 29790 12444 29848 12456
rect 30808 13032 30866 13044
rect 30808 12456 30820 13032
rect 30854 12456 30866 13032
rect 30808 12444 30866 12456
rect 31826 13032 31884 13044
rect 31826 12456 31838 13032
rect 31872 12456 31884 13032
rect 31826 12444 31884 12456
rect 32844 13032 32902 13044
rect 32844 12456 32856 13032
rect 32890 12456 32902 13032
rect 32844 12444 32902 12456
rect 33862 13032 33920 13044
rect 33862 12456 33874 13032
rect 33908 12456 33920 13032
rect 33862 12444 33920 12456
rect 34880 13032 34938 13044
rect 34880 12456 34892 13032
rect 34926 12456 34938 13032
rect 34880 12444 34938 12456
rect 35898 13032 35956 13044
rect 35898 12456 35910 13032
rect 35944 12456 35956 13032
rect 35898 12444 35956 12456
rect 36916 13032 36974 13044
rect 36916 12456 36928 13032
rect 36962 12456 36974 13032
rect 36916 12444 36974 12456
rect 37934 13032 37992 13044
rect 37934 12456 37946 13032
rect 37980 12456 37992 13032
rect 37934 12444 37992 12456
rect 38952 13032 39010 13044
rect 38952 12456 38964 13032
rect 38998 12456 39010 13032
rect 38952 12444 39010 12456
rect 39970 13032 40028 13044
rect 39970 12456 39982 13032
rect 40016 12456 40028 13032
rect 39970 12444 40028 12456
rect 17006 11968 17064 11980
rect 19610 12214 19668 12226
rect 7844 11738 7902 11750
rect 7844 11162 7856 11738
rect 7890 11162 7902 11738
rect 7844 11150 7902 11162
rect 8862 11738 8920 11750
rect 8862 11162 8874 11738
rect 8908 11162 8920 11738
rect 8862 11150 8920 11162
rect 9880 11738 9938 11750
rect 9880 11162 9892 11738
rect 9926 11162 9938 11738
rect 9880 11150 9938 11162
rect 10898 11738 10956 11750
rect 10898 11162 10910 11738
rect 10944 11162 10956 11738
rect 10898 11150 10956 11162
rect 11916 11738 11974 11750
rect 11916 11162 11928 11738
rect 11962 11162 11974 11738
rect 11916 11150 11974 11162
rect 12934 11738 12992 11750
rect 12934 11162 12946 11738
rect 12980 11162 12992 11738
rect 12934 11150 12992 11162
rect 13952 11738 14010 11750
rect 13952 11162 13964 11738
rect 13998 11162 14010 11738
rect 13952 11150 14010 11162
rect 14970 11738 15028 11750
rect 14970 11162 14982 11738
rect 15016 11162 15028 11738
rect 14970 11150 15028 11162
rect 15988 11738 16046 11750
rect 15988 11162 16000 11738
rect 16034 11162 16046 11738
rect 15988 11150 16046 11162
rect 17006 11738 17064 11750
rect 17006 11162 17018 11738
rect 17052 11162 17064 11738
rect 19610 11638 19622 12214
rect 19656 11638 19668 12214
rect 19610 11626 19668 11638
rect 20628 12214 20686 12226
rect 20628 11638 20640 12214
rect 20674 11638 20686 12214
rect 20628 11626 20686 11638
rect 21646 12214 21704 12226
rect 21646 11638 21658 12214
rect 21692 11638 21704 12214
rect 21646 11626 21704 11638
rect 22664 12214 22722 12226
rect 22664 11638 22676 12214
rect 22710 11638 22722 12214
rect 22664 11626 22722 11638
rect 23682 12214 23740 12226
rect 23682 11638 23694 12214
rect 23728 11638 23740 12214
rect 23682 11626 23740 11638
rect 24700 12214 24758 12226
rect 24700 11638 24712 12214
rect 24746 11638 24758 12214
rect 24700 11626 24758 11638
rect 25718 12214 25776 12226
rect 25718 11638 25730 12214
rect 25764 11638 25776 12214
rect 25718 11626 25776 11638
rect 26736 12214 26794 12226
rect 26736 11638 26748 12214
rect 26782 11638 26794 12214
rect 26736 11626 26794 11638
rect 27754 12214 27812 12226
rect 27754 11638 27766 12214
rect 27800 11638 27812 12214
rect 27754 11626 27812 11638
rect 28772 12214 28830 12226
rect 28772 11638 28784 12214
rect 28818 11638 28830 12214
rect 28772 11626 28830 11638
rect 29790 12214 29848 12226
rect 29790 11638 29802 12214
rect 29836 11638 29848 12214
rect 29790 11626 29848 11638
rect 30808 12214 30866 12226
rect 30808 11638 30820 12214
rect 30854 11638 30866 12214
rect 30808 11626 30866 11638
rect 31826 12214 31884 12226
rect 31826 11638 31838 12214
rect 31872 11638 31884 12214
rect 31826 11626 31884 11638
rect 32844 12214 32902 12226
rect 32844 11638 32856 12214
rect 32890 11638 32902 12214
rect 32844 11626 32902 11638
rect 33862 12214 33920 12226
rect 33862 11638 33874 12214
rect 33908 11638 33920 12214
rect 33862 11626 33920 11638
rect 34880 12214 34938 12226
rect 34880 11638 34892 12214
rect 34926 11638 34938 12214
rect 34880 11626 34938 11638
rect 35898 12214 35956 12226
rect 35898 11638 35910 12214
rect 35944 11638 35956 12214
rect 35898 11626 35956 11638
rect 36916 12214 36974 12226
rect 36916 11638 36928 12214
rect 36962 11638 36974 12214
rect 36916 11626 36974 11638
rect 37934 12214 37992 12226
rect 37934 11638 37946 12214
rect 37980 11638 37992 12214
rect 37934 11626 37992 11638
rect 38952 12214 39010 12226
rect 38952 11638 38964 12214
rect 38998 11638 39010 12214
rect 38952 11626 39010 11638
rect 39970 12214 40028 12226
rect 39970 11638 39982 12214
rect 40016 11638 40028 12214
rect 39970 11626 40028 11638
rect 17006 11150 17064 11162
rect 7844 10920 7902 10932
rect 7844 10344 7856 10920
rect 7890 10344 7902 10920
rect 7844 10332 7902 10344
rect 8862 10920 8920 10932
rect 8862 10344 8874 10920
rect 8908 10344 8920 10920
rect 8862 10332 8920 10344
rect 9880 10920 9938 10932
rect 9880 10344 9892 10920
rect 9926 10344 9938 10920
rect 9880 10332 9938 10344
rect 10898 10920 10956 10932
rect 10898 10344 10910 10920
rect 10944 10344 10956 10920
rect 10898 10332 10956 10344
rect 11916 10920 11974 10932
rect 11916 10344 11928 10920
rect 11962 10344 11974 10920
rect 11916 10332 11974 10344
rect 12934 10920 12992 10932
rect 12934 10344 12946 10920
rect 12980 10344 12992 10920
rect 12934 10332 12992 10344
rect 13952 10920 14010 10932
rect 13952 10344 13964 10920
rect 13998 10344 14010 10920
rect 13952 10332 14010 10344
rect 14970 10920 15028 10932
rect 14970 10344 14982 10920
rect 15016 10344 15028 10920
rect 14970 10332 15028 10344
rect 15988 10920 16046 10932
rect 15988 10344 16000 10920
rect 16034 10344 16046 10920
rect 15988 10332 16046 10344
rect 17006 10920 17064 10932
rect 17006 10344 17018 10920
rect 17052 10344 17064 10920
rect 17006 10332 17064 10344
rect 19610 10836 19668 10848
rect 19610 10260 19622 10836
rect 19656 10260 19668 10836
rect 19610 10248 19668 10260
rect 20628 10836 20686 10848
rect 20628 10260 20640 10836
rect 20674 10260 20686 10836
rect 20628 10248 20686 10260
rect 21646 10836 21704 10848
rect 21646 10260 21658 10836
rect 21692 10260 21704 10836
rect 21646 10248 21704 10260
rect 22664 10836 22722 10848
rect 22664 10260 22676 10836
rect 22710 10260 22722 10836
rect 22664 10248 22722 10260
rect 23682 10836 23740 10848
rect 23682 10260 23694 10836
rect 23728 10260 23740 10836
rect 23682 10248 23740 10260
rect 24700 10836 24758 10848
rect 24700 10260 24712 10836
rect 24746 10260 24758 10836
rect 24700 10248 24758 10260
rect 25718 10836 25776 10848
rect 25718 10260 25730 10836
rect 25764 10260 25776 10836
rect 25718 10248 25776 10260
rect 26736 10836 26794 10848
rect 26736 10260 26748 10836
rect 26782 10260 26794 10836
rect 26736 10248 26794 10260
rect 27754 10836 27812 10848
rect 27754 10260 27766 10836
rect 27800 10260 27812 10836
rect 27754 10248 27812 10260
rect 28772 10836 28830 10848
rect 28772 10260 28784 10836
rect 28818 10260 28830 10836
rect 28772 10248 28830 10260
rect 29790 10836 29848 10848
rect 29790 10260 29802 10836
rect 29836 10260 29848 10836
rect 29790 10248 29848 10260
rect 30808 10836 30866 10848
rect 30808 10260 30820 10836
rect 30854 10260 30866 10836
rect 30808 10248 30866 10260
rect 31826 10836 31884 10848
rect 31826 10260 31838 10836
rect 31872 10260 31884 10836
rect 31826 10248 31884 10260
rect 32844 10836 32902 10848
rect 32844 10260 32856 10836
rect 32890 10260 32902 10836
rect 32844 10248 32902 10260
rect 33862 10836 33920 10848
rect 33862 10260 33874 10836
rect 33908 10260 33920 10836
rect 33862 10248 33920 10260
rect 34880 10836 34938 10848
rect 34880 10260 34892 10836
rect 34926 10260 34938 10836
rect 34880 10248 34938 10260
rect 35898 10836 35956 10848
rect 35898 10260 35910 10836
rect 35944 10260 35956 10836
rect 35898 10248 35956 10260
rect 36916 10836 36974 10848
rect 36916 10260 36928 10836
rect 36962 10260 36974 10836
rect 36916 10248 36974 10260
rect 37934 10836 37992 10848
rect 37934 10260 37946 10836
rect 37980 10260 37992 10836
rect 37934 10248 37992 10260
rect 38952 10836 39010 10848
rect 38952 10260 38964 10836
rect 38998 10260 39010 10836
rect 38952 10248 39010 10260
rect 39970 10836 40028 10848
rect 39970 10260 39982 10836
rect 40016 10260 40028 10836
rect 39970 10248 40028 10260
rect 7844 10102 7902 10114
rect 7844 9526 7856 10102
rect 7890 9526 7902 10102
rect 7844 9514 7902 9526
rect 8862 10102 8920 10114
rect 8862 9526 8874 10102
rect 8908 9526 8920 10102
rect 8862 9514 8920 9526
rect 9880 10102 9938 10114
rect 9880 9526 9892 10102
rect 9926 9526 9938 10102
rect 9880 9514 9938 9526
rect 10898 10102 10956 10114
rect 10898 9526 10910 10102
rect 10944 9526 10956 10102
rect 10898 9514 10956 9526
rect 11916 10102 11974 10114
rect 11916 9526 11928 10102
rect 11962 9526 11974 10102
rect 11916 9514 11974 9526
rect 12934 10102 12992 10114
rect 12934 9526 12946 10102
rect 12980 9526 12992 10102
rect 12934 9514 12992 9526
rect 13952 10102 14010 10114
rect 13952 9526 13964 10102
rect 13998 9526 14010 10102
rect 13952 9514 14010 9526
rect 14970 10102 15028 10114
rect 14970 9526 14982 10102
rect 15016 9526 15028 10102
rect 14970 9514 15028 9526
rect 15988 10102 16046 10114
rect 15988 9526 16000 10102
rect 16034 9526 16046 10102
rect 15988 9514 16046 9526
rect 17006 10102 17064 10114
rect 17006 9526 17018 10102
rect 17052 9526 17064 10102
rect 17006 9514 17064 9526
rect 19610 9604 19668 9616
rect 7844 9284 7902 9296
rect 7844 8708 7856 9284
rect 7890 8708 7902 9284
rect 7844 8696 7902 8708
rect 8862 9284 8920 9296
rect 8862 8708 8874 9284
rect 8908 8708 8920 9284
rect 8862 8696 8920 8708
rect 9880 9284 9938 9296
rect 9880 8708 9892 9284
rect 9926 8708 9938 9284
rect 9880 8696 9938 8708
rect 10898 9284 10956 9296
rect 10898 8708 10910 9284
rect 10944 8708 10956 9284
rect 10898 8696 10956 8708
rect 11916 9284 11974 9296
rect 11916 8708 11928 9284
rect 11962 8708 11974 9284
rect 11916 8696 11974 8708
rect 12934 9284 12992 9296
rect 12934 8708 12946 9284
rect 12980 8708 12992 9284
rect 12934 8696 12992 8708
rect 13952 9284 14010 9296
rect 13952 8708 13964 9284
rect 13998 8708 14010 9284
rect 13952 8696 14010 8708
rect 14970 9284 15028 9296
rect 14970 8708 14982 9284
rect 15016 8708 15028 9284
rect 14970 8696 15028 8708
rect 15988 9284 16046 9296
rect 15988 8708 16000 9284
rect 16034 8708 16046 9284
rect 15988 8696 16046 8708
rect 17006 9284 17064 9296
rect 17006 8708 17018 9284
rect 17052 8708 17064 9284
rect 19610 9028 19622 9604
rect 19656 9028 19668 9604
rect 19610 9016 19668 9028
rect 20628 9604 20686 9616
rect 20628 9028 20640 9604
rect 20674 9028 20686 9604
rect 20628 9016 20686 9028
rect 21646 9604 21704 9616
rect 21646 9028 21658 9604
rect 21692 9028 21704 9604
rect 21646 9016 21704 9028
rect 22664 9604 22722 9616
rect 22664 9028 22676 9604
rect 22710 9028 22722 9604
rect 22664 9016 22722 9028
rect 23682 9604 23740 9616
rect 23682 9028 23694 9604
rect 23728 9028 23740 9604
rect 23682 9016 23740 9028
rect 24700 9604 24758 9616
rect 24700 9028 24712 9604
rect 24746 9028 24758 9604
rect 24700 9016 24758 9028
rect 25718 9604 25776 9616
rect 25718 9028 25730 9604
rect 25764 9028 25776 9604
rect 25718 9016 25776 9028
rect 26736 9604 26794 9616
rect 26736 9028 26748 9604
rect 26782 9028 26794 9604
rect 26736 9016 26794 9028
rect 27754 9604 27812 9616
rect 27754 9028 27766 9604
rect 27800 9028 27812 9604
rect 27754 9016 27812 9028
rect 28772 9604 28830 9616
rect 28772 9028 28784 9604
rect 28818 9028 28830 9604
rect 28772 9016 28830 9028
rect 29790 9604 29848 9616
rect 29790 9028 29802 9604
rect 29836 9028 29848 9604
rect 29790 9016 29848 9028
rect 30808 9604 30866 9616
rect 30808 9028 30820 9604
rect 30854 9028 30866 9604
rect 30808 9016 30866 9028
rect 31826 9604 31884 9616
rect 31826 9028 31838 9604
rect 31872 9028 31884 9604
rect 31826 9016 31884 9028
rect 32844 9604 32902 9616
rect 32844 9028 32856 9604
rect 32890 9028 32902 9604
rect 32844 9016 32902 9028
rect 33862 9604 33920 9616
rect 33862 9028 33874 9604
rect 33908 9028 33920 9604
rect 33862 9016 33920 9028
rect 34880 9604 34938 9616
rect 34880 9028 34892 9604
rect 34926 9028 34938 9604
rect 34880 9016 34938 9028
rect 35898 9604 35956 9616
rect 35898 9028 35910 9604
rect 35944 9028 35956 9604
rect 35898 9016 35956 9028
rect 36916 9604 36974 9616
rect 36916 9028 36928 9604
rect 36962 9028 36974 9604
rect 36916 9016 36974 9028
rect 37934 9604 37992 9616
rect 37934 9028 37946 9604
rect 37980 9028 37992 9604
rect 37934 9016 37992 9028
rect 38952 9604 39010 9616
rect 38952 9028 38964 9604
rect 38998 9028 39010 9604
rect 38952 9016 39010 9028
rect 39970 9604 40028 9616
rect 39970 9028 39982 9604
rect 40016 9028 40028 9604
rect 39970 9016 40028 9028
rect 17006 8696 17064 8708
rect 7844 8466 7902 8478
rect 7844 7890 7856 8466
rect 7890 7890 7902 8466
rect 7844 7878 7902 7890
rect 8862 8466 8920 8478
rect 8862 7890 8874 8466
rect 8908 7890 8920 8466
rect 8862 7878 8920 7890
rect 9880 8466 9938 8478
rect 9880 7890 9892 8466
rect 9926 7890 9938 8466
rect 9880 7878 9938 7890
rect 10898 8466 10956 8478
rect 10898 7890 10910 8466
rect 10944 7890 10956 8466
rect 10898 7878 10956 7890
rect 11916 8466 11974 8478
rect 11916 7890 11928 8466
rect 11962 7890 11974 8466
rect 11916 7878 11974 7890
rect 12934 8466 12992 8478
rect 12934 7890 12946 8466
rect 12980 7890 12992 8466
rect 12934 7878 12992 7890
rect 13952 8466 14010 8478
rect 13952 7890 13964 8466
rect 13998 7890 14010 8466
rect 13952 7878 14010 7890
rect 14970 8466 15028 8478
rect 14970 7890 14982 8466
rect 15016 7890 15028 8466
rect 14970 7878 15028 7890
rect 15988 8466 16046 8478
rect 15988 7890 16000 8466
rect 16034 7890 16046 8466
rect 15988 7878 16046 7890
rect 17006 8466 17064 8478
rect 17006 7890 17018 8466
rect 17052 7890 17064 8466
rect 17006 7878 17064 7890
rect 19608 8370 19666 8382
rect 19608 7794 19620 8370
rect 19654 7794 19666 8370
rect 19608 7782 19666 7794
rect 20626 8370 20684 8382
rect 20626 7794 20638 8370
rect 20672 7794 20684 8370
rect 20626 7782 20684 7794
rect 21644 8370 21702 8382
rect 21644 7794 21656 8370
rect 21690 7794 21702 8370
rect 21644 7782 21702 7794
rect 22662 8370 22720 8382
rect 22662 7794 22674 8370
rect 22708 7794 22720 8370
rect 22662 7782 22720 7794
rect 23680 8370 23738 8382
rect 23680 7794 23692 8370
rect 23726 7794 23738 8370
rect 23680 7782 23738 7794
rect 24698 8370 24756 8382
rect 24698 7794 24710 8370
rect 24744 7794 24756 8370
rect 24698 7782 24756 7794
rect 25716 8370 25774 8382
rect 25716 7794 25728 8370
rect 25762 7794 25774 8370
rect 25716 7782 25774 7794
rect 26734 8370 26792 8382
rect 26734 7794 26746 8370
rect 26780 7794 26792 8370
rect 26734 7782 26792 7794
rect 27752 8370 27810 8382
rect 27752 7794 27764 8370
rect 27798 7794 27810 8370
rect 27752 7782 27810 7794
rect 28770 8370 28828 8382
rect 28770 7794 28782 8370
rect 28816 7794 28828 8370
rect 28770 7782 28828 7794
rect 29788 8370 29846 8382
rect 29788 7794 29800 8370
rect 29834 7794 29846 8370
rect 29788 7782 29846 7794
rect 30806 8370 30864 8382
rect 30806 7794 30818 8370
rect 30852 7794 30864 8370
rect 30806 7782 30864 7794
rect 31824 8370 31882 8382
rect 31824 7794 31836 8370
rect 31870 7794 31882 8370
rect 31824 7782 31882 7794
rect 32842 8370 32900 8382
rect 32842 7794 32854 8370
rect 32888 7794 32900 8370
rect 32842 7782 32900 7794
rect 33860 8370 33918 8382
rect 33860 7794 33872 8370
rect 33906 7794 33918 8370
rect 33860 7782 33918 7794
rect 34878 8370 34936 8382
rect 34878 7794 34890 8370
rect 34924 7794 34936 8370
rect 34878 7782 34936 7794
rect 35896 8370 35954 8382
rect 35896 7794 35908 8370
rect 35942 7794 35954 8370
rect 35896 7782 35954 7794
rect 36914 8370 36972 8382
rect 36914 7794 36926 8370
rect 36960 7794 36972 8370
rect 36914 7782 36972 7794
rect 37932 8370 37990 8382
rect 37932 7794 37944 8370
rect 37978 7794 37990 8370
rect 37932 7782 37990 7794
rect 38950 8370 39008 8382
rect 38950 7794 38962 8370
rect 38996 7794 39008 8370
rect 38950 7782 39008 7794
rect 39968 8370 40026 8382
rect 39968 7794 39980 8370
rect 40014 7794 40026 8370
rect 39968 7782 40026 7794
rect 7844 7648 7902 7660
rect 7844 7072 7856 7648
rect 7890 7072 7902 7648
rect 7844 7060 7902 7072
rect 8862 7648 8920 7660
rect 8862 7072 8874 7648
rect 8908 7072 8920 7648
rect 8862 7060 8920 7072
rect 9880 7648 9938 7660
rect 9880 7072 9892 7648
rect 9926 7072 9938 7648
rect 9880 7060 9938 7072
rect 10898 7648 10956 7660
rect 10898 7072 10910 7648
rect 10944 7072 10956 7648
rect 10898 7060 10956 7072
rect 11916 7648 11974 7660
rect 11916 7072 11928 7648
rect 11962 7072 11974 7648
rect 11916 7060 11974 7072
rect 12934 7648 12992 7660
rect 12934 7072 12946 7648
rect 12980 7072 12992 7648
rect 12934 7060 12992 7072
rect 13952 7648 14010 7660
rect 13952 7072 13964 7648
rect 13998 7072 14010 7648
rect 13952 7060 14010 7072
rect 14970 7648 15028 7660
rect 14970 7072 14982 7648
rect 15016 7072 15028 7648
rect 14970 7060 15028 7072
rect 15988 7648 16046 7660
rect 15988 7072 16000 7648
rect 16034 7072 16046 7648
rect 15988 7060 16046 7072
rect 17006 7648 17064 7660
rect 17006 7072 17018 7648
rect 17052 7072 17064 7648
rect 17006 7060 17064 7072
rect 19608 7136 19666 7148
rect 7844 6830 7902 6842
rect 7844 6254 7856 6830
rect 7890 6254 7902 6830
rect 7844 6242 7902 6254
rect 8862 6830 8920 6842
rect 8862 6254 8874 6830
rect 8908 6254 8920 6830
rect 8862 6242 8920 6254
rect 9880 6830 9938 6842
rect 9880 6254 9892 6830
rect 9926 6254 9938 6830
rect 9880 6242 9938 6254
rect 10898 6830 10956 6842
rect 10898 6254 10910 6830
rect 10944 6254 10956 6830
rect 10898 6242 10956 6254
rect 11916 6830 11974 6842
rect 11916 6254 11928 6830
rect 11962 6254 11974 6830
rect 11916 6242 11974 6254
rect 12934 6830 12992 6842
rect 12934 6254 12946 6830
rect 12980 6254 12992 6830
rect 12934 6242 12992 6254
rect 13952 6830 14010 6842
rect 13952 6254 13964 6830
rect 13998 6254 14010 6830
rect 13952 6242 14010 6254
rect 14970 6830 15028 6842
rect 14970 6254 14982 6830
rect 15016 6254 15028 6830
rect 14970 6242 15028 6254
rect 15988 6830 16046 6842
rect 15988 6254 16000 6830
rect 16034 6254 16046 6830
rect 15988 6242 16046 6254
rect 17006 6830 17064 6842
rect 17006 6254 17018 6830
rect 17052 6254 17064 6830
rect 19608 6560 19620 7136
rect 19654 6560 19666 7136
rect 19608 6548 19666 6560
rect 20626 7136 20684 7148
rect 20626 6560 20638 7136
rect 20672 6560 20684 7136
rect 20626 6548 20684 6560
rect 21644 7136 21702 7148
rect 21644 6560 21656 7136
rect 21690 6560 21702 7136
rect 21644 6548 21702 6560
rect 22662 7136 22720 7148
rect 22662 6560 22674 7136
rect 22708 6560 22720 7136
rect 22662 6548 22720 6560
rect 23680 7136 23738 7148
rect 23680 6560 23692 7136
rect 23726 6560 23738 7136
rect 23680 6548 23738 6560
rect 24698 7136 24756 7148
rect 24698 6560 24710 7136
rect 24744 6560 24756 7136
rect 24698 6548 24756 6560
rect 25716 7136 25774 7148
rect 25716 6560 25728 7136
rect 25762 6560 25774 7136
rect 25716 6548 25774 6560
rect 26734 7136 26792 7148
rect 26734 6560 26746 7136
rect 26780 6560 26792 7136
rect 26734 6548 26792 6560
rect 27752 7136 27810 7148
rect 27752 6560 27764 7136
rect 27798 6560 27810 7136
rect 27752 6548 27810 6560
rect 28770 7136 28828 7148
rect 28770 6560 28782 7136
rect 28816 6560 28828 7136
rect 28770 6548 28828 6560
rect 29788 7136 29846 7148
rect 29788 6560 29800 7136
rect 29834 6560 29846 7136
rect 29788 6548 29846 6560
rect 30806 7136 30864 7148
rect 30806 6560 30818 7136
rect 30852 6560 30864 7136
rect 30806 6548 30864 6560
rect 31824 7136 31882 7148
rect 31824 6560 31836 7136
rect 31870 6560 31882 7136
rect 31824 6548 31882 6560
rect 32842 7136 32900 7148
rect 32842 6560 32854 7136
rect 32888 6560 32900 7136
rect 32842 6548 32900 6560
rect 33860 7136 33918 7148
rect 33860 6560 33872 7136
rect 33906 6560 33918 7136
rect 33860 6548 33918 6560
rect 34878 7136 34936 7148
rect 34878 6560 34890 7136
rect 34924 6560 34936 7136
rect 34878 6548 34936 6560
rect 35896 7136 35954 7148
rect 35896 6560 35908 7136
rect 35942 6560 35954 7136
rect 35896 6548 35954 6560
rect 36914 7136 36972 7148
rect 36914 6560 36926 7136
rect 36960 6560 36972 7136
rect 36914 6548 36972 6560
rect 37932 7136 37990 7148
rect 37932 6560 37944 7136
rect 37978 6560 37990 7136
rect 37932 6548 37990 6560
rect 38950 7136 39008 7148
rect 38950 6560 38962 7136
rect 38996 6560 39008 7136
rect 38950 6548 39008 6560
rect 39968 7136 40026 7148
rect 39968 6560 39980 7136
rect 40014 6560 40026 7136
rect 39968 6548 40026 6560
rect 17006 6242 17064 6254
rect 19608 5904 19666 5916
rect 19608 5328 19620 5904
rect 19654 5328 19666 5904
rect 19608 5316 19666 5328
rect 20626 5904 20684 5916
rect 20626 5328 20638 5904
rect 20672 5328 20684 5904
rect 20626 5316 20684 5328
rect 21644 5904 21702 5916
rect 21644 5328 21656 5904
rect 21690 5328 21702 5904
rect 21644 5316 21702 5328
rect 22662 5904 22720 5916
rect 22662 5328 22674 5904
rect 22708 5328 22720 5904
rect 22662 5316 22720 5328
rect 23680 5904 23738 5916
rect 23680 5328 23692 5904
rect 23726 5328 23738 5904
rect 23680 5316 23738 5328
rect 24698 5904 24756 5916
rect 24698 5328 24710 5904
rect 24744 5328 24756 5904
rect 24698 5316 24756 5328
rect 25716 5904 25774 5916
rect 25716 5328 25728 5904
rect 25762 5328 25774 5904
rect 25716 5316 25774 5328
rect 26734 5904 26792 5916
rect 26734 5328 26746 5904
rect 26780 5328 26792 5904
rect 26734 5316 26792 5328
rect 27752 5904 27810 5916
rect 27752 5328 27764 5904
rect 27798 5328 27810 5904
rect 27752 5316 27810 5328
rect 28770 5904 28828 5916
rect 28770 5328 28782 5904
rect 28816 5328 28828 5904
rect 28770 5316 28828 5328
rect 29788 5904 29846 5916
rect 29788 5328 29800 5904
rect 29834 5328 29846 5904
rect 29788 5316 29846 5328
rect 30806 5904 30864 5916
rect 30806 5328 30818 5904
rect 30852 5328 30864 5904
rect 30806 5316 30864 5328
rect 31824 5904 31882 5916
rect 31824 5328 31836 5904
rect 31870 5328 31882 5904
rect 31824 5316 31882 5328
rect 32842 5904 32900 5916
rect 32842 5328 32854 5904
rect 32888 5328 32900 5904
rect 32842 5316 32900 5328
rect 33860 5904 33918 5916
rect 33860 5328 33872 5904
rect 33906 5328 33918 5904
rect 33860 5316 33918 5328
rect 34878 5904 34936 5916
rect 34878 5328 34890 5904
rect 34924 5328 34936 5904
rect 34878 5316 34936 5328
rect 35896 5904 35954 5916
rect 35896 5328 35908 5904
rect 35942 5328 35954 5904
rect 35896 5316 35954 5328
rect 36914 5904 36972 5916
rect 36914 5328 36926 5904
rect 36960 5328 36972 5904
rect 36914 5316 36972 5328
rect 37932 5904 37990 5916
rect 37932 5328 37944 5904
rect 37978 5328 37990 5904
rect 37932 5316 37990 5328
rect 38950 5904 39008 5916
rect 38950 5328 38962 5904
rect 38996 5328 39008 5904
rect 38950 5316 39008 5328
rect 39968 5904 40026 5916
rect 39968 5328 39980 5904
rect 40014 5328 40026 5904
rect 39968 5316 40026 5328
rect 6520 4806 6578 4818
rect 6520 4230 6532 4806
rect 6566 4230 6578 4806
rect 6520 4218 6578 4230
rect 7538 4806 7596 4818
rect 7538 4230 7550 4806
rect 7584 4230 7596 4806
rect 7538 4218 7596 4230
rect 8556 4806 8614 4818
rect 8556 4230 8568 4806
rect 8602 4230 8614 4806
rect 8556 4218 8614 4230
rect 9574 4806 9632 4818
rect 9574 4230 9586 4806
rect 9620 4230 9632 4806
rect 9574 4218 9632 4230
rect 10592 4806 10650 4818
rect 10592 4230 10604 4806
rect 10638 4230 10650 4806
rect 10592 4218 10650 4230
rect 11610 4806 11668 4818
rect 11610 4230 11622 4806
rect 11656 4230 11668 4806
rect 11610 4218 11668 4230
rect 12628 4806 12686 4818
rect 12628 4230 12640 4806
rect 12674 4230 12686 4806
rect 12628 4218 12686 4230
rect 13646 4806 13704 4818
rect 13646 4230 13658 4806
rect 13692 4230 13704 4806
rect 13646 4218 13704 4230
rect 14664 4806 14722 4818
rect 14664 4230 14676 4806
rect 14710 4230 14722 4806
rect 14664 4218 14722 4230
rect 15682 4806 15740 4818
rect 15682 4230 15694 4806
rect 15728 4230 15740 4806
rect 15682 4218 15740 4230
rect 16700 4806 16758 4818
rect 16700 4230 16712 4806
rect 16746 4230 16758 4806
rect 16700 4218 16758 4230
rect 17718 4806 17776 4818
rect 17718 4230 17730 4806
rect 17764 4230 17776 4806
rect 17718 4218 17776 4230
rect 19608 4670 19666 4682
rect 19608 4094 19620 4670
rect 19654 4094 19666 4670
rect 19608 4082 19666 4094
rect 20626 4670 20684 4682
rect 20626 4094 20638 4670
rect 20672 4094 20684 4670
rect 20626 4082 20684 4094
rect 21644 4670 21702 4682
rect 21644 4094 21656 4670
rect 21690 4094 21702 4670
rect 21644 4082 21702 4094
rect 22662 4670 22720 4682
rect 22662 4094 22674 4670
rect 22708 4094 22720 4670
rect 22662 4082 22720 4094
rect 23680 4670 23738 4682
rect 23680 4094 23692 4670
rect 23726 4094 23738 4670
rect 23680 4082 23738 4094
rect 24698 4670 24756 4682
rect 24698 4094 24710 4670
rect 24744 4094 24756 4670
rect 24698 4082 24756 4094
rect 25716 4670 25774 4682
rect 25716 4094 25728 4670
rect 25762 4094 25774 4670
rect 25716 4082 25774 4094
rect 26734 4670 26792 4682
rect 26734 4094 26746 4670
rect 26780 4094 26792 4670
rect 26734 4082 26792 4094
rect 27752 4670 27810 4682
rect 27752 4094 27764 4670
rect 27798 4094 27810 4670
rect 27752 4082 27810 4094
rect 28770 4670 28828 4682
rect 28770 4094 28782 4670
rect 28816 4094 28828 4670
rect 28770 4082 28828 4094
rect 29788 4670 29846 4682
rect 29788 4094 29800 4670
rect 29834 4094 29846 4670
rect 29788 4082 29846 4094
rect 30806 4670 30864 4682
rect 30806 4094 30818 4670
rect 30852 4094 30864 4670
rect 30806 4082 30864 4094
rect 31824 4670 31882 4682
rect 31824 4094 31836 4670
rect 31870 4094 31882 4670
rect 31824 4082 31882 4094
rect 32842 4670 32900 4682
rect 32842 4094 32854 4670
rect 32888 4094 32900 4670
rect 32842 4082 32900 4094
rect 33860 4670 33918 4682
rect 33860 4094 33872 4670
rect 33906 4094 33918 4670
rect 33860 4082 33918 4094
rect 34878 4670 34936 4682
rect 34878 4094 34890 4670
rect 34924 4094 34936 4670
rect 34878 4082 34936 4094
rect 35896 4670 35954 4682
rect 35896 4094 35908 4670
rect 35942 4094 35954 4670
rect 35896 4082 35954 4094
rect 36914 4670 36972 4682
rect 36914 4094 36926 4670
rect 36960 4094 36972 4670
rect 36914 4082 36972 4094
rect 37932 4670 37990 4682
rect 37932 4094 37944 4670
rect 37978 4094 37990 4670
rect 37932 4082 37990 4094
rect 38950 4670 39008 4682
rect 38950 4094 38962 4670
rect 38996 4094 39008 4670
rect 38950 4082 39008 4094
rect 39968 4670 40026 4682
rect 39968 4094 39980 4670
rect 40014 4094 40026 4670
rect 39968 4082 40026 4094
rect 6520 3694 6578 3706
rect 6520 3118 6532 3694
rect 6566 3118 6578 3694
rect 6520 3106 6578 3118
rect 7538 3694 7596 3706
rect 7538 3118 7550 3694
rect 7584 3118 7596 3694
rect 7538 3106 7596 3118
rect 8556 3694 8614 3706
rect 8556 3118 8568 3694
rect 8602 3118 8614 3694
rect 8556 3106 8614 3118
rect 9574 3694 9632 3706
rect 9574 3118 9586 3694
rect 9620 3118 9632 3694
rect 9574 3106 9632 3118
rect 10592 3694 10650 3706
rect 10592 3118 10604 3694
rect 10638 3118 10650 3694
rect 10592 3106 10650 3118
rect 11610 3694 11668 3706
rect 11610 3118 11622 3694
rect 11656 3118 11668 3694
rect 11610 3106 11668 3118
rect 12628 3694 12686 3706
rect 12628 3118 12640 3694
rect 12674 3118 12686 3694
rect 12628 3106 12686 3118
rect 13646 3694 13704 3706
rect 13646 3118 13658 3694
rect 13692 3118 13704 3694
rect 13646 3106 13704 3118
rect 14664 3694 14722 3706
rect 14664 3118 14676 3694
rect 14710 3118 14722 3694
rect 14664 3106 14722 3118
rect 15682 3694 15740 3706
rect 15682 3118 15694 3694
rect 15728 3118 15740 3694
rect 15682 3106 15740 3118
rect 16700 3694 16758 3706
rect 16700 3118 16712 3694
rect 16746 3118 16758 3694
rect 16700 3106 16758 3118
rect 17718 3694 17776 3706
rect 17718 3118 17730 3694
rect 17764 3118 17776 3694
rect 17718 3106 17776 3118
rect 19608 3436 19666 3448
rect 19608 2860 19620 3436
rect 19654 2860 19666 3436
rect 19608 2848 19666 2860
rect 20626 3436 20684 3448
rect 20626 2860 20638 3436
rect 20672 2860 20684 3436
rect 20626 2848 20684 2860
rect 21644 3436 21702 3448
rect 21644 2860 21656 3436
rect 21690 2860 21702 3436
rect 21644 2848 21702 2860
rect 22662 3436 22720 3448
rect 22662 2860 22674 3436
rect 22708 2860 22720 3436
rect 22662 2848 22720 2860
rect 23680 3436 23738 3448
rect 23680 2860 23692 3436
rect 23726 2860 23738 3436
rect 23680 2848 23738 2860
rect 24698 3436 24756 3448
rect 24698 2860 24710 3436
rect 24744 2860 24756 3436
rect 24698 2848 24756 2860
rect 25716 3436 25774 3448
rect 25716 2860 25728 3436
rect 25762 2860 25774 3436
rect 25716 2848 25774 2860
rect 26734 3436 26792 3448
rect 26734 2860 26746 3436
rect 26780 2860 26792 3436
rect 26734 2848 26792 2860
rect 27752 3436 27810 3448
rect 27752 2860 27764 3436
rect 27798 2860 27810 3436
rect 27752 2848 27810 2860
rect 28770 3436 28828 3448
rect 28770 2860 28782 3436
rect 28816 2860 28828 3436
rect 28770 2848 28828 2860
rect 29788 3436 29846 3448
rect 29788 2860 29800 3436
rect 29834 2860 29846 3436
rect 29788 2848 29846 2860
rect 30806 3436 30864 3448
rect 30806 2860 30818 3436
rect 30852 2860 30864 3436
rect 30806 2848 30864 2860
rect 31824 3436 31882 3448
rect 31824 2860 31836 3436
rect 31870 2860 31882 3436
rect 31824 2848 31882 2860
rect 32842 3436 32900 3448
rect 32842 2860 32854 3436
rect 32888 2860 32900 3436
rect 32842 2848 32900 2860
rect 33860 3436 33918 3448
rect 33860 2860 33872 3436
rect 33906 2860 33918 3436
rect 33860 2848 33918 2860
rect 34878 3436 34936 3448
rect 34878 2860 34890 3436
rect 34924 2860 34936 3436
rect 34878 2848 34936 2860
rect 35896 3436 35954 3448
rect 35896 2860 35908 3436
rect 35942 2860 35954 3436
rect 35896 2848 35954 2860
rect 36914 3436 36972 3448
rect 36914 2860 36926 3436
rect 36960 2860 36972 3436
rect 36914 2848 36972 2860
rect 37932 3436 37990 3448
rect 37932 2860 37944 3436
rect 37978 2860 37990 3436
rect 37932 2848 37990 2860
rect 38950 3436 39008 3448
rect 38950 2860 38962 3436
rect 38996 2860 39008 3436
rect 38950 2848 39008 2860
rect 39968 3436 40026 3448
rect 39968 2860 39980 3436
rect 40014 2860 40026 3436
rect 39968 2848 40026 2860
rect 6520 2582 6578 2594
rect 6520 2006 6532 2582
rect 6566 2006 6578 2582
rect 6520 1994 6578 2006
rect 7538 2582 7596 2594
rect 7538 2006 7550 2582
rect 7584 2006 7596 2582
rect 7538 1994 7596 2006
rect 8556 2582 8614 2594
rect 8556 2006 8568 2582
rect 8602 2006 8614 2582
rect 8556 1994 8614 2006
rect 9574 2582 9632 2594
rect 9574 2006 9586 2582
rect 9620 2006 9632 2582
rect 9574 1994 9632 2006
rect 10592 2582 10650 2594
rect 10592 2006 10604 2582
rect 10638 2006 10650 2582
rect 10592 1994 10650 2006
rect 11610 2582 11668 2594
rect 11610 2006 11622 2582
rect 11656 2006 11668 2582
rect 11610 1994 11668 2006
rect 12628 2582 12686 2594
rect 12628 2006 12640 2582
rect 12674 2006 12686 2582
rect 12628 1994 12686 2006
rect 13646 2582 13704 2594
rect 13646 2006 13658 2582
rect 13692 2006 13704 2582
rect 13646 1994 13704 2006
rect 14664 2582 14722 2594
rect 14664 2006 14676 2582
rect 14710 2006 14722 2582
rect 14664 1994 14722 2006
rect 15682 2582 15740 2594
rect 15682 2006 15694 2582
rect 15728 2006 15740 2582
rect 15682 1994 15740 2006
rect 16700 2582 16758 2594
rect 16700 2006 16712 2582
rect 16746 2006 16758 2582
rect 16700 1994 16758 2006
rect 17718 2582 17776 2594
rect 17718 2006 17730 2582
rect 17764 2006 17776 2582
rect 17718 1994 17776 2006
rect 19608 2204 19666 2216
rect 19608 1628 19620 2204
rect 19654 1628 19666 2204
rect 19608 1616 19666 1628
rect 20626 2204 20684 2216
rect 20626 1628 20638 2204
rect 20672 1628 20684 2204
rect 20626 1616 20684 1628
rect 21644 2204 21702 2216
rect 21644 1628 21656 2204
rect 21690 1628 21702 2204
rect 21644 1616 21702 1628
rect 22662 2204 22720 2216
rect 22662 1628 22674 2204
rect 22708 1628 22720 2204
rect 22662 1616 22720 1628
rect 23680 2204 23738 2216
rect 23680 1628 23692 2204
rect 23726 1628 23738 2204
rect 23680 1616 23738 1628
rect 24698 2204 24756 2216
rect 24698 1628 24710 2204
rect 24744 1628 24756 2204
rect 24698 1616 24756 1628
rect 25716 2204 25774 2216
rect 25716 1628 25728 2204
rect 25762 1628 25774 2204
rect 25716 1616 25774 1628
rect 26734 2204 26792 2216
rect 26734 1628 26746 2204
rect 26780 1628 26792 2204
rect 26734 1616 26792 1628
rect 27752 2204 27810 2216
rect 27752 1628 27764 2204
rect 27798 1628 27810 2204
rect 27752 1616 27810 1628
rect 28770 2204 28828 2216
rect 28770 1628 28782 2204
rect 28816 1628 28828 2204
rect 28770 1616 28828 1628
rect 29788 2204 29846 2216
rect 29788 1628 29800 2204
rect 29834 1628 29846 2204
rect 29788 1616 29846 1628
rect 30806 2204 30864 2216
rect 30806 1628 30818 2204
rect 30852 1628 30864 2204
rect 30806 1616 30864 1628
rect 31824 2204 31882 2216
rect 31824 1628 31836 2204
rect 31870 1628 31882 2204
rect 31824 1616 31882 1628
rect 32842 2204 32900 2216
rect 32842 1628 32854 2204
rect 32888 1628 32900 2204
rect 32842 1616 32900 1628
rect 33860 2204 33918 2216
rect 33860 1628 33872 2204
rect 33906 1628 33918 2204
rect 33860 1616 33918 1628
rect 34878 2204 34936 2216
rect 34878 1628 34890 2204
rect 34924 1628 34936 2204
rect 34878 1616 34936 1628
rect 35896 2204 35954 2216
rect 35896 1628 35908 2204
rect 35942 1628 35954 2204
rect 35896 1616 35954 1628
rect 36914 2204 36972 2216
rect 36914 1628 36926 2204
rect 36960 1628 36972 2204
rect 36914 1616 36972 1628
rect 37932 2204 37990 2216
rect 37932 1628 37944 2204
rect 37978 1628 37990 2204
rect 37932 1616 37990 1628
rect 38950 2204 39008 2216
rect 38950 1628 38962 2204
rect 38996 1628 39008 2204
rect 38950 1616 39008 1628
rect 39968 2204 40026 2216
rect 39968 1628 39980 2204
rect 40014 1628 40026 2204
rect 39968 1616 40026 1628
rect 6520 1470 6578 1482
rect 6520 894 6532 1470
rect 6566 894 6578 1470
rect 6520 882 6578 894
rect 7538 1470 7596 1482
rect 7538 894 7550 1470
rect 7584 894 7596 1470
rect 7538 882 7596 894
rect 8556 1470 8614 1482
rect 8556 894 8568 1470
rect 8602 894 8614 1470
rect 8556 882 8614 894
rect 9574 1470 9632 1482
rect 9574 894 9586 1470
rect 9620 894 9632 1470
rect 9574 882 9632 894
rect 10592 1470 10650 1482
rect 10592 894 10604 1470
rect 10638 894 10650 1470
rect 10592 882 10650 894
rect 11610 1470 11668 1482
rect 11610 894 11622 1470
rect 11656 894 11668 1470
rect 11610 882 11668 894
rect 12628 1470 12686 1482
rect 12628 894 12640 1470
rect 12674 894 12686 1470
rect 12628 882 12686 894
rect 13646 1470 13704 1482
rect 13646 894 13658 1470
rect 13692 894 13704 1470
rect 13646 882 13704 894
rect 14664 1470 14722 1482
rect 14664 894 14676 1470
rect 14710 894 14722 1470
rect 14664 882 14722 894
rect 15682 1470 15740 1482
rect 15682 894 15694 1470
rect 15728 894 15740 1470
rect 15682 882 15740 894
rect 16700 1470 16758 1482
rect 16700 894 16712 1470
rect 16746 894 16758 1470
rect 16700 882 16758 894
rect 17718 1470 17776 1482
rect 17718 894 17730 1470
rect 17764 894 17776 1470
rect 17718 882 17776 894
rect 19608 970 19666 982
rect 19608 394 19620 970
rect 19654 394 19666 970
rect 19608 382 19666 394
rect 20626 970 20684 982
rect 20626 394 20638 970
rect 20672 394 20684 970
rect 20626 382 20684 394
rect 21644 970 21702 982
rect 21644 394 21656 970
rect 21690 394 21702 970
rect 21644 382 21702 394
rect 22662 970 22720 982
rect 22662 394 22674 970
rect 22708 394 22720 970
rect 22662 382 22720 394
rect 23680 970 23738 982
rect 23680 394 23692 970
rect 23726 394 23738 970
rect 23680 382 23738 394
rect 24698 970 24756 982
rect 24698 394 24710 970
rect 24744 394 24756 970
rect 24698 382 24756 394
rect 25716 970 25774 982
rect 25716 394 25728 970
rect 25762 394 25774 970
rect 25716 382 25774 394
rect 26734 970 26792 982
rect 26734 394 26746 970
rect 26780 394 26792 970
rect 26734 382 26792 394
rect 27752 970 27810 982
rect 27752 394 27764 970
rect 27798 394 27810 970
rect 27752 382 27810 394
rect 28770 970 28828 982
rect 28770 394 28782 970
rect 28816 394 28828 970
rect 28770 382 28828 394
rect 29788 970 29846 982
rect 29788 394 29800 970
rect 29834 394 29846 970
rect 29788 382 29846 394
rect 30806 970 30864 982
rect 30806 394 30818 970
rect 30852 394 30864 970
rect 30806 382 30864 394
rect 31824 970 31882 982
rect 31824 394 31836 970
rect 31870 394 31882 970
rect 31824 382 31882 394
rect 32842 970 32900 982
rect 32842 394 32854 970
rect 32888 394 32900 970
rect 32842 382 32900 394
rect 33860 970 33918 982
rect 33860 394 33872 970
rect 33906 394 33918 970
rect 33860 382 33918 394
rect 34878 970 34936 982
rect 34878 394 34890 970
rect 34924 394 34936 970
rect 34878 382 34936 394
rect 35896 970 35954 982
rect 35896 394 35908 970
rect 35942 394 35954 970
rect 35896 382 35954 394
rect 36914 970 36972 982
rect 36914 394 36926 970
rect 36960 394 36972 970
rect 36914 382 36972 394
rect 37932 970 37990 982
rect 37932 394 37944 970
rect 37978 394 37990 970
rect 37932 382 37990 394
rect 38950 970 39008 982
rect 38950 394 38962 970
rect 38996 394 39008 970
rect 38950 382 39008 394
rect 39968 970 40026 982
rect 39968 394 39980 970
rect 40014 394 40026 970
rect 39968 382 40026 394
rect 6978 -72 7036 -60
rect 6978 -648 6990 -72
rect 7024 -648 7036 -72
rect 6978 -660 7036 -648
rect 7996 -72 8054 -60
rect 7996 -648 8008 -72
rect 8042 -648 8054 -72
rect 7996 -660 8054 -648
rect 9014 -72 9072 -60
rect 9014 -648 9026 -72
rect 9060 -648 9072 -72
rect 9014 -660 9072 -648
rect 10032 -72 10090 -60
rect 10032 -648 10044 -72
rect 10078 -648 10090 -72
rect 10032 -660 10090 -648
rect 11050 -72 11108 -60
rect 11050 -648 11062 -72
rect 11096 -648 11108 -72
rect 11050 -660 11108 -648
rect 12068 -72 12126 -60
rect 12068 -648 12080 -72
rect 12114 -648 12126 -72
rect 12068 -660 12126 -648
rect 13086 -72 13144 -60
rect 13086 -648 13098 -72
rect 13132 -648 13144 -72
rect 13086 -660 13144 -648
rect 14104 -72 14162 -60
rect 14104 -648 14116 -72
rect 14150 -648 14162 -72
rect 14104 -660 14162 -648
rect 15122 -72 15180 -60
rect 15122 -648 15134 -72
rect 15168 -648 15180 -72
rect 15122 -660 15180 -648
rect 16140 -72 16198 -60
rect 16140 -648 16152 -72
rect 16186 -648 16198 -72
rect 16140 -660 16198 -648
rect 17158 -72 17216 -60
rect 17158 -648 17170 -72
rect 17204 -648 17216 -72
rect 17158 -660 17216 -648
rect 19608 -262 19666 -250
rect 19608 -838 19620 -262
rect 19654 -838 19666 -262
rect 19608 -850 19666 -838
rect 20626 -262 20684 -250
rect 20626 -838 20638 -262
rect 20672 -838 20684 -262
rect 20626 -850 20684 -838
rect 21644 -262 21702 -250
rect 21644 -838 21656 -262
rect 21690 -838 21702 -262
rect 21644 -850 21702 -838
rect 22662 -262 22720 -250
rect 22662 -838 22674 -262
rect 22708 -838 22720 -262
rect 22662 -850 22720 -838
rect 23680 -262 23738 -250
rect 23680 -838 23692 -262
rect 23726 -838 23738 -262
rect 23680 -850 23738 -838
rect 24698 -262 24756 -250
rect 24698 -838 24710 -262
rect 24744 -838 24756 -262
rect 24698 -850 24756 -838
rect 25716 -262 25774 -250
rect 25716 -838 25728 -262
rect 25762 -838 25774 -262
rect 25716 -850 25774 -838
rect 26734 -262 26792 -250
rect 26734 -838 26746 -262
rect 26780 -838 26792 -262
rect 26734 -850 26792 -838
rect 27752 -262 27810 -250
rect 27752 -838 27764 -262
rect 27798 -838 27810 -262
rect 27752 -850 27810 -838
rect 28770 -262 28828 -250
rect 28770 -838 28782 -262
rect 28816 -838 28828 -262
rect 28770 -850 28828 -838
rect 29788 -262 29846 -250
rect 29788 -838 29800 -262
rect 29834 -838 29846 -262
rect 29788 -850 29846 -838
rect 30806 -262 30864 -250
rect 30806 -838 30818 -262
rect 30852 -838 30864 -262
rect 30806 -850 30864 -838
rect 31824 -262 31882 -250
rect 31824 -838 31836 -262
rect 31870 -838 31882 -262
rect 31824 -850 31882 -838
rect 32842 -262 32900 -250
rect 32842 -838 32854 -262
rect 32888 -838 32900 -262
rect 32842 -850 32900 -838
rect 33860 -262 33918 -250
rect 33860 -838 33872 -262
rect 33906 -838 33918 -262
rect 33860 -850 33918 -838
rect 34878 -262 34936 -250
rect 34878 -838 34890 -262
rect 34924 -838 34936 -262
rect 34878 -850 34936 -838
rect 35896 -262 35954 -250
rect 35896 -838 35908 -262
rect 35942 -838 35954 -262
rect 35896 -850 35954 -838
rect 36914 -262 36972 -250
rect 36914 -838 36926 -262
rect 36960 -838 36972 -262
rect 36914 -850 36972 -838
rect 37932 -262 37990 -250
rect 37932 -838 37944 -262
rect 37978 -838 37990 -262
rect 37932 -850 37990 -838
rect 38950 -262 39008 -250
rect 38950 -838 38962 -262
rect 38996 -838 39008 -262
rect 38950 -850 39008 -838
rect 39968 -262 40026 -250
rect 39968 -838 39980 -262
rect 40014 -838 40026 -262
rect 39968 -850 40026 -838
<< pdiff >>
rect 23516 26542 23574 26554
rect 23516 25966 23528 26542
rect 23562 25966 23574 26542
rect 23516 25954 23574 25966
rect 24534 26542 24592 26554
rect 24534 25966 24546 26542
rect 24580 25966 24592 26542
rect 24534 25954 24592 25966
rect 25552 26542 25610 26554
rect 25552 25966 25564 26542
rect 25598 25966 25610 26542
rect 25552 25954 25610 25966
rect 26570 26542 26628 26554
rect 26570 25966 26582 26542
rect 26616 25966 26628 26542
rect 26570 25954 26628 25966
rect 27588 26542 27646 26554
rect 27588 25966 27600 26542
rect 27634 25966 27646 26542
rect 27588 25954 27646 25966
rect 28606 26542 28664 26554
rect 28606 25966 28618 26542
rect 28652 25966 28664 26542
rect 28606 25954 28664 25966
rect 29624 26542 29682 26554
rect 29624 25966 29636 26542
rect 29670 25966 29682 26542
rect 29624 25954 29682 25966
rect 30642 26542 30700 26554
rect 30642 25966 30654 26542
rect 30688 25966 30700 26542
rect 30642 25954 30700 25966
rect 31660 26542 31718 26554
rect 31660 25966 31672 26542
rect 31706 25966 31718 26542
rect 31660 25954 31718 25966
rect 32678 26542 32736 26554
rect 32678 25966 32690 26542
rect 32724 25966 32736 26542
rect 32678 25954 32736 25966
rect 33696 26542 33754 26554
rect 33696 25966 33708 26542
rect 33742 25966 33754 26542
rect 33696 25954 33754 25966
rect 34714 26542 34772 26554
rect 34714 25966 34726 26542
rect 34760 25966 34772 26542
rect 34714 25954 34772 25966
rect 35732 26542 35790 26554
rect 35732 25966 35744 26542
rect 35778 25966 35790 26542
rect 35732 25954 35790 25966
rect 36750 26542 36808 26554
rect 36750 25966 36762 26542
rect 36796 25966 36808 26542
rect 36750 25954 36808 25966
rect 37768 26542 37826 26554
rect 37768 25966 37780 26542
rect 37814 25966 37826 26542
rect 37768 25954 37826 25966
rect 38786 26542 38844 26554
rect 38786 25966 38798 26542
rect 38832 25966 38844 26542
rect 38786 25954 38844 25966
rect 39804 26542 39862 26554
rect 39804 25966 39816 26542
rect 39850 25966 39862 26542
rect 39804 25954 39862 25966
rect 23516 25406 23574 25418
rect 23516 24830 23528 25406
rect 23562 24830 23574 25406
rect 23516 24818 23574 24830
rect 24534 25406 24592 25418
rect 24534 24830 24546 25406
rect 24580 24830 24592 25406
rect 24534 24818 24592 24830
rect 25552 25406 25610 25418
rect 25552 24830 25564 25406
rect 25598 24830 25610 25406
rect 25552 24818 25610 24830
rect 26570 25406 26628 25418
rect 26570 24830 26582 25406
rect 26616 24830 26628 25406
rect 26570 24818 26628 24830
rect 27588 25406 27646 25418
rect 27588 24830 27600 25406
rect 27634 24830 27646 25406
rect 27588 24818 27646 24830
rect 28606 25406 28664 25418
rect 28606 24830 28618 25406
rect 28652 24830 28664 25406
rect 28606 24818 28664 24830
rect 29624 25406 29682 25418
rect 29624 24830 29636 25406
rect 29670 24830 29682 25406
rect 29624 24818 29682 24830
rect 30642 25406 30700 25418
rect 30642 24830 30654 25406
rect 30688 24830 30700 25406
rect 30642 24818 30700 24830
rect 31660 25406 31718 25418
rect 31660 24830 31672 25406
rect 31706 24830 31718 25406
rect 31660 24818 31718 24830
rect 32678 25406 32736 25418
rect 32678 24830 32690 25406
rect 32724 24830 32736 25406
rect 32678 24818 32736 24830
rect 33696 25406 33754 25418
rect 33696 24830 33708 25406
rect 33742 24830 33754 25406
rect 33696 24818 33754 24830
rect 34714 25406 34772 25418
rect 34714 24830 34726 25406
rect 34760 24830 34772 25406
rect 34714 24818 34772 24830
rect 35732 25406 35790 25418
rect 35732 24830 35744 25406
rect 35778 24830 35790 25406
rect 35732 24818 35790 24830
rect 36750 25406 36808 25418
rect 36750 24830 36762 25406
rect 36796 24830 36808 25406
rect 36750 24818 36808 24830
rect 37768 25406 37826 25418
rect 37768 24830 37780 25406
rect 37814 24830 37826 25406
rect 37768 24818 37826 24830
rect 38786 25406 38844 25418
rect 38786 24830 38798 25406
rect 38832 24830 38844 25406
rect 38786 24818 38844 24830
rect 39804 25406 39862 25418
rect 39804 24830 39816 25406
rect 39850 24830 39862 25406
rect 39804 24818 39862 24830
rect 23516 24270 23574 24282
rect 23516 23694 23528 24270
rect 23562 23694 23574 24270
rect 23516 23682 23574 23694
rect 24534 24270 24592 24282
rect 24534 23694 24546 24270
rect 24580 23694 24592 24270
rect 24534 23682 24592 23694
rect 25552 24270 25610 24282
rect 25552 23694 25564 24270
rect 25598 23694 25610 24270
rect 25552 23682 25610 23694
rect 26570 24270 26628 24282
rect 26570 23694 26582 24270
rect 26616 23694 26628 24270
rect 26570 23682 26628 23694
rect 27588 24270 27646 24282
rect 27588 23694 27600 24270
rect 27634 23694 27646 24270
rect 27588 23682 27646 23694
rect 28606 24270 28664 24282
rect 28606 23694 28618 24270
rect 28652 23694 28664 24270
rect 28606 23682 28664 23694
rect 29624 24270 29682 24282
rect 29624 23694 29636 24270
rect 29670 23694 29682 24270
rect 29624 23682 29682 23694
rect 30642 24270 30700 24282
rect 30642 23694 30654 24270
rect 30688 23694 30700 24270
rect 30642 23682 30700 23694
rect 31660 24270 31718 24282
rect 31660 23694 31672 24270
rect 31706 23694 31718 24270
rect 31660 23682 31718 23694
rect 32678 24270 32736 24282
rect 32678 23694 32690 24270
rect 32724 23694 32736 24270
rect 32678 23682 32736 23694
rect 33696 24270 33754 24282
rect 33696 23694 33708 24270
rect 33742 23694 33754 24270
rect 33696 23682 33754 23694
rect 34714 24270 34772 24282
rect 34714 23694 34726 24270
rect 34760 23694 34772 24270
rect 34714 23682 34772 23694
rect 35732 24270 35790 24282
rect 35732 23694 35744 24270
rect 35778 23694 35790 24270
rect 35732 23682 35790 23694
rect 36750 24270 36808 24282
rect 36750 23694 36762 24270
rect 36796 23694 36808 24270
rect 36750 23682 36808 23694
rect 37768 24270 37826 24282
rect 37768 23694 37780 24270
rect 37814 23694 37826 24270
rect 37768 23682 37826 23694
rect 38786 24270 38844 24282
rect 38786 23694 38798 24270
rect 38832 23694 38844 24270
rect 38786 23682 38844 23694
rect 39804 24270 39862 24282
rect 39804 23694 39816 24270
rect 39850 23694 39862 24270
rect 39804 23682 39862 23694
rect 24710 22632 24768 22644
rect 24710 22056 24722 22632
rect 24756 22056 24768 22632
rect 24710 22044 24768 22056
rect 25728 22632 25786 22644
rect 25728 22056 25740 22632
rect 25774 22056 25786 22632
rect 25728 22044 25786 22056
rect 26746 22632 26804 22644
rect 26746 22056 26758 22632
rect 26792 22056 26804 22632
rect 26746 22044 26804 22056
rect 27764 22632 27822 22644
rect 27764 22056 27776 22632
rect 27810 22056 27822 22632
rect 27764 22044 27822 22056
rect 28782 22632 28840 22644
rect 28782 22056 28794 22632
rect 28828 22056 28840 22632
rect 28782 22044 28840 22056
rect 29800 22632 29858 22644
rect 29800 22056 29812 22632
rect 29846 22056 29858 22632
rect 29800 22044 29858 22056
rect 30818 22632 30876 22644
rect 30818 22056 30830 22632
rect 30864 22056 30876 22632
rect 30818 22044 30876 22056
rect 31836 22632 31894 22644
rect 31836 22056 31848 22632
rect 31882 22056 31894 22632
rect 31836 22044 31894 22056
rect 32854 22632 32912 22644
rect 32854 22056 32866 22632
rect 32900 22056 32912 22632
rect 32854 22044 32912 22056
rect 33872 22632 33930 22644
rect 33872 22056 33884 22632
rect 33918 22056 33930 22632
rect 33872 22044 33930 22056
rect 34890 22632 34948 22644
rect 34890 22056 34902 22632
rect 34936 22056 34948 22632
rect 34890 22044 34948 22056
rect 35908 22632 35966 22644
rect 35908 22056 35920 22632
rect 35954 22056 35966 22632
rect 35908 22044 35966 22056
rect 36926 22632 36984 22644
rect 36926 22056 36938 22632
rect 36972 22056 36984 22632
rect 36926 22044 36984 22056
rect 37944 22632 38002 22644
rect 37944 22056 37956 22632
rect 37990 22056 38002 22632
rect 37944 22044 38002 22056
rect 38962 22632 39020 22644
rect 38962 22056 38974 22632
rect 39008 22056 39020 22632
rect 38962 22044 39020 22056
rect 24710 21600 24768 21612
rect 24710 21024 24722 21600
rect 24756 21024 24768 21600
rect 24710 21012 24768 21024
rect 25728 21600 25786 21612
rect 25728 21024 25740 21600
rect 25774 21024 25786 21600
rect 25728 21012 25786 21024
rect 26746 21600 26804 21612
rect 26746 21024 26758 21600
rect 26792 21024 26804 21600
rect 26746 21012 26804 21024
rect 27764 21600 27822 21612
rect 27764 21024 27776 21600
rect 27810 21024 27822 21600
rect 27764 21012 27822 21024
rect 28782 21600 28840 21612
rect 28782 21024 28794 21600
rect 28828 21024 28840 21600
rect 28782 21012 28840 21024
rect 29800 21600 29858 21612
rect 29800 21024 29812 21600
rect 29846 21024 29858 21600
rect 29800 21012 29858 21024
rect 30818 21600 30876 21612
rect 30818 21024 30830 21600
rect 30864 21024 30876 21600
rect 30818 21012 30876 21024
rect 31836 21600 31894 21612
rect 31836 21024 31848 21600
rect 31882 21024 31894 21600
rect 31836 21012 31894 21024
rect 32854 21600 32912 21612
rect 32854 21024 32866 21600
rect 32900 21024 32912 21600
rect 32854 21012 32912 21024
rect 33872 21600 33930 21612
rect 33872 21024 33884 21600
rect 33918 21024 33930 21600
rect 33872 21012 33930 21024
rect 34890 21600 34948 21612
rect 34890 21024 34902 21600
rect 34936 21024 34948 21600
rect 34890 21012 34948 21024
rect 35908 21600 35966 21612
rect 35908 21024 35920 21600
rect 35954 21024 35966 21600
rect 35908 21012 35966 21024
rect 36926 21600 36984 21612
rect 36926 21024 36938 21600
rect 36972 21024 36984 21600
rect 36926 21012 36984 21024
rect 37944 21600 38002 21612
rect 37944 21024 37956 21600
rect 37990 21024 38002 21600
rect 37944 21012 38002 21024
rect 38962 21600 39020 21612
rect 38962 21024 38974 21600
rect 39008 21024 39020 21600
rect 38962 21012 39020 21024
rect 24502 19996 24560 20008
rect 19198 19892 19256 19904
rect 19198 19316 19210 19892
rect 19244 19316 19256 19892
rect 19198 19304 19256 19316
rect 20216 19892 20274 19904
rect 20216 19316 20228 19892
rect 20262 19316 20274 19892
rect 20216 19304 20274 19316
rect 21234 19892 21292 19904
rect 21234 19316 21246 19892
rect 21280 19316 21292 19892
rect 21234 19304 21292 19316
rect 22252 19892 22310 19904
rect 22252 19316 22264 19892
rect 22298 19316 22310 19892
rect 22252 19304 22310 19316
rect 23270 19892 23328 19904
rect 23270 19316 23282 19892
rect 23316 19316 23328 19892
rect 24502 19420 24514 19996
rect 24548 19420 24560 19996
rect 24502 19408 24560 19420
rect 25520 19996 25578 20008
rect 25520 19420 25532 19996
rect 25566 19420 25578 19996
rect 25520 19408 25578 19420
rect 26538 19996 26596 20008
rect 26538 19420 26550 19996
rect 26584 19420 26596 19996
rect 26538 19408 26596 19420
rect 27556 19996 27614 20008
rect 27556 19420 27568 19996
rect 27602 19420 27614 19996
rect 27556 19408 27614 19420
rect 28574 19996 28632 20008
rect 28574 19420 28586 19996
rect 28620 19420 28632 19996
rect 28574 19408 28632 19420
rect 29592 19996 29650 20008
rect 29592 19420 29604 19996
rect 29638 19420 29650 19996
rect 29592 19408 29650 19420
rect 30610 19996 30668 20008
rect 30610 19420 30622 19996
rect 30656 19420 30668 19996
rect 30610 19408 30668 19420
rect 31628 19996 31686 20008
rect 31628 19420 31640 19996
rect 31674 19420 31686 19996
rect 31628 19408 31686 19420
rect 32646 19996 32704 20008
rect 32646 19420 32658 19996
rect 32692 19420 32704 19996
rect 32646 19408 32704 19420
rect 33664 19996 33722 20008
rect 33664 19420 33676 19996
rect 33710 19420 33722 19996
rect 33664 19408 33722 19420
rect 34682 19996 34740 20008
rect 34682 19420 34694 19996
rect 34728 19420 34740 19996
rect 34682 19408 34740 19420
rect 35700 19996 35758 20008
rect 35700 19420 35712 19996
rect 35746 19420 35758 19996
rect 35700 19408 35758 19420
rect 36718 19996 36776 20008
rect 36718 19420 36730 19996
rect 36764 19420 36776 19996
rect 36718 19408 36776 19420
rect 37736 19996 37794 20008
rect 37736 19420 37748 19996
rect 37782 19420 37794 19996
rect 37736 19408 37794 19420
rect 38754 19996 38812 20008
rect 38754 19420 38766 19996
rect 38800 19420 38812 19996
rect 38754 19408 38812 19420
rect 39772 19996 39830 20008
rect 39772 19420 39784 19996
rect 39818 19420 39830 19996
rect 39772 19408 39830 19420
rect 23270 19304 23328 19316
rect 19198 18860 19256 18872
rect 19198 18284 19210 18860
rect 19244 18284 19256 18860
rect 19198 18272 19256 18284
rect 20216 18860 20274 18872
rect 20216 18284 20228 18860
rect 20262 18284 20274 18860
rect 20216 18272 20274 18284
rect 21234 18860 21292 18872
rect 21234 18284 21246 18860
rect 21280 18284 21292 18860
rect 21234 18272 21292 18284
rect 22252 18860 22310 18872
rect 22252 18284 22264 18860
rect 22298 18284 22310 18860
rect 22252 18272 22310 18284
rect 23270 18860 23328 18872
rect 23270 18284 23282 18860
rect 23316 18284 23328 18860
rect 23270 18272 23328 18284
rect 24502 18740 24560 18752
rect 24502 18164 24514 18740
rect 24548 18164 24560 18740
rect 24502 18152 24560 18164
rect 25520 18740 25578 18752
rect 25520 18164 25532 18740
rect 25566 18164 25578 18740
rect 25520 18152 25578 18164
rect 26538 18740 26596 18752
rect 26538 18164 26550 18740
rect 26584 18164 26596 18740
rect 26538 18152 26596 18164
rect 27556 18740 27614 18752
rect 27556 18164 27568 18740
rect 27602 18164 27614 18740
rect 27556 18152 27614 18164
rect 28574 18740 28632 18752
rect 28574 18164 28586 18740
rect 28620 18164 28632 18740
rect 28574 18152 28632 18164
rect 29592 18740 29650 18752
rect 29592 18164 29604 18740
rect 29638 18164 29650 18740
rect 29592 18152 29650 18164
rect 30610 18740 30668 18752
rect 30610 18164 30622 18740
rect 30656 18164 30668 18740
rect 30610 18152 30668 18164
rect 31628 18740 31686 18752
rect 31628 18164 31640 18740
rect 31674 18164 31686 18740
rect 31628 18152 31686 18164
rect 32646 18740 32704 18752
rect 32646 18164 32658 18740
rect 32692 18164 32704 18740
rect 32646 18152 32704 18164
rect 33664 18740 33722 18752
rect 33664 18164 33676 18740
rect 33710 18164 33722 18740
rect 33664 18152 33722 18164
rect 34682 18740 34740 18752
rect 34682 18164 34694 18740
rect 34728 18164 34740 18740
rect 34682 18152 34740 18164
rect 35700 18740 35758 18752
rect 35700 18164 35712 18740
rect 35746 18164 35758 18740
rect 35700 18152 35758 18164
rect 36718 18740 36776 18752
rect 36718 18164 36730 18740
rect 36764 18164 36776 18740
rect 36718 18152 36776 18164
rect 37736 18740 37794 18752
rect 37736 18164 37748 18740
rect 37782 18164 37794 18740
rect 37736 18152 37794 18164
rect 38754 18740 38812 18752
rect 38754 18164 38766 18740
rect 38800 18164 38812 18740
rect 38754 18152 38812 18164
rect 39772 18740 39830 18752
rect 39772 18164 39784 18740
rect 39818 18164 39830 18740
rect 39772 18152 39830 18164
rect 19198 17828 19256 17840
rect 19198 17252 19210 17828
rect 19244 17252 19256 17828
rect 19198 17240 19256 17252
rect 20216 17828 20274 17840
rect 20216 17252 20228 17828
rect 20262 17252 20274 17828
rect 20216 17240 20274 17252
rect 21234 17828 21292 17840
rect 21234 17252 21246 17828
rect 21280 17252 21292 17828
rect 21234 17240 21292 17252
rect 22252 17828 22310 17840
rect 22252 17252 22264 17828
rect 22298 17252 22310 17828
rect 22252 17240 22310 17252
rect 23270 17828 23328 17840
rect 23270 17252 23282 17828
rect 23316 17252 23328 17828
rect 23270 17240 23328 17252
rect 24502 17484 24560 17496
rect 24502 16908 24514 17484
rect 24548 16908 24560 17484
rect 24502 16896 24560 16908
rect 25520 17484 25578 17496
rect 25520 16908 25532 17484
rect 25566 16908 25578 17484
rect 25520 16896 25578 16908
rect 26538 17484 26596 17496
rect 26538 16908 26550 17484
rect 26584 16908 26596 17484
rect 26538 16896 26596 16908
rect 27556 17484 27614 17496
rect 27556 16908 27568 17484
rect 27602 16908 27614 17484
rect 27556 16896 27614 16908
rect 28574 17484 28632 17496
rect 28574 16908 28586 17484
rect 28620 16908 28632 17484
rect 28574 16896 28632 16908
rect 29592 17484 29650 17496
rect 29592 16908 29604 17484
rect 29638 16908 29650 17484
rect 29592 16896 29650 16908
rect 30610 17484 30668 17496
rect 30610 16908 30622 17484
rect 30656 16908 30668 17484
rect 30610 16896 30668 16908
rect 31628 17484 31686 17496
rect 31628 16908 31640 17484
rect 31674 16908 31686 17484
rect 31628 16896 31686 16908
rect 32646 17484 32704 17496
rect 32646 16908 32658 17484
rect 32692 16908 32704 17484
rect 32646 16896 32704 16908
rect 33664 17484 33722 17496
rect 33664 16908 33676 17484
rect 33710 16908 33722 17484
rect 33664 16896 33722 16908
rect 34682 17484 34740 17496
rect 34682 16908 34694 17484
rect 34728 16908 34740 17484
rect 34682 16896 34740 16908
rect 35700 17484 35758 17496
rect 35700 16908 35712 17484
rect 35746 16908 35758 17484
rect 35700 16896 35758 16908
rect 36718 17484 36776 17496
rect 36718 16908 36730 17484
rect 36764 16908 36776 17484
rect 36718 16896 36776 16908
rect 37736 17484 37794 17496
rect 37736 16908 37748 17484
rect 37782 16908 37794 17484
rect 37736 16896 37794 16908
rect 38754 17484 38812 17496
rect 38754 16908 38766 17484
rect 38800 16908 38812 17484
rect 38754 16896 38812 16908
rect 39772 17484 39830 17496
rect 39772 16908 39784 17484
rect 39818 16908 39830 17484
rect 39772 16896 39830 16908
rect 19198 16796 19256 16808
rect 19198 16220 19210 16796
rect 19244 16220 19256 16796
rect 19198 16208 19256 16220
rect 20216 16796 20274 16808
rect 20216 16220 20228 16796
rect 20262 16220 20274 16796
rect 20216 16208 20274 16220
rect 21234 16796 21292 16808
rect 21234 16220 21246 16796
rect 21280 16220 21292 16796
rect 21234 16208 21292 16220
rect 22252 16796 22310 16808
rect 22252 16220 22264 16796
rect 22298 16220 22310 16796
rect 22252 16208 22310 16220
rect 23270 16796 23328 16808
rect 23270 16220 23282 16796
rect 23316 16220 23328 16796
rect 23270 16208 23328 16220
rect 24502 16228 24560 16240
rect 24502 15652 24514 16228
rect 24548 15652 24560 16228
rect 24502 15640 24560 15652
rect 25520 16228 25578 16240
rect 25520 15652 25532 16228
rect 25566 15652 25578 16228
rect 25520 15640 25578 15652
rect 26538 16228 26596 16240
rect 26538 15652 26550 16228
rect 26584 15652 26596 16228
rect 26538 15640 26596 15652
rect 27556 16228 27614 16240
rect 27556 15652 27568 16228
rect 27602 15652 27614 16228
rect 27556 15640 27614 15652
rect 28574 16228 28632 16240
rect 28574 15652 28586 16228
rect 28620 15652 28632 16228
rect 28574 15640 28632 15652
rect 29592 16228 29650 16240
rect 29592 15652 29604 16228
rect 29638 15652 29650 16228
rect 29592 15640 29650 15652
rect 30610 16228 30668 16240
rect 30610 15652 30622 16228
rect 30656 15652 30668 16228
rect 30610 15640 30668 15652
rect 31628 16228 31686 16240
rect 31628 15652 31640 16228
rect 31674 15652 31686 16228
rect 31628 15640 31686 15652
rect 32646 16228 32704 16240
rect 32646 15652 32658 16228
rect 32692 15652 32704 16228
rect 32646 15640 32704 15652
rect 33664 16228 33722 16240
rect 33664 15652 33676 16228
rect 33710 15652 33722 16228
rect 33664 15640 33722 15652
rect 34682 16228 34740 16240
rect 34682 15652 34694 16228
rect 34728 15652 34740 16228
rect 34682 15640 34740 15652
rect 35700 16228 35758 16240
rect 35700 15652 35712 16228
rect 35746 15652 35758 16228
rect 35700 15640 35758 15652
rect 36718 16228 36776 16240
rect 36718 15652 36730 16228
rect 36764 15652 36776 16228
rect 36718 15640 36776 15652
rect 37736 16228 37794 16240
rect 37736 15652 37748 16228
rect 37782 15652 37794 16228
rect 37736 15640 37794 15652
rect 38754 16228 38812 16240
rect 38754 15652 38766 16228
rect 38800 15652 38812 16228
rect 38754 15640 38812 15652
rect 39772 16228 39830 16240
rect 39772 15652 39784 16228
rect 39818 15652 39830 16228
rect 39772 15640 39830 15652
<< ndiffc >>
rect 286 54 320 430
rect 544 54 578 430
rect 802 54 836 430
rect 1060 54 1094 430
rect 1318 54 1352 430
rect 1576 54 1610 430
rect 1834 54 1868 430
rect 2092 54 2126 430
rect 2350 54 2384 430
rect 2608 54 2642 430
rect 2866 54 2900 430
rect 3124 54 3158 430
rect 3382 54 3416 430
rect 3640 54 3674 430
rect 3898 54 3932 430
rect 286 -946 320 -570
rect 544 -946 578 -570
rect 802 -946 836 -570
rect 1060 -946 1094 -570
rect 1318 -946 1352 -570
rect 1576 -946 1610 -570
rect 1834 -946 1868 -570
rect 2092 -946 2126 -570
rect 2350 -946 2384 -570
rect 2608 -946 2642 -570
rect 2866 -946 2900 -570
rect 3124 -946 3158 -570
rect 3382 -946 3416 -570
rect 3640 -946 3674 -570
rect 3898 -946 3932 -570
rect 7856 11980 7890 12556
rect 8874 11980 8908 12556
rect 9892 11980 9926 12556
rect 10910 11980 10944 12556
rect 11928 11980 11962 12556
rect 12946 11980 12980 12556
rect 13964 11980 13998 12556
rect 14982 11980 15016 12556
rect 16000 11980 16034 12556
rect 17018 11980 17052 12556
rect 19622 12456 19656 13032
rect 20640 12456 20674 13032
rect 21658 12456 21692 13032
rect 22676 12456 22710 13032
rect 23694 12456 23728 13032
rect 24712 12456 24746 13032
rect 25730 12456 25764 13032
rect 26748 12456 26782 13032
rect 27766 12456 27800 13032
rect 28784 12456 28818 13032
rect 29802 12456 29836 13032
rect 30820 12456 30854 13032
rect 31838 12456 31872 13032
rect 32856 12456 32890 13032
rect 33874 12456 33908 13032
rect 34892 12456 34926 13032
rect 35910 12456 35944 13032
rect 36928 12456 36962 13032
rect 37946 12456 37980 13032
rect 38964 12456 38998 13032
rect 39982 12456 40016 13032
rect 7856 11162 7890 11738
rect 8874 11162 8908 11738
rect 9892 11162 9926 11738
rect 10910 11162 10944 11738
rect 11928 11162 11962 11738
rect 12946 11162 12980 11738
rect 13964 11162 13998 11738
rect 14982 11162 15016 11738
rect 16000 11162 16034 11738
rect 17018 11162 17052 11738
rect 19622 11638 19656 12214
rect 20640 11638 20674 12214
rect 21658 11638 21692 12214
rect 22676 11638 22710 12214
rect 23694 11638 23728 12214
rect 24712 11638 24746 12214
rect 25730 11638 25764 12214
rect 26748 11638 26782 12214
rect 27766 11638 27800 12214
rect 28784 11638 28818 12214
rect 29802 11638 29836 12214
rect 30820 11638 30854 12214
rect 31838 11638 31872 12214
rect 32856 11638 32890 12214
rect 33874 11638 33908 12214
rect 34892 11638 34926 12214
rect 35910 11638 35944 12214
rect 36928 11638 36962 12214
rect 37946 11638 37980 12214
rect 38964 11638 38998 12214
rect 39982 11638 40016 12214
rect 7856 10344 7890 10920
rect 8874 10344 8908 10920
rect 9892 10344 9926 10920
rect 10910 10344 10944 10920
rect 11928 10344 11962 10920
rect 12946 10344 12980 10920
rect 13964 10344 13998 10920
rect 14982 10344 15016 10920
rect 16000 10344 16034 10920
rect 17018 10344 17052 10920
rect 19622 10260 19656 10836
rect 20640 10260 20674 10836
rect 21658 10260 21692 10836
rect 22676 10260 22710 10836
rect 23694 10260 23728 10836
rect 24712 10260 24746 10836
rect 25730 10260 25764 10836
rect 26748 10260 26782 10836
rect 27766 10260 27800 10836
rect 28784 10260 28818 10836
rect 29802 10260 29836 10836
rect 30820 10260 30854 10836
rect 31838 10260 31872 10836
rect 32856 10260 32890 10836
rect 33874 10260 33908 10836
rect 34892 10260 34926 10836
rect 35910 10260 35944 10836
rect 36928 10260 36962 10836
rect 37946 10260 37980 10836
rect 38964 10260 38998 10836
rect 39982 10260 40016 10836
rect 7856 9526 7890 10102
rect 8874 9526 8908 10102
rect 9892 9526 9926 10102
rect 10910 9526 10944 10102
rect 11928 9526 11962 10102
rect 12946 9526 12980 10102
rect 13964 9526 13998 10102
rect 14982 9526 15016 10102
rect 16000 9526 16034 10102
rect 17018 9526 17052 10102
rect 7856 8708 7890 9284
rect 8874 8708 8908 9284
rect 9892 8708 9926 9284
rect 10910 8708 10944 9284
rect 11928 8708 11962 9284
rect 12946 8708 12980 9284
rect 13964 8708 13998 9284
rect 14982 8708 15016 9284
rect 16000 8708 16034 9284
rect 17018 8708 17052 9284
rect 19622 9028 19656 9604
rect 20640 9028 20674 9604
rect 21658 9028 21692 9604
rect 22676 9028 22710 9604
rect 23694 9028 23728 9604
rect 24712 9028 24746 9604
rect 25730 9028 25764 9604
rect 26748 9028 26782 9604
rect 27766 9028 27800 9604
rect 28784 9028 28818 9604
rect 29802 9028 29836 9604
rect 30820 9028 30854 9604
rect 31838 9028 31872 9604
rect 32856 9028 32890 9604
rect 33874 9028 33908 9604
rect 34892 9028 34926 9604
rect 35910 9028 35944 9604
rect 36928 9028 36962 9604
rect 37946 9028 37980 9604
rect 38964 9028 38998 9604
rect 39982 9028 40016 9604
rect 7856 7890 7890 8466
rect 8874 7890 8908 8466
rect 9892 7890 9926 8466
rect 10910 7890 10944 8466
rect 11928 7890 11962 8466
rect 12946 7890 12980 8466
rect 13964 7890 13998 8466
rect 14982 7890 15016 8466
rect 16000 7890 16034 8466
rect 17018 7890 17052 8466
rect 19620 7794 19654 8370
rect 20638 7794 20672 8370
rect 21656 7794 21690 8370
rect 22674 7794 22708 8370
rect 23692 7794 23726 8370
rect 24710 7794 24744 8370
rect 25728 7794 25762 8370
rect 26746 7794 26780 8370
rect 27764 7794 27798 8370
rect 28782 7794 28816 8370
rect 29800 7794 29834 8370
rect 30818 7794 30852 8370
rect 31836 7794 31870 8370
rect 32854 7794 32888 8370
rect 33872 7794 33906 8370
rect 34890 7794 34924 8370
rect 35908 7794 35942 8370
rect 36926 7794 36960 8370
rect 37944 7794 37978 8370
rect 38962 7794 38996 8370
rect 39980 7794 40014 8370
rect 7856 7072 7890 7648
rect 8874 7072 8908 7648
rect 9892 7072 9926 7648
rect 10910 7072 10944 7648
rect 11928 7072 11962 7648
rect 12946 7072 12980 7648
rect 13964 7072 13998 7648
rect 14982 7072 15016 7648
rect 16000 7072 16034 7648
rect 17018 7072 17052 7648
rect 7856 6254 7890 6830
rect 8874 6254 8908 6830
rect 9892 6254 9926 6830
rect 10910 6254 10944 6830
rect 11928 6254 11962 6830
rect 12946 6254 12980 6830
rect 13964 6254 13998 6830
rect 14982 6254 15016 6830
rect 16000 6254 16034 6830
rect 17018 6254 17052 6830
rect 19620 6560 19654 7136
rect 20638 6560 20672 7136
rect 21656 6560 21690 7136
rect 22674 6560 22708 7136
rect 23692 6560 23726 7136
rect 24710 6560 24744 7136
rect 25728 6560 25762 7136
rect 26746 6560 26780 7136
rect 27764 6560 27798 7136
rect 28782 6560 28816 7136
rect 29800 6560 29834 7136
rect 30818 6560 30852 7136
rect 31836 6560 31870 7136
rect 32854 6560 32888 7136
rect 33872 6560 33906 7136
rect 34890 6560 34924 7136
rect 35908 6560 35942 7136
rect 36926 6560 36960 7136
rect 37944 6560 37978 7136
rect 38962 6560 38996 7136
rect 39980 6560 40014 7136
rect 19620 5328 19654 5904
rect 20638 5328 20672 5904
rect 21656 5328 21690 5904
rect 22674 5328 22708 5904
rect 23692 5328 23726 5904
rect 24710 5328 24744 5904
rect 25728 5328 25762 5904
rect 26746 5328 26780 5904
rect 27764 5328 27798 5904
rect 28782 5328 28816 5904
rect 29800 5328 29834 5904
rect 30818 5328 30852 5904
rect 31836 5328 31870 5904
rect 32854 5328 32888 5904
rect 33872 5328 33906 5904
rect 34890 5328 34924 5904
rect 35908 5328 35942 5904
rect 36926 5328 36960 5904
rect 37944 5328 37978 5904
rect 38962 5328 38996 5904
rect 39980 5328 40014 5904
rect 6532 4230 6566 4806
rect 7550 4230 7584 4806
rect 8568 4230 8602 4806
rect 9586 4230 9620 4806
rect 10604 4230 10638 4806
rect 11622 4230 11656 4806
rect 12640 4230 12674 4806
rect 13658 4230 13692 4806
rect 14676 4230 14710 4806
rect 15694 4230 15728 4806
rect 16712 4230 16746 4806
rect 17730 4230 17764 4806
rect 19620 4094 19654 4670
rect 20638 4094 20672 4670
rect 21656 4094 21690 4670
rect 22674 4094 22708 4670
rect 23692 4094 23726 4670
rect 24710 4094 24744 4670
rect 25728 4094 25762 4670
rect 26746 4094 26780 4670
rect 27764 4094 27798 4670
rect 28782 4094 28816 4670
rect 29800 4094 29834 4670
rect 30818 4094 30852 4670
rect 31836 4094 31870 4670
rect 32854 4094 32888 4670
rect 33872 4094 33906 4670
rect 34890 4094 34924 4670
rect 35908 4094 35942 4670
rect 36926 4094 36960 4670
rect 37944 4094 37978 4670
rect 38962 4094 38996 4670
rect 39980 4094 40014 4670
rect 6532 3118 6566 3694
rect 7550 3118 7584 3694
rect 8568 3118 8602 3694
rect 9586 3118 9620 3694
rect 10604 3118 10638 3694
rect 11622 3118 11656 3694
rect 12640 3118 12674 3694
rect 13658 3118 13692 3694
rect 14676 3118 14710 3694
rect 15694 3118 15728 3694
rect 16712 3118 16746 3694
rect 17730 3118 17764 3694
rect 19620 2860 19654 3436
rect 20638 2860 20672 3436
rect 21656 2860 21690 3436
rect 22674 2860 22708 3436
rect 23692 2860 23726 3436
rect 24710 2860 24744 3436
rect 25728 2860 25762 3436
rect 26746 2860 26780 3436
rect 27764 2860 27798 3436
rect 28782 2860 28816 3436
rect 29800 2860 29834 3436
rect 30818 2860 30852 3436
rect 31836 2860 31870 3436
rect 32854 2860 32888 3436
rect 33872 2860 33906 3436
rect 34890 2860 34924 3436
rect 35908 2860 35942 3436
rect 36926 2860 36960 3436
rect 37944 2860 37978 3436
rect 38962 2860 38996 3436
rect 39980 2860 40014 3436
rect 6532 2006 6566 2582
rect 7550 2006 7584 2582
rect 8568 2006 8602 2582
rect 9586 2006 9620 2582
rect 10604 2006 10638 2582
rect 11622 2006 11656 2582
rect 12640 2006 12674 2582
rect 13658 2006 13692 2582
rect 14676 2006 14710 2582
rect 15694 2006 15728 2582
rect 16712 2006 16746 2582
rect 17730 2006 17764 2582
rect 19620 1628 19654 2204
rect 20638 1628 20672 2204
rect 21656 1628 21690 2204
rect 22674 1628 22708 2204
rect 23692 1628 23726 2204
rect 24710 1628 24744 2204
rect 25728 1628 25762 2204
rect 26746 1628 26780 2204
rect 27764 1628 27798 2204
rect 28782 1628 28816 2204
rect 29800 1628 29834 2204
rect 30818 1628 30852 2204
rect 31836 1628 31870 2204
rect 32854 1628 32888 2204
rect 33872 1628 33906 2204
rect 34890 1628 34924 2204
rect 35908 1628 35942 2204
rect 36926 1628 36960 2204
rect 37944 1628 37978 2204
rect 38962 1628 38996 2204
rect 39980 1628 40014 2204
rect 6532 894 6566 1470
rect 7550 894 7584 1470
rect 8568 894 8602 1470
rect 9586 894 9620 1470
rect 10604 894 10638 1470
rect 11622 894 11656 1470
rect 12640 894 12674 1470
rect 13658 894 13692 1470
rect 14676 894 14710 1470
rect 15694 894 15728 1470
rect 16712 894 16746 1470
rect 17730 894 17764 1470
rect 19620 394 19654 970
rect 20638 394 20672 970
rect 21656 394 21690 970
rect 22674 394 22708 970
rect 23692 394 23726 970
rect 24710 394 24744 970
rect 25728 394 25762 970
rect 26746 394 26780 970
rect 27764 394 27798 970
rect 28782 394 28816 970
rect 29800 394 29834 970
rect 30818 394 30852 970
rect 31836 394 31870 970
rect 32854 394 32888 970
rect 33872 394 33906 970
rect 34890 394 34924 970
rect 35908 394 35942 970
rect 36926 394 36960 970
rect 37944 394 37978 970
rect 38962 394 38996 970
rect 39980 394 40014 970
rect 6990 -648 7024 -72
rect 8008 -648 8042 -72
rect 9026 -648 9060 -72
rect 10044 -648 10078 -72
rect 11062 -648 11096 -72
rect 12080 -648 12114 -72
rect 13098 -648 13132 -72
rect 14116 -648 14150 -72
rect 15134 -648 15168 -72
rect 16152 -648 16186 -72
rect 17170 -648 17204 -72
rect 19620 -838 19654 -262
rect 20638 -838 20672 -262
rect 21656 -838 21690 -262
rect 22674 -838 22708 -262
rect 23692 -838 23726 -262
rect 24710 -838 24744 -262
rect 25728 -838 25762 -262
rect 26746 -838 26780 -262
rect 27764 -838 27798 -262
rect 28782 -838 28816 -262
rect 29800 -838 29834 -262
rect 30818 -838 30852 -262
rect 31836 -838 31870 -262
rect 32854 -838 32888 -262
rect 33872 -838 33906 -262
rect 34890 -838 34924 -262
rect 35908 -838 35942 -262
rect 36926 -838 36960 -262
rect 37944 -838 37978 -262
rect 38962 -838 38996 -262
rect 39980 -838 40014 -262
<< pdiffc >>
rect 23528 25966 23562 26542
rect 24546 25966 24580 26542
rect 25564 25966 25598 26542
rect 26582 25966 26616 26542
rect 27600 25966 27634 26542
rect 28618 25966 28652 26542
rect 29636 25966 29670 26542
rect 30654 25966 30688 26542
rect 31672 25966 31706 26542
rect 32690 25966 32724 26542
rect 33708 25966 33742 26542
rect 34726 25966 34760 26542
rect 35744 25966 35778 26542
rect 36762 25966 36796 26542
rect 37780 25966 37814 26542
rect 38798 25966 38832 26542
rect 39816 25966 39850 26542
rect 23528 24830 23562 25406
rect 24546 24830 24580 25406
rect 25564 24830 25598 25406
rect 26582 24830 26616 25406
rect 27600 24830 27634 25406
rect 28618 24830 28652 25406
rect 29636 24830 29670 25406
rect 30654 24830 30688 25406
rect 31672 24830 31706 25406
rect 32690 24830 32724 25406
rect 33708 24830 33742 25406
rect 34726 24830 34760 25406
rect 35744 24830 35778 25406
rect 36762 24830 36796 25406
rect 37780 24830 37814 25406
rect 38798 24830 38832 25406
rect 39816 24830 39850 25406
rect 23528 23694 23562 24270
rect 24546 23694 24580 24270
rect 25564 23694 25598 24270
rect 26582 23694 26616 24270
rect 27600 23694 27634 24270
rect 28618 23694 28652 24270
rect 29636 23694 29670 24270
rect 30654 23694 30688 24270
rect 31672 23694 31706 24270
rect 32690 23694 32724 24270
rect 33708 23694 33742 24270
rect 34726 23694 34760 24270
rect 35744 23694 35778 24270
rect 36762 23694 36796 24270
rect 37780 23694 37814 24270
rect 38798 23694 38832 24270
rect 39816 23694 39850 24270
rect 24722 22056 24756 22632
rect 25740 22056 25774 22632
rect 26758 22056 26792 22632
rect 27776 22056 27810 22632
rect 28794 22056 28828 22632
rect 29812 22056 29846 22632
rect 30830 22056 30864 22632
rect 31848 22056 31882 22632
rect 32866 22056 32900 22632
rect 33884 22056 33918 22632
rect 34902 22056 34936 22632
rect 35920 22056 35954 22632
rect 36938 22056 36972 22632
rect 37956 22056 37990 22632
rect 38974 22056 39008 22632
rect 24722 21024 24756 21600
rect 25740 21024 25774 21600
rect 26758 21024 26792 21600
rect 27776 21024 27810 21600
rect 28794 21024 28828 21600
rect 29812 21024 29846 21600
rect 30830 21024 30864 21600
rect 31848 21024 31882 21600
rect 32866 21024 32900 21600
rect 33884 21024 33918 21600
rect 34902 21024 34936 21600
rect 35920 21024 35954 21600
rect 36938 21024 36972 21600
rect 37956 21024 37990 21600
rect 38974 21024 39008 21600
rect 19210 19316 19244 19892
rect 20228 19316 20262 19892
rect 21246 19316 21280 19892
rect 22264 19316 22298 19892
rect 23282 19316 23316 19892
rect 24514 19420 24548 19996
rect 25532 19420 25566 19996
rect 26550 19420 26584 19996
rect 27568 19420 27602 19996
rect 28586 19420 28620 19996
rect 29604 19420 29638 19996
rect 30622 19420 30656 19996
rect 31640 19420 31674 19996
rect 32658 19420 32692 19996
rect 33676 19420 33710 19996
rect 34694 19420 34728 19996
rect 35712 19420 35746 19996
rect 36730 19420 36764 19996
rect 37748 19420 37782 19996
rect 38766 19420 38800 19996
rect 39784 19420 39818 19996
rect 19210 18284 19244 18860
rect 20228 18284 20262 18860
rect 21246 18284 21280 18860
rect 22264 18284 22298 18860
rect 23282 18284 23316 18860
rect 24514 18164 24548 18740
rect 25532 18164 25566 18740
rect 26550 18164 26584 18740
rect 27568 18164 27602 18740
rect 28586 18164 28620 18740
rect 29604 18164 29638 18740
rect 30622 18164 30656 18740
rect 31640 18164 31674 18740
rect 32658 18164 32692 18740
rect 33676 18164 33710 18740
rect 34694 18164 34728 18740
rect 35712 18164 35746 18740
rect 36730 18164 36764 18740
rect 37748 18164 37782 18740
rect 38766 18164 38800 18740
rect 39784 18164 39818 18740
rect 19210 17252 19244 17828
rect 20228 17252 20262 17828
rect 21246 17252 21280 17828
rect 22264 17252 22298 17828
rect 23282 17252 23316 17828
rect 24514 16908 24548 17484
rect 25532 16908 25566 17484
rect 26550 16908 26584 17484
rect 27568 16908 27602 17484
rect 28586 16908 28620 17484
rect 29604 16908 29638 17484
rect 30622 16908 30656 17484
rect 31640 16908 31674 17484
rect 32658 16908 32692 17484
rect 33676 16908 33710 17484
rect 34694 16908 34728 17484
rect 35712 16908 35746 17484
rect 36730 16908 36764 17484
rect 37748 16908 37782 17484
rect 38766 16908 38800 17484
rect 39784 16908 39818 17484
rect 19210 16220 19244 16796
rect 20228 16220 20262 16796
rect 21246 16220 21280 16796
rect 22264 16220 22298 16796
rect 23282 16220 23316 16796
rect 24514 15652 24548 16228
rect 25532 15652 25566 16228
rect 26550 15652 26584 16228
rect 27568 15652 27602 16228
rect 28586 15652 28620 16228
rect 29604 15652 29638 16228
rect 30622 15652 30656 16228
rect 31640 15652 31674 16228
rect 32658 15652 32692 16228
rect 33676 15652 33710 16228
rect 34694 15652 34728 16228
rect 35712 15652 35746 16228
rect 36730 15652 36764 16228
rect 37748 15652 37782 16228
rect 38766 15652 38800 16228
rect 39784 15652 39818 16228
<< psubdiff >>
rect 4718 13802 4880 13902
rect 41800 13802 41962 13902
rect 4718 13740 4818 13802
rect -202 842 -40 942
rect 4240 842 4402 942
rect -202 780 -102 842
rect 4302 780 4402 842
rect -202 -1942 -102 -1880
rect 4302 -1942 4402 -1880
rect -202 -2042 -40 -1942
rect 4240 -2042 4402 -1942
rect 41862 13740 41962 13802
rect 20126 13296 20208 13320
rect 20126 13262 20150 13296
rect 20184 13262 20208 13296
rect 20126 13238 20208 13262
rect 21144 13296 21226 13320
rect 21144 13262 21168 13296
rect 21202 13262 21226 13296
rect 21144 13238 21226 13262
rect 22162 13296 22244 13320
rect 22162 13262 22186 13296
rect 22220 13262 22244 13296
rect 22162 13238 22244 13262
rect 23180 13296 23262 13320
rect 23180 13262 23204 13296
rect 23238 13262 23262 13296
rect 23180 13238 23262 13262
rect 24198 13296 24280 13320
rect 24198 13262 24222 13296
rect 24256 13262 24280 13296
rect 24198 13238 24280 13262
rect 25216 13296 25298 13320
rect 25216 13262 25240 13296
rect 25274 13262 25298 13296
rect 25216 13238 25298 13262
rect 26234 13296 26316 13320
rect 26234 13262 26258 13296
rect 26292 13262 26316 13296
rect 26234 13238 26316 13262
rect 27252 13296 27334 13320
rect 27252 13262 27276 13296
rect 27310 13262 27334 13296
rect 27252 13238 27334 13262
rect 28270 13296 28352 13320
rect 28270 13262 28294 13296
rect 28328 13262 28352 13296
rect 28270 13238 28352 13262
rect 29288 13296 29370 13320
rect 29288 13262 29312 13296
rect 29346 13262 29370 13296
rect 29288 13238 29370 13262
rect 30306 13296 30388 13320
rect 30306 13262 30330 13296
rect 30364 13262 30388 13296
rect 30306 13238 30388 13262
rect 31324 13296 31406 13320
rect 31324 13262 31348 13296
rect 31382 13262 31406 13296
rect 31324 13238 31406 13262
rect 32342 13296 32424 13320
rect 32342 13262 32366 13296
rect 32400 13262 32424 13296
rect 32342 13238 32424 13262
rect 33360 13296 33442 13320
rect 33360 13262 33384 13296
rect 33418 13262 33442 13296
rect 33360 13238 33442 13262
rect 34378 13296 34460 13320
rect 34378 13262 34402 13296
rect 34436 13262 34460 13296
rect 34378 13238 34460 13262
rect 35396 13296 35478 13320
rect 35396 13262 35420 13296
rect 35454 13262 35478 13296
rect 35396 13238 35478 13262
rect 36414 13296 36496 13320
rect 36414 13262 36438 13296
rect 36472 13262 36496 13296
rect 36414 13238 36496 13262
rect 37432 13296 37514 13320
rect 37432 13262 37456 13296
rect 37490 13262 37514 13296
rect 37432 13238 37514 13262
rect 38450 13296 38532 13320
rect 38450 13262 38474 13296
rect 38508 13262 38532 13296
rect 38450 13238 38532 13262
rect 39468 13296 39550 13320
rect 39468 13262 39492 13296
rect 39526 13262 39550 13296
rect 39468 13238 39550 13262
rect 7832 12694 7914 12718
rect 7832 12660 7856 12694
rect 7890 12660 7914 12694
rect 7832 12636 7914 12660
rect 8850 12694 8932 12718
rect 8850 12660 8874 12694
rect 8908 12660 8932 12694
rect 8850 12636 8932 12660
rect 9868 12694 9950 12718
rect 9868 12660 9892 12694
rect 9926 12660 9950 12694
rect 9868 12636 9950 12660
rect 10886 12694 10968 12718
rect 10886 12660 10910 12694
rect 10944 12660 10968 12694
rect 10886 12636 10968 12660
rect 11904 12694 11986 12718
rect 11904 12660 11928 12694
rect 11962 12660 11986 12694
rect 11904 12636 11986 12660
rect 12922 12694 13004 12718
rect 12922 12660 12946 12694
rect 12980 12660 13004 12694
rect 12922 12636 13004 12660
rect 13940 12694 14022 12718
rect 13940 12660 13964 12694
rect 13998 12660 14022 12694
rect 13940 12636 14022 12660
rect 14958 12694 15040 12718
rect 14958 12660 14982 12694
rect 15016 12660 15040 12694
rect 14958 12636 15040 12660
rect 15976 12694 16058 12718
rect 15976 12660 16000 12694
rect 16034 12660 16058 12694
rect 15976 12636 16058 12660
rect 17004 12694 17086 12718
rect 17004 12660 17028 12694
rect 17062 12660 17086 12694
rect 17004 12636 17086 12660
rect 7832 11876 7914 11900
rect 7832 11842 7856 11876
rect 7890 11842 7914 11876
rect 7832 11818 7914 11842
rect 8850 11876 8932 11900
rect 8850 11842 8874 11876
rect 8908 11842 8932 11876
rect 8850 11818 8932 11842
rect 9868 11876 9950 11900
rect 9868 11842 9892 11876
rect 9926 11842 9950 11876
rect 9868 11818 9950 11842
rect 10886 11876 10968 11900
rect 10886 11842 10910 11876
rect 10944 11842 10968 11876
rect 10886 11818 10968 11842
rect 11904 11876 11986 11900
rect 11904 11842 11928 11876
rect 11962 11842 11986 11876
rect 11904 11818 11986 11842
rect 12922 11876 13004 11900
rect 12922 11842 12946 11876
rect 12980 11842 13004 11876
rect 12922 11818 13004 11842
rect 13940 11876 14022 11900
rect 13940 11842 13964 11876
rect 13998 11842 14022 11876
rect 13940 11818 14022 11842
rect 14958 11876 15040 11900
rect 14958 11842 14982 11876
rect 15016 11842 15040 11876
rect 14958 11818 15040 11842
rect 15976 11876 16058 11900
rect 15976 11842 16000 11876
rect 16034 11842 16058 11876
rect 15976 11818 16058 11842
rect 17004 11876 17086 11900
rect 17004 11842 17028 11876
rect 17062 11842 17086 11876
rect 17004 11818 17086 11842
rect 20138 11270 20220 11294
rect 20138 11236 20162 11270
rect 20196 11236 20220 11270
rect 20138 11212 20220 11236
rect 21156 11270 21238 11294
rect 21156 11236 21180 11270
rect 21214 11236 21238 11270
rect 21156 11212 21238 11236
rect 22174 11270 22256 11294
rect 22174 11236 22198 11270
rect 22232 11236 22256 11270
rect 22174 11212 22256 11236
rect 23192 11270 23274 11294
rect 23192 11236 23216 11270
rect 23250 11236 23274 11270
rect 23192 11212 23274 11236
rect 24210 11270 24292 11294
rect 24210 11236 24234 11270
rect 24268 11236 24292 11270
rect 24210 11212 24292 11236
rect 25228 11270 25310 11294
rect 25228 11236 25252 11270
rect 25286 11236 25310 11270
rect 25228 11212 25310 11236
rect 26246 11270 26328 11294
rect 26246 11236 26270 11270
rect 26304 11236 26328 11270
rect 26246 11212 26328 11236
rect 27264 11270 27346 11294
rect 27264 11236 27288 11270
rect 27322 11236 27346 11270
rect 27264 11212 27346 11236
rect 28282 11270 28364 11294
rect 28282 11236 28306 11270
rect 28340 11236 28364 11270
rect 28282 11212 28364 11236
rect 29300 11270 29382 11294
rect 29300 11236 29324 11270
rect 29358 11236 29382 11270
rect 29300 11212 29382 11236
rect 30318 11270 30400 11294
rect 30318 11236 30342 11270
rect 30376 11236 30400 11270
rect 30318 11212 30400 11236
rect 31336 11270 31418 11294
rect 31336 11236 31360 11270
rect 31394 11236 31418 11270
rect 31336 11212 31418 11236
rect 32354 11270 32436 11294
rect 32354 11236 32378 11270
rect 32412 11236 32436 11270
rect 32354 11212 32436 11236
rect 33372 11270 33454 11294
rect 33372 11236 33396 11270
rect 33430 11236 33454 11270
rect 33372 11212 33454 11236
rect 34390 11270 34472 11294
rect 34390 11236 34414 11270
rect 34448 11236 34472 11270
rect 34390 11212 34472 11236
rect 35408 11270 35490 11294
rect 35408 11236 35432 11270
rect 35466 11236 35490 11270
rect 35408 11212 35490 11236
rect 36426 11270 36508 11294
rect 36426 11236 36450 11270
rect 36484 11236 36508 11270
rect 36426 11212 36508 11236
rect 37444 11270 37526 11294
rect 37444 11236 37468 11270
rect 37502 11236 37526 11270
rect 37444 11212 37526 11236
rect 38462 11270 38544 11294
rect 38462 11236 38486 11270
rect 38520 11236 38544 11270
rect 38462 11212 38544 11236
rect 39480 11270 39562 11294
rect 39480 11236 39504 11270
rect 39538 11236 39562 11270
rect 39480 11212 39562 11236
rect 7832 11058 7914 11082
rect 7832 11024 7856 11058
rect 7890 11024 7914 11058
rect 7832 11000 7914 11024
rect 8850 11058 8932 11082
rect 8850 11024 8874 11058
rect 8908 11024 8932 11058
rect 8850 11000 8932 11024
rect 9868 11058 9950 11082
rect 9868 11024 9892 11058
rect 9926 11024 9950 11058
rect 9868 11000 9950 11024
rect 10886 11058 10968 11082
rect 10886 11024 10910 11058
rect 10944 11024 10968 11058
rect 10886 11000 10968 11024
rect 11904 11058 11986 11082
rect 11904 11024 11928 11058
rect 11962 11024 11986 11058
rect 11904 11000 11986 11024
rect 12922 11058 13004 11082
rect 12922 11024 12946 11058
rect 12980 11024 13004 11058
rect 12922 11000 13004 11024
rect 13940 11058 14022 11082
rect 13940 11024 13964 11058
rect 13998 11024 14022 11058
rect 13940 11000 14022 11024
rect 14958 11058 15040 11082
rect 14958 11024 14982 11058
rect 15016 11024 15040 11058
rect 14958 11000 15040 11024
rect 15976 11058 16058 11082
rect 15976 11024 16000 11058
rect 16034 11024 16058 11058
rect 15976 11000 16058 11024
rect 17004 11058 17086 11082
rect 17004 11024 17028 11058
rect 17062 11024 17086 11058
rect 17004 11000 17086 11024
rect 7832 10240 7914 10264
rect 7832 10206 7856 10240
rect 7890 10206 7914 10240
rect 7832 10182 7914 10206
rect 8850 10240 8932 10264
rect 8850 10206 8874 10240
rect 8908 10206 8932 10240
rect 8850 10182 8932 10206
rect 9868 10240 9950 10264
rect 9868 10206 9892 10240
rect 9926 10206 9950 10240
rect 9868 10182 9950 10206
rect 10886 10240 10968 10264
rect 10886 10206 10910 10240
rect 10944 10206 10968 10240
rect 10886 10182 10968 10206
rect 11904 10240 11986 10264
rect 11904 10206 11928 10240
rect 11962 10206 11986 10240
rect 11904 10182 11986 10206
rect 12922 10240 13004 10264
rect 12922 10206 12946 10240
rect 12980 10206 13004 10240
rect 12922 10182 13004 10206
rect 13940 10240 14022 10264
rect 13940 10206 13964 10240
rect 13998 10206 14022 10240
rect 13940 10182 14022 10206
rect 14958 10240 15040 10264
rect 14958 10206 14982 10240
rect 15016 10206 15040 10240
rect 14958 10182 15040 10206
rect 15976 10240 16058 10264
rect 15976 10206 16000 10240
rect 16034 10206 16058 10240
rect 15976 10182 16058 10206
rect 17004 10240 17086 10264
rect 17004 10206 17028 10240
rect 17062 10206 17086 10240
rect 17004 10182 17086 10206
rect 20126 9964 20208 9988
rect 20126 9930 20150 9964
rect 20184 9930 20208 9964
rect 20126 9906 20208 9930
rect 21144 9964 21226 9988
rect 21144 9930 21168 9964
rect 21202 9930 21226 9964
rect 21144 9906 21226 9930
rect 22162 9964 22244 9988
rect 22162 9930 22186 9964
rect 22220 9930 22244 9964
rect 22162 9906 22244 9930
rect 23180 9964 23262 9988
rect 23180 9930 23204 9964
rect 23238 9930 23262 9964
rect 23180 9906 23262 9930
rect 24198 9964 24280 9988
rect 24198 9930 24222 9964
rect 24256 9930 24280 9964
rect 24198 9906 24280 9930
rect 25216 9964 25298 9988
rect 25216 9930 25240 9964
rect 25274 9930 25298 9964
rect 25216 9906 25298 9930
rect 26234 9964 26316 9988
rect 26234 9930 26258 9964
rect 26292 9930 26316 9964
rect 26234 9906 26316 9930
rect 27252 9964 27334 9988
rect 27252 9930 27276 9964
rect 27310 9930 27334 9964
rect 27252 9906 27334 9930
rect 28270 9964 28352 9988
rect 28270 9930 28294 9964
rect 28328 9930 28352 9964
rect 28270 9906 28352 9930
rect 29288 9964 29370 9988
rect 29288 9930 29312 9964
rect 29346 9930 29370 9964
rect 29288 9906 29370 9930
rect 30306 9964 30388 9988
rect 30306 9930 30330 9964
rect 30364 9930 30388 9964
rect 30306 9906 30388 9930
rect 31324 9964 31406 9988
rect 31324 9930 31348 9964
rect 31382 9930 31406 9964
rect 31324 9906 31406 9930
rect 32342 9964 32424 9988
rect 32342 9930 32366 9964
rect 32400 9930 32424 9964
rect 32342 9906 32424 9930
rect 33360 9964 33442 9988
rect 33360 9930 33384 9964
rect 33418 9930 33442 9964
rect 33360 9906 33442 9930
rect 34378 9964 34460 9988
rect 34378 9930 34402 9964
rect 34436 9930 34460 9964
rect 34378 9906 34460 9930
rect 35396 9964 35478 9988
rect 35396 9930 35420 9964
rect 35454 9930 35478 9964
rect 35396 9906 35478 9930
rect 36414 9964 36496 9988
rect 36414 9930 36438 9964
rect 36472 9930 36496 9964
rect 36414 9906 36496 9930
rect 37432 9964 37514 9988
rect 37432 9930 37456 9964
rect 37490 9930 37514 9964
rect 37432 9906 37514 9930
rect 38450 9964 38532 9988
rect 38450 9930 38474 9964
rect 38508 9930 38532 9964
rect 38450 9906 38532 9930
rect 39468 9964 39550 9988
rect 39468 9930 39492 9964
rect 39526 9930 39550 9964
rect 39468 9906 39550 9930
rect 7832 9422 7914 9446
rect 7832 9388 7856 9422
rect 7890 9388 7914 9422
rect 7832 9364 7914 9388
rect 8850 9422 8932 9446
rect 8850 9388 8874 9422
rect 8908 9388 8932 9422
rect 8850 9364 8932 9388
rect 9868 9422 9950 9446
rect 9868 9388 9892 9422
rect 9926 9388 9950 9422
rect 9868 9364 9950 9388
rect 10886 9422 10968 9446
rect 10886 9388 10910 9422
rect 10944 9388 10968 9422
rect 10886 9364 10968 9388
rect 11904 9422 11986 9446
rect 11904 9388 11928 9422
rect 11962 9388 11986 9422
rect 11904 9364 11986 9388
rect 12922 9422 13004 9446
rect 12922 9388 12946 9422
rect 12980 9388 13004 9422
rect 12922 9364 13004 9388
rect 13940 9422 14022 9446
rect 13940 9388 13964 9422
rect 13998 9388 14022 9422
rect 13940 9364 14022 9388
rect 14958 9422 15040 9446
rect 14958 9388 14982 9422
rect 15016 9388 15040 9422
rect 14958 9364 15040 9388
rect 15976 9422 16058 9446
rect 15976 9388 16000 9422
rect 16034 9388 16058 9422
rect 15976 9364 16058 9388
rect 17004 9422 17086 9446
rect 17004 9388 17028 9422
rect 17062 9388 17086 9422
rect 17004 9364 17086 9388
rect 20114 8728 20196 8752
rect 7832 8604 7914 8628
rect 7832 8570 7856 8604
rect 7890 8570 7914 8604
rect 7832 8546 7914 8570
rect 8850 8604 8932 8628
rect 8850 8570 8874 8604
rect 8908 8570 8932 8604
rect 8850 8546 8932 8570
rect 9868 8604 9950 8628
rect 9868 8570 9892 8604
rect 9926 8570 9950 8604
rect 9868 8546 9950 8570
rect 10886 8604 10968 8628
rect 10886 8570 10910 8604
rect 10944 8570 10968 8604
rect 10886 8546 10968 8570
rect 11904 8604 11986 8628
rect 11904 8570 11928 8604
rect 11962 8570 11986 8604
rect 11904 8546 11986 8570
rect 12922 8604 13004 8628
rect 12922 8570 12946 8604
rect 12980 8570 13004 8604
rect 12922 8546 13004 8570
rect 13940 8604 14022 8628
rect 13940 8570 13964 8604
rect 13998 8570 14022 8604
rect 13940 8546 14022 8570
rect 14958 8604 15040 8628
rect 20114 8694 20138 8728
rect 20172 8694 20196 8728
rect 20114 8670 20196 8694
rect 21132 8728 21214 8752
rect 21132 8694 21156 8728
rect 21190 8694 21214 8728
rect 21132 8670 21214 8694
rect 22150 8728 22232 8752
rect 22150 8694 22174 8728
rect 22208 8694 22232 8728
rect 22150 8670 22232 8694
rect 23168 8728 23250 8752
rect 23168 8694 23192 8728
rect 23226 8694 23250 8728
rect 23168 8670 23250 8694
rect 24186 8728 24268 8752
rect 24186 8694 24210 8728
rect 24244 8694 24268 8728
rect 24186 8670 24268 8694
rect 25204 8728 25286 8752
rect 25204 8694 25228 8728
rect 25262 8694 25286 8728
rect 25204 8670 25286 8694
rect 26222 8728 26304 8752
rect 26222 8694 26246 8728
rect 26280 8694 26304 8728
rect 26222 8670 26304 8694
rect 27240 8728 27322 8752
rect 27240 8694 27264 8728
rect 27298 8694 27322 8728
rect 27240 8670 27322 8694
rect 28258 8728 28340 8752
rect 28258 8694 28282 8728
rect 28316 8694 28340 8728
rect 28258 8670 28340 8694
rect 29276 8728 29358 8752
rect 29276 8694 29300 8728
rect 29334 8694 29358 8728
rect 29276 8670 29358 8694
rect 30294 8728 30376 8752
rect 30294 8694 30318 8728
rect 30352 8694 30376 8728
rect 30294 8670 30376 8694
rect 31312 8728 31394 8752
rect 31312 8694 31336 8728
rect 31370 8694 31394 8728
rect 31312 8670 31394 8694
rect 32330 8728 32412 8752
rect 32330 8694 32354 8728
rect 32388 8694 32412 8728
rect 32330 8670 32412 8694
rect 33348 8728 33430 8752
rect 33348 8694 33372 8728
rect 33406 8694 33430 8728
rect 33348 8670 33430 8694
rect 34366 8728 34448 8752
rect 34366 8694 34390 8728
rect 34424 8694 34448 8728
rect 34366 8670 34448 8694
rect 35384 8728 35466 8752
rect 35384 8694 35408 8728
rect 35442 8694 35466 8728
rect 35384 8670 35466 8694
rect 36402 8728 36484 8752
rect 36402 8694 36426 8728
rect 36460 8694 36484 8728
rect 36402 8670 36484 8694
rect 37420 8728 37502 8752
rect 37420 8694 37444 8728
rect 37478 8694 37502 8728
rect 37420 8670 37502 8694
rect 38438 8728 38520 8752
rect 38438 8694 38462 8728
rect 38496 8694 38520 8728
rect 38438 8670 38520 8694
rect 39456 8728 39538 8752
rect 39456 8694 39480 8728
rect 39514 8694 39538 8728
rect 39456 8670 39538 8694
rect 14958 8570 14982 8604
rect 15016 8570 15040 8604
rect 14958 8546 15040 8570
rect 15976 8604 16058 8628
rect 15976 8570 16000 8604
rect 16034 8570 16058 8604
rect 15976 8546 16058 8570
rect 17004 8604 17086 8628
rect 17004 8570 17028 8604
rect 17062 8570 17086 8604
rect 17004 8546 17086 8570
rect 7832 7786 7914 7810
rect 7832 7752 7856 7786
rect 7890 7752 7914 7786
rect 7832 7728 7914 7752
rect 8850 7786 8932 7810
rect 8850 7752 8874 7786
rect 8908 7752 8932 7786
rect 8850 7728 8932 7752
rect 9868 7786 9950 7810
rect 9868 7752 9892 7786
rect 9926 7752 9950 7786
rect 9868 7728 9950 7752
rect 10886 7786 10968 7810
rect 10886 7752 10910 7786
rect 10944 7752 10968 7786
rect 10886 7728 10968 7752
rect 11904 7786 11986 7810
rect 11904 7752 11928 7786
rect 11962 7752 11986 7786
rect 11904 7728 11986 7752
rect 12922 7786 13004 7810
rect 12922 7752 12946 7786
rect 12980 7752 13004 7786
rect 12922 7728 13004 7752
rect 13940 7786 14022 7810
rect 13940 7752 13964 7786
rect 13998 7752 14022 7786
rect 13940 7728 14022 7752
rect 14958 7786 15040 7810
rect 14958 7752 14982 7786
rect 15016 7752 15040 7786
rect 14958 7728 15040 7752
rect 15976 7786 16058 7810
rect 15976 7752 16000 7786
rect 16034 7752 16058 7786
rect 15976 7728 16058 7752
rect 17004 7786 17086 7810
rect 17004 7752 17028 7786
rect 17062 7752 17086 7786
rect 17004 7728 17086 7752
rect 20114 7504 20196 7528
rect 20114 7470 20138 7504
rect 20172 7470 20196 7504
rect 20114 7446 20196 7470
rect 21132 7504 21214 7528
rect 21132 7470 21156 7504
rect 21190 7470 21214 7504
rect 21132 7446 21214 7470
rect 22150 7504 22232 7528
rect 22150 7470 22174 7504
rect 22208 7470 22232 7504
rect 22150 7446 22232 7470
rect 23168 7504 23250 7528
rect 23168 7470 23192 7504
rect 23226 7470 23250 7504
rect 23168 7446 23250 7470
rect 24186 7504 24268 7528
rect 24186 7470 24210 7504
rect 24244 7470 24268 7504
rect 24186 7446 24268 7470
rect 25204 7504 25286 7528
rect 25204 7470 25228 7504
rect 25262 7470 25286 7504
rect 25204 7446 25286 7470
rect 26222 7504 26304 7528
rect 26222 7470 26246 7504
rect 26280 7470 26304 7504
rect 26222 7446 26304 7470
rect 27240 7504 27322 7528
rect 27240 7470 27264 7504
rect 27298 7470 27322 7504
rect 27240 7446 27322 7470
rect 28258 7504 28340 7528
rect 28258 7470 28282 7504
rect 28316 7470 28340 7504
rect 28258 7446 28340 7470
rect 29276 7504 29358 7528
rect 29276 7470 29300 7504
rect 29334 7470 29358 7504
rect 29276 7446 29358 7470
rect 30294 7504 30376 7528
rect 30294 7470 30318 7504
rect 30352 7470 30376 7504
rect 30294 7446 30376 7470
rect 31312 7504 31394 7528
rect 31312 7470 31336 7504
rect 31370 7470 31394 7504
rect 31312 7446 31394 7470
rect 32330 7504 32412 7528
rect 32330 7470 32354 7504
rect 32388 7470 32412 7504
rect 32330 7446 32412 7470
rect 33348 7504 33430 7528
rect 33348 7470 33372 7504
rect 33406 7470 33430 7504
rect 33348 7446 33430 7470
rect 34366 7504 34448 7528
rect 34366 7470 34390 7504
rect 34424 7470 34448 7504
rect 34366 7446 34448 7470
rect 35384 7504 35466 7528
rect 35384 7470 35408 7504
rect 35442 7470 35466 7504
rect 35384 7446 35466 7470
rect 36402 7504 36484 7528
rect 36402 7470 36426 7504
rect 36460 7470 36484 7504
rect 36402 7446 36484 7470
rect 37420 7504 37502 7528
rect 37420 7470 37444 7504
rect 37478 7470 37502 7504
rect 37420 7446 37502 7470
rect 38438 7504 38520 7528
rect 38438 7470 38462 7504
rect 38496 7470 38520 7504
rect 38438 7446 38520 7470
rect 39456 7504 39538 7528
rect 39456 7470 39480 7504
rect 39514 7470 39538 7504
rect 39456 7446 39538 7470
rect 7832 6968 7914 6992
rect 7832 6934 7856 6968
rect 7890 6934 7914 6968
rect 7832 6910 7914 6934
rect 8850 6968 8932 6992
rect 8850 6934 8874 6968
rect 8908 6934 8932 6968
rect 8850 6910 8932 6934
rect 9868 6968 9950 6992
rect 9868 6934 9892 6968
rect 9926 6934 9950 6968
rect 9868 6910 9950 6934
rect 10886 6968 10968 6992
rect 10886 6934 10910 6968
rect 10944 6934 10968 6968
rect 10886 6910 10968 6934
rect 11904 6968 11986 6992
rect 11904 6934 11928 6968
rect 11962 6934 11986 6968
rect 11904 6910 11986 6934
rect 12922 6968 13004 6992
rect 12922 6934 12946 6968
rect 12980 6934 13004 6968
rect 12922 6910 13004 6934
rect 13940 6968 14022 6992
rect 13940 6934 13964 6968
rect 13998 6934 14022 6968
rect 13940 6910 14022 6934
rect 14958 6968 15040 6992
rect 14958 6934 14982 6968
rect 15016 6934 15040 6968
rect 14958 6910 15040 6934
rect 15976 6968 16058 6992
rect 15976 6934 16000 6968
rect 16034 6934 16058 6968
rect 15976 6910 16058 6934
rect 17004 6968 17086 6992
rect 17004 6934 17028 6968
rect 17062 6934 17086 6968
rect 17004 6910 17086 6934
rect 20126 6268 20208 6292
rect 20126 6234 20150 6268
rect 20184 6234 20208 6268
rect 20126 6210 20208 6234
rect 21144 6268 21226 6292
rect 21144 6234 21168 6268
rect 21202 6234 21226 6268
rect 21144 6210 21226 6234
rect 22162 6268 22244 6292
rect 22162 6234 22186 6268
rect 22220 6234 22244 6268
rect 22162 6210 22244 6234
rect 23180 6268 23262 6292
rect 23180 6234 23204 6268
rect 23238 6234 23262 6268
rect 23180 6210 23262 6234
rect 24198 6268 24280 6292
rect 24198 6234 24222 6268
rect 24256 6234 24280 6268
rect 24198 6210 24280 6234
rect 25216 6268 25298 6292
rect 25216 6234 25240 6268
rect 25274 6234 25298 6268
rect 25216 6210 25298 6234
rect 26234 6268 26316 6292
rect 26234 6234 26258 6268
rect 26292 6234 26316 6268
rect 26234 6210 26316 6234
rect 27252 6268 27334 6292
rect 27252 6234 27276 6268
rect 27310 6234 27334 6268
rect 27252 6210 27334 6234
rect 28270 6268 28352 6292
rect 28270 6234 28294 6268
rect 28328 6234 28352 6268
rect 28270 6210 28352 6234
rect 29288 6268 29370 6292
rect 29288 6234 29312 6268
rect 29346 6234 29370 6268
rect 29288 6210 29370 6234
rect 30306 6268 30388 6292
rect 30306 6234 30330 6268
rect 30364 6234 30388 6268
rect 30306 6210 30388 6234
rect 31324 6268 31406 6292
rect 31324 6234 31348 6268
rect 31382 6234 31406 6268
rect 31324 6210 31406 6234
rect 32342 6268 32424 6292
rect 32342 6234 32366 6268
rect 32400 6234 32424 6268
rect 32342 6210 32424 6234
rect 33360 6268 33442 6292
rect 33360 6234 33384 6268
rect 33418 6234 33442 6268
rect 33360 6210 33442 6234
rect 34378 6268 34460 6292
rect 34378 6234 34402 6268
rect 34436 6234 34460 6268
rect 34378 6210 34460 6234
rect 35396 6268 35478 6292
rect 35396 6234 35420 6268
rect 35454 6234 35478 6268
rect 35396 6210 35478 6234
rect 36414 6268 36496 6292
rect 36414 6234 36438 6268
rect 36472 6234 36496 6268
rect 36414 6210 36496 6234
rect 37432 6268 37514 6292
rect 37432 6234 37456 6268
rect 37490 6234 37514 6268
rect 37432 6210 37514 6234
rect 38450 6268 38532 6292
rect 38450 6234 38474 6268
rect 38508 6234 38532 6268
rect 38450 6210 38532 6234
rect 39468 6268 39550 6292
rect 39468 6234 39492 6268
rect 39526 6234 39550 6268
rect 39468 6210 39550 6234
rect 7820 6074 7902 6098
rect 7820 6040 7844 6074
rect 7878 6040 7902 6074
rect 7820 6016 7902 6040
rect 8838 6074 8920 6098
rect 8838 6040 8862 6074
rect 8896 6040 8920 6074
rect 8838 6016 8920 6040
rect 9856 6074 9938 6098
rect 9856 6040 9880 6074
rect 9914 6040 9938 6074
rect 9856 6016 9938 6040
rect 10874 6074 10956 6098
rect 10874 6040 10898 6074
rect 10932 6040 10956 6074
rect 10874 6016 10956 6040
rect 11892 6074 11974 6098
rect 11892 6040 11916 6074
rect 11950 6040 11974 6074
rect 11892 6016 11974 6040
rect 12910 6074 12992 6098
rect 12910 6040 12934 6074
rect 12968 6040 12992 6074
rect 12910 6016 12992 6040
rect 13928 6074 14010 6098
rect 13928 6040 13952 6074
rect 13986 6040 14010 6074
rect 13928 6016 14010 6040
rect 14946 6074 15028 6098
rect 14946 6040 14970 6074
rect 15004 6040 15028 6074
rect 14946 6016 15028 6040
rect 15964 6074 16046 6098
rect 15964 6040 15988 6074
rect 16022 6040 16046 6074
rect 15964 6016 16046 6040
rect 16992 6074 17074 6098
rect 16992 6040 17016 6074
rect 17050 6040 17074 6074
rect 16992 6016 17074 6040
rect 7024 5126 7106 5150
rect 7024 5092 7048 5126
rect 7082 5092 7106 5126
rect 7024 5068 7106 5092
rect 8042 5126 8124 5150
rect 8042 5092 8066 5126
rect 8100 5092 8124 5126
rect 8042 5068 8124 5092
rect 9060 5126 9142 5150
rect 9060 5092 9084 5126
rect 9118 5092 9142 5126
rect 9060 5068 9142 5092
rect 10078 5126 10160 5150
rect 10078 5092 10102 5126
rect 10136 5092 10160 5126
rect 10078 5068 10160 5092
rect 11096 5126 11178 5150
rect 11096 5092 11120 5126
rect 11154 5092 11178 5126
rect 11096 5068 11178 5092
rect 12114 5126 12196 5150
rect 12114 5092 12138 5126
rect 12172 5092 12196 5126
rect 12114 5068 12196 5092
rect 13132 5126 13214 5150
rect 13132 5092 13156 5126
rect 13190 5092 13214 5126
rect 13132 5068 13214 5092
rect 14150 5126 14232 5150
rect 14150 5092 14174 5126
rect 14208 5092 14232 5126
rect 14150 5068 14232 5092
rect 15168 5126 15250 5150
rect 15168 5092 15192 5126
rect 15226 5092 15250 5126
rect 15168 5068 15250 5092
rect 16186 5126 16268 5150
rect 16186 5092 16210 5126
rect 16244 5092 16268 5126
rect 16186 5068 16268 5092
rect 17204 5126 17286 5150
rect 17204 5092 17228 5126
rect 17262 5092 17286 5126
rect 17204 5068 17286 5092
rect 20126 5020 20208 5044
rect 20126 4986 20150 5020
rect 20184 4986 20208 5020
rect 20126 4962 20208 4986
rect 21144 5020 21226 5044
rect 21144 4986 21168 5020
rect 21202 4986 21226 5020
rect 21144 4962 21226 4986
rect 22162 5020 22244 5044
rect 22162 4986 22186 5020
rect 22220 4986 22244 5020
rect 22162 4962 22244 4986
rect 23180 5020 23262 5044
rect 23180 4986 23204 5020
rect 23238 4986 23262 5020
rect 23180 4962 23262 4986
rect 24198 5020 24280 5044
rect 24198 4986 24222 5020
rect 24256 4986 24280 5020
rect 24198 4962 24280 4986
rect 25216 5020 25298 5044
rect 25216 4986 25240 5020
rect 25274 4986 25298 5020
rect 25216 4962 25298 4986
rect 26234 5020 26316 5044
rect 26234 4986 26258 5020
rect 26292 4986 26316 5020
rect 26234 4962 26316 4986
rect 27252 5020 27334 5044
rect 27252 4986 27276 5020
rect 27310 4986 27334 5020
rect 27252 4962 27334 4986
rect 28270 5020 28352 5044
rect 28270 4986 28294 5020
rect 28328 4986 28352 5020
rect 28270 4962 28352 4986
rect 29288 5020 29370 5044
rect 29288 4986 29312 5020
rect 29346 4986 29370 5020
rect 29288 4962 29370 4986
rect 30306 5020 30388 5044
rect 30306 4986 30330 5020
rect 30364 4986 30388 5020
rect 30306 4962 30388 4986
rect 31324 5020 31406 5044
rect 31324 4986 31348 5020
rect 31382 4986 31406 5020
rect 31324 4962 31406 4986
rect 32342 5020 32424 5044
rect 32342 4986 32366 5020
rect 32400 4986 32424 5020
rect 32342 4962 32424 4986
rect 33360 5020 33442 5044
rect 33360 4986 33384 5020
rect 33418 4986 33442 5020
rect 33360 4962 33442 4986
rect 34378 5020 34460 5044
rect 34378 4986 34402 5020
rect 34436 4986 34460 5020
rect 34378 4962 34460 4986
rect 35396 5020 35478 5044
rect 35396 4986 35420 5020
rect 35454 4986 35478 5020
rect 35396 4962 35478 4986
rect 36414 5020 36496 5044
rect 36414 4986 36438 5020
rect 36472 4986 36496 5020
rect 36414 4962 36496 4986
rect 37432 5020 37514 5044
rect 37432 4986 37456 5020
rect 37490 4986 37514 5020
rect 37432 4962 37514 4986
rect 38450 5020 38532 5044
rect 38450 4986 38474 5020
rect 38508 4986 38532 5020
rect 38450 4962 38532 4986
rect 39468 5020 39550 5044
rect 39468 4986 39492 5020
rect 39526 4986 39550 5020
rect 39468 4962 39550 4986
rect 7036 3984 7118 4008
rect 7036 3950 7060 3984
rect 7094 3950 7118 3984
rect 7036 3926 7118 3950
rect 8054 3984 8136 4008
rect 8054 3950 8078 3984
rect 8112 3950 8136 3984
rect 8054 3926 8136 3950
rect 9072 3984 9154 4008
rect 9072 3950 9096 3984
rect 9130 3950 9154 3984
rect 9072 3926 9154 3950
rect 10090 3984 10172 4008
rect 10090 3950 10114 3984
rect 10148 3950 10172 3984
rect 10090 3926 10172 3950
rect 11108 3984 11190 4008
rect 11108 3950 11132 3984
rect 11166 3950 11190 3984
rect 11108 3926 11190 3950
rect 12126 3984 12208 4008
rect 12126 3950 12150 3984
rect 12184 3950 12208 3984
rect 12126 3926 12208 3950
rect 13144 3984 13226 4008
rect 13144 3950 13168 3984
rect 13202 3950 13226 3984
rect 13144 3926 13226 3950
rect 14162 3984 14244 4008
rect 14162 3950 14186 3984
rect 14220 3950 14244 3984
rect 14162 3926 14244 3950
rect 15180 3984 15262 4008
rect 15180 3950 15204 3984
rect 15238 3950 15262 3984
rect 15180 3926 15262 3950
rect 16198 3984 16280 4008
rect 16198 3950 16222 3984
rect 16256 3950 16280 3984
rect 16198 3926 16280 3950
rect 17216 3984 17298 4008
rect 17216 3950 17240 3984
rect 17274 3950 17298 3984
rect 17216 3926 17298 3950
rect 20102 3784 20184 3808
rect 20102 3750 20126 3784
rect 20160 3750 20184 3784
rect 20102 3726 20184 3750
rect 21120 3784 21202 3808
rect 21120 3750 21144 3784
rect 21178 3750 21202 3784
rect 21120 3726 21202 3750
rect 22138 3784 22220 3808
rect 22138 3750 22162 3784
rect 22196 3750 22220 3784
rect 22138 3726 22220 3750
rect 23156 3784 23238 3808
rect 23156 3750 23180 3784
rect 23214 3750 23238 3784
rect 23156 3726 23238 3750
rect 24174 3784 24256 3808
rect 24174 3750 24198 3784
rect 24232 3750 24256 3784
rect 24174 3726 24256 3750
rect 25192 3784 25274 3808
rect 25192 3750 25216 3784
rect 25250 3750 25274 3784
rect 25192 3726 25274 3750
rect 26210 3784 26292 3808
rect 26210 3750 26234 3784
rect 26268 3750 26292 3784
rect 26210 3726 26292 3750
rect 27228 3784 27310 3808
rect 27228 3750 27252 3784
rect 27286 3750 27310 3784
rect 27228 3726 27310 3750
rect 28246 3784 28328 3808
rect 28246 3750 28270 3784
rect 28304 3750 28328 3784
rect 28246 3726 28328 3750
rect 29264 3784 29346 3808
rect 29264 3750 29288 3784
rect 29322 3750 29346 3784
rect 29264 3726 29346 3750
rect 30282 3784 30364 3808
rect 30282 3750 30306 3784
rect 30340 3750 30364 3784
rect 30282 3726 30364 3750
rect 31300 3784 31382 3808
rect 31300 3750 31324 3784
rect 31358 3750 31382 3784
rect 31300 3726 31382 3750
rect 32318 3784 32400 3808
rect 32318 3750 32342 3784
rect 32376 3750 32400 3784
rect 32318 3726 32400 3750
rect 33336 3784 33418 3808
rect 33336 3750 33360 3784
rect 33394 3750 33418 3784
rect 33336 3726 33418 3750
rect 34354 3784 34436 3808
rect 34354 3750 34378 3784
rect 34412 3750 34436 3784
rect 34354 3726 34436 3750
rect 35372 3784 35454 3808
rect 35372 3750 35396 3784
rect 35430 3750 35454 3784
rect 35372 3726 35454 3750
rect 36390 3784 36472 3808
rect 36390 3750 36414 3784
rect 36448 3750 36472 3784
rect 36390 3726 36472 3750
rect 37408 3784 37490 3808
rect 37408 3750 37432 3784
rect 37466 3750 37490 3784
rect 37408 3726 37490 3750
rect 38426 3784 38508 3808
rect 38426 3750 38450 3784
rect 38484 3750 38508 3784
rect 38426 3726 38508 3750
rect 39444 3784 39526 3808
rect 39444 3750 39468 3784
rect 39502 3750 39526 3784
rect 39444 3726 39526 3750
rect 7014 2876 7096 2900
rect 7014 2842 7038 2876
rect 7072 2842 7096 2876
rect 7014 2818 7096 2842
rect 8032 2876 8114 2900
rect 8032 2842 8056 2876
rect 8090 2842 8114 2876
rect 8032 2818 8114 2842
rect 9050 2876 9132 2900
rect 9050 2842 9074 2876
rect 9108 2842 9132 2876
rect 9050 2818 9132 2842
rect 10068 2876 10150 2900
rect 10068 2842 10092 2876
rect 10126 2842 10150 2876
rect 10068 2818 10150 2842
rect 11086 2876 11168 2900
rect 11086 2842 11110 2876
rect 11144 2842 11168 2876
rect 11086 2818 11168 2842
rect 12104 2876 12186 2900
rect 12104 2842 12128 2876
rect 12162 2842 12186 2876
rect 12104 2818 12186 2842
rect 13122 2876 13204 2900
rect 13122 2842 13146 2876
rect 13180 2842 13204 2876
rect 13122 2818 13204 2842
rect 14140 2876 14222 2900
rect 14140 2842 14164 2876
rect 14198 2842 14222 2876
rect 14140 2818 14222 2842
rect 15158 2876 15240 2900
rect 15158 2842 15182 2876
rect 15216 2842 15240 2876
rect 15158 2818 15240 2842
rect 16176 2876 16258 2900
rect 16176 2842 16200 2876
rect 16234 2842 16258 2876
rect 16176 2818 16258 2842
rect 17194 2876 17276 2900
rect 17194 2842 17218 2876
rect 17252 2842 17276 2876
rect 17194 2818 17276 2842
rect 20114 2560 20196 2584
rect 20114 2526 20138 2560
rect 20172 2526 20196 2560
rect 20114 2502 20196 2526
rect 21132 2560 21214 2584
rect 21132 2526 21156 2560
rect 21190 2526 21214 2560
rect 21132 2502 21214 2526
rect 22150 2560 22232 2584
rect 22150 2526 22174 2560
rect 22208 2526 22232 2560
rect 22150 2502 22232 2526
rect 23168 2560 23250 2584
rect 23168 2526 23192 2560
rect 23226 2526 23250 2560
rect 23168 2502 23250 2526
rect 24186 2560 24268 2584
rect 24186 2526 24210 2560
rect 24244 2526 24268 2560
rect 24186 2502 24268 2526
rect 25204 2560 25286 2584
rect 25204 2526 25228 2560
rect 25262 2526 25286 2560
rect 25204 2502 25286 2526
rect 26222 2560 26304 2584
rect 26222 2526 26246 2560
rect 26280 2526 26304 2560
rect 26222 2502 26304 2526
rect 27240 2560 27322 2584
rect 27240 2526 27264 2560
rect 27298 2526 27322 2560
rect 27240 2502 27322 2526
rect 28258 2560 28340 2584
rect 28258 2526 28282 2560
rect 28316 2526 28340 2560
rect 28258 2502 28340 2526
rect 29276 2560 29358 2584
rect 29276 2526 29300 2560
rect 29334 2526 29358 2560
rect 29276 2502 29358 2526
rect 30294 2560 30376 2584
rect 30294 2526 30318 2560
rect 30352 2526 30376 2560
rect 30294 2502 30376 2526
rect 31312 2560 31394 2584
rect 31312 2526 31336 2560
rect 31370 2526 31394 2560
rect 31312 2502 31394 2526
rect 32330 2560 32412 2584
rect 32330 2526 32354 2560
rect 32388 2526 32412 2560
rect 32330 2502 32412 2526
rect 33348 2560 33430 2584
rect 33348 2526 33372 2560
rect 33406 2526 33430 2560
rect 33348 2502 33430 2526
rect 34366 2560 34448 2584
rect 34366 2526 34390 2560
rect 34424 2526 34448 2560
rect 34366 2502 34448 2526
rect 35384 2560 35466 2584
rect 35384 2526 35408 2560
rect 35442 2526 35466 2560
rect 35384 2502 35466 2526
rect 36402 2560 36484 2584
rect 36402 2526 36426 2560
rect 36460 2526 36484 2560
rect 36402 2502 36484 2526
rect 37420 2560 37502 2584
rect 37420 2526 37444 2560
rect 37478 2526 37502 2560
rect 37420 2502 37502 2526
rect 38438 2560 38520 2584
rect 38438 2526 38462 2560
rect 38496 2526 38520 2560
rect 38438 2502 38520 2526
rect 39456 2560 39538 2584
rect 39456 2526 39480 2560
rect 39514 2526 39538 2560
rect 39456 2502 39538 2526
rect 7014 1770 7096 1794
rect 7014 1736 7038 1770
rect 7072 1736 7096 1770
rect 7014 1712 7096 1736
rect 8032 1770 8114 1794
rect 8032 1736 8056 1770
rect 8090 1736 8114 1770
rect 8032 1712 8114 1736
rect 9050 1770 9132 1794
rect 9050 1736 9074 1770
rect 9108 1736 9132 1770
rect 9050 1712 9132 1736
rect 10068 1770 10150 1794
rect 10068 1736 10092 1770
rect 10126 1736 10150 1770
rect 10068 1712 10150 1736
rect 11086 1770 11168 1794
rect 11086 1736 11110 1770
rect 11144 1736 11168 1770
rect 11086 1712 11168 1736
rect 12104 1770 12186 1794
rect 12104 1736 12128 1770
rect 12162 1736 12186 1770
rect 12104 1712 12186 1736
rect 13122 1770 13204 1794
rect 13122 1736 13146 1770
rect 13180 1736 13204 1770
rect 13122 1712 13204 1736
rect 14140 1770 14222 1794
rect 14140 1736 14164 1770
rect 14198 1736 14222 1770
rect 14140 1712 14222 1736
rect 15158 1770 15240 1794
rect 15158 1736 15182 1770
rect 15216 1736 15240 1770
rect 15158 1712 15240 1736
rect 16176 1770 16258 1794
rect 16176 1736 16200 1770
rect 16234 1736 16258 1770
rect 16176 1712 16258 1736
rect 17194 1770 17276 1794
rect 17194 1736 17218 1770
rect 17252 1736 17276 1770
rect 17194 1712 17276 1736
rect 20114 1324 20196 1348
rect 20114 1290 20138 1324
rect 20172 1290 20196 1324
rect 20114 1266 20196 1290
rect 21132 1324 21214 1348
rect 21132 1290 21156 1324
rect 21190 1290 21214 1324
rect 21132 1266 21214 1290
rect 22150 1324 22232 1348
rect 22150 1290 22174 1324
rect 22208 1290 22232 1324
rect 22150 1266 22232 1290
rect 23168 1324 23250 1348
rect 23168 1290 23192 1324
rect 23226 1290 23250 1324
rect 23168 1266 23250 1290
rect 24186 1324 24268 1348
rect 24186 1290 24210 1324
rect 24244 1290 24268 1324
rect 24186 1266 24268 1290
rect 25204 1324 25286 1348
rect 25204 1290 25228 1324
rect 25262 1290 25286 1324
rect 25204 1266 25286 1290
rect 26222 1324 26304 1348
rect 26222 1290 26246 1324
rect 26280 1290 26304 1324
rect 26222 1266 26304 1290
rect 27240 1324 27322 1348
rect 27240 1290 27264 1324
rect 27298 1290 27322 1324
rect 27240 1266 27322 1290
rect 28258 1324 28340 1348
rect 28258 1290 28282 1324
rect 28316 1290 28340 1324
rect 28258 1266 28340 1290
rect 29276 1324 29358 1348
rect 29276 1290 29300 1324
rect 29334 1290 29358 1324
rect 29276 1266 29358 1290
rect 30294 1324 30376 1348
rect 30294 1290 30318 1324
rect 30352 1290 30376 1324
rect 30294 1266 30376 1290
rect 31312 1324 31394 1348
rect 31312 1290 31336 1324
rect 31370 1290 31394 1324
rect 31312 1266 31394 1290
rect 32330 1324 32412 1348
rect 32330 1290 32354 1324
rect 32388 1290 32412 1324
rect 32330 1266 32412 1290
rect 33348 1324 33430 1348
rect 33348 1290 33372 1324
rect 33406 1290 33430 1324
rect 33348 1266 33430 1290
rect 34366 1324 34448 1348
rect 34366 1290 34390 1324
rect 34424 1290 34448 1324
rect 34366 1266 34448 1290
rect 35384 1324 35466 1348
rect 35384 1290 35408 1324
rect 35442 1290 35466 1324
rect 35384 1266 35466 1290
rect 36402 1324 36484 1348
rect 36402 1290 36426 1324
rect 36460 1290 36484 1324
rect 36402 1266 36484 1290
rect 37420 1324 37502 1348
rect 37420 1290 37444 1324
rect 37478 1290 37502 1324
rect 37420 1266 37502 1290
rect 38438 1324 38520 1348
rect 38438 1290 38462 1324
rect 38496 1290 38520 1324
rect 38438 1266 38520 1290
rect 39456 1324 39538 1348
rect 39456 1290 39480 1324
rect 39514 1290 39538 1324
rect 39456 1266 39538 1290
rect 7014 428 7096 452
rect 7014 394 7038 428
rect 7072 394 7096 428
rect 7014 370 7096 394
rect 8032 428 8114 452
rect 8032 394 8056 428
rect 8090 394 8114 428
rect 8032 370 8114 394
rect 9050 428 9132 452
rect 9050 394 9074 428
rect 9108 394 9132 428
rect 9050 370 9132 394
rect 10068 428 10150 452
rect 10068 394 10092 428
rect 10126 394 10150 428
rect 10068 370 10150 394
rect 11086 428 11168 452
rect 11086 394 11110 428
rect 11144 394 11168 428
rect 11086 370 11168 394
rect 12104 428 12186 452
rect 12104 394 12128 428
rect 12162 394 12186 428
rect 12104 370 12186 394
rect 13122 428 13204 452
rect 13122 394 13146 428
rect 13180 394 13204 428
rect 13122 370 13204 394
rect 14140 428 14222 452
rect 14140 394 14164 428
rect 14198 394 14222 428
rect 14140 370 14222 394
rect 15158 428 15240 452
rect 15158 394 15182 428
rect 15216 394 15240 428
rect 15158 370 15240 394
rect 16176 428 16258 452
rect 16176 394 16200 428
rect 16234 394 16258 428
rect 16176 370 16258 394
rect 17194 428 17276 452
rect 17194 394 17218 428
rect 17252 394 17276 428
rect 17194 370 17276 394
rect 20126 78 20208 102
rect 20126 44 20150 78
rect 20184 44 20208 78
rect 20126 20 20208 44
rect 21144 78 21226 102
rect 21144 44 21168 78
rect 21202 44 21226 78
rect 21144 20 21226 44
rect 22162 78 22244 102
rect 22162 44 22186 78
rect 22220 44 22244 78
rect 22162 20 22244 44
rect 23180 78 23262 102
rect 23180 44 23204 78
rect 23238 44 23262 78
rect 23180 20 23262 44
rect 24198 78 24280 102
rect 24198 44 24222 78
rect 24256 44 24280 78
rect 24198 20 24280 44
rect 25216 78 25298 102
rect 25216 44 25240 78
rect 25274 44 25298 78
rect 25216 20 25298 44
rect 26234 78 26316 102
rect 26234 44 26258 78
rect 26292 44 26316 78
rect 26234 20 26316 44
rect 27252 78 27334 102
rect 27252 44 27276 78
rect 27310 44 27334 78
rect 27252 20 27334 44
rect 28270 78 28352 102
rect 28270 44 28294 78
rect 28328 44 28352 78
rect 28270 20 28352 44
rect 29288 78 29370 102
rect 29288 44 29312 78
rect 29346 44 29370 78
rect 29288 20 29370 44
rect 30306 78 30388 102
rect 30306 44 30330 78
rect 30364 44 30388 78
rect 30306 20 30388 44
rect 31324 78 31406 102
rect 31324 44 31348 78
rect 31382 44 31406 78
rect 31324 20 31406 44
rect 32342 78 32424 102
rect 32342 44 32366 78
rect 32400 44 32424 78
rect 32342 20 32424 44
rect 33360 78 33442 102
rect 33360 44 33384 78
rect 33418 44 33442 78
rect 33360 20 33442 44
rect 34378 78 34460 102
rect 34378 44 34402 78
rect 34436 44 34460 78
rect 34378 20 34460 44
rect 35396 78 35478 102
rect 35396 44 35420 78
rect 35454 44 35478 78
rect 35396 20 35478 44
rect 36414 78 36496 102
rect 36414 44 36438 78
rect 36472 44 36496 78
rect 36414 20 36496 44
rect 37432 78 37514 102
rect 37432 44 37456 78
rect 37490 44 37514 78
rect 37432 20 37514 44
rect 38450 78 38532 102
rect 38450 44 38474 78
rect 38508 44 38532 78
rect 38450 20 38532 44
rect 39468 78 39550 102
rect 39468 44 39492 78
rect 39526 44 39550 78
rect 39468 20 39550 44
rect 6824 -1018 6906 -994
rect 6824 -1052 6848 -1018
rect 6882 -1052 6906 -1018
rect 6824 -1076 6906 -1052
rect 7842 -1018 7924 -994
rect 7842 -1052 7866 -1018
rect 7900 -1052 7924 -1018
rect 7842 -1076 7924 -1052
rect 8860 -1018 8942 -994
rect 8860 -1052 8884 -1018
rect 8918 -1052 8942 -1018
rect 8860 -1076 8942 -1052
rect 9878 -1018 9960 -994
rect 9878 -1052 9902 -1018
rect 9936 -1052 9960 -1018
rect 9878 -1076 9960 -1052
rect 10896 -1018 10978 -994
rect 10896 -1052 10920 -1018
rect 10954 -1052 10978 -1018
rect 10896 -1076 10978 -1052
rect 11914 -1018 11996 -994
rect 11914 -1052 11938 -1018
rect 11972 -1052 11996 -1018
rect 11914 -1076 11996 -1052
rect 12932 -1018 13014 -994
rect 12932 -1052 12956 -1018
rect 12990 -1052 13014 -1018
rect 12932 -1076 13014 -1052
rect 13950 -1018 14032 -994
rect 13950 -1052 13974 -1018
rect 14008 -1052 14032 -1018
rect 13950 -1076 14032 -1052
rect 14968 -1018 15050 -994
rect 14968 -1052 14992 -1018
rect 15026 -1052 15050 -1018
rect 14968 -1076 15050 -1052
rect 15986 -1018 16068 -994
rect 15986 -1052 16010 -1018
rect 16044 -1052 16068 -1018
rect 15986 -1076 16068 -1052
rect 17004 -1018 17086 -994
rect 17004 -1052 17028 -1018
rect 17062 -1052 17086 -1018
rect 17004 -1076 17086 -1052
rect 20114 -1100 20196 -1076
rect 20114 -1134 20138 -1100
rect 20172 -1134 20196 -1100
rect 20114 -1158 20196 -1134
rect 21132 -1100 21214 -1076
rect 21132 -1134 21156 -1100
rect 21190 -1134 21214 -1100
rect 21132 -1158 21214 -1134
rect 22150 -1100 22232 -1076
rect 22150 -1134 22174 -1100
rect 22208 -1134 22232 -1100
rect 22150 -1158 22232 -1134
rect 23168 -1100 23250 -1076
rect 23168 -1134 23192 -1100
rect 23226 -1134 23250 -1100
rect 23168 -1158 23250 -1134
rect 24186 -1100 24268 -1076
rect 24186 -1134 24210 -1100
rect 24244 -1134 24268 -1100
rect 24186 -1158 24268 -1134
rect 25204 -1100 25286 -1076
rect 25204 -1134 25228 -1100
rect 25262 -1134 25286 -1100
rect 25204 -1158 25286 -1134
rect 26222 -1100 26304 -1076
rect 26222 -1134 26246 -1100
rect 26280 -1134 26304 -1100
rect 26222 -1158 26304 -1134
rect 27240 -1100 27322 -1076
rect 27240 -1134 27264 -1100
rect 27298 -1134 27322 -1100
rect 27240 -1158 27322 -1134
rect 28258 -1100 28340 -1076
rect 28258 -1134 28282 -1100
rect 28316 -1134 28340 -1100
rect 28258 -1158 28340 -1134
rect 29276 -1100 29358 -1076
rect 29276 -1134 29300 -1100
rect 29334 -1134 29358 -1100
rect 29276 -1158 29358 -1134
rect 30294 -1100 30376 -1076
rect 30294 -1134 30318 -1100
rect 30352 -1134 30376 -1100
rect 30294 -1158 30376 -1134
rect 31312 -1100 31394 -1076
rect 31312 -1134 31336 -1100
rect 31370 -1134 31394 -1100
rect 31312 -1158 31394 -1134
rect 32330 -1100 32412 -1076
rect 32330 -1134 32354 -1100
rect 32388 -1134 32412 -1100
rect 32330 -1158 32412 -1134
rect 33348 -1100 33430 -1076
rect 33348 -1134 33372 -1100
rect 33406 -1134 33430 -1100
rect 33348 -1158 33430 -1134
rect 34366 -1100 34448 -1076
rect 34366 -1134 34390 -1100
rect 34424 -1134 34448 -1100
rect 34366 -1158 34448 -1134
rect 35384 -1100 35466 -1076
rect 35384 -1134 35408 -1100
rect 35442 -1134 35466 -1100
rect 35384 -1158 35466 -1134
rect 36402 -1100 36484 -1076
rect 36402 -1134 36426 -1100
rect 36460 -1134 36484 -1100
rect 36402 -1158 36484 -1134
rect 37420 -1100 37502 -1076
rect 37420 -1134 37444 -1100
rect 37478 -1134 37502 -1100
rect 37420 -1158 37502 -1134
rect 38438 -1100 38520 -1076
rect 38438 -1134 38462 -1100
rect 38496 -1134 38520 -1100
rect 38438 -1158 38520 -1134
rect 39456 -1100 39538 -1076
rect 39456 -1134 39480 -1100
rect 39514 -1134 39538 -1100
rect 39456 -1158 39538 -1134
rect 4718 -2042 4818 -1980
rect 41862 -2042 41962 -1980
rect 4718 -2142 4880 -2042
rect 41800 -2142 41962 -2042
<< nsubdiff >>
rect 17418 29302 17580 29402
rect 41700 29302 41862 29402
rect 17418 29240 17518 29302
rect 41762 29240 41862 29302
rect 24012 26858 24094 26884
rect 24012 26824 24036 26858
rect 24070 26824 24094 26858
rect 24012 26800 24094 26824
rect 25030 26858 25112 26884
rect 25030 26824 25054 26858
rect 25088 26824 25112 26858
rect 25030 26800 25112 26824
rect 26048 26858 26130 26884
rect 26048 26824 26072 26858
rect 26106 26824 26130 26858
rect 26048 26800 26130 26824
rect 27066 26858 27148 26884
rect 27066 26824 27090 26858
rect 27124 26824 27148 26858
rect 27066 26800 27148 26824
rect 28084 26858 28166 26884
rect 28084 26824 28108 26858
rect 28142 26824 28166 26858
rect 28084 26800 28166 26824
rect 29102 26858 29184 26884
rect 29102 26824 29126 26858
rect 29160 26824 29184 26858
rect 29102 26800 29184 26824
rect 30120 26858 30202 26884
rect 30120 26824 30144 26858
rect 30178 26824 30202 26858
rect 30120 26800 30202 26824
rect 31138 26858 31220 26884
rect 31138 26824 31162 26858
rect 31196 26824 31220 26858
rect 31138 26800 31220 26824
rect 32156 26858 32238 26884
rect 32156 26824 32180 26858
rect 32214 26824 32238 26858
rect 32156 26800 32238 26824
rect 33174 26858 33256 26884
rect 33174 26824 33198 26858
rect 33232 26824 33256 26858
rect 33174 26800 33256 26824
rect 34192 26858 34274 26884
rect 34192 26824 34216 26858
rect 34250 26824 34274 26858
rect 34192 26800 34274 26824
rect 35210 26858 35292 26884
rect 35210 26824 35234 26858
rect 35268 26824 35292 26858
rect 35210 26800 35292 26824
rect 36228 26858 36310 26884
rect 36228 26824 36252 26858
rect 36286 26824 36310 26858
rect 36228 26800 36310 26824
rect 37246 26858 37328 26884
rect 37246 26824 37270 26858
rect 37304 26824 37328 26858
rect 37246 26800 37328 26824
rect 38264 26858 38346 26884
rect 38264 26824 38288 26858
rect 38322 26824 38346 26858
rect 38264 26800 38346 26824
rect 39282 26858 39364 26884
rect 39282 26824 39306 26858
rect 39340 26824 39364 26858
rect 39282 26800 39364 26824
rect 24034 25704 24116 25730
rect 24034 25670 24058 25704
rect 24092 25670 24116 25704
rect 24034 25646 24116 25670
rect 25052 25704 25134 25730
rect 25052 25670 25076 25704
rect 25110 25670 25134 25704
rect 25052 25646 25134 25670
rect 26070 25704 26152 25730
rect 26070 25670 26094 25704
rect 26128 25670 26152 25704
rect 26070 25646 26152 25670
rect 27088 25704 27170 25730
rect 27088 25670 27112 25704
rect 27146 25670 27170 25704
rect 27088 25646 27170 25670
rect 28106 25704 28188 25730
rect 28106 25670 28130 25704
rect 28164 25670 28188 25704
rect 28106 25646 28188 25670
rect 29124 25704 29206 25730
rect 29124 25670 29148 25704
rect 29182 25670 29206 25704
rect 29124 25646 29206 25670
rect 30142 25704 30224 25730
rect 30142 25670 30166 25704
rect 30200 25670 30224 25704
rect 30142 25646 30224 25670
rect 31160 25704 31242 25730
rect 31160 25670 31184 25704
rect 31218 25670 31242 25704
rect 31160 25646 31242 25670
rect 32178 25704 32260 25730
rect 32178 25670 32202 25704
rect 32236 25670 32260 25704
rect 32178 25646 32260 25670
rect 33196 25704 33278 25730
rect 33196 25670 33220 25704
rect 33254 25670 33278 25704
rect 33196 25646 33278 25670
rect 34214 25704 34296 25730
rect 34214 25670 34238 25704
rect 34272 25670 34296 25704
rect 34214 25646 34296 25670
rect 35232 25704 35314 25730
rect 35232 25670 35256 25704
rect 35290 25670 35314 25704
rect 35232 25646 35314 25670
rect 36250 25704 36332 25730
rect 36250 25670 36274 25704
rect 36308 25670 36332 25704
rect 36250 25646 36332 25670
rect 37268 25704 37350 25730
rect 37268 25670 37292 25704
rect 37326 25670 37350 25704
rect 37268 25646 37350 25670
rect 38286 25704 38368 25730
rect 38286 25670 38310 25704
rect 38344 25670 38368 25704
rect 38286 25646 38368 25670
rect 39304 25704 39386 25730
rect 39304 25670 39328 25704
rect 39362 25670 39386 25704
rect 39304 25646 39386 25670
rect 24012 24572 24094 24598
rect 24012 24538 24036 24572
rect 24070 24538 24094 24572
rect 24012 24514 24094 24538
rect 25030 24572 25112 24598
rect 25030 24538 25054 24572
rect 25088 24538 25112 24572
rect 25030 24514 25112 24538
rect 26048 24572 26130 24598
rect 26048 24538 26072 24572
rect 26106 24538 26130 24572
rect 26048 24514 26130 24538
rect 27066 24572 27148 24598
rect 27066 24538 27090 24572
rect 27124 24538 27148 24572
rect 27066 24514 27148 24538
rect 28084 24572 28166 24598
rect 28084 24538 28108 24572
rect 28142 24538 28166 24572
rect 28084 24514 28166 24538
rect 29102 24572 29184 24598
rect 29102 24538 29126 24572
rect 29160 24538 29184 24572
rect 29102 24514 29184 24538
rect 30120 24572 30202 24598
rect 30120 24538 30144 24572
rect 30178 24538 30202 24572
rect 30120 24514 30202 24538
rect 31138 24572 31220 24598
rect 31138 24538 31162 24572
rect 31196 24538 31220 24572
rect 31138 24514 31220 24538
rect 32156 24572 32238 24598
rect 32156 24538 32180 24572
rect 32214 24538 32238 24572
rect 32156 24514 32238 24538
rect 33174 24572 33256 24598
rect 33174 24538 33198 24572
rect 33232 24538 33256 24572
rect 33174 24514 33256 24538
rect 34192 24572 34274 24598
rect 34192 24538 34216 24572
rect 34250 24538 34274 24572
rect 34192 24514 34274 24538
rect 35210 24572 35292 24598
rect 35210 24538 35234 24572
rect 35268 24538 35292 24572
rect 35210 24514 35292 24538
rect 36228 24572 36310 24598
rect 36228 24538 36252 24572
rect 36286 24538 36310 24572
rect 36228 24514 36310 24538
rect 37246 24572 37328 24598
rect 37246 24538 37270 24572
rect 37304 24538 37328 24572
rect 37246 24514 37328 24538
rect 38264 24572 38346 24598
rect 38264 24538 38288 24572
rect 38322 24538 38346 24572
rect 38264 24514 38346 24538
rect 39282 24572 39364 24598
rect 39282 24538 39306 24572
rect 39340 24538 39364 24572
rect 39282 24514 39364 24538
rect 24012 23190 24094 23216
rect 24012 23156 24036 23190
rect 24070 23156 24094 23190
rect 24012 23132 24094 23156
rect 25030 23190 25112 23216
rect 25030 23156 25054 23190
rect 25088 23156 25112 23190
rect 25030 23132 25112 23156
rect 26048 23190 26130 23216
rect 26048 23156 26072 23190
rect 26106 23156 26130 23190
rect 26048 23132 26130 23156
rect 27066 23190 27148 23216
rect 27066 23156 27090 23190
rect 27124 23156 27148 23190
rect 27066 23132 27148 23156
rect 28084 23190 28166 23216
rect 28084 23156 28108 23190
rect 28142 23156 28166 23190
rect 28084 23132 28166 23156
rect 29102 23190 29184 23216
rect 29102 23156 29126 23190
rect 29160 23156 29184 23190
rect 29102 23132 29184 23156
rect 30120 23190 30202 23216
rect 30120 23156 30144 23190
rect 30178 23156 30202 23190
rect 30120 23132 30202 23156
rect 31138 23190 31220 23216
rect 31138 23156 31162 23190
rect 31196 23156 31220 23190
rect 31138 23132 31220 23156
rect 32156 23190 32238 23216
rect 32156 23156 32180 23190
rect 32214 23156 32238 23190
rect 32156 23132 32238 23156
rect 33174 23190 33256 23216
rect 33174 23156 33198 23190
rect 33232 23156 33256 23190
rect 33174 23132 33256 23156
rect 34192 23190 34274 23216
rect 34192 23156 34216 23190
rect 34250 23156 34274 23190
rect 34192 23132 34274 23156
rect 35210 23190 35292 23216
rect 35210 23156 35234 23190
rect 35268 23156 35292 23190
rect 35210 23132 35292 23156
rect 36228 23190 36310 23216
rect 36228 23156 36252 23190
rect 36286 23156 36310 23190
rect 36228 23132 36310 23156
rect 37246 23190 37328 23216
rect 37246 23156 37270 23190
rect 37304 23156 37328 23190
rect 37246 23132 37328 23156
rect 38264 23190 38346 23216
rect 38264 23156 38288 23190
rect 38322 23156 38346 23190
rect 38264 23132 38346 23156
rect 39282 23190 39364 23216
rect 39282 23156 39306 23190
rect 39340 23156 39364 23190
rect 39282 23132 39364 23156
rect 24700 21842 24782 21868
rect 24700 21808 24724 21842
rect 24758 21808 24782 21842
rect 24700 21784 24782 21808
rect 25718 21842 25800 21868
rect 25718 21808 25742 21842
rect 25776 21808 25800 21842
rect 25718 21784 25800 21808
rect 26736 21842 26818 21868
rect 26736 21808 26760 21842
rect 26794 21808 26818 21842
rect 26736 21784 26818 21808
rect 27754 21842 27836 21868
rect 27754 21808 27778 21842
rect 27812 21808 27836 21842
rect 27754 21784 27836 21808
rect 28772 21842 28854 21868
rect 28772 21808 28796 21842
rect 28830 21808 28854 21842
rect 28772 21784 28854 21808
rect 29790 21842 29872 21868
rect 29790 21808 29814 21842
rect 29848 21808 29872 21842
rect 29790 21784 29872 21808
rect 30808 21842 30890 21868
rect 30808 21808 30832 21842
rect 30866 21808 30890 21842
rect 30808 21784 30890 21808
rect 31826 21842 31908 21868
rect 31826 21808 31850 21842
rect 31884 21808 31908 21842
rect 31826 21784 31908 21808
rect 32844 21842 32926 21868
rect 32844 21808 32868 21842
rect 32902 21808 32926 21842
rect 32844 21784 32926 21808
rect 33862 21842 33944 21868
rect 33862 21808 33886 21842
rect 33920 21808 33944 21842
rect 33862 21784 33944 21808
rect 34880 21842 34962 21868
rect 34880 21808 34904 21842
rect 34938 21808 34962 21842
rect 34880 21784 34962 21808
rect 35898 21842 35980 21868
rect 35898 21808 35922 21842
rect 35956 21808 35980 21842
rect 35898 21784 35980 21808
rect 36916 21842 36998 21868
rect 36916 21808 36940 21842
rect 36974 21808 36998 21842
rect 36916 21784 36998 21808
rect 37934 21842 38016 21868
rect 37934 21808 37958 21842
rect 37992 21808 38016 21842
rect 37934 21784 38016 21808
rect 38952 21842 39034 21868
rect 38952 21808 38976 21842
rect 39010 21808 39034 21842
rect 38952 21784 39034 21808
rect 24306 20564 24388 20590
rect 24306 20530 24330 20564
rect 24364 20530 24388 20564
rect 24306 20506 24388 20530
rect 25324 20564 25406 20590
rect 25324 20530 25348 20564
rect 25382 20530 25406 20564
rect 25324 20506 25406 20530
rect 26342 20564 26424 20590
rect 26342 20530 26366 20564
rect 26400 20530 26424 20564
rect 26342 20506 26424 20530
rect 27360 20564 27442 20590
rect 27360 20530 27384 20564
rect 27418 20530 27442 20564
rect 27360 20506 27442 20530
rect 28378 20564 28460 20590
rect 28378 20530 28402 20564
rect 28436 20530 28460 20564
rect 28378 20506 28460 20530
rect 29396 20564 29478 20590
rect 29396 20530 29420 20564
rect 29454 20530 29478 20564
rect 29396 20506 29478 20530
rect 30414 20564 30496 20590
rect 30414 20530 30438 20564
rect 30472 20530 30496 20564
rect 30414 20506 30496 20530
rect 31432 20564 31514 20590
rect 31432 20530 31456 20564
rect 31490 20530 31514 20564
rect 31432 20506 31514 20530
rect 32450 20564 32532 20590
rect 32450 20530 32474 20564
rect 32508 20530 32532 20564
rect 32450 20506 32532 20530
rect 33468 20564 33550 20590
rect 33468 20530 33492 20564
rect 33526 20530 33550 20564
rect 33468 20506 33550 20530
rect 34486 20564 34568 20590
rect 34486 20530 34510 20564
rect 34544 20530 34568 20564
rect 34486 20506 34568 20530
rect 35504 20564 35586 20590
rect 35504 20530 35528 20564
rect 35562 20530 35586 20564
rect 35504 20506 35586 20530
rect 36522 20564 36604 20590
rect 36522 20530 36546 20564
rect 36580 20530 36604 20564
rect 36522 20506 36604 20530
rect 37540 20564 37622 20590
rect 37540 20530 37564 20564
rect 37598 20530 37622 20564
rect 37540 20506 37622 20530
rect 38558 20564 38640 20590
rect 38558 20530 38582 20564
rect 38616 20530 38640 20564
rect 38558 20506 38640 20530
rect 39576 20564 39658 20590
rect 39576 20530 39600 20564
rect 39634 20530 39658 20564
rect 39576 20506 39658 20530
rect 19708 20254 19790 20280
rect 19708 20220 19732 20254
rect 19766 20220 19790 20254
rect 19708 20196 19790 20220
rect 20726 20254 20808 20280
rect 20726 20220 20750 20254
rect 20784 20220 20808 20254
rect 20726 20196 20808 20220
rect 21744 20254 21826 20280
rect 21744 20220 21768 20254
rect 21802 20220 21826 20254
rect 21744 20196 21826 20220
rect 22762 20254 22844 20280
rect 22762 20220 22786 20254
rect 22820 20220 22844 20254
rect 22762 20196 22844 20220
rect 19184 19100 19266 19126
rect 19184 19066 19208 19100
rect 19242 19066 19266 19100
rect 19184 19042 19266 19066
rect 20202 19100 20284 19126
rect 20202 19066 20226 19100
rect 20260 19066 20284 19100
rect 20202 19042 20284 19066
rect 21220 19100 21302 19126
rect 21220 19066 21244 19100
rect 21278 19066 21302 19100
rect 21220 19042 21302 19066
rect 22238 19100 22320 19126
rect 22238 19066 22262 19100
rect 22296 19066 22320 19100
rect 22238 19042 22320 19066
rect 24396 19116 24478 19142
rect 24396 19082 24420 19116
rect 24454 19082 24478 19116
rect 24396 19058 24478 19082
rect 25414 19116 25496 19142
rect 25414 19082 25438 19116
rect 25472 19082 25496 19116
rect 25414 19058 25496 19082
rect 26432 19116 26514 19142
rect 26432 19082 26456 19116
rect 26490 19082 26514 19116
rect 26432 19058 26514 19082
rect 27450 19116 27532 19142
rect 27450 19082 27474 19116
rect 27508 19082 27532 19116
rect 27450 19058 27532 19082
rect 28468 19116 28550 19142
rect 28468 19082 28492 19116
rect 28526 19082 28550 19116
rect 28468 19058 28550 19082
rect 29486 19116 29568 19142
rect 29486 19082 29510 19116
rect 29544 19082 29568 19116
rect 29486 19058 29568 19082
rect 30504 19116 30586 19142
rect 30504 19082 30528 19116
rect 30562 19082 30586 19116
rect 30504 19058 30586 19082
rect 31522 19116 31604 19142
rect 31522 19082 31546 19116
rect 31580 19082 31604 19116
rect 31522 19058 31604 19082
rect 32540 19116 32622 19142
rect 32540 19082 32564 19116
rect 32598 19082 32622 19116
rect 32540 19058 32622 19082
rect 33558 19116 33640 19142
rect 33558 19082 33582 19116
rect 33616 19082 33640 19116
rect 33558 19058 33640 19082
rect 34576 19116 34658 19142
rect 34576 19082 34600 19116
rect 34634 19082 34658 19116
rect 34576 19058 34658 19082
rect 35594 19116 35676 19142
rect 35594 19082 35618 19116
rect 35652 19082 35676 19116
rect 35594 19058 35676 19082
rect 36612 19116 36694 19142
rect 36612 19082 36636 19116
rect 36670 19082 36694 19116
rect 36612 19058 36694 19082
rect 37630 19116 37712 19142
rect 37630 19082 37654 19116
rect 37688 19082 37712 19116
rect 37630 19058 37712 19082
rect 38648 19116 38730 19142
rect 38648 19082 38672 19116
rect 38706 19082 38730 19116
rect 38648 19058 38730 19082
rect 39666 19116 39748 19142
rect 39666 19082 39690 19116
rect 39724 19082 39748 19116
rect 39666 19058 39748 19082
rect 19194 18072 19276 18098
rect 19194 18038 19218 18072
rect 19252 18038 19276 18072
rect 19194 18014 19276 18038
rect 20212 18072 20294 18098
rect 20212 18038 20236 18072
rect 20270 18038 20294 18072
rect 20212 18014 20294 18038
rect 21230 18072 21312 18098
rect 21230 18038 21254 18072
rect 21288 18038 21312 18072
rect 21230 18014 21312 18038
rect 22248 18072 22330 18098
rect 22248 18038 22272 18072
rect 22306 18038 22330 18072
rect 22248 18014 22330 18038
rect 24420 17848 24502 17874
rect 24420 17814 24444 17848
rect 24478 17814 24502 17848
rect 24420 17790 24502 17814
rect 25438 17848 25520 17874
rect 25438 17814 25462 17848
rect 25496 17814 25520 17848
rect 25438 17790 25520 17814
rect 26456 17848 26538 17874
rect 26456 17814 26480 17848
rect 26514 17814 26538 17848
rect 26456 17790 26538 17814
rect 27474 17848 27556 17874
rect 27474 17814 27498 17848
rect 27532 17814 27556 17848
rect 27474 17790 27556 17814
rect 28492 17848 28574 17874
rect 28492 17814 28516 17848
rect 28550 17814 28574 17848
rect 28492 17790 28574 17814
rect 29510 17848 29592 17874
rect 29510 17814 29534 17848
rect 29568 17814 29592 17848
rect 29510 17790 29592 17814
rect 30528 17848 30610 17874
rect 30528 17814 30552 17848
rect 30586 17814 30610 17848
rect 30528 17790 30610 17814
rect 31546 17848 31628 17874
rect 31546 17814 31570 17848
rect 31604 17814 31628 17848
rect 31546 17790 31628 17814
rect 32564 17848 32646 17874
rect 32564 17814 32588 17848
rect 32622 17814 32646 17848
rect 32564 17790 32646 17814
rect 33582 17848 33664 17874
rect 33582 17814 33606 17848
rect 33640 17814 33664 17848
rect 33582 17790 33664 17814
rect 34600 17848 34682 17874
rect 34600 17814 34624 17848
rect 34658 17814 34682 17848
rect 34600 17790 34682 17814
rect 35618 17848 35700 17874
rect 35618 17814 35642 17848
rect 35676 17814 35700 17848
rect 35618 17790 35700 17814
rect 36636 17848 36718 17874
rect 36636 17814 36660 17848
rect 36694 17814 36718 17848
rect 36636 17790 36718 17814
rect 37654 17848 37736 17874
rect 37654 17814 37678 17848
rect 37712 17814 37736 17848
rect 37654 17790 37736 17814
rect 38672 17848 38754 17874
rect 38672 17814 38696 17848
rect 38730 17814 38754 17848
rect 38672 17790 38754 17814
rect 39690 17848 39772 17874
rect 39690 17814 39714 17848
rect 39748 17814 39772 17848
rect 39690 17790 39772 17814
rect 19184 17044 19266 17070
rect 19184 17010 19208 17044
rect 19242 17010 19266 17044
rect 19184 16986 19266 17010
rect 20202 17044 20284 17070
rect 20202 17010 20226 17044
rect 20260 17010 20284 17044
rect 20202 16986 20284 17010
rect 21220 17044 21302 17070
rect 21220 17010 21244 17044
rect 21278 17010 21302 17044
rect 21220 16986 21302 17010
rect 22238 17044 22320 17070
rect 22238 17010 22262 17044
rect 22296 17010 22320 17044
rect 22238 16986 22320 17010
rect 24284 16604 24366 16630
rect 24284 16570 24308 16604
rect 24342 16570 24366 16604
rect 24284 16546 24366 16570
rect 25302 16604 25384 16630
rect 25302 16570 25326 16604
rect 25360 16570 25384 16604
rect 25302 16546 25384 16570
rect 26320 16604 26402 16630
rect 26320 16570 26344 16604
rect 26378 16570 26402 16604
rect 26320 16546 26402 16570
rect 27338 16604 27420 16630
rect 27338 16570 27362 16604
rect 27396 16570 27420 16604
rect 27338 16546 27420 16570
rect 28356 16604 28438 16630
rect 28356 16570 28380 16604
rect 28414 16570 28438 16604
rect 28356 16546 28438 16570
rect 29374 16604 29456 16630
rect 29374 16570 29398 16604
rect 29432 16570 29456 16604
rect 29374 16546 29456 16570
rect 30392 16604 30474 16630
rect 30392 16570 30416 16604
rect 30450 16570 30474 16604
rect 30392 16546 30474 16570
rect 31410 16604 31492 16630
rect 31410 16570 31434 16604
rect 31468 16570 31492 16604
rect 31410 16546 31492 16570
rect 32428 16604 32510 16630
rect 32428 16570 32452 16604
rect 32486 16570 32510 16604
rect 32428 16546 32510 16570
rect 33446 16604 33528 16630
rect 33446 16570 33470 16604
rect 33504 16570 33528 16604
rect 33446 16546 33528 16570
rect 34464 16604 34546 16630
rect 34464 16570 34488 16604
rect 34522 16570 34546 16604
rect 34464 16546 34546 16570
rect 35482 16604 35564 16630
rect 35482 16570 35506 16604
rect 35540 16570 35564 16604
rect 35482 16546 35564 16570
rect 36500 16604 36582 16630
rect 36500 16570 36524 16604
rect 36558 16570 36582 16604
rect 36500 16546 36582 16570
rect 37518 16604 37600 16630
rect 37518 16570 37542 16604
rect 37576 16570 37600 16604
rect 37518 16546 37600 16570
rect 38536 16604 38618 16630
rect 38536 16570 38560 16604
rect 38594 16570 38618 16604
rect 38536 16546 38618 16570
rect 39554 16604 39636 16630
rect 39554 16570 39578 16604
rect 39612 16570 39636 16604
rect 39554 16546 39636 16570
rect 19708 15892 19790 15918
rect 19708 15858 19732 15892
rect 19766 15858 19790 15892
rect 19708 15834 19790 15858
rect 20726 15892 20808 15918
rect 20726 15858 20750 15892
rect 20784 15858 20808 15892
rect 20726 15834 20808 15858
rect 21744 15892 21826 15918
rect 21744 15858 21768 15892
rect 21802 15858 21826 15892
rect 21744 15834 21826 15858
rect 22762 15892 22844 15918
rect 22762 15858 22786 15892
rect 22820 15858 22844 15892
rect 22762 15834 22844 15858
rect 17418 14832 17518 14894
rect 41762 14832 41862 14894
rect 17418 14732 17580 14832
rect 41700 14732 41862 14832
<< psubdiffcont >>
rect 4880 13802 41800 13902
rect -40 842 4240 942
rect -202 -1880 -102 780
rect 4302 -1880 4402 780
rect -40 -2042 4240 -1942
rect 4718 -1980 4818 13740
rect 20150 13262 20184 13296
rect 21168 13262 21202 13296
rect 22186 13262 22220 13296
rect 23204 13262 23238 13296
rect 24222 13262 24256 13296
rect 25240 13262 25274 13296
rect 26258 13262 26292 13296
rect 27276 13262 27310 13296
rect 28294 13262 28328 13296
rect 29312 13262 29346 13296
rect 30330 13262 30364 13296
rect 31348 13262 31382 13296
rect 32366 13262 32400 13296
rect 33384 13262 33418 13296
rect 34402 13262 34436 13296
rect 35420 13262 35454 13296
rect 36438 13262 36472 13296
rect 37456 13262 37490 13296
rect 38474 13262 38508 13296
rect 39492 13262 39526 13296
rect 7856 12660 7890 12694
rect 8874 12660 8908 12694
rect 9892 12660 9926 12694
rect 10910 12660 10944 12694
rect 11928 12660 11962 12694
rect 12946 12660 12980 12694
rect 13964 12660 13998 12694
rect 14982 12660 15016 12694
rect 16000 12660 16034 12694
rect 17028 12660 17062 12694
rect 7856 11842 7890 11876
rect 8874 11842 8908 11876
rect 9892 11842 9926 11876
rect 10910 11842 10944 11876
rect 11928 11842 11962 11876
rect 12946 11842 12980 11876
rect 13964 11842 13998 11876
rect 14982 11842 15016 11876
rect 16000 11842 16034 11876
rect 17028 11842 17062 11876
rect 20162 11236 20196 11270
rect 21180 11236 21214 11270
rect 22198 11236 22232 11270
rect 23216 11236 23250 11270
rect 24234 11236 24268 11270
rect 25252 11236 25286 11270
rect 26270 11236 26304 11270
rect 27288 11236 27322 11270
rect 28306 11236 28340 11270
rect 29324 11236 29358 11270
rect 30342 11236 30376 11270
rect 31360 11236 31394 11270
rect 32378 11236 32412 11270
rect 33396 11236 33430 11270
rect 34414 11236 34448 11270
rect 35432 11236 35466 11270
rect 36450 11236 36484 11270
rect 37468 11236 37502 11270
rect 38486 11236 38520 11270
rect 39504 11236 39538 11270
rect 7856 11024 7890 11058
rect 8874 11024 8908 11058
rect 9892 11024 9926 11058
rect 10910 11024 10944 11058
rect 11928 11024 11962 11058
rect 12946 11024 12980 11058
rect 13964 11024 13998 11058
rect 14982 11024 15016 11058
rect 16000 11024 16034 11058
rect 17028 11024 17062 11058
rect 7856 10206 7890 10240
rect 8874 10206 8908 10240
rect 9892 10206 9926 10240
rect 10910 10206 10944 10240
rect 11928 10206 11962 10240
rect 12946 10206 12980 10240
rect 13964 10206 13998 10240
rect 14982 10206 15016 10240
rect 16000 10206 16034 10240
rect 17028 10206 17062 10240
rect 20150 9930 20184 9964
rect 21168 9930 21202 9964
rect 22186 9930 22220 9964
rect 23204 9930 23238 9964
rect 24222 9930 24256 9964
rect 25240 9930 25274 9964
rect 26258 9930 26292 9964
rect 27276 9930 27310 9964
rect 28294 9930 28328 9964
rect 29312 9930 29346 9964
rect 30330 9930 30364 9964
rect 31348 9930 31382 9964
rect 32366 9930 32400 9964
rect 33384 9930 33418 9964
rect 34402 9930 34436 9964
rect 35420 9930 35454 9964
rect 36438 9930 36472 9964
rect 37456 9930 37490 9964
rect 38474 9930 38508 9964
rect 39492 9930 39526 9964
rect 7856 9388 7890 9422
rect 8874 9388 8908 9422
rect 9892 9388 9926 9422
rect 10910 9388 10944 9422
rect 11928 9388 11962 9422
rect 12946 9388 12980 9422
rect 13964 9388 13998 9422
rect 14982 9388 15016 9422
rect 16000 9388 16034 9422
rect 17028 9388 17062 9422
rect 7856 8570 7890 8604
rect 8874 8570 8908 8604
rect 9892 8570 9926 8604
rect 10910 8570 10944 8604
rect 11928 8570 11962 8604
rect 12946 8570 12980 8604
rect 13964 8570 13998 8604
rect 20138 8694 20172 8728
rect 21156 8694 21190 8728
rect 22174 8694 22208 8728
rect 23192 8694 23226 8728
rect 24210 8694 24244 8728
rect 25228 8694 25262 8728
rect 26246 8694 26280 8728
rect 27264 8694 27298 8728
rect 28282 8694 28316 8728
rect 29300 8694 29334 8728
rect 30318 8694 30352 8728
rect 31336 8694 31370 8728
rect 32354 8694 32388 8728
rect 33372 8694 33406 8728
rect 34390 8694 34424 8728
rect 35408 8694 35442 8728
rect 36426 8694 36460 8728
rect 37444 8694 37478 8728
rect 38462 8694 38496 8728
rect 39480 8694 39514 8728
rect 14982 8570 15016 8604
rect 16000 8570 16034 8604
rect 17028 8570 17062 8604
rect 7856 7752 7890 7786
rect 8874 7752 8908 7786
rect 9892 7752 9926 7786
rect 10910 7752 10944 7786
rect 11928 7752 11962 7786
rect 12946 7752 12980 7786
rect 13964 7752 13998 7786
rect 14982 7752 15016 7786
rect 16000 7752 16034 7786
rect 17028 7752 17062 7786
rect 20138 7470 20172 7504
rect 21156 7470 21190 7504
rect 22174 7470 22208 7504
rect 23192 7470 23226 7504
rect 24210 7470 24244 7504
rect 25228 7470 25262 7504
rect 26246 7470 26280 7504
rect 27264 7470 27298 7504
rect 28282 7470 28316 7504
rect 29300 7470 29334 7504
rect 30318 7470 30352 7504
rect 31336 7470 31370 7504
rect 32354 7470 32388 7504
rect 33372 7470 33406 7504
rect 34390 7470 34424 7504
rect 35408 7470 35442 7504
rect 36426 7470 36460 7504
rect 37444 7470 37478 7504
rect 38462 7470 38496 7504
rect 39480 7470 39514 7504
rect 7856 6934 7890 6968
rect 8874 6934 8908 6968
rect 9892 6934 9926 6968
rect 10910 6934 10944 6968
rect 11928 6934 11962 6968
rect 12946 6934 12980 6968
rect 13964 6934 13998 6968
rect 14982 6934 15016 6968
rect 16000 6934 16034 6968
rect 17028 6934 17062 6968
rect 20150 6234 20184 6268
rect 21168 6234 21202 6268
rect 22186 6234 22220 6268
rect 23204 6234 23238 6268
rect 24222 6234 24256 6268
rect 25240 6234 25274 6268
rect 26258 6234 26292 6268
rect 27276 6234 27310 6268
rect 28294 6234 28328 6268
rect 29312 6234 29346 6268
rect 30330 6234 30364 6268
rect 31348 6234 31382 6268
rect 32366 6234 32400 6268
rect 33384 6234 33418 6268
rect 34402 6234 34436 6268
rect 35420 6234 35454 6268
rect 36438 6234 36472 6268
rect 37456 6234 37490 6268
rect 38474 6234 38508 6268
rect 39492 6234 39526 6268
rect 7844 6040 7878 6074
rect 8862 6040 8896 6074
rect 9880 6040 9914 6074
rect 10898 6040 10932 6074
rect 11916 6040 11950 6074
rect 12934 6040 12968 6074
rect 13952 6040 13986 6074
rect 14970 6040 15004 6074
rect 15988 6040 16022 6074
rect 17016 6040 17050 6074
rect 7048 5092 7082 5126
rect 8066 5092 8100 5126
rect 9084 5092 9118 5126
rect 10102 5092 10136 5126
rect 11120 5092 11154 5126
rect 12138 5092 12172 5126
rect 13156 5092 13190 5126
rect 14174 5092 14208 5126
rect 15192 5092 15226 5126
rect 16210 5092 16244 5126
rect 17228 5092 17262 5126
rect 20150 4986 20184 5020
rect 21168 4986 21202 5020
rect 22186 4986 22220 5020
rect 23204 4986 23238 5020
rect 24222 4986 24256 5020
rect 25240 4986 25274 5020
rect 26258 4986 26292 5020
rect 27276 4986 27310 5020
rect 28294 4986 28328 5020
rect 29312 4986 29346 5020
rect 30330 4986 30364 5020
rect 31348 4986 31382 5020
rect 32366 4986 32400 5020
rect 33384 4986 33418 5020
rect 34402 4986 34436 5020
rect 35420 4986 35454 5020
rect 36438 4986 36472 5020
rect 37456 4986 37490 5020
rect 38474 4986 38508 5020
rect 39492 4986 39526 5020
rect 7060 3950 7094 3984
rect 8078 3950 8112 3984
rect 9096 3950 9130 3984
rect 10114 3950 10148 3984
rect 11132 3950 11166 3984
rect 12150 3950 12184 3984
rect 13168 3950 13202 3984
rect 14186 3950 14220 3984
rect 15204 3950 15238 3984
rect 16222 3950 16256 3984
rect 17240 3950 17274 3984
rect 20126 3750 20160 3784
rect 21144 3750 21178 3784
rect 22162 3750 22196 3784
rect 23180 3750 23214 3784
rect 24198 3750 24232 3784
rect 25216 3750 25250 3784
rect 26234 3750 26268 3784
rect 27252 3750 27286 3784
rect 28270 3750 28304 3784
rect 29288 3750 29322 3784
rect 30306 3750 30340 3784
rect 31324 3750 31358 3784
rect 32342 3750 32376 3784
rect 33360 3750 33394 3784
rect 34378 3750 34412 3784
rect 35396 3750 35430 3784
rect 36414 3750 36448 3784
rect 37432 3750 37466 3784
rect 38450 3750 38484 3784
rect 39468 3750 39502 3784
rect 7038 2842 7072 2876
rect 8056 2842 8090 2876
rect 9074 2842 9108 2876
rect 10092 2842 10126 2876
rect 11110 2842 11144 2876
rect 12128 2842 12162 2876
rect 13146 2842 13180 2876
rect 14164 2842 14198 2876
rect 15182 2842 15216 2876
rect 16200 2842 16234 2876
rect 17218 2842 17252 2876
rect 20138 2526 20172 2560
rect 21156 2526 21190 2560
rect 22174 2526 22208 2560
rect 23192 2526 23226 2560
rect 24210 2526 24244 2560
rect 25228 2526 25262 2560
rect 26246 2526 26280 2560
rect 27264 2526 27298 2560
rect 28282 2526 28316 2560
rect 29300 2526 29334 2560
rect 30318 2526 30352 2560
rect 31336 2526 31370 2560
rect 32354 2526 32388 2560
rect 33372 2526 33406 2560
rect 34390 2526 34424 2560
rect 35408 2526 35442 2560
rect 36426 2526 36460 2560
rect 37444 2526 37478 2560
rect 38462 2526 38496 2560
rect 39480 2526 39514 2560
rect 7038 1736 7072 1770
rect 8056 1736 8090 1770
rect 9074 1736 9108 1770
rect 10092 1736 10126 1770
rect 11110 1736 11144 1770
rect 12128 1736 12162 1770
rect 13146 1736 13180 1770
rect 14164 1736 14198 1770
rect 15182 1736 15216 1770
rect 16200 1736 16234 1770
rect 17218 1736 17252 1770
rect 20138 1290 20172 1324
rect 21156 1290 21190 1324
rect 22174 1290 22208 1324
rect 23192 1290 23226 1324
rect 24210 1290 24244 1324
rect 25228 1290 25262 1324
rect 26246 1290 26280 1324
rect 27264 1290 27298 1324
rect 28282 1290 28316 1324
rect 29300 1290 29334 1324
rect 30318 1290 30352 1324
rect 31336 1290 31370 1324
rect 32354 1290 32388 1324
rect 33372 1290 33406 1324
rect 34390 1290 34424 1324
rect 35408 1290 35442 1324
rect 36426 1290 36460 1324
rect 37444 1290 37478 1324
rect 38462 1290 38496 1324
rect 39480 1290 39514 1324
rect 7038 394 7072 428
rect 8056 394 8090 428
rect 9074 394 9108 428
rect 10092 394 10126 428
rect 11110 394 11144 428
rect 12128 394 12162 428
rect 13146 394 13180 428
rect 14164 394 14198 428
rect 15182 394 15216 428
rect 16200 394 16234 428
rect 17218 394 17252 428
rect 20150 44 20184 78
rect 21168 44 21202 78
rect 22186 44 22220 78
rect 23204 44 23238 78
rect 24222 44 24256 78
rect 25240 44 25274 78
rect 26258 44 26292 78
rect 27276 44 27310 78
rect 28294 44 28328 78
rect 29312 44 29346 78
rect 30330 44 30364 78
rect 31348 44 31382 78
rect 32366 44 32400 78
rect 33384 44 33418 78
rect 34402 44 34436 78
rect 35420 44 35454 78
rect 36438 44 36472 78
rect 37456 44 37490 78
rect 38474 44 38508 78
rect 39492 44 39526 78
rect 6848 -1052 6882 -1018
rect 7866 -1052 7900 -1018
rect 8884 -1052 8918 -1018
rect 9902 -1052 9936 -1018
rect 10920 -1052 10954 -1018
rect 11938 -1052 11972 -1018
rect 12956 -1052 12990 -1018
rect 13974 -1052 14008 -1018
rect 14992 -1052 15026 -1018
rect 16010 -1052 16044 -1018
rect 17028 -1052 17062 -1018
rect 20138 -1134 20172 -1100
rect 21156 -1134 21190 -1100
rect 22174 -1134 22208 -1100
rect 23192 -1134 23226 -1100
rect 24210 -1134 24244 -1100
rect 25228 -1134 25262 -1100
rect 26246 -1134 26280 -1100
rect 27264 -1134 27298 -1100
rect 28282 -1134 28316 -1100
rect 29300 -1134 29334 -1100
rect 30318 -1134 30352 -1100
rect 31336 -1134 31370 -1100
rect 32354 -1134 32388 -1100
rect 33372 -1134 33406 -1100
rect 34390 -1134 34424 -1100
rect 35408 -1134 35442 -1100
rect 36426 -1134 36460 -1100
rect 37444 -1134 37478 -1100
rect 38462 -1134 38496 -1100
rect 39480 -1134 39514 -1100
rect 41862 -1980 41962 13740
rect 4880 -2142 41800 -2042
<< nsubdiffcont >>
rect 17580 29302 41700 29402
rect 17418 14894 17518 29240
rect 24036 26824 24070 26858
rect 25054 26824 25088 26858
rect 26072 26824 26106 26858
rect 27090 26824 27124 26858
rect 28108 26824 28142 26858
rect 29126 26824 29160 26858
rect 30144 26824 30178 26858
rect 31162 26824 31196 26858
rect 32180 26824 32214 26858
rect 33198 26824 33232 26858
rect 34216 26824 34250 26858
rect 35234 26824 35268 26858
rect 36252 26824 36286 26858
rect 37270 26824 37304 26858
rect 38288 26824 38322 26858
rect 39306 26824 39340 26858
rect 24058 25670 24092 25704
rect 25076 25670 25110 25704
rect 26094 25670 26128 25704
rect 27112 25670 27146 25704
rect 28130 25670 28164 25704
rect 29148 25670 29182 25704
rect 30166 25670 30200 25704
rect 31184 25670 31218 25704
rect 32202 25670 32236 25704
rect 33220 25670 33254 25704
rect 34238 25670 34272 25704
rect 35256 25670 35290 25704
rect 36274 25670 36308 25704
rect 37292 25670 37326 25704
rect 38310 25670 38344 25704
rect 39328 25670 39362 25704
rect 24036 24538 24070 24572
rect 25054 24538 25088 24572
rect 26072 24538 26106 24572
rect 27090 24538 27124 24572
rect 28108 24538 28142 24572
rect 29126 24538 29160 24572
rect 30144 24538 30178 24572
rect 31162 24538 31196 24572
rect 32180 24538 32214 24572
rect 33198 24538 33232 24572
rect 34216 24538 34250 24572
rect 35234 24538 35268 24572
rect 36252 24538 36286 24572
rect 37270 24538 37304 24572
rect 38288 24538 38322 24572
rect 39306 24538 39340 24572
rect 24036 23156 24070 23190
rect 25054 23156 25088 23190
rect 26072 23156 26106 23190
rect 27090 23156 27124 23190
rect 28108 23156 28142 23190
rect 29126 23156 29160 23190
rect 30144 23156 30178 23190
rect 31162 23156 31196 23190
rect 32180 23156 32214 23190
rect 33198 23156 33232 23190
rect 34216 23156 34250 23190
rect 35234 23156 35268 23190
rect 36252 23156 36286 23190
rect 37270 23156 37304 23190
rect 38288 23156 38322 23190
rect 39306 23156 39340 23190
rect 24724 21808 24758 21842
rect 25742 21808 25776 21842
rect 26760 21808 26794 21842
rect 27778 21808 27812 21842
rect 28796 21808 28830 21842
rect 29814 21808 29848 21842
rect 30832 21808 30866 21842
rect 31850 21808 31884 21842
rect 32868 21808 32902 21842
rect 33886 21808 33920 21842
rect 34904 21808 34938 21842
rect 35922 21808 35956 21842
rect 36940 21808 36974 21842
rect 37958 21808 37992 21842
rect 38976 21808 39010 21842
rect 24330 20530 24364 20564
rect 25348 20530 25382 20564
rect 26366 20530 26400 20564
rect 27384 20530 27418 20564
rect 28402 20530 28436 20564
rect 29420 20530 29454 20564
rect 30438 20530 30472 20564
rect 31456 20530 31490 20564
rect 32474 20530 32508 20564
rect 33492 20530 33526 20564
rect 34510 20530 34544 20564
rect 35528 20530 35562 20564
rect 36546 20530 36580 20564
rect 37564 20530 37598 20564
rect 38582 20530 38616 20564
rect 39600 20530 39634 20564
rect 19732 20220 19766 20254
rect 20750 20220 20784 20254
rect 21768 20220 21802 20254
rect 22786 20220 22820 20254
rect 19208 19066 19242 19100
rect 20226 19066 20260 19100
rect 21244 19066 21278 19100
rect 22262 19066 22296 19100
rect 24420 19082 24454 19116
rect 25438 19082 25472 19116
rect 26456 19082 26490 19116
rect 27474 19082 27508 19116
rect 28492 19082 28526 19116
rect 29510 19082 29544 19116
rect 30528 19082 30562 19116
rect 31546 19082 31580 19116
rect 32564 19082 32598 19116
rect 33582 19082 33616 19116
rect 34600 19082 34634 19116
rect 35618 19082 35652 19116
rect 36636 19082 36670 19116
rect 37654 19082 37688 19116
rect 38672 19082 38706 19116
rect 39690 19082 39724 19116
rect 19218 18038 19252 18072
rect 20236 18038 20270 18072
rect 21254 18038 21288 18072
rect 22272 18038 22306 18072
rect 24444 17814 24478 17848
rect 25462 17814 25496 17848
rect 26480 17814 26514 17848
rect 27498 17814 27532 17848
rect 28516 17814 28550 17848
rect 29534 17814 29568 17848
rect 30552 17814 30586 17848
rect 31570 17814 31604 17848
rect 32588 17814 32622 17848
rect 33606 17814 33640 17848
rect 34624 17814 34658 17848
rect 35642 17814 35676 17848
rect 36660 17814 36694 17848
rect 37678 17814 37712 17848
rect 38696 17814 38730 17848
rect 39714 17814 39748 17848
rect 19208 17010 19242 17044
rect 20226 17010 20260 17044
rect 21244 17010 21278 17044
rect 22262 17010 22296 17044
rect 24308 16570 24342 16604
rect 25326 16570 25360 16604
rect 26344 16570 26378 16604
rect 27362 16570 27396 16604
rect 28380 16570 28414 16604
rect 29398 16570 29432 16604
rect 30416 16570 30450 16604
rect 31434 16570 31468 16604
rect 32452 16570 32486 16604
rect 33470 16570 33504 16604
rect 34488 16570 34522 16604
rect 35506 16570 35540 16604
rect 36524 16570 36558 16604
rect 37542 16570 37576 16604
rect 38560 16570 38594 16604
rect 39578 16570 39612 16604
rect 19732 15858 19766 15892
rect 20750 15858 20784 15892
rect 21768 15858 21802 15892
rect 22786 15858 22820 15892
rect 41762 14894 41862 29240
rect 17580 14732 41700 14832
<< poly >>
rect 23760 26635 24348 26651
rect 23760 26618 23776 26635
rect 23574 26601 23776 26618
rect 24332 26618 24348 26635
rect 24778 26635 25366 26651
rect 24778 26618 24794 26635
rect 24332 26601 24534 26618
rect 23574 26554 24534 26601
rect 24592 26601 24794 26618
rect 25350 26618 25366 26635
rect 25796 26635 26384 26651
rect 25796 26618 25812 26635
rect 25350 26601 25552 26618
rect 24592 26554 25552 26601
rect 25610 26601 25812 26618
rect 26368 26618 26384 26635
rect 26814 26635 27402 26651
rect 26814 26618 26830 26635
rect 26368 26601 26570 26618
rect 25610 26554 26570 26601
rect 26628 26601 26830 26618
rect 27386 26618 27402 26635
rect 27832 26635 28420 26651
rect 27832 26618 27848 26635
rect 27386 26601 27588 26618
rect 26628 26554 27588 26601
rect 27646 26601 27848 26618
rect 28404 26618 28420 26635
rect 28850 26635 29438 26651
rect 28850 26618 28866 26635
rect 28404 26601 28606 26618
rect 27646 26554 28606 26601
rect 28664 26601 28866 26618
rect 29422 26618 29438 26635
rect 29868 26635 30456 26651
rect 29868 26618 29884 26635
rect 29422 26601 29624 26618
rect 28664 26554 29624 26601
rect 29682 26601 29884 26618
rect 30440 26618 30456 26635
rect 30886 26635 31474 26651
rect 30886 26618 30902 26635
rect 30440 26601 30642 26618
rect 29682 26554 30642 26601
rect 30700 26601 30902 26618
rect 31458 26618 31474 26635
rect 31904 26635 32492 26651
rect 31904 26618 31920 26635
rect 31458 26601 31660 26618
rect 30700 26554 31660 26601
rect 31718 26601 31920 26618
rect 32476 26618 32492 26635
rect 32922 26635 33510 26651
rect 32922 26618 32938 26635
rect 32476 26601 32678 26618
rect 31718 26554 32678 26601
rect 32736 26601 32938 26618
rect 33494 26618 33510 26635
rect 33940 26635 34528 26651
rect 33940 26618 33956 26635
rect 33494 26601 33696 26618
rect 32736 26554 33696 26601
rect 33754 26601 33956 26618
rect 34512 26618 34528 26635
rect 34958 26635 35546 26651
rect 34958 26618 34974 26635
rect 34512 26601 34714 26618
rect 33754 26554 34714 26601
rect 34772 26601 34974 26618
rect 35530 26618 35546 26635
rect 35976 26635 36564 26651
rect 35976 26618 35992 26635
rect 35530 26601 35732 26618
rect 34772 26554 35732 26601
rect 35790 26601 35992 26618
rect 36548 26618 36564 26635
rect 36994 26635 37582 26651
rect 36994 26618 37010 26635
rect 36548 26601 36750 26618
rect 35790 26554 36750 26601
rect 36808 26601 37010 26618
rect 37566 26618 37582 26635
rect 38012 26635 38600 26651
rect 38012 26618 38028 26635
rect 37566 26601 37768 26618
rect 36808 26554 37768 26601
rect 37826 26601 38028 26618
rect 38584 26618 38600 26635
rect 39030 26635 39618 26651
rect 39030 26618 39046 26635
rect 38584 26601 38786 26618
rect 37826 26554 38786 26601
rect 38844 26601 39046 26618
rect 39602 26618 39618 26635
rect 39602 26601 39804 26618
rect 38844 26554 39804 26601
rect 23574 25907 24534 25954
rect 23574 25890 23776 25907
rect 23760 25873 23776 25890
rect 24332 25890 24534 25907
rect 24592 25907 25552 25954
rect 24592 25890 24794 25907
rect 24332 25873 24348 25890
rect 23760 25857 24348 25873
rect 24778 25873 24794 25890
rect 25350 25890 25552 25907
rect 25610 25907 26570 25954
rect 25610 25890 25812 25907
rect 25350 25873 25366 25890
rect 24778 25857 25366 25873
rect 25796 25873 25812 25890
rect 26368 25890 26570 25907
rect 26628 25907 27588 25954
rect 26628 25890 26830 25907
rect 26368 25873 26384 25890
rect 25796 25857 26384 25873
rect 26814 25873 26830 25890
rect 27386 25890 27588 25907
rect 27646 25907 28606 25954
rect 27646 25890 27848 25907
rect 27386 25873 27402 25890
rect 26814 25857 27402 25873
rect 27832 25873 27848 25890
rect 28404 25890 28606 25907
rect 28664 25907 29624 25954
rect 28664 25890 28866 25907
rect 28404 25873 28420 25890
rect 27832 25857 28420 25873
rect 28850 25873 28866 25890
rect 29422 25890 29624 25907
rect 29682 25907 30642 25954
rect 29682 25890 29884 25907
rect 29422 25873 29438 25890
rect 28850 25857 29438 25873
rect 29868 25873 29884 25890
rect 30440 25890 30642 25907
rect 30700 25907 31660 25954
rect 30700 25890 30902 25907
rect 30440 25873 30456 25890
rect 29868 25857 30456 25873
rect 30886 25873 30902 25890
rect 31458 25890 31660 25907
rect 31718 25907 32678 25954
rect 31718 25890 31920 25907
rect 31458 25873 31474 25890
rect 30886 25857 31474 25873
rect 31904 25873 31920 25890
rect 32476 25890 32678 25907
rect 32736 25907 33696 25954
rect 32736 25890 32938 25907
rect 32476 25873 32492 25890
rect 31904 25857 32492 25873
rect 32922 25873 32938 25890
rect 33494 25890 33696 25907
rect 33754 25907 34714 25954
rect 33754 25890 33956 25907
rect 33494 25873 33510 25890
rect 32922 25857 33510 25873
rect 33940 25873 33956 25890
rect 34512 25890 34714 25907
rect 34772 25907 35732 25954
rect 34772 25890 34974 25907
rect 34512 25873 34528 25890
rect 33940 25857 34528 25873
rect 34958 25873 34974 25890
rect 35530 25890 35732 25907
rect 35790 25907 36750 25954
rect 35790 25890 35992 25907
rect 35530 25873 35546 25890
rect 34958 25857 35546 25873
rect 35976 25873 35992 25890
rect 36548 25890 36750 25907
rect 36808 25907 37768 25954
rect 36808 25890 37010 25907
rect 36548 25873 36564 25890
rect 35976 25857 36564 25873
rect 36994 25873 37010 25890
rect 37566 25890 37768 25907
rect 37826 25907 38786 25954
rect 37826 25890 38028 25907
rect 37566 25873 37582 25890
rect 36994 25857 37582 25873
rect 38012 25873 38028 25890
rect 38584 25890 38786 25907
rect 38844 25907 39804 25954
rect 38844 25890 39046 25907
rect 38584 25873 38600 25890
rect 38012 25857 38600 25873
rect 39030 25873 39046 25890
rect 39602 25890 39804 25907
rect 39602 25873 39618 25890
rect 39030 25857 39618 25873
rect 23760 25499 24348 25515
rect 23760 25482 23776 25499
rect 23574 25465 23776 25482
rect 24332 25482 24348 25499
rect 24778 25499 25366 25515
rect 24778 25482 24794 25499
rect 24332 25465 24534 25482
rect 23574 25418 24534 25465
rect 24592 25465 24794 25482
rect 25350 25482 25366 25499
rect 25796 25499 26384 25515
rect 25796 25482 25812 25499
rect 25350 25465 25552 25482
rect 24592 25418 25552 25465
rect 25610 25465 25812 25482
rect 26368 25482 26384 25499
rect 26814 25499 27402 25515
rect 26814 25482 26830 25499
rect 26368 25465 26570 25482
rect 25610 25418 26570 25465
rect 26628 25465 26830 25482
rect 27386 25482 27402 25499
rect 27832 25499 28420 25515
rect 27832 25482 27848 25499
rect 27386 25465 27588 25482
rect 26628 25418 27588 25465
rect 27646 25465 27848 25482
rect 28404 25482 28420 25499
rect 28850 25499 29438 25515
rect 28850 25482 28866 25499
rect 28404 25465 28606 25482
rect 27646 25418 28606 25465
rect 28664 25465 28866 25482
rect 29422 25482 29438 25499
rect 29868 25499 30456 25515
rect 29868 25482 29884 25499
rect 29422 25465 29624 25482
rect 28664 25418 29624 25465
rect 29682 25465 29884 25482
rect 30440 25482 30456 25499
rect 30886 25499 31474 25515
rect 30886 25482 30902 25499
rect 30440 25465 30642 25482
rect 29682 25418 30642 25465
rect 30700 25465 30902 25482
rect 31458 25482 31474 25499
rect 31904 25499 32492 25515
rect 31904 25482 31920 25499
rect 31458 25465 31660 25482
rect 30700 25418 31660 25465
rect 31718 25465 31920 25482
rect 32476 25482 32492 25499
rect 32922 25499 33510 25515
rect 32922 25482 32938 25499
rect 32476 25465 32678 25482
rect 31718 25418 32678 25465
rect 32736 25465 32938 25482
rect 33494 25482 33510 25499
rect 33940 25499 34528 25515
rect 33940 25482 33956 25499
rect 33494 25465 33696 25482
rect 32736 25418 33696 25465
rect 33754 25465 33956 25482
rect 34512 25482 34528 25499
rect 34958 25499 35546 25515
rect 34958 25482 34974 25499
rect 34512 25465 34714 25482
rect 33754 25418 34714 25465
rect 34772 25465 34974 25482
rect 35530 25482 35546 25499
rect 35976 25499 36564 25515
rect 35976 25482 35992 25499
rect 35530 25465 35732 25482
rect 34772 25418 35732 25465
rect 35790 25465 35992 25482
rect 36548 25482 36564 25499
rect 36994 25499 37582 25515
rect 36994 25482 37010 25499
rect 36548 25465 36750 25482
rect 35790 25418 36750 25465
rect 36808 25465 37010 25482
rect 37566 25482 37582 25499
rect 38012 25499 38600 25515
rect 38012 25482 38028 25499
rect 37566 25465 37768 25482
rect 36808 25418 37768 25465
rect 37826 25465 38028 25482
rect 38584 25482 38600 25499
rect 39030 25499 39618 25515
rect 39030 25482 39046 25499
rect 38584 25465 38786 25482
rect 37826 25418 38786 25465
rect 38844 25465 39046 25482
rect 39602 25482 39618 25499
rect 39602 25465 39804 25482
rect 38844 25418 39804 25465
rect 23574 24771 24534 24818
rect 23574 24754 23776 24771
rect 23760 24737 23776 24754
rect 24332 24754 24534 24771
rect 24592 24771 25552 24818
rect 24592 24754 24794 24771
rect 24332 24737 24348 24754
rect 23760 24721 24348 24737
rect 24778 24737 24794 24754
rect 25350 24754 25552 24771
rect 25610 24771 26570 24818
rect 25610 24754 25812 24771
rect 25350 24737 25366 24754
rect 24778 24721 25366 24737
rect 25796 24737 25812 24754
rect 26368 24754 26570 24771
rect 26628 24771 27588 24818
rect 26628 24754 26830 24771
rect 26368 24737 26384 24754
rect 25796 24721 26384 24737
rect 26814 24737 26830 24754
rect 27386 24754 27588 24771
rect 27646 24771 28606 24818
rect 27646 24754 27848 24771
rect 27386 24737 27402 24754
rect 26814 24721 27402 24737
rect 27832 24737 27848 24754
rect 28404 24754 28606 24771
rect 28664 24771 29624 24818
rect 28664 24754 28866 24771
rect 28404 24737 28420 24754
rect 27832 24721 28420 24737
rect 28850 24737 28866 24754
rect 29422 24754 29624 24771
rect 29682 24771 30642 24818
rect 29682 24754 29884 24771
rect 29422 24737 29438 24754
rect 28850 24721 29438 24737
rect 29868 24737 29884 24754
rect 30440 24754 30642 24771
rect 30700 24771 31660 24818
rect 30700 24754 30902 24771
rect 30440 24737 30456 24754
rect 29868 24721 30456 24737
rect 30886 24737 30902 24754
rect 31458 24754 31660 24771
rect 31718 24771 32678 24818
rect 31718 24754 31920 24771
rect 31458 24737 31474 24754
rect 30886 24721 31474 24737
rect 31904 24737 31920 24754
rect 32476 24754 32678 24771
rect 32736 24771 33696 24818
rect 32736 24754 32938 24771
rect 32476 24737 32492 24754
rect 31904 24721 32492 24737
rect 32922 24737 32938 24754
rect 33494 24754 33696 24771
rect 33754 24771 34714 24818
rect 33754 24754 33956 24771
rect 33494 24737 33510 24754
rect 32922 24721 33510 24737
rect 33940 24737 33956 24754
rect 34512 24754 34714 24771
rect 34772 24771 35732 24818
rect 34772 24754 34974 24771
rect 34512 24737 34528 24754
rect 33940 24721 34528 24737
rect 34958 24737 34974 24754
rect 35530 24754 35732 24771
rect 35790 24771 36750 24818
rect 35790 24754 35992 24771
rect 35530 24737 35546 24754
rect 34958 24721 35546 24737
rect 35976 24737 35992 24754
rect 36548 24754 36750 24771
rect 36808 24771 37768 24818
rect 36808 24754 37010 24771
rect 36548 24737 36564 24754
rect 35976 24721 36564 24737
rect 36994 24737 37010 24754
rect 37566 24754 37768 24771
rect 37826 24771 38786 24818
rect 37826 24754 38028 24771
rect 37566 24737 37582 24754
rect 36994 24721 37582 24737
rect 38012 24737 38028 24754
rect 38584 24754 38786 24771
rect 38844 24771 39804 24818
rect 38844 24754 39046 24771
rect 38584 24737 38600 24754
rect 38012 24721 38600 24737
rect 39030 24737 39046 24754
rect 39602 24754 39804 24771
rect 39602 24737 39618 24754
rect 39030 24721 39618 24737
rect 23760 24363 24348 24379
rect 23760 24346 23776 24363
rect 23574 24329 23776 24346
rect 24332 24346 24348 24363
rect 24778 24363 25366 24379
rect 24778 24346 24794 24363
rect 24332 24329 24534 24346
rect 23574 24282 24534 24329
rect 24592 24329 24794 24346
rect 25350 24346 25366 24363
rect 25796 24363 26384 24379
rect 25796 24346 25812 24363
rect 25350 24329 25552 24346
rect 24592 24282 25552 24329
rect 25610 24329 25812 24346
rect 26368 24346 26384 24363
rect 26814 24363 27402 24379
rect 26814 24346 26830 24363
rect 26368 24329 26570 24346
rect 25610 24282 26570 24329
rect 26628 24329 26830 24346
rect 27386 24346 27402 24363
rect 27832 24363 28420 24379
rect 27832 24346 27848 24363
rect 27386 24329 27588 24346
rect 26628 24282 27588 24329
rect 27646 24329 27848 24346
rect 28404 24346 28420 24363
rect 28850 24363 29438 24379
rect 28850 24346 28866 24363
rect 28404 24329 28606 24346
rect 27646 24282 28606 24329
rect 28664 24329 28866 24346
rect 29422 24346 29438 24363
rect 29868 24363 30456 24379
rect 29868 24346 29884 24363
rect 29422 24329 29624 24346
rect 28664 24282 29624 24329
rect 29682 24329 29884 24346
rect 30440 24346 30456 24363
rect 30886 24363 31474 24379
rect 30886 24346 30902 24363
rect 30440 24329 30642 24346
rect 29682 24282 30642 24329
rect 30700 24329 30902 24346
rect 31458 24346 31474 24363
rect 31904 24363 32492 24379
rect 31904 24346 31920 24363
rect 31458 24329 31660 24346
rect 30700 24282 31660 24329
rect 31718 24329 31920 24346
rect 32476 24346 32492 24363
rect 32922 24363 33510 24379
rect 32922 24346 32938 24363
rect 32476 24329 32678 24346
rect 31718 24282 32678 24329
rect 32736 24329 32938 24346
rect 33494 24346 33510 24363
rect 33940 24363 34528 24379
rect 33940 24346 33956 24363
rect 33494 24329 33696 24346
rect 32736 24282 33696 24329
rect 33754 24329 33956 24346
rect 34512 24346 34528 24363
rect 34958 24363 35546 24379
rect 34958 24346 34974 24363
rect 34512 24329 34714 24346
rect 33754 24282 34714 24329
rect 34772 24329 34974 24346
rect 35530 24346 35546 24363
rect 35976 24363 36564 24379
rect 35976 24346 35992 24363
rect 35530 24329 35732 24346
rect 34772 24282 35732 24329
rect 35790 24329 35992 24346
rect 36548 24346 36564 24363
rect 36994 24363 37582 24379
rect 36994 24346 37010 24363
rect 36548 24329 36750 24346
rect 35790 24282 36750 24329
rect 36808 24329 37010 24346
rect 37566 24346 37582 24363
rect 38012 24363 38600 24379
rect 38012 24346 38028 24363
rect 37566 24329 37768 24346
rect 36808 24282 37768 24329
rect 37826 24329 38028 24346
rect 38584 24346 38600 24363
rect 39030 24363 39618 24379
rect 39030 24346 39046 24363
rect 38584 24329 38786 24346
rect 37826 24282 38786 24329
rect 38844 24329 39046 24346
rect 39602 24346 39618 24363
rect 39602 24329 39804 24346
rect 38844 24282 39804 24329
rect 23574 23635 24534 23682
rect 23574 23618 23776 23635
rect 23760 23601 23776 23618
rect 24332 23618 24534 23635
rect 24592 23635 25552 23682
rect 24592 23618 24794 23635
rect 24332 23601 24348 23618
rect 23760 23585 24348 23601
rect 24778 23601 24794 23618
rect 25350 23618 25552 23635
rect 25610 23635 26570 23682
rect 25610 23618 25812 23635
rect 25350 23601 25366 23618
rect 24778 23585 25366 23601
rect 25796 23601 25812 23618
rect 26368 23618 26570 23635
rect 26628 23635 27588 23682
rect 26628 23618 26830 23635
rect 26368 23601 26384 23618
rect 25796 23585 26384 23601
rect 26814 23601 26830 23618
rect 27386 23618 27588 23635
rect 27646 23635 28606 23682
rect 27646 23618 27848 23635
rect 27386 23601 27402 23618
rect 26814 23585 27402 23601
rect 27832 23601 27848 23618
rect 28404 23618 28606 23635
rect 28664 23635 29624 23682
rect 28664 23618 28866 23635
rect 28404 23601 28420 23618
rect 27832 23585 28420 23601
rect 28850 23601 28866 23618
rect 29422 23618 29624 23635
rect 29682 23635 30642 23682
rect 29682 23618 29884 23635
rect 29422 23601 29438 23618
rect 28850 23585 29438 23601
rect 29868 23601 29884 23618
rect 30440 23618 30642 23635
rect 30700 23635 31660 23682
rect 30700 23618 30902 23635
rect 30440 23601 30456 23618
rect 29868 23585 30456 23601
rect 30886 23601 30902 23618
rect 31458 23618 31660 23635
rect 31718 23635 32678 23682
rect 31718 23618 31920 23635
rect 31458 23601 31474 23618
rect 30886 23585 31474 23601
rect 31904 23601 31920 23618
rect 32476 23618 32678 23635
rect 32736 23635 33696 23682
rect 32736 23618 32938 23635
rect 32476 23601 32492 23618
rect 31904 23585 32492 23601
rect 32922 23601 32938 23618
rect 33494 23618 33696 23635
rect 33754 23635 34714 23682
rect 33754 23618 33956 23635
rect 33494 23601 33510 23618
rect 32922 23585 33510 23601
rect 33940 23601 33956 23618
rect 34512 23618 34714 23635
rect 34772 23635 35732 23682
rect 34772 23618 34974 23635
rect 34512 23601 34528 23618
rect 33940 23585 34528 23601
rect 34958 23601 34974 23618
rect 35530 23618 35732 23635
rect 35790 23635 36750 23682
rect 35790 23618 35992 23635
rect 35530 23601 35546 23618
rect 34958 23585 35546 23601
rect 35976 23601 35992 23618
rect 36548 23618 36750 23635
rect 36808 23635 37768 23682
rect 36808 23618 37010 23635
rect 36548 23601 36564 23618
rect 35976 23585 36564 23601
rect 36994 23601 37010 23618
rect 37566 23618 37768 23635
rect 37826 23635 38786 23682
rect 37826 23618 38028 23635
rect 37566 23601 37582 23618
rect 36994 23585 37582 23601
rect 38012 23601 38028 23618
rect 38584 23618 38786 23635
rect 38844 23635 39804 23682
rect 38844 23618 39046 23635
rect 38584 23601 38600 23618
rect 38012 23585 38600 23601
rect 39030 23601 39046 23618
rect 39602 23618 39804 23635
rect 39602 23601 39618 23618
rect 39030 23585 39618 23601
rect 24954 22725 25542 22741
rect 24954 22708 24970 22725
rect 24768 22691 24970 22708
rect 25526 22708 25542 22725
rect 25972 22725 26560 22741
rect 25972 22708 25988 22725
rect 25526 22691 25728 22708
rect 24768 22644 25728 22691
rect 25786 22691 25988 22708
rect 26544 22708 26560 22725
rect 26990 22725 27578 22741
rect 26990 22708 27006 22725
rect 26544 22691 26746 22708
rect 25786 22644 26746 22691
rect 26804 22691 27006 22708
rect 27562 22708 27578 22725
rect 28008 22725 28596 22741
rect 28008 22708 28024 22725
rect 27562 22691 27764 22708
rect 26804 22644 27764 22691
rect 27822 22691 28024 22708
rect 28580 22708 28596 22725
rect 29026 22725 29614 22741
rect 29026 22708 29042 22725
rect 28580 22691 28782 22708
rect 27822 22644 28782 22691
rect 28840 22691 29042 22708
rect 29598 22708 29614 22725
rect 30044 22725 30632 22741
rect 30044 22708 30060 22725
rect 29598 22691 29800 22708
rect 28840 22644 29800 22691
rect 29858 22691 30060 22708
rect 30616 22708 30632 22725
rect 31062 22725 31650 22741
rect 31062 22708 31078 22725
rect 30616 22691 30818 22708
rect 29858 22644 30818 22691
rect 30876 22691 31078 22708
rect 31634 22708 31650 22725
rect 32080 22725 32668 22741
rect 32080 22708 32096 22725
rect 31634 22691 31836 22708
rect 30876 22644 31836 22691
rect 31894 22691 32096 22708
rect 32652 22708 32668 22725
rect 33098 22725 33686 22741
rect 33098 22708 33114 22725
rect 32652 22691 32854 22708
rect 31894 22644 32854 22691
rect 32912 22691 33114 22708
rect 33670 22708 33686 22725
rect 34116 22725 34704 22741
rect 34116 22708 34132 22725
rect 33670 22691 33872 22708
rect 32912 22644 33872 22691
rect 33930 22691 34132 22708
rect 34688 22708 34704 22725
rect 35134 22725 35722 22741
rect 35134 22708 35150 22725
rect 34688 22691 34890 22708
rect 33930 22644 34890 22691
rect 34948 22691 35150 22708
rect 35706 22708 35722 22725
rect 36152 22725 36740 22741
rect 36152 22708 36168 22725
rect 35706 22691 35908 22708
rect 34948 22644 35908 22691
rect 35966 22691 36168 22708
rect 36724 22708 36740 22725
rect 37170 22725 37758 22741
rect 37170 22708 37186 22725
rect 36724 22691 36926 22708
rect 35966 22644 36926 22691
rect 36984 22691 37186 22708
rect 37742 22708 37758 22725
rect 38188 22725 38776 22741
rect 38188 22708 38204 22725
rect 37742 22691 37944 22708
rect 36984 22644 37944 22691
rect 38002 22691 38204 22708
rect 38760 22708 38776 22725
rect 38760 22691 38962 22708
rect 38002 22644 38962 22691
rect 24768 21997 25728 22044
rect 24768 21980 24970 21997
rect 24954 21963 24970 21980
rect 25526 21980 25728 21997
rect 25786 21997 26746 22044
rect 25786 21980 25988 21997
rect 25526 21963 25542 21980
rect 24954 21947 25542 21963
rect 25972 21963 25988 21980
rect 26544 21980 26746 21997
rect 26804 21997 27764 22044
rect 26804 21980 27006 21997
rect 26544 21963 26560 21980
rect 25972 21947 26560 21963
rect 26990 21963 27006 21980
rect 27562 21980 27764 21997
rect 27822 21997 28782 22044
rect 27822 21980 28024 21997
rect 27562 21963 27578 21980
rect 26990 21947 27578 21963
rect 28008 21963 28024 21980
rect 28580 21980 28782 21997
rect 28840 21997 29800 22044
rect 28840 21980 29042 21997
rect 28580 21963 28596 21980
rect 28008 21947 28596 21963
rect 29026 21963 29042 21980
rect 29598 21980 29800 21997
rect 29858 21997 30818 22044
rect 29858 21980 30060 21997
rect 29598 21963 29614 21980
rect 29026 21947 29614 21963
rect 30044 21963 30060 21980
rect 30616 21980 30818 21997
rect 30876 21997 31836 22044
rect 30876 21980 31078 21997
rect 30616 21963 30632 21980
rect 30044 21947 30632 21963
rect 31062 21963 31078 21980
rect 31634 21980 31836 21997
rect 31894 21997 32854 22044
rect 31894 21980 32096 21997
rect 31634 21963 31650 21980
rect 31062 21947 31650 21963
rect 32080 21963 32096 21980
rect 32652 21980 32854 21997
rect 32912 21997 33872 22044
rect 32912 21980 33114 21997
rect 32652 21963 32668 21980
rect 32080 21947 32668 21963
rect 33098 21963 33114 21980
rect 33670 21980 33872 21997
rect 33930 21997 34890 22044
rect 33930 21980 34132 21997
rect 33670 21963 33686 21980
rect 33098 21947 33686 21963
rect 34116 21963 34132 21980
rect 34688 21980 34890 21997
rect 34948 21997 35908 22044
rect 34948 21980 35150 21997
rect 34688 21963 34704 21980
rect 34116 21947 34704 21963
rect 35134 21963 35150 21980
rect 35706 21980 35908 21997
rect 35966 21997 36926 22044
rect 35966 21980 36168 21997
rect 35706 21963 35722 21980
rect 35134 21947 35722 21963
rect 36152 21963 36168 21980
rect 36724 21980 36926 21997
rect 36984 21997 37944 22044
rect 36984 21980 37186 21997
rect 36724 21963 36740 21980
rect 36152 21947 36740 21963
rect 37170 21963 37186 21980
rect 37742 21980 37944 21997
rect 38002 21997 38962 22044
rect 38002 21980 38204 21997
rect 37742 21963 37758 21980
rect 37170 21947 37758 21963
rect 38188 21963 38204 21980
rect 38760 21980 38962 21997
rect 38760 21963 38776 21980
rect 38188 21947 38776 21963
rect 24954 21693 25542 21709
rect 24954 21676 24970 21693
rect 24768 21659 24970 21676
rect 25526 21676 25542 21693
rect 25972 21693 26560 21709
rect 25972 21676 25988 21693
rect 25526 21659 25728 21676
rect 24768 21612 25728 21659
rect 25786 21659 25988 21676
rect 26544 21676 26560 21693
rect 26990 21693 27578 21709
rect 26990 21676 27006 21693
rect 26544 21659 26746 21676
rect 25786 21612 26746 21659
rect 26804 21659 27006 21676
rect 27562 21676 27578 21693
rect 28008 21693 28596 21709
rect 28008 21676 28024 21693
rect 27562 21659 27764 21676
rect 26804 21612 27764 21659
rect 27822 21659 28024 21676
rect 28580 21676 28596 21693
rect 29026 21693 29614 21709
rect 29026 21676 29042 21693
rect 28580 21659 28782 21676
rect 27822 21612 28782 21659
rect 28840 21659 29042 21676
rect 29598 21676 29614 21693
rect 30044 21693 30632 21709
rect 30044 21676 30060 21693
rect 29598 21659 29800 21676
rect 28840 21612 29800 21659
rect 29858 21659 30060 21676
rect 30616 21676 30632 21693
rect 31062 21693 31650 21709
rect 31062 21676 31078 21693
rect 30616 21659 30818 21676
rect 29858 21612 30818 21659
rect 30876 21659 31078 21676
rect 31634 21676 31650 21693
rect 32080 21693 32668 21709
rect 32080 21676 32096 21693
rect 31634 21659 31836 21676
rect 30876 21612 31836 21659
rect 31894 21659 32096 21676
rect 32652 21676 32668 21693
rect 33098 21693 33686 21709
rect 33098 21676 33114 21693
rect 32652 21659 32854 21676
rect 31894 21612 32854 21659
rect 32912 21659 33114 21676
rect 33670 21676 33686 21693
rect 34116 21693 34704 21709
rect 34116 21676 34132 21693
rect 33670 21659 33872 21676
rect 32912 21612 33872 21659
rect 33930 21659 34132 21676
rect 34688 21676 34704 21693
rect 35134 21693 35722 21709
rect 35134 21676 35150 21693
rect 34688 21659 34890 21676
rect 33930 21612 34890 21659
rect 34948 21659 35150 21676
rect 35706 21676 35722 21693
rect 36152 21693 36740 21709
rect 36152 21676 36168 21693
rect 35706 21659 35908 21676
rect 34948 21612 35908 21659
rect 35966 21659 36168 21676
rect 36724 21676 36740 21693
rect 37170 21693 37758 21709
rect 37170 21676 37186 21693
rect 36724 21659 36926 21676
rect 35966 21612 36926 21659
rect 36984 21659 37186 21676
rect 37742 21676 37758 21693
rect 38188 21693 38776 21709
rect 38188 21676 38204 21693
rect 37742 21659 37944 21676
rect 36984 21612 37944 21659
rect 38002 21659 38204 21676
rect 38760 21676 38776 21693
rect 38760 21659 38962 21676
rect 38002 21612 38962 21659
rect 24768 20965 25728 21012
rect 24768 20948 24970 20965
rect 24954 20931 24970 20948
rect 25526 20948 25728 20965
rect 25786 20965 26746 21012
rect 25786 20948 25988 20965
rect 25526 20931 25542 20948
rect 24954 20915 25542 20931
rect 25972 20931 25988 20948
rect 26544 20948 26746 20965
rect 26804 20965 27764 21012
rect 26804 20948 27006 20965
rect 26544 20931 26560 20948
rect 25972 20915 26560 20931
rect 26990 20931 27006 20948
rect 27562 20948 27764 20965
rect 27822 20965 28782 21012
rect 27822 20948 28024 20965
rect 27562 20931 27578 20948
rect 26990 20915 27578 20931
rect 28008 20931 28024 20948
rect 28580 20948 28782 20965
rect 28840 20965 29800 21012
rect 28840 20948 29042 20965
rect 28580 20931 28596 20948
rect 28008 20915 28596 20931
rect 29026 20931 29042 20948
rect 29598 20948 29800 20965
rect 29858 20965 30818 21012
rect 29858 20948 30060 20965
rect 29598 20931 29614 20948
rect 29026 20915 29614 20931
rect 30044 20931 30060 20948
rect 30616 20948 30818 20965
rect 30876 20965 31836 21012
rect 30876 20948 31078 20965
rect 30616 20931 30632 20948
rect 30044 20915 30632 20931
rect 31062 20931 31078 20948
rect 31634 20948 31836 20965
rect 31894 20965 32854 21012
rect 31894 20948 32096 20965
rect 31634 20931 31650 20948
rect 31062 20915 31650 20931
rect 32080 20931 32096 20948
rect 32652 20948 32854 20965
rect 32912 20965 33872 21012
rect 32912 20948 33114 20965
rect 32652 20931 32668 20948
rect 32080 20915 32668 20931
rect 33098 20931 33114 20948
rect 33670 20948 33872 20965
rect 33930 20965 34890 21012
rect 33930 20948 34132 20965
rect 33670 20931 33686 20948
rect 33098 20915 33686 20931
rect 34116 20931 34132 20948
rect 34688 20948 34890 20965
rect 34948 20965 35908 21012
rect 34948 20948 35150 20965
rect 34688 20931 34704 20948
rect 34116 20915 34704 20931
rect 35134 20931 35150 20948
rect 35706 20948 35908 20965
rect 35966 20965 36926 21012
rect 35966 20948 36168 20965
rect 35706 20931 35722 20948
rect 35134 20915 35722 20931
rect 36152 20931 36168 20948
rect 36724 20948 36926 20965
rect 36984 20965 37944 21012
rect 36984 20948 37186 20965
rect 36724 20931 36740 20948
rect 36152 20915 36740 20931
rect 37170 20931 37186 20948
rect 37742 20948 37944 20965
rect 38002 20965 38962 21012
rect 38002 20948 38204 20965
rect 37742 20931 37758 20948
rect 37170 20915 37758 20931
rect 38188 20931 38204 20948
rect 38760 20948 38962 20965
rect 38760 20931 38776 20948
rect 38188 20915 38776 20931
rect 24746 20089 25334 20105
rect 24746 20072 24762 20089
rect 24560 20055 24762 20072
rect 25318 20072 25334 20089
rect 25764 20089 26352 20105
rect 25764 20072 25780 20089
rect 25318 20055 25520 20072
rect 24560 20008 25520 20055
rect 25578 20055 25780 20072
rect 26336 20072 26352 20089
rect 26782 20089 27370 20105
rect 26782 20072 26798 20089
rect 26336 20055 26538 20072
rect 25578 20008 26538 20055
rect 26596 20055 26798 20072
rect 27354 20072 27370 20089
rect 27800 20089 28388 20105
rect 27800 20072 27816 20089
rect 27354 20055 27556 20072
rect 26596 20008 27556 20055
rect 27614 20055 27816 20072
rect 28372 20072 28388 20089
rect 28818 20089 29406 20105
rect 28818 20072 28834 20089
rect 28372 20055 28574 20072
rect 27614 20008 28574 20055
rect 28632 20055 28834 20072
rect 29390 20072 29406 20089
rect 29836 20089 30424 20105
rect 29836 20072 29852 20089
rect 29390 20055 29592 20072
rect 28632 20008 29592 20055
rect 29650 20055 29852 20072
rect 30408 20072 30424 20089
rect 30854 20089 31442 20105
rect 30854 20072 30870 20089
rect 30408 20055 30610 20072
rect 29650 20008 30610 20055
rect 30668 20055 30870 20072
rect 31426 20072 31442 20089
rect 31872 20089 32460 20105
rect 31872 20072 31888 20089
rect 31426 20055 31628 20072
rect 30668 20008 31628 20055
rect 31686 20055 31888 20072
rect 32444 20072 32460 20089
rect 32890 20089 33478 20105
rect 32890 20072 32906 20089
rect 32444 20055 32646 20072
rect 31686 20008 32646 20055
rect 32704 20055 32906 20072
rect 33462 20072 33478 20089
rect 33908 20089 34496 20105
rect 33908 20072 33924 20089
rect 33462 20055 33664 20072
rect 32704 20008 33664 20055
rect 33722 20055 33924 20072
rect 34480 20072 34496 20089
rect 34926 20089 35514 20105
rect 34926 20072 34942 20089
rect 34480 20055 34682 20072
rect 33722 20008 34682 20055
rect 34740 20055 34942 20072
rect 35498 20072 35514 20089
rect 35944 20089 36532 20105
rect 35944 20072 35960 20089
rect 35498 20055 35700 20072
rect 34740 20008 35700 20055
rect 35758 20055 35960 20072
rect 36516 20072 36532 20089
rect 36962 20089 37550 20105
rect 36962 20072 36978 20089
rect 36516 20055 36718 20072
rect 35758 20008 36718 20055
rect 36776 20055 36978 20072
rect 37534 20072 37550 20089
rect 37980 20089 38568 20105
rect 37980 20072 37996 20089
rect 37534 20055 37736 20072
rect 36776 20008 37736 20055
rect 37794 20055 37996 20072
rect 38552 20072 38568 20089
rect 38998 20089 39586 20105
rect 38998 20072 39014 20089
rect 38552 20055 38754 20072
rect 37794 20008 38754 20055
rect 38812 20055 39014 20072
rect 39570 20072 39586 20089
rect 39570 20055 39772 20072
rect 38812 20008 39772 20055
rect 19442 19985 20030 20001
rect 19442 19968 19458 19985
rect 19256 19951 19458 19968
rect 20014 19968 20030 19985
rect 20460 19985 21048 20001
rect 20460 19968 20476 19985
rect 20014 19951 20216 19968
rect 19256 19904 20216 19951
rect 20274 19951 20476 19968
rect 21032 19968 21048 19985
rect 21478 19985 22066 20001
rect 21478 19968 21494 19985
rect 21032 19951 21234 19968
rect 20274 19904 21234 19951
rect 21292 19951 21494 19968
rect 22050 19968 22066 19985
rect 22496 19985 23084 20001
rect 22496 19968 22512 19985
rect 22050 19951 22252 19968
rect 21292 19904 22252 19951
rect 22310 19951 22512 19968
rect 23068 19968 23084 19985
rect 23068 19951 23270 19968
rect 22310 19904 23270 19951
rect 24560 19361 25520 19408
rect 24560 19344 24762 19361
rect 24746 19327 24762 19344
rect 25318 19344 25520 19361
rect 25578 19361 26538 19408
rect 25578 19344 25780 19361
rect 25318 19327 25334 19344
rect 24746 19311 25334 19327
rect 25764 19327 25780 19344
rect 26336 19344 26538 19361
rect 26596 19361 27556 19408
rect 26596 19344 26798 19361
rect 26336 19327 26352 19344
rect 25764 19311 26352 19327
rect 26782 19327 26798 19344
rect 27354 19344 27556 19361
rect 27614 19361 28574 19408
rect 27614 19344 27816 19361
rect 27354 19327 27370 19344
rect 26782 19311 27370 19327
rect 27800 19327 27816 19344
rect 28372 19344 28574 19361
rect 28632 19361 29592 19408
rect 28632 19344 28834 19361
rect 28372 19327 28388 19344
rect 27800 19311 28388 19327
rect 28818 19327 28834 19344
rect 29390 19344 29592 19361
rect 29650 19361 30610 19408
rect 29650 19344 29852 19361
rect 29390 19327 29406 19344
rect 28818 19311 29406 19327
rect 29836 19327 29852 19344
rect 30408 19344 30610 19361
rect 30668 19361 31628 19408
rect 30668 19344 30870 19361
rect 30408 19327 30424 19344
rect 29836 19311 30424 19327
rect 30854 19327 30870 19344
rect 31426 19344 31628 19361
rect 31686 19361 32646 19408
rect 31686 19344 31888 19361
rect 31426 19327 31442 19344
rect 30854 19311 31442 19327
rect 31872 19327 31888 19344
rect 32444 19344 32646 19361
rect 32704 19361 33664 19408
rect 32704 19344 32906 19361
rect 32444 19327 32460 19344
rect 31872 19311 32460 19327
rect 32890 19327 32906 19344
rect 33462 19344 33664 19361
rect 33722 19361 34682 19408
rect 33722 19344 33924 19361
rect 33462 19327 33478 19344
rect 32890 19311 33478 19327
rect 33908 19327 33924 19344
rect 34480 19344 34682 19361
rect 34740 19361 35700 19408
rect 34740 19344 34942 19361
rect 34480 19327 34496 19344
rect 33908 19311 34496 19327
rect 34926 19327 34942 19344
rect 35498 19344 35700 19361
rect 35758 19361 36718 19408
rect 35758 19344 35960 19361
rect 35498 19327 35514 19344
rect 34926 19311 35514 19327
rect 35944 19327 35960 19344
rect 36516 19344 36718 19361
rect 36776 19361 37736 19408
rect 36776 19344 36978 19361
rect 36516 19327 36532 19344
rect 35944 19311 36532 19327
rect 36962 19327 36978 19344
rect 37534 19344 37736 19361
rect 37794 19361 38754 19408
rect 37794 19344 37996 19361
rect 37534 19327 37550 19344
rect 36962 19311 37550 19327
rect 37980 19327 37996 19344
rect 38552 19344 38754 19361
rect 38812 19361 39772 19408
rect 38812 19344 39014 19361
rect 38552 19327 38568 19344
rect 37980 19311 38568 19327
rect 38998 19327 39014 19344
rect 39570 19344 39772 19361
rect 39570 19327 39586 19344
rect 38998 19311 39586 19327
rect 19256 19257 20216 19304
rect 19256 19240 19458 19257
rect 19442 19223 19458 19240
rect 20014 19240 20216 19257
rect 20274 19257 21234 19304
rect 20274 19240 20476 19257
rect 20014 19223 20030 19240
rect 19442 19207 20030 19223
rect 20460 19223 20476 19240
rect 21032 19240 21234 19257
rect 21292 19257 22252 19304
rect 21292 19240 21494 19257
rect 21032 19223 21048 19240
rect 20460 19207 21048 19223
rect 21478 19223 21494 19240
rect 22050 19240 22252 19257
rect 22310 19257 23270 19304
rect 22310 19240 22512 19257
rect 22050 19223 22066 19240
rect 21478 19207 22066 19223
rect 22496 19223 22512 19240
rect 23068 19240 23270 19257
rect 23068 19223 23084 19240
rect 22496 19207 23084 19223
rect 19442 18953 20030 18969
rect 19442 18936 19458 18953
rect 19256 18919 19458 18936
rect 20014 18936 20030 18953
rect 20460 18953 21048 18969
rect 20460 18936 20476 18953
rect 20014 18919 20216 18936
rect 19256 18872 20216 18919
rect 20274 18919 20476 18936
rect 21032 18936 21048 18953
rect 21478 18953 22066 18969
rect 21478 18936 21494 18953
rect 21032 18919 21234 18936
rect 20274 18872 21234 18919
rect 21292 18919 21494 18936
rect 22050 18936 22066 18953
rect 22496 18953 23084 18969
rect 22496 18936 22512 18953
rect 22050 18919 22252 18936
rect 21292 18872 22252 18919
rect 22310 18919 22512 18936
rect 23068 18936 23084 18953
rect 23068 18919 23270 18936
rect 22310 18872 23270 18919
rect 24746 18833 25334 18849
rect 24746 18816 24762 18833
rect 24560 18799 24762 18816
rect 25318 18816 25334 18833
rect 25764 18833 26352 18849
rect 25764 18816 25780 18833
rect 25318 18799 25520 18816
rect 24560 18752 25520 18799
rect 25578 18799 25780 18816
rect 26336 18816 26352 18833
rect 26782 18833 27370 18849
rect 26782 18816 26798 18833
rect 26336 18799 26538 18816
rect 25578 18752 26538 18799
rect 26596 18799 26798 18816
rect 27354 18816 27370 18833
rect 27800 18833 28388 18849
rect 27800 18816 27816 18833
rect 27354 18799 27556 18816
rect 26596 18752 27556 18799
rect 27614 18799 27816 18816
rect 28372 18816 28388 18833
rect 28818 18833 29406 18849
rect 28818 18816 28834 18833
rect 28372 18799 28574 18816
rect 27614 18752 28574 18799
rect 28632 18799 28834 18816
rect 29390 18816 29406 18833
rect 29836 18833 30424 18849
rect 29836 18816 29852 18833
rect 29390 18799 29592 18816
rect 28632 18752 29592 18799
rect 29650 18799 29852 18816
rect 30408 18816 30424 18833
rect 30854 18833 31442 18849
rect 30854 18816 30870 18833
rect 30408 18799 30610 18816
rect 29650 18752 30610 18799
rect 30668 18799 30870 18816
rect 31426 18816 31442 18833
rect 31872 18833 32460 18849
rect 31872 18816 31888 18833
rect 31426 18799 31628 18816
rect 30668 18752 31628 18799
rect 31686 18799 31888 18816
rect 32444 18816 32460 18833
rect 32890 18833 33478 18849
rect 32890 18816 32906 18833
rect 32444 18799 32646 18816
rect 31686 18752 32646 18799
rect 32704 18799 32906 18816
rect 33462 18816 33478 18833
rect 33908 18833 34496 18849
rect 33908 18816 33924 18833
rect 33462 18799 33664 18816
rect 32704 18752 33664 18799
rect 33722 18799 33924 18816
rect 34480 18816 34496 18833
rect 34926 18833 35514 18849
rect 34926 18816 34942 18833
rect 34480 18799 34682 18816
rect 33722 18752 34682 18799
rect 34740 18799 34942 18816
rect 35498 18816 35514 18833
rect 35944 18833 36532 18849
rect 35944 18816 35960 18833
rect 35498 18799 35700 18816
rect 34740 18752 35700 18799
rect 35758 18799 35960 18816
rect 36516 18816 36532 18833
rect 36962 18833 37550 18849
rect 36962 18816 36978 18833
rect 36516 18799 36718 18816
rect 35758 18752 36718 18799
rect 36776 18799 36978 18816
rect 37534 18816 37550 18833
rect 37980 18833 38568 18849
rect 37980 18816 37996 18833
rect 37534 18799 37736 18816
rect 36776 18752 37736 18799
rect 37794 18799 37996 18816
rect 38552 18816 38568 18833
rect 38998 18833 39586 18849
rect 38998 18816 39014 18833
rect 38552 18799 38754 18816
rect 37794 18752 38754 18799
rect 38812 18799 39014 18816
rect 39570 18816 39586 18833
rect 39570 18799 39772 18816
rect 38812 18752 39772 18799
rect 19256 18225 20216 18272
rect 19256 18208 19458 18225
rect 19442 18191 19458 18208
rect 20014 18208 20216 18225
rect 20274 18225 21234 18272
rect 20274 18208 20476 18225
rect 20014 18191 20030 18208
rect 19442 18175 20030 18191
rect 20460 18191 20476 18208
rect 21032 18208 21234 18225
rect 21292 18225 22252 18272
rect 21292 18208 21494 18225
rect 21032 18191 21048 18208
rect 20460 18175 21048 18191
rect 21478 18191 21494 18208
rect 22050 18208 22252 18225
rect 22310 18225 23270 18272
rect 22310 18208 22512 18225
rect 22050 18191 22066 18208
rect 21478 18175 22066 18191
rect 22496 18191 22512 18208
rect 23068 18208 23270 18225
rect 23068 18191 23084 18208
rect 22496 18175 23084 18191
rect 24560 18105 25520 18152
rect 24560 18088 24762 18105
rect 24746 18071 24762 18088
rect 25318 18088 25520 18105
rect 25578 18105 26538 18152
rect 25578 18088 25780 18105
rect 25318 18071 25334 18088
rect 24746 18055 25334 18071
rect 25764 18071 25780 18088
rect 26336 18088 26538 18105
rect 26596 18105 27556 18152
rect 26596 18088 26798 18105
rect 26336 18071 26352 18088
rect 25764 18055 26352 18071
rect 26782 18071 26798 18088
rect 27354 18088 27556 18105
rect 27614 18105 28574 18152
rect 27614 18088 27816 18105
rect 27354 18071 27370 18088
rect 26782 18055 27370 18071
rect 27800 18071 27816 18088
rect 28372 18088 28574 18105
rect 28632 18105 29592 18152
rect 28632 18088 28834 18105
rect 28372 18071 28388 18088
rect 27800 18055 28388 18071
rect 28818 18071 28834 18088
rect 29390 18088 29592 18105
rect 29650 18105 30610 18152
rect 29650 18088 29852 18105
rect 29390 18071 29406 18088
rect 28818 18055 29406 18071
rect 29836 18071 29852 18088
rect 30408 18088 30610 18105
rect 30668 18105 31628 18152
rect 30668 18088 30870 18105
rect 30408 18071 30424 18088
rect 29836 18055 30424 18071
rect 30854 18071 30870 18088
rect 31426 18088 31628 18105
rect 31686 18105 32646 18152
rect 31686 18088 31888 18105
rect 31426 18071 31442 18088
rect 30854 18055 31442 18071
rect 31872 18071 31888 18088
rect 32444 18088 32646 18105
rect 32704 18105 33664 18152
rect 32704 18088 32906 18105
rect 32444 18071 32460 18088
rect 31872 18055 32460 18071
rect 32890 18071 32906 18088
rect 33462 18088 33664 18105
rect 33722 18105 34682 18152
rect 33722 18088 33924 18105
rect 33462 18071 33478 18088
rect 32890 18055 33478 18071
rect 33908 18071 33924 18088
rect 34480 18088 34682 18105
rect 34740 18105 35700 18152
rect 34740 18088 34942 18105
rect 34480 18071 34496 18088
rect 33908 18055 34496 18071
rect 34926 18071 34942 18088
rect 35498 18088 35700 18105
rect 35758 18105 36718 18152
rect 35758 18088 35960 18105
rect 35498 18071 35514 18088
rect 34926 18055 35514 18071
rect 35944 18071 35960 18088
rect 36516 18088 36718 18105
rect 36776 18105 37736 18152
rect 36776 18088 36978 18105
rect 36516 18071 36532 18088
rect 35944 18055 36532 18071
rect 36962 18071 36978 18088
rect 37534 18088 37736 18105
rect 37794 18105 38754 18152
rect 37794 18088 37996 18105
rect 37534 18071 37550 18088
rect 36962 18055 37550 18071
rect 37980 18071 37996 18088
rect 38552 18088 38754 18105
rect 38812 18105 39772 18152
rect 38812 18088 39014 18105
rect 38552 18071 38568 18088
rect 37980 18055 38568 18071
rect 38998 18071 39014 18088
rect 39570 18088 39772 18105
rect 39570 18071 39586 18088
rect 38998 18055 39586 18071
rect 19442 17921 20030 17937
rect 19442 17904 19458 17921
rect 19256 17887 19458 17904
rect 20014 17904 20030 17921
rect 20460 17921 21048 17937
rect 20460 17904 20476 17921
rect 20014 17887 20216 17904
rect 19256 17840 20216 17887
rect 20274 17887 20476 17904
rect 21032 17904 21048 17921
rect 21478 17921 22066 17937
rect 21478 17904 21494 17921
rect 21032 17887 21234 17904
rect 20274 17840 21234 17887
rect 21292 17887 21494 17904
rect 22050 17904 22066 17921
rect 22496 17921 23084 17937
rect 22496 17904 22512 17921
rect 22050 17887 22252 17904
rect 21292 17840 22252 17887
rect 22310 17887 22512 17904
rect 23068 17904 23084 17921
rect 23068 17887 23270 17904
rect 22310 17840 23270 17887
rect 24746 17577 25334 17593
rect 24746 17560 24762 17577
rect 24560 17543 24762 17560
rect 25318 17560 25334 17577
rect 25764 17577 26352 17593
rect 25764 17560 25780 17577
rect 25318 17543 25520 17560
rect 24560 17496 25520 17543
rect 25578 17543 25780 17560
rect 26336 17560 26352 17577
rect 26782 17577 27370 17593
rect 26782 17560 26798 17577
rect 26336 17543 26538 17560
rect 25578 17496 26538 17543
rect 26596 17543 26798 17560
rect 27354 17560 27370 17577
rect 27800 17577 28388 17593
rect 27800 17560 27816 17577
rect 27354 17543 27556 17560
rect 26596 17496 27556 17543
rect 27614 17543 27816 17560
rect 28372 17560 28388 17577
rect 28818 17577 29406 17593
rect 28818 17560 28834 17577
rect 28372 17543 28574 17560
rect 27614 17496 28574 17543
rect 28632 17543 28834 17560
rect 29390 17560 29406 17577
rect 29836 17577 30424 17593
rect 29836 17560 29852 17577
rect 29390 17543 29592 17560
rect 28632 17496 29592 17543
rect 29650 17543 29852 17560
rect 30408 17560 30424 17577
rect 30854 17577 31442 17593
rect 30854 17560 30870 17577
rect 30408 17543 30610 17560
rect 29650 17496 30610 17543
rect 30668 17543 30870 17560
rect 31426 17560 31442 17577
rect 31872 17577 32460 17593
rect 31872 17560 31888 17577
rect 31426 17543 31628 17560
rect 30668 17496 31628 17543
rect 31686 17543 31888 17560
rect 32444 17560 32460 17577
rect 32890 17577 33478 17593
rect 32890 17560 32906 17577
rect 32444 17543 32646 17560
rect 31686 17496 32646 17543
rect 32704 17543 32906 17560
rect 33462 17560 33478 17577
rect 33908 17577 34496 17593
rect 33908 17560 33924 17577
rect 33462 17543 33664 17560
rect 32704 17496 33664 17543
rect 33722 17543 33924 17560
rect 34480 17560 34496 17577
rect 34926 17577 35514 17593
rect 34926 17560 34942 17577
rect 34480 17543 34682 17560
rect 33722 17496 34682 17543
rect 34740 17543 34942 17560
rect 35498 17560 35514 17577
rect 35944 17577 36532 17593
rect 35944 17560 35960 17577
rect 35498 17543 35700 17560
rect 34740 17496 35700 17543
rect 35758 17543 35960 17560
rect 36516 17560 36532 17577
rect 36962 17577 37550 17593
rect 36962 17560 36978 17577
rect 36516 17543 36718 17560
rect 35758 17496 36718 17543
rect 36776 17543 36978 17560
rect 37534 17560 37550 17577
rect 37980 17577 38568 17593
rect 37980 17560 37996 17577
rect 37534 17543 37736 17560
rect 36776 17496 37736 17543
rect 37794 17543 37996 17560
rect 38552 17560 38568 17577
rect 38998 17577 39586 17593
rect 38998 17560 39014 17577
rect 38552 17543 38754 17560
rect 37794 17496 38754 17543
rect 38812 17543 39014 17560
rect 39570 17560 39586 17577
rect 39570 17543 39772 17560
rect 38812 17496 39772 17543
rect 19256 17193 20216 17240
rect 19256 17176 19458 17193
rect 19442 17159 19458 17176
rect 20014 17176 20216 17193
rect 20274 17193 21234 17240
rect 20274 17176 20476 17193
rect 20014 17159 20030 17176
rect 19442 17143 20030 17159
rect 20460 17159 20476 17176
rect 21032 17176 21234 17193
rect 21292 17193 22252 17240
rect 21292 17176 21494 17193
rect 21032 17159 21048 17176
rect 20460 17143 21048 17159
rect 21478 17159 21494 17176
rect 22050 17176 22252 17193
rect 22310 17193 23270 17240
rect 22310 17176 22512 17193
rect 22050 17159 22066 17176
rect 21478 17143 22066 17159
rect 22496 17159 22512 17176
rect 23068 17176 23270 17193
rect 23068 17159 23084 17176
rect 22496 17143 23084 17159
rect 19442 16889 20030 16905
rect 19442 16872 19458 16889
rect 19256 16855 19458 16872
rect 20014 16872 20030 16889
rect 20460 16889 21048 16905
rect 20460 16872 20476 16889
rect 20014 16855 20216 16872
rect 19256 16808 20216 16855
rect 20274 16855 20476 16872
rect 21032 16872 21048 16889
rect 21478 16889 22066 16905
rect 21478 16872 21494 16889
rect 21032 16855 21234 16872
rect 20274 16808 21234 16855
rect 21292 16855 21494 16872
rect 22050 16872 22066 16889
rect 22496 16889 23084 16905
rect 22496 16872 22512 16889
rect 22050 16855 22252 16872
rect 21292 16808 22252 16855
rect 22310 16855 22512 16872
rect 23068 16872 23084 16889
rect 23068 16855 23270 16872
rect 22310 16808 23270 16855
rect 24560 16849 25520 16896
rect 24560 16832 24762 16849
rect 24746 16815 24762 16832
rect 25318 16832 25520 16849
rect 25578 16849 26538 16896
rect 25578 16832 25780 16849
rect 25318 16815 25334 16832
rect 24746 16799 25334 16815
rect 25764 16815 25780 16832
rect 26336 16832 26538 16849
rect 26596 16849 27556 16896
rect 26596 16832 26798 16849
rect 26336 16815 26352 16832
rect 25764 16799 26352 16815
rect 26782 16815 26798 16832
rect 27354 16832 27556 16849
rect 27614 16849 28574 16896
rect 27614 16832 27816 16849
rect 27354 16815 27370 16832
rect 26782 16799 27370 16815
rect 27800 16815 27816 16832
rect 28372 16832 28574 16849
rect 28632 16849 29592 16896
rect 28632 16832 28834 16849
rect 28372 16815 28388 16832
rect 27800 16799 28388 16815
rect 28818 16815 28834 16832
rect 29390 16832 29592 16849
rect 29650 16849 30610 16896
rect 29650 16832 29852 16849
rect 29390 16815 29406 16832
rect 28818 16799 29406 16815
rect 29836 16815 29852 16832
rect 30408 16832 30610 16849
rect 30668 16849 31628 16896
rect 30668 16832 30870 16849
rect 30408 16815 30424 16832
rect 29836 16799 30424 16815
rect 30854 16815 30870 16832
rect 31426 16832 31628 16849
rect 31686 16849 32646 16896
rect 31686 16832 31888 16849
rect 31426 16815 31442 16832
rect 30854 16799 31442 16815
rect 31872 16815 31888 16832
rect 32444 16832 32646 16849
rect 32704 16849 33664 16896
rect 32704 16832 32906 16849
rect 32444 16815 32460 16832
rect 31872 16799 32460 16815
rect 32890 16815 32906 16832
rect 33462 16832 33664 16849
rect 33722 16849 34682 16896
rect 33722 16832 33924 16849
rect 33462 16815 33478 16832
rect 32890 16799 33478 16815
rect 33908 16815 33924 16832
rect 34480 16832 34682 16849
rect 34740 16849 35700 16896
rect 34740 16832 34942 16849
rect 34480 16815 34496 16832
rect 33908 16799 34496 16815
rect 34926 16815 34942 16832
rect 35498 16832 35700 16849
rect 35758 16849 36718 16896
rect 35758 16832 35960 16849
rect 35498 16815 35514 16832
rect 34926 16799 35514 16815
rect 35944 16815 35960 16832
rect 36516 16832 36718 16849
rect 36776 16849 37736 16896
rect 36776 16832 36978 16849
rect 36516 16815 36532 16832
rect 35944 16799 36532 16815
rect 36962 16815 36978 16832
rect 37534 16832 37736 16849
rect 37794 16849 38754 16896
rect 37794 16832 37996 16849
rect 37534 16815 37550 16832
rect 36962 16799 37550 16815
rect 37980 16815 37996 16832
rect 38552 16832 38754 16849
rect 38812 16849 39772 16896
rect 38812 16832 39014 16849
rect 38552 16815 38568 16832
rect 37980 16799 38568 16815
rect 38998 16815 39014 16832
rect 39570 16832 39772 16849
rect 39570 16815 39586 16832
rect 38998 16799 39586 16815
rect 24746 16321 25334 16337
rect 24746 16304 24762 16321
rect 24560 16287 24762 16304
rect 25318 16304 25334 16321
rect 25764 16321 26352 16337
rect 25764 16304 25780 16321
rect 25318 16287 25520 16304
rect 24560 16240 25520 16287
rect 25578 16287 25780 16304
rect 26336 16304 26352 16321
rect 26782 16321 27370 16337
rect 26782 16304 26798 16321
rect 26336 16287 26538 16304
rect 25578 16240 26538 16287
rect 26596 16287 26798 16304
rect 27354 16304 27370 16321
rect 27800 16321 28388 16337
rect 27800 16304 27816 16321
rect 27354 16287 27556 16304
rect 26596 16240 27556 16287
rect 27614 16287 27816 16304
rect 28372 16304 28388 16321
rect 28818 16321 29406 16337
rect 28818 16304 28834 16321
rect 28372 16287 28574 16304
rect 27614 16240 28574 16287
rect 28632 16287 28834 16304
rect 29390 16304 29406 16321
rect 29836 16321 30424 16337
rect 29836 16304 29852 16321
rect 29390 16287 29592 16304
rect 28632 16240 29592 16287
rect 29650 16287 29852 16304
rect 30408 16304 30424 16321
rect 30854 16321 31442 16337
rect 30854 16304 30870 16321
rect 30408 16287 30610 16304
rect 29650 16240 30610 16287
rect 30668 16287 30870 16304
rect 31426 16304 31442 16321
rect 31872 16321 32460 16337
rect 31872 16304 31888 16321
rect 31426 16287 31628 16304
rect 30668 16240 31628 16287
rect 31686 16287 31888 16304
rect 32444 16304 32460 16321
rect 32890 16321 33478 16337
rect 32890 16304 32906 16321
rect 32444 16287 32646 16304
rect 31686 16240 32646 16287
rect 32704 16287 32906 16304
rect 33462 16304 33478 16321
rect 33908 16321 34496 16337
rect 33908 16304 33924 16321
rect 33462 16287 33664 16304
rect 32704 16240 33664 16287
rect 33722 16287 33924 16304
rect 34480 16304 34496 16321
rect 34926 16321 35514 16337
rect 34926 16304 34942 16321
rect 34480 16287 34682 16304
rect 33722 16240 34682 16287
rect 34740 16287 34942 16304
rect 35498 16304 35514 16321
rect 35944 16321 36532 16337
rect 35944 16304 35960 16321
rect 35498 16287 35700 16304
rect 34740 16240 35700 16287
rect 35758 16287 35960 16304
rect 36516 16304 36532 16321
rect 36962 16321 37550 16337
rect 36962 16304 36978 16321
rect 36516 16287 36718 16304
rect 35758 16240 36718 16287
rect 36776 16287 36978 16304
rect 37534 16304 37550 16321
rect 37980 16321 38568 16337
rect 37980 16304 37996 16321
rect 37534 16287 37736 16304
rect 36776 16240 37736 16287
rect 37794 16287 37996 16304
rect 38552 16304 38568 16321
rect 38998 16321 39586 16337
rect 38998 16304 39014 16321
rect 38552 16287 38754 16304
rect 37794 16240 38754 16287
rect 38812 16287 39014 16304
rect 39570 16304 39586 16321
rect 39570 16287 39772 16304
rect 38812 16240 39772 16287
rect 19256 16161 20216 16208
rect 19256 16144 19458 16161
rect 19442 16127 19458 16144
rect 20014 16144 20216 16161
rect 20274 16161 21234 16208
rect 20274 16144 20476 16161
rect 20014 16127 20030 16144
rect 19442 16111 20030 16127
rect 20460 16127 20476 16144
rect 21032 16144 21234 16161
rect 21292 16161 22252 16208
rect 21292 16144 21494 16161
rect 21032 16127 21048 16144
rect 20460 16111 21048 16127
rect 21478 16127 21494 16144
rect 22050 16144 22252 16161
rect 22310 16161 23270 16208
rect 22310 16144 22512 16161
rect 22050 16127 22066 16144
rect 21478 16111 22066 16127
rect 22496 16127 22512 16144
rect 23068 16144 23270 16161
rect 23068 16127 23084 16144
rect 22496 16111 23084 16127
rect 24560 15593 25520 15640
rect 24560 15576 24762 15593
rect 24746 15559 24762 15576
rect 25318 15576 25520 15593
rect 25578 15593 26538 15640
rect 25578 15576 25780 15593
rect 25318 15559 25334 15576
rect 24746 15543 25334 15559
rect 25764 15559 25780 15576
rect 26336 15576 26538 15593
rect 26596 15593 27556 15640
rect 26596 15576 26798 15593
rect 26336 15559 26352 15576
rect 25764 15543 26352 15559
rect 26782 15559 26798 15576
rect 27354 15576 27556 15593
rect 27614 15593 28574 15640
rect 27614 15576 27816 15593
rect 27354 15559 27370 15576
rect 26782 15543 27370 15559
rect 27800 15559 27816 15576
rect 28372 15576 28574 15593
rect 28632 15593 29592 15640
rect 28632 15576 28834 15593
rect 28372 15559 28388 15576
rect 27800 15543 28388 15559
rect 28818 15559 28834 15576
rect 29390 15576 29592 15593
rect 29650 15593 30610 15640
rect 29650 15576 29852 15593
rect 29390 15559 29406 15576
rect 28818 15543 29406 15559
rect 29836 15559 29852 15576
rect 30408 15576 30610 15593
rect 30668 15593 31628 15640
rect 30668 15576 30870 15593
rect 30408 15559 30424 15576
rect 29836 15543 30424 15559
rect 30854 15559 30870 15576
rect 31426 15576 31628 15593
rect 31686 15593 32646 15640
rect 31686 15576 31888 15593
rect 31426 15559 31442 15576
rect 30854 15543 31442 15559
rect 31872 15559 31888 15576
rect 32444 15576 32646 15593
rect 32704 15593 33664 15640
rect 32704 15576 32906 15593
rect 32444 15559 32460 15576
rect 31872 15543 32460 15559
rect 32890 15559 32906 15576
rect 33462 15576 33664 15593
rect 33722 15593 34682 15640
rect 33722 15576 33924 15593
rect 33462 15559 33478 15576
rect 32890 15543 33478 15559
rect 33908 15559 33924 15576
rect 34480 15576 34682 15593
rect 34740 15593 35700 15640
rect 34740 15576 34942 15593
rect 34480 15559 34496 15576
rect 33908 15543 34496 15559
rect 34926 15559 34942 15576
rect 35498 15576 35700 15593
rect 35758 15593 36718 15640
rect 35758 15576 35960 15593
rect 35498 15559 35514 15576
rect 34926 15543 35514 15559
rect 35944 15559 35960 15576
rect 36516 15576 36718 15593
rect 36776 15593 37736 15640
rect 36776 15576 36978 15593
rect 36516 15559 36532 15576
rect 35944 15543 36532 15559
rect 36962 15559 36978 15576
rect 37534 15576 37736 15593
rect 37794 15593 38754 15640
rect 37794 15576 37996 15593
rect 37534 15559 37550 15576
rect 36962 15543 37550 15559
rect 37980 15559 37996 15576
rect 38552 15576 38754 15593
rect 38812 15593 39772 15640
rect 38812 15576 39014 15593
rect 38552 15559 38568 15576
rect 37980 15543 38568 15559
rect 38998 15559 39014 15576
rect 39570 15576 39772 15593
rect 39570 15559 39586 15576
rect 38998 15543 39586 15559
rect 366 514 498 530
rect 366 497 382 514
rect 332 480 382 497
rect 482 497 498 514
rect 624 514 756 530
rect 624 497 640 514
rect 482 480 532 497
rect 332 442 532 480
rect 590 480 640 497
rect 740 497 756 514
rect 882 514 1014 530
rect 882 497 898 514
rect 740 480 790 497
rect 590 442 790 480
rect 848 480 898 497
rect 998 497 1014 514
rect 1140 514 1272 530
rect 1140 497 1156 514
rect 998 480 1048 497
rect 848 442 1048 480
rect 1106 480 1156 497
rect 1256 497 1272 514
rect 1398 514 1530 530
rect 1398 497 1414 514
rect 1256 480 1306 497
rect 1106 442 1306 480
rect 1364 480 1414 497
rect 1514 497 1530 514
rect 1656 514 1788 530
rect 1656 497 1672 514
rect 1514 480 1564 497
rect 1364 442 1564 480
rect 1622 480 1672 497
rect 1772 497 1788 514
rect 1914 514 2046 530
rect 1914 497 1930 514
rect 1772 480 1822 497
rect 1622 442 1822 480
rect 1880 480 1930 497
rect 2030 497 2046 514
rect 2172 514 2304 530
rect 2172 497 2188 514
rect 2030 480 2080 497
rect 1880 442 2080 480
rect 2138 480 2188 497
rect 2288 497 2304 514
rect 2430 514 2562 530
rect 2430 497 2446 514
rect 2288 480 2338 497
rect 2138 442 2338 480
rect 2396 480 2446 497
rect 2546 497 2562 514
rect 2688 514 2820 530
rect 2688 497 2704 514
rect 2546 480 2596 497
rect 2396 442 2596 480
rect 2654 480 2704 497
rect 2804 497 2820 514
rect 2946 514 3078 530
rect 2946 497 2962 514
rect 2804 480 2854 497
rect 2654 442 2854 480
rect 2912 480 2962 497
rect 3062 497 3078 514
rect 3204 514 3336 530
rect 3204 497 3220 514
rect 3062 480 3112 497
rect 2912 442 3112 480
rect 3170 480 3220 497
rect 3320 497 3336 514
rect 3462 514 3594 530
rect 3462 497 3478 514
rect 3320 480 3370 497
rect 3170 442 3370 480
rect 3428 480 3478 497
rect 3578 497 3594 514
rect 3720 514 3852 530
rect 3720 497 3736 514
rect 3578 480 3628 497
rect 3428 442 3628 480
rect 3686 480 3736 497
rect 3836 497 3852 514
rect 3836 480 3886 497
rect 3686 442 3886 480
rect 332 4 532 42
rect 332 -13 382 4
rect 366 -30 382 -13
rect 482 -13 532 4
rect 590 4 790 42
rect 590 -13 640 4
rect 482 -30 498 -13
rect 366 -46 498 -30
rect 624 -30 640 -13
rect 740 -13 790 4
rect 848 4 1048 42
rect 848 -13 898 4
rect 740 -30 756 -13
rect 624 -46 756 -30
rect 882 -30 898 -13
rect 998 -13 1048 4
rect 1106 4 1306 42
rect 1106 -13 1156 4
rect 998 -30 1014 -13
rect 882 -46 1014 -30
rect 1140 -30 1156 -13
rect 1256 -13 1306 4
rect 1364 4 1564 42
rect 1364 -13 1414 4
rect 1256 -30 1272 -13
rect 1140 -46 1272 -30
rect 1398 -30 1414 -13
rect 1514 -13 1564 4
rect 1622 4 1822 42
rect 1622 -13 1672 4
rect 1514 -30 1530 -13
rect 1398 -46 1530 -30
rect 1656 -30 1672 -13
rect 1772 -13 1822 4
rect 1880 4 2080 42
rect 1880 -13 1930 4
rect 1772 -30 1788 -13
rect 1656 -46 1788 -30
rect 1914 -30 1930 -13
rect 2030 -13 2080 4
rect 2138 4 2338 42
rect 2138 -13 2188 4
rect 2030 -30 2046 -13
rect 1914 -46 2046 -30
rect 2172 -30 2188 -13
rect 2288 -13 2338 4
rect 2396 4 2596 42
rect 2396 -13 2446 4
rect 2288 -30 2304 -13
rect 2172 -46 2304 -30
rect 2430 -30 2446 -13
rect 2546 -13 2596 4
rect 2654 4 2854 42
rect 2654 -13 2704 4
rect 2546 -30 2562 -13
rect 2430 -46 2562 -30
rect 2688 -30 2704 -13
rect 2804 -13 2854 4
rect 2912 4 3112 42
rect 2912 -13 2962 4
rect 2804 -30 2820 -13
rect 2688 -46 2820 -30
rect 2946 -30 2962 -13
rect 3062 -13 3112 4
rect 3170 4 3370 42
rect 3170 -13 3220 4
rect 3062 -30 3078 -13
rect 2946 -46 3078 -30
rect 3204 -30 3220 -13
rect 3320 -13 3370 4
rect 3428 4 3628 42
rect 3428 -13 3478 4
rect 3320 -30 3336 -13
rect 3204 -46 3336 -30
rect 3462 -30 3478 -13
rect 3578 -13 3628 4
rect 3686 4 3886 42
rect 3686 -13 3736 4
rect 3578 -30 3594 -13
rect 3462 -46 3594 -30
rect 3720 -30 3736 -13
rect 3836 -13 3886 4
rect 3836 -30 3852 -13
rect 3720 -46 3852 -30
rect 366 -486 498 -470
rect 366 -503 382 -486
rect 332 -520 382 -503
rect 482 -503 498 -486
rect 624 -486 756 -470
rect 624 -503 640 -486
rect 482 -520 532 -503
rect 332 -558 532 -520
rect 590 -520 640 -503
rect 740 -503 756 -486
rect 882 -486 1014 -470
rect 882 -503 898 -486
rect 740 -520 790 -503
rect 590 -558 790 -520
rect 848 -520 898 -503
rect 998 -503 1014 -486
rect 1140 -486 1272 -470
rect 1140 -503 1156 -486
rect 998 -520 1048 -503
rect 848 -558 1048 -520
rect 1106 -520 1156 -503
rect 1256 -503 1272 -486
rect 1398 -486 1530 -470
rect 1398 -503 1414 -486
rect 1256 -520 1306 -503
rect 1106 -558 1306 -520
rect 1364 -520 1414 -503
rect 1514 -503 1530 -486
rect 1656 -486 1788 -470
rect 1656 -503 1672 -486
rect 1514 -520 1564 -503
rect 1364 -558 1564 -520
rect 1622 -520 1672 -503
rect 1772 -503 1788 -486
rect 1914 -486 2046 -470
rect 1914 -503 1930 -486
rect 1772 -520 1822 -503
rect 1622 -558 1822 -520
rect 1880 -520 1930 -503
rect 2030 -503 2046 -486
rect 2172 -486 2304 -470
rect 2172 -503 2188 -486
rect 2030 -520 2080 -503
rect 1880 -558 2080 -520
rect 2138 -520 2188 -503
rect 2288 -503 2304 -486
rect 2430 -486 2562 -470
rect 2430 -503 2446 -486
rect 2288 -520 2338 -503
rect 2138 -558 2338 -520
rect 2396 -520 2446 -503
rect 2546 -503 2562 -486
rect 2688 -486 2820 -470
rect 2688 -503 2704 -486
rect 2546 -520 2596 -503
rect 2396 -558 2596 -520
rect 2654 -520 2704 -503
rect 2804 -503 2820 -486
rect 2946 -486 3078 -470
rect 2946 -503 2962 -486
rect 2804 -520 2854 -503
rect 2654 -558 2854 -520
rect 2912 -520 2962 -503
rect 3062 -503 3078 -486
rect 3204 -486 3336 -470
rect 3204 -503 3220 -486
rect 3062 -520 3112 -503
rect 2912 -558 3112 -520
rect 3170 -520 3220 -503
rect 3320 -503 3336 -486
rect 3462 -486 3594 -470
rect 3462 -503 3478 -486
rect 3320 -520 3370 -503
rect 3170 -558 3370 -520
rect 3428 -520 3478 -503
rect 3578 -503 3594 -486
rect 3720 -486 3852 -470
rect 3720 -503 3736 -486
rect 3578 -520 3628 -503
rect 3428 -558 3628 -520
rect 3686 -520 3736 -503
rect 3836 -503 3852 -486
rect 3836 -520 3886 -503
rect 3686 -558 3886 -520
rect 332 -996 532 -958
rect 332 -1013 382 -996
rect 366 -1030 382 -1013
rect 482 -1013 532 -996
rect 590 -996 790 -958
rect 590 -1013 640 -996
rect 482 -1030 498 -1013
rect 366 -1046 498 -1030
rect 624 -1030 640 -1013
rect 740 -1013 790 -996
rect 848 -996 1048 -958
rect 848 -1013 898 -996
rect 740 -1030 756 -1013
rect 624 -1046 756 -1030
rect 882 -1030 898 -1013
rect 998 -1013 1048 -996
rect 1106 -996 1306 -958
rect 1106 -1013 1156 -996
rect 998 -1030 1014 -1013
rect 882 -1046 1014 -1030
rect 1140 -1030 1156 -1013
rect 1256 -1013 1306 -996
rect 1364 -996 1564 -958
rect 1364 -1013 1414 -996
rect 1256 -1030 1272 -1013
rect 1140 -1046 1272 -1030
rect 1398 -1030 1414 -1013
rect 1514 -1013 1564 -996
rect 1622 -996 1822 -958
rect 1622 -1013 1672 -996
rect 1514 -1030 1530 -1013
rect 1398 -1046 1530 -1030
rect 1656 -1030 1672 -1013
rect 1772 -1013 1822 -996
rect 1880 -996 2080 -958
rect 1880 -1013 1930 -996
rect 1772 -1030 1788 -1013
rect 1656 -1046 1788 -1030
rect 1914 -1030 1930 -1013
rect 2030 -1013 2080 -996
rect 2138 -996 2338 -958
rect 2138 -1013 2188 -996
rect 2030 -1030 2046 -1013
rect 1914 -1046 2046 -1030
rect 2172 -1030 2188 -1013
rect 2288 -1013 2338 -996
rect 2396 -996 2596 -958
rect 2396 -1013 2446 -996
rect 2288 -1030 2304 -1013
rect 2172 -1046 2304 -1030
rect 2430 -1030 2446 -1013
rect 2546 -1013 2596 -996
rect 2654 -996 2854 -958
rect 2654 -1013 2704 -996
rect 2546 -1030 2562 -1013
rect 2430 -1046 2562 -1030
rect 2688 -1030 2704 -1013
rect 2804 -1013 2854 -996
rect 2912 -996 3112 -958
rect 2912 -1013 2962 -996
rect 2804 -1030 2820 -1013
rect 2688 -1046 2820 -1030
rect 2946 -1030 2962 -1013
rect 3062 -1013 3112 -996
rect 3170 -996 3370 -958
rect 3170 -1013 3220 -996
rect 3062 -1030 3078 -1013
rect 2946 -1046 3078 -1030
rect 3204 -1030 3220 -1013
rect 3320 -1013 3370 -996
rect 3428 -996 3628 -958
rect 3428 -1013 3478 -996
rect 3320 -1030 3336 -1013
rect 3204 -1046 3336 -1030
rect 3462 -1030 3478 -1013
rect 3578 -1013 3628 -996
rect 3686 -996 3886 -958
rect 3686 -1013 3736 -996
rect 3578 -1030 3594 -1013
rect 3462 -1046 3594 -1030
rect 3720 -1030 3736 -1013
rect 3836 -1013 3886 -996
rect 3836 -1030 3852 -1013
rect 3720 -1046 3852 -1030
rect 19854 13116 20442 13132
rect 19854 13099 19870 13116
rect 19668 13082 19870 13099
rect 20426 13099 20442 13116
rect 20872 13116 21460 13132
rect 20872 13099 20888 13116
rect 20426 13082 20628 13099
rect 19668 13044 20628 13082
rect 20686 13082 20888 13099
rect 21444 13099 21460 13116
rect 21890 13116 22478 13132
rect 21890 13099 21906 13116
rect 21444 13082 21646 13099
rect 20686 13044 21646 13082
rect 21704 13082 21906 13099
rect 22462 13099 22478 13116
rect 22908 13116 23496 13132
rect 22908 13099 22924 13116
rect 22462 13082 22664 13099
rect 21704 13044 22664 13082
rect 22722 13082 22924 13099
rect 23480 13099 23496 13116
rect 23926 13116 24514 13132
rect 23926 13099 23942 13116
rect 23480 13082 23682 13099
rect 22722 13044 23682 13082
rect 23740 13082 23942 13099
rect 24498 13099 24514 13116
rect 24944 13116 25532 13132
rect 24944 13099 24960 13116
rect 24498 13082 24700 13099
rect 23740 13044 24700 13082
rect 24758 13082 24960 13099
rect 25516 13099 25532 13116
rect 25962 13116 26550 13132
rect 25962 13099 25978 13116
rect 25516 13082 25718 13099
rect 24758 13044 25718 13082
rect 25776 13082 25978 13099
rect 26534 13099 26550 13116
rect 26980 13116 27568 13132
rect 26980 13099 26996 13116
rect 26534 13082 26736 13099
rect 25776 13044 26736 13082
rect 26794 13082 26996 13099
rect 27552 13099 27568 13116
rect 27998 13116 28586 13132
rect 27998 13099 28014 13116
rect 27552 13082 27754 13099
rect 26794 13044 27754 13082
rect 27812 13082 28014 13099
rect 28570 13099 28586 13116
rect 29016 13116 29604 13132
rect 29016 13099 29032 13116
rect 28570 13082 28772 13099
rect 27812 13044 28772 13082
rect 28830 13082 29032 13099
rect 29588 13099 29604 13116
rect 30034 13116 30622 13132
rect 30034 13099 30050 13116
rect 29588 13082 29790 13099
rect 28830 13044 29790 13082
rect 29848 13082 30050 13099
rect 30606 13099 30622 13116
rect 31052 13116 31640 13132
rect 31052 13099 31068 13116
rect 30606 13082 30808 13099
rect 29848 13044 30808 13082
rect 30866 13082 31068 13099
rect 31624 13099 31640 13116
rect 32070 13116 32658 13132
rect 32070 13099 32086 13116
rect 31624 13082 31826 13099
rect 30866 13044 31826 13082
rect 31884 13082 32086 13099
rect 32642 13099 32658 13116
rect 33088 13116 33676 13132
rect 33088 13099 33104 13116
rect 32642 13082 32844 13099
rect 31884 13044 32844 13082
rect 32902 13082 33104 13099
rect 33660 13099 33676 13116
rect 34106 13116 34694 13132
rect 34106 13099 34122 13116
rect 33660 13082 33862 13099
rect 32902 13044 33862 13082
rect 33920 13082 34122 13099
rect 34678 13099 34694 13116
rect 35124 13116 35712 13132
rect 35124 13099 35140 13116
rect 34678 13082 34880 13099
rect 33920 13044 34880 13082
rect 34938 13082 35140 13099
rect 35696 13099 35712 13116
rect 36142 13116 36730 13132
rect 36142 13099 36158 13116
rect 35696 13082 35898 13099
rect 34938 13044 35898 13082
rect 35956 13082 36158 13099
rect 36714 13099 36730 13116
rect 37160 13116 37748 13132
rect 37160 13099 37176 13116
rect 36714 13082 36916 13099
rect 35956 13044 36916 13082
rect 36974 13082 37176 13099
rect 37732 13099 37748 13116
rect 38178 13116 38766 13132
rect 38178 13099 38194 13116
rect 37732 13082 37934 13099
rect 36974 13044 37934 13082
rect 37992 13082 38194 13099
rect 38750 13099 38766 13116
rect 39196 13116 39784 13132
rect 39196 13099 39212 13116
rect 38750 13082 38952 13099
rect 37992 13044 38952 13082
rect 39010 13082 39212 13099
rect 39768 13099 39784 13116
rect 39768 13082 39970 13099
rect 39010 13044 39970 13082
rect 8088 12640 8676 12656
rect 8088 12623 8104 12640
rect 7902 12606 8104 12623
rect 8660 12623 8676 12640
rect 9106 12640 9694 12656
rect 9106 12623 9122 12640
rect 8660 12606 8862 12623
rect 7902 12568 8862 12606
rect 8920 12606 9122 12623
rect 9678 12623 9694 12640
rect 10124 12640 10712 12656
rect 10124 12623 10140 12640
rect 9678 12606 9880 12623
rect 8920 12568 9880 12606
rect 9938 12606 10140 12623
rect 10696 12623 10712 12640
rect 11142 12640 11730 12656
rect 11142 12623 11158 12640
rect 10696 12606 10898 12623
rect 9938 12568 10898 12606
rect 10956 12606 11158 12623
rect 11714 12623 11730 12640
rect 12160 12640 12748 12656
rect 12160 12623 12176 12640
rect 11714 12606 11916 12623
rect 10956 12568 11916 12606
rect 11974 12606 12176 12623
rect 12732 12623 12748 12640
rect 13178 12640 13766 12656
rect 13178 12623 13194 12640
rect 12732 12606 12934 12623
rect 11974 12568 12934 12606
rect 12992 12606 13194 12623
rect 13750 12623 13766 12640
rect 14196 12640 14784 12656
rect 14196 12623 14212 12640
rect 13750 12606 13952 12623
rect 12992 12568 13952 12606
rect 14010 12606 14212 12623
rect 14768 12623 14784 12640
rect 15214 12640 15802 12656
rect 15214 12623 15230 12640
rect 14768 12606 14970 12623
rect 14010 12568 14970 12606
rect 15028 12606 15230 12623
rect 15786 12623 15802 12640
rect 16232 12640 16820 12656
rect 16232 12623 16248 12640
rect 15786 12606 15988 12623
rect 15028 12568 15988 12606
rect 16046 12606 16248 12623
rect 16804 12623 16820 12640
rect 16804 12606 17006 12623
rect 16046 12568 17006 12606
rect 19668 12406 20628 12444
rect 19668 12389 19870 12406
rect 19854 12372 19870 12389
rect 20426 12389 20628 12406
rect 20686 12406 21646 12444
rect 20686 12389 20888 12406
rect 20426 12372 20442 12389
rect 19854 12356 20442 12372
rect 20872 12372 20888 12389
rect 21444 12389 21646 12406
rect 21704 12406 22664 12444
rect 21704 12389 21906 12406
rect 21444 12372 21460 12389
rect 20872 12356 21460 12372
rect 21890 12372 21906 12389
rect 22462 12389 22664 12406
rect 22722 12406 23682 12444
rect 22722 12389 22924 12406
rect 22462 12372 22478 12389
rect 21890 12356 22478 12372
rect 22908 12372 22924 12389
rect 23480 12389 23682 12406
rect 23740 12406 24700 12444
rect 23740 12389 23942 12406
rect 23480 12372 23496 12389
rect 22908 12356 23496 12372
rect 23926 12372 23942 12389
rect 24498 12389 24700 12406
rect 24758 12406 25718 12444
rect 24758 12389 24960 12406
rect 24498 12372 24514 12389
rect 23926 12356 24514 12372
rect 24944 12372 24960 12389
rect 25516 12389 25718 12406
rect 25776 12406 26736 12444
rect 25776 12389 25978 12406
rect 25516 12372 25532 12389
rect 24944 12356 25532 12372
rect 25962 12372 25978 12389
rect 26534 12389 26736 12406
rect 26794 12406 27754 12444
rect 26794 12389 26996 12406
rect 26534 12372 26550 12389
rect 25962 12356 26550 12372
rect 26980 12372 26996 12389
rect 27552 12389 27754 12406
rect 27812 12406 28772 12444
rect 27812 12389 28014 12406
rect 27552 12372 27568 12389
rect 26980 12356 27568 12372
rect 27998 12372 28014 12389
rect 28570 12389 28772 12406
rect 28830 12406 29790 12444
rect 28830 12389 29032 12406
rect 28570 12372 28586 12389
rect 27998 12356 28586 12372
rect 29016 12372 29032 12389
rect 29588 12389 29790 12406
rect 29848 12406 30808 12444
rect 29848 12389 30050 12406
rect 29588 12372 29604 12389
rect 29016 12356 29604 12372
rect 30034 12372 30050 12389
rect 30606 12389 30808 12406
rect 30866 12406 31826 12444
rect 30866 12389 31068 12406
rect 30606 12372 30622 12389
rect 30034 12356 30622 12372
rect 31052 12372 31068 12389
rect 31624 12389 31826 12406
rect 31884 12406 32844 12444
rect 31884 12389 32086 12406
rect 31624 12372 31640 12389
rect 31052 12356 31640 12372
rect 32070 12372 32086 12389
rect 32642 12389 32844 12406
rect 32902 12406 33862 12444
rect 32902 12389 33104 12406
rect 32642 12372 32658 12389
rect 32070 12356 32658 12372
rect 33088 12372 33104 12389
rect 33660 12389 33862 12406
rect 33920 12406 34880 12444
rect 33920 12389 34122 12406
rect 33660 12372 33676 12389
rect 33088 12356 33676 12372
rect 34106 12372 34122 12389
rect 34678 12389 34880 12406
rect 34938 12406 35898 12444
rect 34938 12389 35140 12406
rect 34678 12372 34694 12389
rect 34106 12356 34694 12372
rect 35124 12372 35140 12389
rect 35696 12389 35898 12406
rect 35956 12406 36916 12444
rect 35956 12389 36158 12406
rect 35696 12372 35712 12389
rect 35124 12356 35712 12372
rect 36142 12372 36158 12389
rect 36714 12389 36916 12406
rect 36974 12406 37934 12444
rect 36974 12389 37176 12406
rect 36714 12372 36730 12389
rect 36142 12356 36730 12372
rect 37160 12372 37176 12389
rect 37732 12389 37934 12406
rect 37992 12406 38952 12444
rect 37992 12389 38194 12406
rect 37732 12372 37748 12389
rect 37160 12356 37748 12372
rect 38178 12372 38194 12389
rect 38750 12389 38952 12406
rect 39010 12406 39970 12444
rect 39010 12389 39212 12406
rect 38750 12372 38766 12389
rect 38178 12356 38766 12372
rect 39196 12372 39212 12389
rect 39768 12389 39970 12406
rect 39768 12372 39784 12389
rect 39196 12356 39784 12372
rect 19854 12298 20442 12314
rect 19854 12281 19870 12298
rect 19668 12264 19870 12281
rect 20426 12281 20442 12298
rect 20872 12298 21460 12314
rect 20872 12281 20888 12298
rect 20426 12264 20628 12281
rect 19668 12226 20628 12264
rect 20686 12264 20888 12281
rect 21444 12281 21460 12298
rect 21890 12298 22478 12314
rect 21890 12281 21906 12298
rect 21444 12264 21646 12281
rect 20686 12226 21646 12264
rect 21704 12264 21906 12281
rect 22462 12281 22478 12298
rect 22908 12298 23496 12314
rect 22908 12281 22924 12298
rect 22462 12264 22664 12281
rect 21704 12226 22664 12264
rect 22722 12264 22924 12281
rect 23480 12281 23496 12298
rect 23926 12298 24514 12314
rect 23926 12281 23942 12298
rect 23480 12264 23682 12281
rect 22722 12226 23682 12264
rect 23740 12264 23942 12281
rect 24498 12281 24514 12298
rect 24944 12298 25532 12314
rect 24944 12281 24960 12298
rect 24498 12264 24700 12281
rect 23740 12226 24700 12264
rect 24758 12264 24960 12281
rect 25516 12281 25532 12298
rect 25962 12298 26550 12314
rect 25962 12281 25978 12298
rect 25516 12264 25718 12281
rect 24758 12226 25718 12264
rect 25776 12264 25978 12281
rect 26534 12281 26550 12298
rect 26980 12298 27568 12314
rect 26980 12281 26996 12298
rect 26534 12264 26736 12281
rect 25776 12226 26736 12264
rect 26794 12264 26996 12281
rect 27552 12281 27568 12298
rect 27998 12298 28586 12314
rect 27998 12281 28014 12298
rect 27552 12264 27754 12281
rect 26794 12226 27754 12264
rect 27812 12264 28014 12281
rect 28570 12281 28586 12298
rect 29016 12298 29604 12314
rect 29016 12281 29032 12298
rect 28570 12264 28772 12281
rect 27812 12226 28772 12264
rect 28830 12264 29032 12281
rect 29588 12281 29604 12298
rect 30034 12298 30622 12314
rect 30034 12281 30050 12298
rect 29588 12264 29790 12281
rect 28830 12226 29790 12264
rect 29848 12264 30050 12281
rect 30606 12281 30622 12298
rect 31052 12298 31640 12314
rect 31052 12281 31068 12298
rect 30606 12264 30808 12281
rect 29848 12226 30808 12264
rect 30866 12264 31068 12281
rect 31624 12281 31640 12298
rect 32070 12298 32658 12314
rect 32070 12281 32086 12298
rect 31624 12264 31826 12281
rect 30866 12226 31826 12264
rect 31884 12264 32086 12281
rect 32642 12281 32658 12298
rect 33088 12298 33676 12314
rect 33088 12281 33104 12298
rect 32642 12264 32844 12281
rect 31884 12226 32844 12264
rect 32902 12264 33104 12281
rect 33660 12281 33676 12298
rect 34106 12298 34694 12314
rect 34106 12281 34122 12298
rect 33660 12264 33862 12281
rect 32902 12226 33862 12264
rect 33920 12264 34122 12281
rect 34678 12281 34694 12298
rect 35124 12298 35712 12314
rect 35124 12281 35140 12298
rect 34678 12264 34880 12281
rect 33920 12226 34880 12264
rect 34938 12264 35140 12281
rect 35696 12281 35712 12298
rect 36142 12298 36730 12314
rect 36142 12281 36158 12298
rect 35696 12264 35898 12281
rect 34938 12226 35898 12264
rect 35956 12264 36158 12281
rect 36714 12281 36730 12298
rect 37160 12298 37748 12314
rect 37160 12281 37176 12298
rect 36714 12264 36916 12281
rect 35956 12226 36916 12264
rect 36974 12264 37176 12281
rect 37732 12281 37748 12298
rect 38178 12298 38766 12314
rect 38178 12281 38194 12298
rect 37732 12264 37934 12281
rect 36974 12226 37934 12264
rect 37992 12264 38194 12281
rect 38750 12281 38766 12298
rect 39196 12298 39784 12314
rect 39196 12281 39212 12298
rect 38750 12264 38952 12281
rect 37992 12226 38952 12264
rect 39010 12264 39212 12281
rect 39768 12281 39784 12298
rect 39768 12264 39970 12281
rect 39010 12226 39970 12264
rect 7902 11930 8862 11968
rect 7902 11913 8104 11930
rect 8088 11896 8104 11913
rect 8660 11913 8862 11930
rect 8920 11930 9880 11968
rect 8920 11913 9122 11930
rect 8660 11896 8676 11913
rect 8088 11880 8676 11896
rect 9106 11896 9122 11913
rect 9678 11913 9880 11930
rect 9938 11930 10898 11968
rect 9938 11913 10140 11930
rect 9678 11896 9694 11913
rect 9106 11880 9694 11896
rect 8088 11822 8676 11838
rect 8088 11805 8104 11822
rect 7902 11788 8104 11805
rect 8660 11805 8676 11822
rect 10124 11896 10140 11913
rect 10696 11913 10898 11930
rect 10956 11930 11916 11968
rect 10956 11913 11158 11930
rect 10696 11896 10712 11913
rect 10124 11880 10712 11896
rect 9106 11822 9694 11838
rect 9106 11805 9122 11822
rect 8660 11788 8862 11805
rect 7902 11750 8862 11788
rect 8920 11788 9122 11805
rect 9678 11805 9694 11822
rect 11142 11896 11158 11913
rect 11714 11913 11916 11930
rect 11974 11930 12934 11968
rect 11974 11913 12176 11930
rect 11714 11896 11730 11913
rect 11142 11880 11730 11896
rect 10124 11822 10712 11838
rect 10124 11805 10140 11822
rect 9678 11788 9880 11805
rect 8920 11750 9880 11788
rect 9938 11788 10140 11805
rect 10696 11805 10712 11822
rect 12160 11896 12176 11913
rect 12732 11913 12934 11930
rect 12992 11930 13952 11968
rect 12992 11913 13194 11930
rect 12732 11896 12748 11913
rect 12160 11880 12748 11896
rect 11142 11822 11730 11838
rect 11142 11805 11158 11822
rect 10696 11788 10898 11805
rect 9938 11750 10898 11788
rect 10956 11788 11158 11805
rect 11714 11805 11730 11822
rect 13178 11896 13194 11913
rect 13750 11913 13952 11930
rect 14010 11930 14970 11968
rect 14010 11913 14212 11930
rect 13750 11896 13766 11913
rect 13178 11880 13766 11896
rect 12160 11822 12748 11838
rect 12160 11805 12176 11822
rect 11714 11788 11916 11805
rect 10956 11750 11916 11788
rect 11974 11788 12176 11805
rect 12732 11805 12748 11822
rect 14196 11896 14212 11913
rect 14768 11913 14970 11930
rect 15028 11930 15988 11968
rect 15028 11913 15230 11930
rect 14768 11896 14784 11913
rect 14196 11880 14784 11896
rect 13178 11822 13766 11838
rect 13178 11805 13194 11822
rect 12732 11788 12934 11805
rect 11974 11750 12934 11788
rect 12992 11788 13194 11805
rect 13750 11805 13766 11822
rect 15214 11896 15230 11913
rect 15786 11913 15988 11930
rect 16046 11930 17006 11968
rect 16046 11913 16248 11930
rect 15786 11896 15802 11913
rect 15214 11880 15802 11896
rect 14196 11822 14784 11838
rect 14196 11805 14212 11822
rect 13750 11788 13952 11805
rect 12992 11750 13952 11788
rect 14010 11788 14212 11805
rect 14768 11805 14784 11822
rect 16232 11896 16248 11913
rect 16804 11913 17006 11930
rect 16804 11896 16820 11913
rect 16232 11880 16820 11896
rect 15214 11822 15802 11838
rect 15214 11805 15230 11822
rect 14768 11788 14970 11805
rect 14010 11750 14970 11788
rect 15028 11788 15230 11805
rect 15786 11805 15802 11822
rect 16232 11822 16820 11838
rect 16232 11805 16248 11822
rect 15786 11788 15988 11805
rect 15028 11750 15988 11788
rect 16046 11788 16248 11805
rect 16804 11805 16820 11822
rect 16804 11788 17006 11805
rect 16046 11750 17006 11788
rect 19668 11588 20628 11626
rect 19668 11571 19870 11588
rect 19854 11554 19870 11571
rect 20426 11571 20628 11588
rect 20686 11588 21646 11626
rect 20686 11571 20888 11588
rect 20426 11554 20442 11571
rect 19854 11538 20442 11554
rect 20872 11554 20888 11571
rect 21444 11571 21646 11588
rect 21704 11588 22664 11626
rect 21704 11571 21906 11588
rect 21444 11554 21460 11571
rect 20872 11538 21460 11554
rect 21890 11554 21906 11571
rect 22462 11571 22664 11588
rect 22722 11588 23682 11626
rect 22722 11571 22924 11588
rect 22462 11554 22478 11571
rect 21890 11538 22478 11554
rect 22908 11554 22924 11571
rect 23480 11571 23682 11588
rect 23740 11588 24700 11626
rect 23740 11571 23942 11588
rect 23480 11554 23496 11571
rect 22908 11538 23496 11554
rect 23926 11554 23942 11571
rect 24498 11571 24700 11588
rect 24758 11588 25718 11626
rect 24758 11571 24960 11588
rect 24498 11554 24514 11571
rect 23926 11538 24514 11554
rect 24944 11554 24960 11571
rect 25516 11571 25718 11588
rect 25776 11588 26736 11626
rect 25776 11571 25978 11588
rect 25516 11554 25532 11571
rect 24944 11538 25532 11554
rect 25962 11554 25978 11571
rect 26534 11571 26736 11588
rect 26794 11588 27754 11626
rect 26794 11571 26996 11588
rect 26534 11554 26550 11571
rect 25962 11538 26550 11554
rect 26980 11554 26996 11571
rect 27552 11571 27754 11588
rect 27812 11588 28772 11626
rect 27812 11571 28014 11588
rect 27552 11554 27568 11571
rect 26980 11538 27568 11554
rect 27998 11554 28014 11571
rect 28570 11571 28772 11588
rect 28830 11588 29790 11626
rect 28830 11571 29032 11588
rect 28570 11554 28586 11571
rect 27998 11538 28586 11554
rect 29016 11554 29032 11571
rect 29588 11571 29790 11588
rect 29848 11588 30808 11626
rect 29848 11571 30050 11588
rect 29588 11554 29604 11571
rect 29016 11538 29604 11554
rect 30034 11554 30050 11571
rect 30606 11571 30808 11588
rect 30866 11588 31826 11626
rect 30866 11571 31068 11588
rect 30606 11554 30622 11571
rect 30034 11538 30622 11554
rect 31052 11554 31068 11571
rect 31624 11571 31826 11588
rect 31884 11588 32844 11626
rect 31884 11571 32086 11588
rect 31624 11554 31640 11571
rect 31052 11538 31640 11554
rect 32070 11554 32086 11571
rect 32642 11571 32844 11588
rect 32902 11588 33862 11626
rect 32902 11571 33104 11588
rect 32642 11554 32658 11571
rect 32070 11538 32658 11554
rect 33088 11554 33104 11571
rect 33660 11571 33862 11588
rect 33920 11588 34880 11626
rect 33920 11571 34122 11588
rect 33660 11554 33676 11571
rect 33088 11538 33676 11554
rect 34106 11554 34122 11571
rect 34678 11571 34880 11588
rect 34938 11588 35898 11626
rect 34938 11571 35140 11588
rect 34678 11554 34694 11571
rect 34106 11538 34694 11554
rect 35124 11554 35140 11571
rect 35696 11571 35898 11588
rect 35956 11588 36916 11626
rect 35956 11571 36158 11588
rect 35696 11554 35712 11571
rect 35124 11538 35712 11554
rect 36142 11554 36158 11571
rect 36714 11571 36916 11588
rect 36974 11588 37934 11626
rect 36974 11571 37176 11588
rect 36714 11554 36730 11571
rect 36142 11538 36730 11554
rect 37160 11554 37176 11571
rect 37732 11571 37934 11588
rect 37992 11588 38952 11626
rect 37992 11571 38194 11588
rect 37732 11554 37748 11571
rect 37160 11538 37748 11554
rect 38178 11554 38194 11571
rect 38750 11571 38952 11588
rect 39010 11588 39970 11626
rect 39010 11571 39212 11588
rect 38750 11554 38766 11571
rect 38178 11538 38766 11554
rect 39196 11554 39212 11571
rect 39768 11571 39970 11588
rect 39768 11554 39784 11571
rect 39196 11538 39784 11554
rect 7902 11112 8862 11150
rect 7902 11095 8104 11112
rect 8088 11078 8104 11095
rect 8660 11095 8862 11112
rect 8920 11112 9880 11150
rect 8920 11095 9122 11112
rect 8660 11078 8676 11095
rect 8088 11062 8676 11078
rect 9106 11078 9122 11095
rect 9678 11095 9880 11112
rect 9938 11112 10898 11150
rect 9938 11095 10140 11112
rect 9678 11078 9694 11095
rect 9106 11062 9694 11078
rect 8088 11004 8676 11020
rect 8088 10987 8104 11004
rect 7902 10970 8104 10987
rect 8660 10987 8676 11004
rect 10124 11078 10140 11095
rect 10696 11095 10898 11112
rect 10956 11112 11916 11150
rect 10956 11095 11158 11112
rect 10696 11078 10712 11095
rect 10124 11062 10712 11078
rect 9106 11004 9694 11020
rect 9106 10987 9122 11004
rect 8660 10970 8862 10987
rect 7902 10932 8862 10970
rect 8920 10970 9122 10987
rect 9678 10987 9694 11004
rect 11142 11078 11158 11095
rect 11714 11095 11916 11112
rect 11974 11112 12934 11150
rect 11974 11095 12176 11112
rect 11714 11078 11730 11095
rect 11142 11062 11730 11078
rect 10124 11004 10712 11020
rect 10124 10987 10140 11004
rect 9678 10970 9880 10987
rect 8920 10932 9880 10970
rect 9938 10970 10140 10987
rect 10696 10987 10712 11004
rect 12160 11078 12176 11095
rect 12732 11095 12934 11112
rect 12992 11112 13952 11150
rect 12992 11095 13194 11112
rect 12732 11078 12748 11095
rect 12160 11062 12748 11078
rect 11142 11004 11730 11020
rect 11142 10987 11158 11004
rect 10696 10970 10898 10987
rect 9938 10932 10898 10970
rect 10956 10970 11158 10987
rect 11714 10987 11730 11004
rect 13178 11078 13194 11095
rect 13750 11095 13952 11112
rect 14010 11112 14970 11150
rect 14010 11095 14212 11112
rect 13750 11078 13766 11095
rect 13178 11062 13766 11078
rect 12160 11004 12748 11020
rect 12160 10987 12176 11004
rect 11714 10970 11916 10987
rect 10956 10932 11916 10970
rect 11974 10970 12176 10987
rect 12732 10987 12748 11004
rect 14196 11078 14212 11095
rect 14768 11095 14970 11112
rect 15028 11112 15988 11150
rect 15028 11095 15230 11112
rect 14768 11078 14784 11095
rect 14196 11062 14784 11078
rect 13178 11004 13766 11020
rect 13178 10987 13194 11004
rect 12732 10970 12934 10987
rect 11974 10932 12934 10970
rect 12992 10970 13194 10987
rect 13750 10987 13766 11004
rect 15214 11078 15230 11095
rect 15786 11095 15988 11112
rect 16046 11112 17006 11150
rect 16046 11095 16248 11112
rect 15786 11078 15802 11095
rect 15214 11062 15802 11078
rect 14196 11004 14784 11020
rect 14196 10987 14212 11004
rect 13750 10970 13952 10987
rect 12992 10932 13952 10970
rect 14010 10970 14212 10987
rect 14768 10987 14784 11004
rect 16232 11078 16248 11095
rect 16804 11095 17006 11112
rect 16804 11078 16820 11095
rect 16232 11062 16820 11078
rect 15214 11004 15802 11020
rect 15214 10987 15230 11004
rect 14768 10970 14970 10987
rect 14010 10932 14970 10970
rect 15028 10970 15230 10987
rect 15786 10987 15802 11004
rect 16232 11004 16820 11020
rect 16232 10987 16248 11004
rect 15786 10970 15988 10987
rect 15028 10932 15988 10970
rect 16046 10970 16248 10987
rect 16804 10987 16820 11004
rect 16804 10970 17006 10987
rect 16046 10932 17006 10970
rect 19854 10920 20442 10936
rect 19854 10903 19870 10920
rect 19668 10886 19870 10903
rect 20426 10903 20442 10920
rect 20872 10920 21460 10936
rect 20872 10903 20888 10920
rect 20426 10886 20628 10903
rect 19668 10848 20628 10886
rect 20686 10886 20888 10903
rect 21444 10903 21460 10920
rect 21890 10920 22478 10936
rect 21890 10903 21906 10920
rect 21444 10886 21646 10903
rect 20686 10848 21646 10886
rect 21704 10886 21906 10903
rect 22462 10903 22478 10920
rect 22908 10920 23496 10936
rect 22908 10903 22924 10920
rect 22462 10886 22664 10903
rect 21704 10848 22664 10886
rect 22722 10886 22924 10903
rect 23480 10903 23496 10920
rect 23926 10920 24514 10936
rect 23926 10903 23942 10920
rect 23480 10886 23682 10903
rect 22722 10848 23682 10886
rect 23740 10886 23942 10903
rect 24498 10903 24514 10920
rect 24944 10920 25532 10936
rect 24944 10903 24960 10920
rect 24498 10886 24700 10903
rect 23740 10848 24700 10886
rect 24758 10886 24960 10903
rect 25516 10903 25532 10920
rect 25962 10920 26550 10936
rect 25962 10903 25978 10920
rect 25516 10886 25718 10903
rect 24758 10848 25718 10886
rect 25776 10886 25978 10903
rect 26534 10903 26550 10920
rect 26980 10920 27568 10936
rect 26980 10903 26996 10920
rect 26534 10886 26736 10903
rect 25776 10848 26736 10886
rect 26794 10886 26996 10903
rect 27552 10903 27568 10920
rect 27998 10920 28586 10936
rect 27998 10903 28014 10920
rect 27552 10886 27754 10903
rect 26794 10848 27754 10886
rect 27812 10886 28014 10903
rect 28570 10903 28586 10920
rect 29016 10920 29604 10936
rect 29016 10903 29032 10920
rect 28570 10886 28772 10903
rect 27812 10848 28772 10886
rect 28830 10886 29032 10903
rect 29588 10903 29604 10920
rect 30034 10920 30622 10936
rect 30034 10903 30050 10920
rect 29588 10886 29790 10903
rect 28830 10848 29790 10886
rect 29848 10886 30050 10903
rect 30606 10903 30622 10920
rect 31052 10920 31640 10936
rect 31052 10903 31068 10920
rect 30606 10886 30808 10903
rect 29848 10848 30808 10886
rect 30866 10886 31068 10903
rect 31624 10903 31640 10920
rect 32070 10920 32658 10936
rect 32070 10903 32086 10920
rect 31624 10886 31826 10903
rect 30866 10848 31826 10886
rect 31884 10886 32086 10903
rect 32642 10903 32658 10920
rect 33088 10920 33676 10936
rect 33088 10903 33104 10920
rect 32642 10886 32844 10903
rect 31884 10848 32844 10886
rect 32902 10886 33104 10903
rect 33660 10903 33676 10920
rect 34106 10920 34694 10936
rect 34106 10903 34122 10920
rect 33660 10886 33862 10903
rect 32902 10848 33862 10886
rect 33920 10886 34122 10903
rect 34678 10903 34694 10920
rect 35124 10920 35712 10936
rect 35124 10903 35140 10920
rect 34678 10886 34880 10903
rect 33920 10848 34880 10886
rect 34938 10886 35140 10903
rect 35696 10903 35712 10920
rect 36142 10920 36730 10936
rect 36142 10903 36158 10920
rect 35696 10886 35898 10903
rect 34938 10848 35898 10886
rect 35956 10886 36158 10903
rect 36714 10903 36730 10920
rect 37160 10920 37748 10936
rect 37160 10903 37176 10920
rect 36714 10886 36916 10903
rect 35956 10848 36916 10886
rect 36974 10886 37176 10903
rect 37732 10903 37748 10920
rect 38178 10920 38766 10936
rect 38178 10903 38194 10920
rect 37732 10886 37934 10903
rect 36974 10848 37934 10886
rect 37992 10886 38194 10903
rect 38750 10903 38766 10920
rect 39196 10920 39784 10936
rect 39196 10903 39212 10920
rect 38750 10886 38952 10903
rect 37992 10848 38952 10886
rect 39010 10886 39212 10903
rect 39768 10903 39784 10920
rect 39768 10886 39970 10903
rect 39010 10848 39970 10886
rect 7902 10294 8862 10332
rect 7902 10277 8104 10294
rect 8088 10260 8104 10277
rect 8660 10277 8862 10294
rect 8920 10294 9880 10332
rect 8920 10277 9122 10294
rect 8660 10260 8676 10277
rect 8088 10244 8676 10260
rect 9106 10260 9122 10277
rect 9678 10277 9880 10294
rect 9938 10294 10898 10332
rect 9938 10277 10140 10294
rect 9678 10260 9694 10277
rect 9106 10244 9694 10260
rect 8088 10186 8676 10202
rect 8088 10169 8104 10186
rect 7902 10152 8104 10169
rect 8660 10169 8676 10186
rect 10124 10260 10140 10277
rect 10696 10277 10898 10294
rect 10956 10294 11916 10332
rect 10956 10277 11158 10294
rect 10696 10260 10712 10277
rect 10124 10244 10712 10260
rect 9106 10186 9694 10202
rect 9106 10169 9122 10186
rect 8660 10152 8862 10169
rect 7902 10114 8862 10152
rect 8920 10152 9122 10169
rect 9678 10169 9694 10186
rect 11142 10260 11158 10277
rect 11714 10277 11916 10294
rect 11974 10294 12934 10332
rect 11974 10277 12176 10294
rect 11714 10260 11730 10277
rect 11142 10244 11730 10260
rect 10124 10186 10712 10202
rect 10124 10169 10140 10186
rect 9678 10152 9880 10169
rect 8920 10114 9880 10152
rect 9938 10152 10140 10169
rect 10696 10169 10712 10186
rect 12160 10260 12176 10277
rect 12732 10277 12934 10294
rect 12992 10294 13952 10332
rect 12992 10277 13194 10294
rect 12732 10260 12748 10277
rect 12160 10244 12748 10260
rect 11142 10186 11730 10202
rect 11142 10169 11158 10186
rect 10696 10152 10898 10169
rect 9938 10114 10898 10152
rect 10956 10152 11158 10169
rect 11714 10169 11730 10186
rect 13178 10260 13194 10277
rect 13750 10277 13952 10294
rect 14010 10294 14970 10332
rect 14010 10277 14212 10294
rect 13750 10260 13766 10277
rect 13178 10244 13766 10260
rect 12160 10186 12748 10202
rect 12160 10169 12176 10186
rect 11714 10152 11916 10169
rect 10956 10114 11916 10152
rect 11974 10152 12176 10169
rect 12732 10169 12748 10186
rect 14196 10260 14212 10277
rect 14768 10277 14970 10294
rect 15028 10294 15988 10332
rect 15028 10277 15230 10294
rect 14768 10260 14784 10277
rect 14196 10244 14784 10260
rect 13178 10186 13766 10202
rect 13178 10169 13194 10186
rect 12732 10152 12934 10169
rect 11974 10114 12934 10152
rect 12992 10152 13194 10169
rect 13750 10169 13766 10186
rect 15214 10260 15230 10277
rect 15786 10277 15988 10294
rect 16046 10294 17006 10332
rect 16046 10277 16248 10294
rect 15786 10260 15802 10277
rect 15214 10244 15802 10260
rect 14196 10186 14784 10202
rect 14196 10169 14212 10186
rect 13750 10152 13952 10169
rect 12992 10114 13952 10152
rect 14010 10152 14212 10169
rect 14768 10169 14784 10186
rect 16232 10260 16248 10277
rect 16804 10277 17006 10294
rect 16804 10260 16820 10277
rect 16232 10244 16820 10260
rect 15214 10186 15802 10202
rect 15214 10169 15230 10186
rect 14768 10152 14970 10169
rect 14010 10114 14970 10152
rect 15028 10152 15230 10169
rect 15786 10169 15802 10186
rect 16232 10186 16820 10202
rect 16232 10169 16248 10186
rect 15786 10152 15988 10169
rect 15028 10114 15988 10152
rect 16046 10152 16248 10169
rect 16804 10169 16820 10186
rect 19668 10210 20628 10248
rect 19668 10193 19870 10210
rect 19854 10176 19870 10193
rect 20426 10193 20628 10210
rect 20686 10210 21646 10248
rect 20686 10193 20888 10210
rect 20426 10176 20442 10193
rect 16804 10152 17006 10169
rect 19854 10160 20442 10176
rect 20872 10176 20888 10193
rect 21444 10193 21646 10210
rect 21704 10210 22664 10248
rect 21704 10193 21906 10210
rect 21444 10176 21460 10193
rect 20872 10160 21460 10176
rect 21890 10176 21906 10193
rect 22462 10193 22664 10210
rect 22722 10210 23682 10248
rect 22722 10193 22924 10210
rect 22462 10176 22478 10193
rect 21890 10160 22478 10176
rect 22908 10176 22924 10193
rect 23480 10193 23682 10210
rect 23740 10210 24700 10248
rect 23740 10193 23942 10210
rect 23480 10176 23496 10193
rect 22908 10160 23496 10176
rect 23926 10176 23942 10193
rect 24498 10193 24700 10210
rect 24758 10210 25718 10248
rect 24758 10193 24960 10210
rect 24498 10176 24514 10193
rect 23926 10160 24514 10176
rect 24944 10176 24960 10193
rect 25516 10193 25718 10210
rect 25776 10210 26736 10248
rect 25776 10193 25978 10210
rect 25516 10176 25532 10193
rect 24944 10160 25532 10176
rect 25962 10176 25978 10193
rect 26534 10193 26736 10210
rect 26794 10210 27754 10248
rect 26794 10193 26996 10210
rect 26534 10176 26550 10193
rect 25962 10160 26550 10176
rect 26980 10176 26996 10193
rect 27552 10193 27754 10210
rect 27812 10210 28772 10248
rect 27812 10193 28014 10210
rect 27552 10176 27568 10193
rect 26980 10160 27568 10176
rect 27998 10176 28014 10193
rect 28570 10193 28772 10210
rect 28830 10210 29790 10248
rect 28830 10193 29032 10210
rect 28570 10176 28586 10193
rect 27998 10160 28586 10176
rect 29016 10176 29032 10193
rect 29588 10193 29790 10210
rect 29848 10210 30808 10248
rect 29848 10193 30050 10210
rect 29588 10176 29604 10193
rect 29016 10160 29604 10176
rect 30034 10176 30050 10193
rect 30606 10193 30808 10210
rect 30866 10210 31826 10248
rect 30866 10193 31068 10210
rect 30606 10176 30622 10193
rect 30034 10160 30622 10176
rect 31052 10176 31068 10193
rect 31624 10193 31826 10210
rect 31884 10210 32844 10248
rect 31884 10193 32086 10210
rect 31624 10176 31640 10193
rect 31052 10160 31640 10176
rect 32070 10176 32086 10193
rect 32642 10193 32844 10210
rect 32902 10210 33862 10248
rect 32902 10193 33104 10210
rect 32642 10176 32658 10193
rect 32070 10160 32658 10176
rect 33088 10176 33104 10193
rect 33660 10193 33862 10210
rect 33920 10210 34880 10248
rect 33920 10193 34122 10210
rect 33660 10176 33676 10193
rect 33088 10160 33676 10176
rect 34106 10176 34122 10193
rect 34678 10193 34880 10210
rect 34938 10210 35898 10248
rect 34938 10193 35140 10210
rect 34678 10176 34694 10193
rect 34106 10160 34694 10176
rect 35124 10176 35140 10193
rect 35696 10193 35898 10210
rect 35956 10210 36916 10248
rect 35956 10193 36158 10210
rect 35696 10176 35712 10193
rect 35124 10160 35712 10176
rect 36142 10176 36158 10193
rect 36714 10193 36916 10210
rect 36974 10210 37934 10248
rect 36974 10193 37176 10210
rect 36714 10176 36730 10193
rect 36142 10160 36730 10176
rect 37160 10176 37176 10193
rect 37732 10193 37934 10210
rect 37992 10210 38952 10248
rect 37992 10193 38194 10210
rect 37732 10176 37748 10193
rect 37160 10160 37748 10176
rect 38178 10176 38194 10193
rect 38750 10193 38952 10210
rect 39010 10210 39970 10248
rect 39010 10193 39212 10210
rect 38750 10176 38766 10193
rect 38178 10160 38766 10176
rect 39196 10176 39212 10193
rect 39768 10193 39970 10210
rect 39768 10176 39784 10193
rect 39196 10160 39784 10176
rect 16046 10114 17006 10152
rect 19854 9688 20442 9704
rect 19854 9671 19870 9688
rect 19668 9654 19870 9671
rect 20426 9671 20442 9688
rect 20872 9688 21460 9704
rect 20872 9671 20888 9688
rect 20426 9654 20628 9671
rect 19668 9616 20628 9654
rect 20686 9654 20888 9671
rect 21444 9671 21460 9688
rect 21890 9688 22478 9704
rect 21890 9671 21906 9688
rect 21444 9654 21646 9671
rect 20686 9616 21646 9654
rect 21704 9654 21906 9671
rect 22462 9671 22478 9688
rect 22908 9688 23496 9704
rect 22908 9671 22924 9688
rect 22462 9654 22664 9671
rect 21704 9616 22664 9654
rect 22722 9654 22924 9671
rect 23480 9671 23496 9688
rect 23926 9688 24514 9704
rect 23926 9671 23942 9688
rect 23480 9654 23682 9671
rect 22722 9616 23682 9654
rect 23740 9654 23942 9671
rect 24498 9671 24514 9688
rect 24944 9688 25532 9704
rect 24944 9671 24960 9688
rect 24498 9654 24700 9671
rect 23740 9616 24700 9654
rect 24758 9654 24960 9671
rect 25516 9671 25532 9688
rect 25962 9688 26550 9704
rect 25962 9671 25978 9688
rect 25516 9654 25718 9671
rect 24758 9616 25718 9654
rect 25776 9654 25978 9671
rect 26534 9671 26550 9688
rect 26980 9688 27568 9704
rect 26980 9671 26996 9688
rect 26534 9654 26736 9671
rect 25776 9616 26736 9654
rect 26794 9654 26996 9671
rect 27552 9671 27568 9688
rect 27998 9688 28586 9704
rect 27998 9671 28014 9688
rect 27552 9654 27754 9671
rect 26794 9616 27754 9654
rect 27812 9654 28014 9671
rect 28570 9671 28586 9688
rect 29016 9688 29604 9704
rect 29016 9671 29032 9688
rect 28570 9654 28772 9671
rect 27812 9616 28772 9654
rect 28830 9654 29032 9671
rect 29588 9671 29604 9688
rect 30034 9688 30622 9704
rect 30034 9671 30050 9688
rect 29588 9654 29790 9671
rect 28830 9616 29790 9654
rect 29848 9654 30050 9671
rect 30606 9671 30622 9688
rect 31052 9688 31640 9704
rect 31052 9671 31068 9688
rect 30606 9654 30808 9671
rect 29848 9616 30808 9654
rect 30866 9654 31068 9671
rect 31624 9671 31640 9688
rect 32070 9688 32658 9704
rect 32070 9671 32086 9688
rect 31624 9654 31826 9671
rect 30866 9616 31826 9654
rect 31884 9654 32086 9671
rect 32642 9671 32658 9688
rect 33088 9688 33676 9704
rect 33088 9671 33104 9688
rect 32642 9654 32844 9671
rect 31884 9616 32844 9654
rect 32902 9654 33104 9671
rect 33660 9671 33676 9688
rect 34106 9688 34694 9704
rect 34106 9671 34122 9688
rect 33660 9654 33862 9671
rect 32902 9616 33862 9654
rect 33920 9654 34122 9671
rect 34678 9671 34694 9688
rect 35124 9688 35712 9704
rect 35124 9671 35140 9688
rect 34678 9654 34880 9671
rect 33920 9616 34880 9654
rect 34938 9654 35140 9671
rect 35696 9671 35712 9688
rect 36142 9688 36730 9704
rect 36142 9671 36158 9688
rect 35696 9654 35898 9671
rect 34938 9616 35898 9654
rect 35956 9654 36158 9671
rect 36714 9671 36730 9688
rect 37160 9688 37748 9704
rect 37160 9671 37176 9688
rect 36714 9654 36916 9671
rect 35956 9616 36916 9654
rect 36974 9654 37176 9671
rect 37732 9671 37748 9688
rect 38178 9688 38766 9704
rect 38178 9671 38194 9688
rect 37732 9654 37934 9671
rect 36974 9616 37934 9654
rect 37992 9654 38194 9671
rect 38750 9671 38766 9688
rect 39196 9688 39784 9704
rect 39196 9671 39212 9688
rect 38750 9654 38952 9671
rect 37992 9616 38952 9654
rect 39010 9654 39212 9671
rect 39768 9671 39784 9688
rect 39768 9654 39970 9671
rect 39010 9616 39970 9654
rect 7902 9476 8862 9514
rect 7902 9459 8104 9476
rect 8088 9442 8104 9459
rect 8660 9459 8862 9476
rect 8920 9476 9880 9514
rect 8920 9459 9122 9476
rect 8660 9442 8676 9459
rect 8088 9426 8676 9442
rect 9106 9442 9122 9459
rect 9678 9459 9880 9476
rect 9938 9476 10898 9514
rect 9938 9459 10140 9476
rect 9678 9442 9694 9459
rect 9106 9426 9694 9442
rect 8088 9368 8676 9384
rect 8088 9351 8104 9368
rect 7902 9334 8104 9351
rect 8660 9351 8676 9368
rect 10124 9442 10140 9459
rect 10696 9459 10898 9476
rect 10956 9476 11916 9514
rect 10956 9459 11158 9476
rect 10696 9442 10712 9459
rect 10124 9426 10712 9442
rect 9106 9368 9694 9384
rect 9106 9351 9122 9368
rect 8660 9334 8862 9351
rect 7902 9296 8862 9334
rect 8920 9334 9122 9351
rect 9678 9351 9694 9368
rect 11142 9442 11158 9459
rect 11714 9459 11916 9476
rect 11974 9476 12934 9514
rect 11974 9459 12176 9476
rect 11714 9442 11730 9459
rect 11142 9426 11730 9442
rect 10124 9368 10712 9384
rect 10124 9351 10140 9368
rect 9678 9334 9880 9351
rect 8920 9296 9880 9334
rect 9938 9334 10140 9351
rect 10696 9351 10712 9368
rect 12160 9442 12176 9459
rect 12732 9459 12934 9476
rect 12992 9476 13952 9514
rect 12992 9459 13194 9476
rect 12732 9442 12748 9459
rect 12160 9426 12748 9442
rect 11142 9368 11730 9384
rect 11142 9351 11158 9368
rect 10696 9334 10898 9351
rect 9938 9296 10898 9334
rect 10956 9334 11158 9351
rect 11714 9351 11730 9368
rect 13178 9442 13194 9459
rect 13750 9459 13952 9476
rect 14010 9476 14970 9514
rect 14010 9459 14212 9476
rect 13750 9442 13766 9459
rect 13178 9426 13766 9442
rect 12160 9368 12748 9384
rect 12160 9351 12176 9368
rect 11714 9334 11916 9351
rect 10956 9296 11916 9334
rect 11974 9334 12176 9351
rect 12732 9351 12748 9368
rect 14196 9442 14212 9459
rect 14768 9459 14970 9476
rect 15028 9476 15988 9514
rect 15028 9459 15230 9476
rect 14768 9442 14784 9459
rect 14196 9426 14784 9442
rect 13178 9368 13766 9384
rect 13178 9351 13194 9368
rect 12732 9334 12934 9351
rect 11974 9296 12934 9334
rect 12992 9334 13194 9351
rect 13750 9351 13766 9368
rect 15214 9442 15230 9459
rect 15786 9459 15988 9476
rect 16046 9476 17006 9514
rect 16046 9459 16248 9476
rect 15786 9442 15802 9459
rect 15214 9426 15802 9442
rect 14196 9368 14784 9384
rect 14196 9351 14212 9368
rect 13750 9334 13952 9351
rect 12992 9296 13952 9334
rect 14010 9334 14212 9351
rect 14768 9351 14784 9368
rect 16232 9442 16248 9459
rect 16804 9459 17006 9476
rect 16804 9442 16820 9459
rect 16232 9426 16820 9442
rect 15214 9368 15802 9384
rect 15214 9351 15230 9368
rect 14768 9334 14970 9351
rect 14010 9296 14970 9334
rect 15028 9334 15230 9351
rect 15786 9351 15802 9368
rect 16232 9368 16820 9384
rect 16232 9351 16248 9368
rect 15786 9334 15988 9351
rect 15028 9296 15988 9334
rect 16046 9334 16248 9351
rect 16804 9351 16820 9368
rect 16804 9334 17006 9351
rect 16046 9296 17006 9334
rect 19668 8978 20628 9016
rect 19668 8961 19870 8978
rect 19854 8944 19870 8961
rect 20426 8961 20628 8978
rect 20686 8978 21646 9016
rect 20686 8961 20888 8978
rect 20426 8944 20442 8961
rect 19854 8928 20442 8944
rect 20872 8944 20888 8961
rect 21444 8961 21646 8978
rect 21704 8978 22664 9016
rect 21704 8961 21906 8978
rect 21444 8944 21460 8961
rect 20872 8928 21460 8944
rect 21890 8944 21906 8961
rect 22462 8961 22664 8978
rect 22722 8978 23682 9016
rect 22722 8961 22924 8978
rect 22462 8944 22478 8961
rect 21890 8928 22478 8944
rect 22908 8944 22924 8961
rect 23480 8961 23682 8978
rect 23740 8978 24700 9016
rect 23740 8961 23942 8978
rect 23480 8944 23496 8961
rect 22908 8928 23496 8944
rect 23926 8944 23942 8961
rect 24498 8961 24700 8978
rect 24758 8978 25718 9016
rect 24758 8961 24960 8978
rect 24498 8944 24514 8961
rect 23926 8928 24514 8944
rect 24944 8944 24960 8961
rect 25516 8961 25718 8978
rect 25776 8978 26736 9016
rect 25776 8961 25978 8978
rect 25516 8944 25532 8961
rect 24944 8928 25532 8944
rect 25962 8944 25978 8961
rect 26534 8961 26736 8978
rect 26794 8978 27754 9016
rect 26794 8961 26996 8978
rect 26534 8944 26550 8961
rect 25962 8928 26550 8944
rect 26980 8944 26996 8961
rect 27552 8961 27754 8978
rect 27812 8978 28772 9016
rect 27812 8961 28014 8978
rect 27552 8944 27568 8961
rect 26980 8928 27568 8944
rect 27998 8944 28014 8961
rect 28570 8961 28772 8978
rect 28830 8978 29790 9016
rect 28830 8961 29032 8978
rect 28570 8944 28586 8961
rect 27998 8928 28586 8944
rect 29016 8944 29032 8961
rect 29588 8961 29790 8978
rect 29848 8978 30808 9016
rect 29848 8961 30050 8978
rect 29588 8944 29604 8961
rect 29016 8928 29604 8944
rect 30034 8944 30050 8961
rect 30606 8961 30808 8978
rect 30866 8978 31826 9016
rect 30866 8961 31068 8978
rect 30606 8944 30622 8961
rect 30034 8928 30622 8944
rect 31052 8944 31068 8961
rect 31624 8961 31826 8978
rect 31884 8978 32844 9016
rect 31884 8961 32086 8978
rect 31624 8944 31640 8961
rect 31052 8928 31640 8944
rect 32070 8944 32086 8961
rect 32642 8961 32844 8978
rect 32902 8978 33862 9016
rect 32902 8961 33104 8978
rect 32642 8944 32658 8961
rect 32070 8928 32658 8944
rect 33088 8944 33104 8961
rect 33660 8961 33862 8978
rect 33920 8978 34880 9016
rect 33920 8961 34122 8978
rect 33660 8944 33676 8961
rect 33088 8928 33676 8944
rect 34106 8944 34122 8961
rect 34678 8961 34880 8978
rect 34938 8978 35898 9016
rect 34938 8961 35140 8978
rect 34678 8944 34694 8961
rect 34106 8928 34694 8944
rect 35124 8944 35140 8961
rect 35696 8961 35898 8978
rect 35956 8978 36916 9016
rect 35956 8961 36158 8978
rect 35696 8944 35712 8961
rect 35124 8928 35712 8944
rect 36142 8944 36158 8961
rect 36714 8961 36916 8978
rect 36974 8978 37934 9016
rect 36974 8961 37176 8978
rect 36714 8944 36730 8961
rect 36142 8928 36730 8944
rect 37160 8944 37176 8961
rect 37732 8961 37934 8978
rect 37992 8978 38952 9016
rect 37992 8961 38194 8978
rect 37732 8944 37748 8961
rect 37160 8928 37748 8944
rect 38178 8944 38194 8961
rect 38750 8961 38952 8978
rect 39010 8978 39970 9016
rect 39010 8961 39212 8978
rect 38750 8944 38766 8961
rect 38178 8928 38766 8944
rect 39196 8944 39212 8961
rect 39768 8961 39970 8978
rect 39768 8944 39784 8961
rect 39196 8928 39784 8944
rect 7902 8658 8862 8696
rect 7902 8641 8104 8658
rect 8088 8624 8104 8641
rect 8660 8641 8862 8658
rect 8920 8658 9880 8696
rect 8920 8641 9122 8658
rect 8660 8624 8676 8641
rect 8088 8608 8676 8624
rect 9106 8624 9122 8641
rect 9678 8641 9880 8658
rect 9938 8658 10898 8696
rect 9938 8641 10140 8658
rect 9678 8624 9694 8641
rect 9106 8608 9694 8624
rect 8088 8550 8676 8566
rect 8088 8533 8104 8550
rect 7902 8516 8104 8533
rect 8660 8533 8676 8550
rect 10124 8624 10140 8641
rect 10696 8641 10898 8658
rect 10956 8658 11916 8696
rect 10956 8641 11158 8658
rect 10696 8624 10712 8641
rect 10124 8608 10712 8624
rect 9106 8550 9694 8566
rect 9106 8533 9122 8550
rect 8660 8516 8862 8533
rect 7902 8478 8862 8516
rect 8920 8516 9122 8533
rect 9678 8533 9694 8550
rect 11142 8624 11158 8641
rect 11714 8641 11916 8658
rect 11974 8658 12934 8696
rect 11974 8641 12176 8658
rect 11714 8624 11730 8641
rect 11142 8608 11730 8624
rect 10124 8550 10712 8566
rect 10124 8533 10140 8550
rect 9678 8516 9880 8533
rect 8920 8478 9880 8516
rect 9938 8516 10140 8533
rect 10696 8533 10712 8550
rect 12160 8624 12176 8641
rect 12732 8641 12934 8658
rect 12992 8658 13952 8696
rect 12992 8641 13194 8658
rect 12732 8624 12748 8641
rect 12160 8608 12748 8624
rect 11142 8550 11730 8566
rect 11142 8533 11158 8550
rect 10696 8516 10898 8533
rect 9938 8478 10898 8516
rect 10956 8516 11158 8533
rect 11714 8533 11730 8550
rect 13178 8624 13194 8641
rect 13750 8641 13952 8658
rect 14010 8658 14970 8696
rect 14010 8641 14212 8658
rect 13750 8624 13766 8641
rect 13178 8608 13766 8624
rect 12160 8550 12748 8566
rect 12160 8533 12176 8550
rect 11714 8516 11916 8533
rect 10956 8478 11916 8516
rect 11974 8516 12176 8533
rect 12732 8533 12748 8550
rect 14196 8624 14212 8641
rect 14768 8641 14970 8658
rect 15028 8658 15988 8696
rect 15028 8641 15230 8658
rect 14768 8624 14784 8641
rect 14196 8608 14784 8624
rect 13178 8550 13766 8566
rect 13178 8533 13194 8550
rect 12732 8516 12934 8533
rect 11974 8478 12934 8516
rect 12992 8516 13194 8533
rect 13750 8533 13766 8550
rect 15214 8624 15230 8641
rect 15786 8641 15988 8658
rect 16046 8658 17006 8696
rect 16046 8641 16248 8658
rect 15786 8624 15802 8641
rect 15214 8608 15802 8624
rect 14196 8550 14784 8566
rect 14196 8533 14212 8550
rect 13750 8516 13952 8533
rect 12992 8478 13952 8516
rect 14010 8516 14212 8533
rect 14768 8533 14784 8550
rect 16232 8624 16248 8641
rect 16804 8641 17006 8658
rect 16804 8624 16820 8641
rect 16232 8608 16820 8624
rect 15214 8550 15802 8566
rect 15214 8533 15230 8550
rect 14768 8516 14970 8533
rect 14010 8478 14970 8516
rect 15028 8516 15230 8533
rect 15786 8533 15802 8550
rect 16232 8550 16820 8566
rect 16232 8533 16248 8550
rect 15786 8516 15988 8533
rect 15028 8478 15988 8516
rect 16046 8516 16248 8533
rect 16804 8533 16820 8550
rect 16804 8516 17006 8533
rect 16046 8478 17006 8516
rect 19852 8454 20440 8470
rect 19852 8437 19868 8454
rect 19666 8420 19868 8437
rect 20424 8437 20440 8454
rect 20870 8454 21458 8470
rect 20870 8437 20886 8454
rect 20424 8420 20626 8437
rect 19666 8382 20626 8420
rect 20684 8420 20886 8437
rect 21442 8437 21458 8454
rect 21888 8454 22476 8470
rect 21888 8437 21904 8454
rect 21442 8420 21644 8437
rect 20684 8382 21644 8420
rect 21702 8420 21904 8437
rect 22460 8437 22476 8454
rect 22906 8454 23494 8470
rect 22906 8437 22922 8454
rect 22460 8420 22662 8437
rect 21702 8382 22662 8420
rect 22720 8420 22922 8437
rect 23478 8437 23494 8454
rect 23924 8454 24512 8470
rect 23924 8437 23940 8454
rect 23478 8420 23680 8437
rect 22720 8382 23680 8420
rect 23738 8420 23940 8437
rect 24496 8437 24512 8454
rect 24942 8454 25530 8470
rect 24942 8437 24958 8454
rect 24496 8420 24698 8437
rect 23738 8382 24698 8420
rect 24756 8420 24958 8437
rect 25514 8437 25530 8454
rect 25960 8454 26548 8470
rect 25960 8437 25976 8454
rect 25514 8420 25716 8437
rect 24756 8382 25716 8420
rect 25774 8420 25976 8437
rect 26532 8437 26548 8454
rect 26978 8454 27566 8470
rect 26978 8437 26994 8454
rect 26532 8420 26734 8437
rect 25774 8382 26734 8420
rect 26792 8420 26994 8437
rect 27550 8437 27566 8454
rect 27996 8454 28584 8470
rect 27996 8437 28012 8454
rect 27550 8420 27752 8437
rect 26792 8382 27752 8420
rect 27810 8420 28012 8437
rect 28568 8437 28584 8454
rect 29014 8454 29602 8470
rect 29014 8437 29030 8454
rect 28568 8420 28770 8437
rect 27810 8382 28770 8420
rect 28828 8420 29030 8437
rect 29586 8437 29602 8454
rect 30032 8454 30620 8470
rect 30032 8437 30048 8454
rect 29586 8420 29788 8437
rect 28828 8382 29788 8420
rect 29846 8420 30048 8437
rect 30604 8437 30620 8454
rect 31050 8454 31638 8470
rect 31050 8437 31066 8454
rect 30604 8420 30806 8437
rect 29846 8382 30806 8420
rect 30864 8420 31066 8437
rect 31622 8437 31638 8454
rect 32068 8454 32656 8470
rect 32068 8437 32084 8454
rect 31622 8420 31824 8437
rect 30864 8382 31824 8420
rect 31882 8420 32084 8437
rect 32640 8437 32656 8454
rect 33086 8454 33674 8470
rect 33086 8437 33102 8454
rect 32640 8420 32842 8437
rect 31882 8382 32842 8420
rect 32900 8420 33102 8437
rect 33658 8437 33674 8454
rect 34104 8454 34692 8470
rect 34104 8437 34120 8454
rect 33658 8420 33860 8437
rect 32900 8382 33860 8420
rect 33918 8420 34120 8437
rect 34676 8437 34692 8454
rect 35122 8454 35710 8470
rect 35122 8437 35138 8454
rect 34676 8420 34878 8437
rect 33918 8382 34878 8420
rect 34936 8420 35138 8437
rect 35694 8437 35710 8454
rect 36140 8454 36728 8470
rect 36140 8437 36156 8454
rect 35694 8420 35896 8437
rect 34936 8382 35896 8420
rect 35954 8420 36156 8437
rect 36712 8437 36728 8454
rect 37158 8454 37746 8470
rect 37158 8437 37174 8454
rect 36712 8420 36914 8437
rect 35954 8382 36914 8420
rect 36972 8420 37174 8437
rect 37730 8437 37746 8454
rect 38176 8454 38764 8470
rect 38176 8437 38192 8454
rect 37730 8420 37932 8437
rect 36972 8382 37932 8420
rect 37990 8420 38192 8437
rect 38748 8437 38764 8454
rect 39194 8454 39782 8470
rect 39194 8437 39210 8454
rect 38748 8420 38950 8437
rect 37990 8382 38950 8420
rect 39008 8420 39210 8437
rect 39766 8437 39782 8454
rect 39766 8420 39968 8437
rect 39008 8382 39968 8420
rect 7902 7840 8862 7878
rect 7902 7823 8104 7840
rect 8088 7806 8104 7823
rect 8660 7823 8862 7840
rect 8920 7840 9880 7878
rect 8920 7823 9122 7840
rect 8660 7806 8676 7823
rect 8088 7790 8676 7806
rect 9106 7806 9122 7823
rect 9678 7823 9880 7840
rect 9938 7840 10898 7878
rect 9938 7823 10140 7840
rect 9678 7806 9694 7823
rect 9106 7790 9694 7806
rect 8088 7732 8676 7748
rect 8088 7715 8104 7732
rect 7902 7698 8104 7715
rect 8660 7715 8676 7732
rect 10124 7806 10140 7823
rect 10696 7823 10898 7840
rect 10956 7840 11916 7878
rect 10956 7823 11158 7840
rect 10696 7806 10712 7823
rect 10124 7790 10712 7806
rect 9106 7732 9694 7748
rect 9106 7715 9122 7732
rect 8660 7698 8862 7715
rect 7902 7660 8862 7698
rect 8920 7698 9122 7715
rect 9678 7715 9694 7732
rect 11142 7806 11158 7823
rect 11714 7823 11916 7840
rect 11974 7840 12934 7878
rect 11974 7823 12176 7840
rect 11714 7806 11730 7823
rect 11142 7790 11730 7806
rect 10124 7732 10712 7748
rect 10124 7715 10140 7732
rect 9678 7698 9880 7715
rect 8920 7660 9880 7698
rect 9938 7698 10140 7715
rect 10696 7715 10712 7732
rect 12160 7806 12176 7823
rect 12732 7823 12934 7840
rect 12992 7840 13952 7878
rect 12992 7823 13194 7840
rect 12732 7806 12748 7823
rect 12160 7790 12748 7806
rect 11142 7732 11730 7748
rect 11142 7715 11158 7732
rect 10696 7698 10898 7715
rect 9938 7660 10898 7698
rect 10956 7698 11158 7715
rect 11714 7715 11730 7732
rect 13178 7806 13194 7823
rect 13750 7823 13952 7840
rect 14010 7840 14970 7878
rect 14010 7823 14212 7840
rect 13750 7806 13766 7823
rect 13178 7790 13766 7806
rect 12160 7732 12748 7748
rect 12160 7715 12176 7732
rect 11714 7698 11916 7715
rect 10956 7660 11916 7698
rect 11974 7698 12176 7715
rect 12732 7715 12748 7732
rect 14196 7806 14212 7823
rect 14768 7823 14970 7840
rect 15028 7840 15988 7878
rect 15028 7823 15230 7840
rect 14768 7806 14784 7823
rect 14196 7790 14784 7806
rect 13178 7732 13766 7748
rect 13178 7715 13194 7732
rect 12732 7698 12934 7715
rect 11974 7660 12934 7698
rect 12992 7698 13194 7715
rect 13750 7715 13766 7732
rect 15214 7806 15230 7823
rect 15786 7823 15988 7840
rect 16046 7840 17006 7878
rect 16046 7823 16248 7840
rect 15786 7806 15802 7823
rect 15214 7790 15802 7806
rect 14196 7732 14784 7748
rect 14196 7715 14212 7732
rect 13750 7698 13952 7715
rect 12992 7660 13952 7698
rect 14010 7698 14212 7715
rect 14768 7715 14784 7732
rect 16232 7806 16248 7823
rect 16804 7823 17006 7840
rect 16804 7806 16820 7823
rect 16232 7790 16820 7806
rect 15214 7732 15802 7748
rect 15214 7715 15230 7732
rect 14768 7698 14970 7715
rect 14010 7660 14970 7698
rect 15028 7698 15230 7715
rect 15786 7715 15802 7732
rect 16232 7732 16820 7748
rect 16232 7715 16248 7732
rect 15786 7698 15988 7715
rect 15028 7660 15988 7698
rect 16046 7698 16248 7715
rect 16804 7715 16820 7732
rect 19666 7744 20626 7782
rect 19666 7727 19868 7744
rect 16804 7698 17006 7715
rect 16046 7660 17006 7698
rect 19852 7710 19868 7727
rect 20424 7727 20626 7744
rect 20684 7744 21644 7782
rect 20684 7727 20886 7744
rect 20424 7710 20440 7727
rect 19852 7694 20440 7710
rect 20870 7710 20886 7727
rect 21442 7727 21644 7744
rect 21702 7744 22662 7782
rect 21702 7727 21904 7744
rect 21442 7710 21458 7727
rect 20870 7694 21458 7710
rect 21888 7710 21904 7727
rect 22460 7727 22662 7744
rect 22720 7744 23680 7782
rect 22720 7727 22922 7744
rect 22460 7710 22476 7727
rect 21888 7694 22476 7710
rect 22906 7710 22922 7727
rect 23478 7727 23680 7744
rect 23738 7744 24698 7782
rect 23738 7727 23940 7744
rect 23478 7710 23494 7727
rect 22906 7694 23494 7710
rect 23924 7710 23940 7727
rect 24496 7727 24698 7744
rect 24756 7744 25716 7782
rect 24756 7727 24958 7744
rect 24496 7710 24512 7727
rect 23924 7694 24512 7710
rect 24942 7710 24958 7727
rect 25514 7727 25716 7744
rect 25774 7744 26734 7782
rect 25774 7727 25976 7744
rect 25514 7710 25530 7727
rect 24942 7694 25530 7710
rect 25960 7710 25976 7727
rect 26532 7727 26734 7744
rect 26792 7744 27752 7782
rect 26792 7727 26994 7744
rect 26532 7710 26548 7727
rect 25960 7694 26548 7710
rect 26978 7710 26994 7727
rect 27550 7727 27752 7744
rect 27810 7744 28770 7782
rect 27810 7727 28012 7744
rect 27550 7710 27566 7727
rect 26978 7694 27566 7710
rect 27996 7710 28012 7727
rect 28568 7727 28770 7744
rect 28828 7744 29788 7782
rect 28828 7727 29030 7744
rect 28568 7710 28584 7727
rect 27996 7694 28584 7710
rect 29014 7710 29030 7727
rect 29586 7727 29788 7744
rect 29846 7744 30806 7782
rect 29846 7727 30048 7744
rect 29586 7710 29602 7727
rect 29014 7694 29602 7710
rect 30032 7710 30048 7727
rect 30604 7727 30806 7744
rect 30864 7744 31824 7782
rect 30864 7727 31066 7744
rect 30604 7710 30620 7727
rect 30032 7694 30620 7710
rect 31050 7710 31066 7727
rect 31622 7727 31824 7744
rect 31882 7744 32842 7782
rect 31882 7727 32084 7744
rect 31622 7710 31638 7727
rect 31050 7694 31638 7710
rect 32068 7710 32084 7727
rect 32640 7727 32842 7744
rect 32900 7744 33860 7782
rect 32900 7727 33102 7744
rect 32640 7710 32656 7727
rect 32068 7694 32656 7710
rect 33086 7710 33102 7727
rect 33658 7727 33860 7744
rect 33918 7744 34878 7782
rect 33918 7727 34120 7744
rect 33658 7710 33674 7727
rect 33086 7694 33674 7710
rect 34104 7710 34120 7727
rect 34676 7727 34878 7744
rect 34936 7744 35896 7782
rect 34936 7727 35138 7744
rect 34676 7710 34692 7727
rect 34104 7694 34692 7710
rect 35122 7710 35138 7727
rect 35694 7727 35896 7744
rect 35954 7744 36914 7782
rect 35954 7727 36156 7744
rect 35694 7710 35710 7727
rect 35122 7694 35710 7710
rect 36140 7710 36156 7727
rect 36712 7727 36914 7744
rect 36972 7744 37932 7782
rect 36972 7727 37174 7744
rect 36712 7710 36728 7727
rect 36140 7694 36728 7710
rect 37158 7710 37174 7727
rect 37730 7727 37932 7744
rect 37990 7744 38950 7782
rect 37990 7727 38192 7744
rect 37730 7710 37746 7727
rect 37158 7694 37746 7710
rect 38176 7710 38192 7727
rect 38748 7727 38950 7744
rect 39008 7744 39968 7782
rect 39008 7727 39210 7744
rect 38748 7710 38764 7727
rect 38176 7694 38764 7710
rect 39194 7710 39210 7727
rect 39766 7727 39968 7744
rect 39766 7710 39782 7727
rect 39194 7694 39782 7710
rect 19852 7220 20440 7236
rect 19852 7203 19868 7220
rect 19666 7186 19868 7203
rect 20424 7203 20440 7220
rect 20870 7220 21458 7236
rect 20870 7203 20886 7220
rect 20424 7186 20626 7203
rect 19666 7148 20626 7186
rect 20684 7186 20886 7203
rect 21442 7203 21458 7220
rect 21888 7220 22476 7236
rect 21888 7203 21904 7220
rect 21442 7186 21644 7203
rect 20684 7148 21644 7186
rect 21702 7186 21904 7203
rect 22460 7203 22476 7220
rect 22906 7220 23494 7236
rect 22906 7203 22922 7220
rect 22460 7186 22662 7203
rect 21702 7148 22662 7186
rect 22720 7186 22922 7203
rect 23478 7203 23494 7220
rect 23924 7220 24512 7236
rect 23924 7203 23940 7220
rect 23478 7186 23680 7203
rect 22720 7148 23680 7186
rect 23738 7186 23940 7203
rect 24496 7203 24512 7220
rect 24942 7220 25530 7236
rect 24942 7203 24958 7220
rect 24496 7186 24698 7203
rect 23738 7148 24698 7186
rect 24756 7186 24958 7203
rect 25514 7203 25530 7220
rect 25960 7220 26548 7236
rect 25960 7203 25976 7220
rect 25514 7186 25716 7203
rect 24756 7148 25716 7186
rect 25774 7186 25976 7203
rect 26532 7203 26548 7220
rect 26978 7220 27566 7236
rect 26978 7203 26994 7220
rect 26532 7186 26734 7203
rect 25774 7148 26734 7186
rect 26792 7186 26994 7203
rect 27550 7203 27566 7220
rect 27996 7220 28584 7236
rect 27996 7203 28012 7220
rect 27550 7186 27752 7203
rect 26792 7148 27752 7186
rect 27810 7186 28012 7203
rect 28568 7203 28584 7220
rect 29014 7220 29602 7236
rect 29014 7203 29030 7220
rect 28568 7186 28770 7203
rect 27810 7148 28770 7186
rect 28828 7186 29030 7203
rect 29586 7203 29602 7220
rect 30032 7220 30620 7236
rect 30032 7203 30048 7220
rect 29586 7186 29788 7203
rect 28828 7148 29788 7186
rect 29846 7186 30048 7203
rect 30604 7203 30620 7220
rect 31050 7220 31638 7236
rect 31050 7203 31066 7220
rect 30604 7186 30806 7203
rect 29846 7148 30806 7186
rect 30864 7186 31066 7203
rect 31622 7203 31638 7220
rect 32068 7220 32656 7236
rect 32068 7203 32084 7220
rect 31622 7186 31824 7203
rect 30864 7148 31824 7186
rect 31882 7186 32084 7203
rect 32640 7203 32656 7220
rect 33086 7220 33674 7236
rect 33086 7203 33102 7220
rect 32640 7186 32842 7203
rect 31882 7148 32842 7186
rect 32900 7186 33102 7203
rect 33658 7203 33674 7220
rect 34104 7220 34692 7236
rect 34104 7203 34120 7220
rect 33658 7186 33860 7203
rect 32900 7148 33860 7186
rect 33918 7186 34120 7203
rect 34676 7203 34692 7220
rect 35122 7220 35710 7236
rect 35122 7203 35138 7220
rect 34676 7186 34878 7203
rect 33918 7148 34878 7186
rect 34936 7186 35138 7203
rect 35694 7203 35710 7220
rect 36140 7220 36728 7236
rect 36140 7203 36156 7220
rect 35694 7186 35896 7203
rect 34936 7148 35896 7186
rect 35954 7186 36156 7203
rect 36712 7203 36728 7220
rect 37158 7220 37746 7236
rect 37158 7203 37174 7220
rect 36712 7186 36914 7203
rect 35954 7148 36914 7186
rect 36972 7186 37174 7203
rect 37730 7203 37746 7220
rect 38176 7220 38764 7236
rect 38176 7203 38192 7220
rect 37730 7186 37932 7203
rect 36972 7148 37932 7186
rect 37990 7186 38192 7203
rect 38748 7203 38764 7220
rect 39194 7220 39782 7236
rect 39194 7203 39210 7220
rect 38748 7186 38950 7203
rect 37990 7148 38950 7186
rect 39008 7186 39210 7203
rect 39766 7203 39782 7220
rect 39766 7186 39968 7203
rect 39008 7148 39968 7186
rect 7902 7022 8862 7060
rect 7902 7005 8104 7022
rect 8088 6988 8104 7005
rect 8660 7005 8862 7022
rect 8920 7022 9880 7060
rect 8920 7005 9122 7022
rect 8660 6988 8676 7005
rect 8088 6972 8676 6988
rect 9106 6988 9122 7005
rect 9678 7005 9880 7022
rect 9938 7022 10898 7060
rect 9938 7005 10140 7022
rect 9678 6988 9694 7005
rect 9106 6972 9694 6988
rect 8088 6914 8676 6930
rect 8088 6897 8104 6914
rect 7902 6880 8104 6897
rect 8660 6897 8676 6914
rect 10124 6988 10140 7005
rect 10696 7005 10898 7022
rect 10956 7022 11916 7060
rect 10956 7005 11158 7022
rect 10696 6988 10712 7005
rect 10124 6972 10712 6988
rect 9106 6914 9694 6930
rect 9106 6897 9122 6914
rect 8660 6880 8862 6897
rect 7902 6842 8862 6880
rect 8920 6880 9122 6897
rect 9678 6897 9694 6914
rect 11142 6988 11158 7005
rect 11714 7005 11916 7022
rect 11974 7022 12934 7060
rect 11974 7005 12176 7022
rect 11714 6988 11730 7005
rect 11142 6972 11730 6988
rect 10124 6914 10712 6930
rect 10124 6897 10140 6914
rect 9678 6880 9880 6897
rect 8920 6842 9880 6880
rect 9938 6880 10140 6897
rect 10696 6897 10712 6914
rect 12160 6988 12176 7005
rect 12732 7005 12934 7022
rect 12992 7022 13952 7060
rect 12992 7005 13194 7022
rect 12732 6988 12748 7005
rect 12160 6972 12748 6988
rect 11142 6914 11730 6930
rect 11142 6897 11158 6914
rect 10696 6880 10898 6897
rect 9938 6842 10898 6880
rect 10956 6880 11158 6897
rect 11714 6897 11730 6914
rect 13178 6988 13194 7005
rect 13750 7005 13952 7022
rect 14010 7022 14970 7060
rect 14010 7005 14212 7022
rect 13750 6988 13766 7005
rect 13178 6972 13766 6988
rect 12160 6914 12748 6930
rect 12160 6897 12176 6914
rect 11714 6880 11916 6897
rect 10956 6842 11916 6880
rect 11974 6880 12176 6897
rect 12732 6897 12748 6914
rect 14196 6988 14212 7005
rect 14768 7005 14970 7022
rect 15028 7022 15988 7060
rect 15028 7005 15230 7022
rect 14768 6988 14784 7005
rect 14196 6972 14784 6988
rect 13178 6914 13766 6930
rect 13178 6897 13194 6914
rect 12732 6880 12934 6897
rect 11974 6842 12934 6880
rect 12992 6880 13194 6897
rect 13750 6897 13766 6914
rect 15214 6988 15230 7005
rect 15786 7005 15988 7022
rect 16046 7022 17006 7060
rect 16046 7005 16248 7022
rect 15786 6988 15802 7005
rect 15214 6972 15802 6988
rect 14196 6914 14784 6930
rect 14196 6897 14212 6914
rect 13750 6880 13952 6897
rect 12992 6842 13952 6880
rect 14010 6880 14212 6897
rect 14768 6897 14784 6914
rect 16232 6988 16248 7005
rect 16804 7005 17006 7022
rect 16804 6988 16820 7005
rect 16232 6972 16820 6988
rect 15214 6914 15802 6930
rect 15214 6897 15230 6914
rect 14768 6880 14970 6897
rect 14010 6842 14970 6880
rect 15028 6880 15230 6897
rect 15786 6897 15802 6914
rect 16232 6914 16820 6930
rect 16232 6897 16248 6914
rect 15786 6880 15988 6897
rect 15028 6842 15988 6880
rect 16046 6880 16248 6897
rect 16804 6897 16820 6914
rect 16804 6880 17006 6897
rect 16046 6842 17006 6880
rect 19666 6510 20626 6548
rect 19666 6493 19868 6510
rect 19852 6476 19868 6493
rect 20424 6493 20626 6510
rect 20684 6510 21644 6548
rect 20684 6493 20886 6510
rect 20424 6476 20440 6493
rect 19852 6460 20440 6476
rect 20870 6476 20886 6493
rect 21442 6493 21644 6510
rect 21702 6510 22662 6548
rect 21702 6493 21904 6510
rect 21442 6476 21458 6493
rect 20870 6460 21458 6476
rect 21888 6476 21904 6493
rect 22460 6493 22662 6510
rect 22720 6510 23680 6548
rect 22720 6493 22922 6510
rect 22460 6476 22476 6493
rect 21888 6460 22476 6476
rect 22906 6476 22922 6493
rect 23478 6493 23680 6510
rect 23738 6510 24698 6548
rect 23738 6493 23940 6510
rect 23478 6476 23494 6493
rect 22906 6460 23494 6476
rect 23924 6476 23940 6493
rect 24496 6493 24698 6510
rect 24756 6510 25716 6548
rect 24756 6493 24958 6510
rect 24496 6476 24512 6493
rect 23924 6460 24512 6476
rect 24942 6476 24958 6493
rect 25514 6493 25716 6510
rect 25774 6510 26734 6548
rect 25774 6493 25976 6510
rect 25514 6476 25530 6493
rect 24942 6460 25530 6476
rect 25960 6476 25976 6493
rect 26532 6493 26734 6510
rect 26792 6510 27752 6548
rect 26792 6493 26994 6510
rect 26532 6476 26548 6493
rect 25960 6460 26548 6476
rect 26978 6476 26994 6493
rect 27550 6493 27752 6510
rect 27810 6510 28770 6548
rect 27810 6493 28012 6510
rect 27550 6476 27566 6493
rect 26978 6460 27566 6476
rect 27996 6476 28012 6493
rect 28568 6493 28770 6510
rect 28828 6510 29788 6548
rect 28828 6493 29030 6510
rect 28568 6476 28584 6493
rect 27996 6460 28584 6476
rect 29014 6476 29030 6493
rect 29586 6493 29788 6510
rect 29846 6510 30806 6548
rect 29846 6493 30048 6510
rect 29586 6476 29602 6493
rect 29014 6460 29602 6476
rect 30032 6476 30048 6493
rect 30604 6493 30806 6510
rect 30864 6510 31824 6548
rect 30864 6493 31066 6510
rect 30604 6476 30620 6493
rect 30032 6460 30620 6476
rect 31050 6476 31066 6493
rect 31622 6493 31824 6510
rect 31882 6510 32842 6548
rect 31882 6493 32084 6510
rect 31622 6476 31638 6493
rect 31050 6460 31638 6476
rect 32068 6476 32084 6493
rect 32640 6493 32842 6510
rect 32900 6510 33860 6548
rect 32900 6493 33102 6510
rect 32640 6476 32656 6493
rect 32068 6460 32656 6476
rect 33086 6476 33102 6493
rect 33658 6493 33860 6510
rect 33918 6510 34878 6548
rect 33918 6493 34120 6510
rect 33658 6476 33674 6493
rect 33086 6460 33674 6476
rect 34104 6476 34120 6493
rect 34676 6493 34878 6510
rect 34936 6510 35896 6548
rect 34936 6493 35138 6510
rect 34676 6476 34692 6493
rect 34104 6460 34692 6476
rect 35122 6476 35138 6493
rect 35694 6493 35896 6510
rect 35954 6510 36914 6548
rect 35954 6493 36156 6510
rect 35694 6476 35710 6493
rect 35122 6460 35710 6476
rect 36140 6476 36156 6493
rect 36712 6493 36914 6510
rect 36972 6510 37932 6548
rect 36972 6493 37174 6510
rect 36712 6476 36728 6493
rect 36140 6460 36728 6476
rect 37158 6476 37174 6493
rect 37730 6493 37932 6510
rect 37990 6510 38950 6548
rect 37990 6493 38192 6510
rect 37730 6476 37746 6493
rect 37158 6460 37746 6476
rect 38176 6476 38192 6493
rect 38748 6493 38950 6510
rect 39008 6510 39968 6548
rect 39008 6493 39210 6510
rect 38748 6476 38764 6493
rect 38176 6460 38764 6476
rect 39194 6476 39210 6493
rect 39766 6493 39968 6510
rect 39766 6476 39782 6493
rect 39194 6460 39782 6476
rect 7902 6204 8862 6242
rect 7902 6187 8104 6204
rect 8088 6170 8104 6187
rect 8660 6187 8862 6204
rect 8920 6204 9880 6242
rect 8920 6187 9122 6204
rect 8660 6170 8676 6187
rect 8088 6154 8676 6170
rect 9106 6170 9122 6187
rect 9678 6187 9880 6204
rect 9938 6204 10898 6242
rect 9938 6187 10140 6204
rect 9678 6170 9694 6187
rect 9106 6154 9694 6170
rect 10124 6170 10140 6187
rect 10696 6187 10898 6204
rect 10956 6204 11916 6242
rect 10956 6187 11158 6204
rect 10696 6170 10712 6187
rect 10124 6154 10712 6170
rect 11142 6170 11158 6187
rect 11714 6187 11916 6204
rect 11974 6204 12934 6242
rect 11974 6187 12176 6204
rect 11714 6170 11730 6187
rect 11142 6154 11730 6170
rect 12160 6170 12176 6187
rect 12732 6187 12934 6204
rect 12992 6204 13952 6242
rect 12992 6187 13194 6204
rect 12732 6170 12748 6187
rect 12160 6154 12748 6170
rect 13178 6170 13194 6187
rect 13750 6187 13952 6204
rect 14010 6204 14970 6242
rect 14010 6187 14212 6204
rect 13750 6170 13766 6187
rect 13178 6154 13766 6170
rect 14196 6170 14212 6187
rect 14768 6187 14970 6204
rect 15028 6204 15988 6242
rect 15028 6187 15230 6204
rect 14768 6170 14784 6187
rect 14196 6154 14784 6170
rect 15214 6170 15230 6187
rect 15786 6187 15988 6204
rect 16046 6204 17006 6242
rect 16046 6187 16248 6204
rect 15786 6170 15802 6187
rect 15214 6154 15802 6170
rect 16232 6170 16248 6187
rect 16804 6187 17006 6204
rect 16804 6170 16820 6187
rect 16232 6154 16820 6170
rect 19852 5988 20440 6004
rect 19852 5971 19868 5988
rect 19666 5954 19868 5971
rect 20424 5971 20440 5988
rect 20870 5988 21458 6004
rect 20870 5971 20886 5988
rect 20424 5954 20626 5971
rect 19666 5916 20626 5954
rect 20684 5954 20886 5971
rect 21442 5971 21458 5988
rect 21888 5988 22476 6004
rect 21888 5971 21904 5988
rect 21442 5954 21644 5971
rect 20684 5916 21644 5954
rect 21702 5954 21904 5971
rect 22460 5971 22476 5988
rect 22906 5988 23494 6004
rect 22906 5971 22922 5988
rect 22460 5954 22662 5971
rect 21702 5916 22662 5954
rect 22720 5954 22922 5971
rect 23478 5971 23494 5988
rect 23924 5988 24512 6004
rect 23924 5971 23940 5988
rect 23478 5954 23680 5971
rect 22720 5916 23680 5954
rect 23738 5954 23940 5971
rect 24496 5971 24512 5988
rect 24942 5988 25530 6004
rect 24942 5971 24958 5988
rect 24496 5954 24698 5971
rect 23738 5916 24698 5954
rect 24756 5954 24958 5971
rect 25514 5971 25530 5988
rect 25960 5988 26548 6004
rect 25960 5971 25976 5988
rect 25514 5954 25716 5971
rect 24756 5916 25716 5954
rect 25774 5954 25976 5971
rect 26532 5971 26548 5988
rect 26978 5988 27566 6004
rect 26978 5971 26994 5988
rect 26532 5954 26734 5971
rect 25774 5916 26734 5954
rect 26792 5954 26994 5971
rect 27550 5971 27566 5988
rect 27996 5988 28584 6004
rect 27996 5971 28012 5988
rect 27550 5954 27752 5971
rect 26792 5916 27752 5954
rect 27810 5954 28012 5971
rect 28568 5971 28584 5988
rect 29014 5988 29602 6004
rect 29014 5971 29030 5988
rect 28568 5954 28770 5971
rect 27810 5916 28770 5954
rect 28828 5954 29030 5971
rect 29586 5971 29602 5988
rect 30032 5988 30620 6004
rect 30032 5971 30048 5988
rect 29586 5954 29788 5971
rect 28828 5916 29788 5954
rect 29846 5954 30048 5971
rect 30604 5971 30620 5988
rect 31050 5988 31638 6004
rect 31050 5971 31066 5988
rect 30604 5954 30806 5971
rect 29846 5916 30806 5954
rect 30864 5954 31066 5971
rect 31622 5971 31638 5988
rect 32068 5988 32656 6004
rect 32068 5971 32084 5988
rect 31622 5954 31824 5971
rect 30864 5916 31824 5954
rect 31882 5954 32084 5971
rect 32640 5971 32656 5988
rect 33086 5988 33674 6004
rect 33086 5971 33102 5988
rect 32640 5954 32842 5971
rect 31882 5916 32842 5954
rect 32900 5954 33102 5971
rect 33658 5971 33674 5988
rect 34104 5988 34692 6004
rect 34104 5971 34120 5988
rect 33658 5954 33860 5971
rect 32900 5916 33860 5954
rect 33918 5954 34120 5971
rect 34676 5971 34692 5988
rect 35122 5988 35710 6004
rect 35122 5971 35138 5988
rect 34676 5954 34878 5971
rect 33918 5916 34878 5954
rect 34936 5954 35138 5971
rect 35694 5971 35710 5988
rect 36140 5988 36728 6004
rect 36140 5971 36156 5988
rect 35694 5954 35896 5971
rect 34936 5916 35896 5954
rect 35954 5954 36156 5971
rect 36712 5971 36728 5988
rect 37158 5988 37746 6004
rect 37158 5971 37174 5988
rect 36712 5954 36914 5971
rect 35954 5916 36914 5954
rect 36972 5954 37174 5971
rect 37730 5971 37746 5988
rect 38176 5988 38764 6004
rect 38176 5971 38192 5988
rect 37730 5954 37932 5971
rect 36972 5916 37932 5954
rect 37990 5954 38192 5971
rect 38748 5971 38764 5988
rect 39194 5988 39782 6004
rect 39194 5971 39210 5988
rect 38748 5954 38950 5971
rect 37990 5916 38950 5954
rect 39008 5954 39210 5971
rect 39766 5971 39782 5988
rect 39766 5954 39968 5971
rect 39008 5916 39968 5954
rect 19666 5278 20626 5316
rect 19666 5261 19868 5278
rect 19852 5244 19868 5261
rect 20424 5261 20626 5278
rect 20684 5278 21644 5316
rect 20684 5261 20886 5278
rect 20424 5244 20440 5261
rect 19852 5228 20440 5244
rect 20870 5244 20886 5261
rect 21442 5261 21644 5278
rect 21702 5278 22662 5316
rect 21702 5261 21904 5278
rect 21442 5244 21458 5261
rect 20870 5228 21458 5244
rect 21888 5244 21904 5261
rect 22460 5261 22662 5278
rect 22720 5278 23680 5316
rect 22720 5261 22922 5278
rect 22460 5244 22476 5261
rect 21888 5228 22476 5244
rect 22906 5244 22922 5261
rect 23478 5261 23680 5278
rect 23738 5278 24698 5316
rect 23738 5261 23940 5278
rect 23478 5244 23494 5261
rect 22906 5228 23494 5244
rect 23924 5244 23940 5261
rect 24496 5261 24698 5278
rect 24756 5278 25716 5316
rect 24756 5261 24958 5278
rect 24496 5244 24512 5261
rect 23924 5228 24512 5244
rect 24942 5244 24958 5261
rect 25514 5261 25716 5278
rect 25774 5278 26734 5316
rect 25774 5261 25976 5278
rect 25514 5244 25530 5261
rect 24942 5228 25530 5244
rect 25960 5244 25976 5261
rect 26532 5261 26734 5278
rect 26792 5278 27752 5316
rect 26792 5261 26994 5278
rect 26532 5244 26548 5261
rect 25960 5228 26548 5244
rect 26978 5244 26994 5261
rect 27550 5261 27752 5278
rect 27810 5278 28770 5316
rect 27810 5261 28012 5278
rect 27550 5244 27566 5261
rect 26978 5228 27566 5244
rect 27996 5244 28012 5261
rect 28568 5261 28770 5278
rect 28828 5278 29788 5316
rect 28828 5261 29030 5278
rect 28568 5244 28584 5261
rect 27996 5228 28584 5244
rect 29014 5244 29030 5261
rect 29586 5261 29788 5278
rect 29846 5278 30806 5316
rect 29846 5261 30048 5278
rect 29586 5244 29602 5261
rect 29014 5228 29602 5244
rect 30032 5244 30048 5261
rect 30604 5261 30806 5278
rect 30864 5278 31824 5316
rect 30864 5261 31066 5278
rect 30604 5244 30620 5261
rect 30032 5228 30620 5244
rect 31050 5244 31066 5261
rect 31622 5261 31824 5278
rect 31882 5278 32842 5316
rect 31882 5261 32084 5278
rect 31622 5244 31638 5261
rect 31050 5228 31638 5244
rect 32068 5244 32084 5261
rect 32640 5261 32842 5278
rect 32900 5278 33860 5316
rect 32900 5261 33102 5278
rect 32640 5244 32656 5261
rect 32068 5228 32656 5244
rect 33086 5244 33102 5261
rect 33658 5261 33860 5278
rect 33918 5278 34878 5316
rect 33918 5261 34120 5278
rect 33658 5244 33674 5261
rect 33086 5228 33674 5244
rect 34104 5244 34120 5261
rect 34676 5261 34878 5278
rect 34936 5278 35896 5316
rect 34936 5261 35138 5278
rect 34676 5244 34692 5261
rect 34104 5228 34692 5244
rect 35122 5244 35138 5261
rect 35694 5261 35896 5278
rect 35954 5278 36914 5316
rect 35954 5261 36156 5278
rect 35694 5244 35710 5261
rect 35122 5228 35710 5244
rect 36140 5244 36156 5261
rect 36712 5261 36914 5278
rect 36972 5278 37932 5316
rect 36972 5261 37174 5278
rect 36712 5244 36728 5261
rect 36140 5228 36728 5244
rect 37158 5244 37174 5261
rect 37730 5261 37932 5278
rect 37990 5278 38950 5316
rect 37990 5261 38192 5278
rect 37730 5244 37746 5261
rect 37158 5228 37746 5244
rect 38176 5244 38192 5261
rect 38748 5261 38950 5278
rect 39008 5278 39968 5316
rect 39008 5261 39210 5278
rect 38748 5244 38764 5261
rect 38176 5228 38764 5244
rect 39194 5244 39210 5261
rect 39766 5261 39968 5278
rect 39766 5244 39782 5261
rect 39194 5228 39782 5244
rect 6764 4890 7352 4906
rect 6764 4873 6780 4890
rect 6578 4856 6780 4873
rect 7336 4873 7352 4890
rect 7782 4890 8370 4906
rect 7782 4873 7798 4890
rect 7336 4856 7538 4873
rect 6578 4818 7538 4856
rect 7596 4856 7798 4873
rect 8354 4873 8370 4890
rect 8800 4890 9388 4906
rect 8800 4873 8816 4890
rect 8354 4856 8556 4873
rect 7596 4818 8556 4856
rect 8614 4856 8816 4873
rect 9372 4873 9388 4890
rect 9818 4890 10406 4906
rect 9818 4873 9834 4890
rect 9372 4856 9574 4873
rect 8614 4818 9574 4856
rect 9632 4856 9834 4873
rect 10390 4873 10406 4890
rect 10836 4890 11424 4906
rect 10836 4873 10852 4890
rect 10390 4856 10592 4873
rect 9632 4818 10592 4856
rect 10650 4856 10852 4873
rect 11408 4873 11424 4890
rect 11854 4890 12442 4906
rect 11854 4873 11870 4890
rect 11408 4856 11610 4873
rect 10650 4818 11610 4856
rect 11668 4856 11870 4873
rect 12426 4873 12442 4890
rect 12872 4890 13460 4906
rect 12872 4873 12888 4890
rect 12426 4856 12628 4873
rect 11668 4818 12628 4856
rect 12686 4856 12888 4873
rect 13444 4873 13460 4890
rect 13890 4890 14478 4906
rect 13890 4873 13906 4890
rect 13444 4856 13646 4873
rect 12686 4818 13646 4856
rect 13704 4856 13906 4873
rect 14462 4873 14478 4890
rect 14908 4890 15496 4906
rect 14908 4873 14924 4890
rect 14462 4856 14664 4873
rect 13704 4818 14664 4856
rect 14722 4856 14924 4873
rect 15480 4873 15496 4890
rect 15926 4890 16514 4906
rect 15926 4873 15942 4890
rect 15480 4856 15682 4873
rect 14722 4818 15682 4856
rect 15740 4856 15942 4873
rect 16498 4873 16514 4890
rect 16944 4890 17532 4906
rect 16944 4873 16960 4890
rect 16498 4856 16700 4873
rect 15740 4818 16700 4856
rect 16758 4856 16960 4873
rect 17516 4873 17532 4890
rect 17516 4856 17718 4873
rect 16758 4818 17718 4856
rect 19852 4754 20440 4770
rect 19852 4737 19868 4754
rect 19666 4720 19868 4737
rect 20424 4737 20440 4754
rect 20870 4754 21458 4770
rect 20870 4737 20886 4754
rect 20424 4720 20626 4737
rect 19666 4682 20626 4720
rect 20684 4720 20886 4737
rect 21442 4737 21458 4754
rect 21888 4754 22476 4770
rect 21888 4737 21904 4754
rect 21442 4720 21644 4737
rect 20684 4682 21644 4720
rect 21702 4720 21904 4737
rect 22460 4737 22476 4754
rect 22906 4754 23494 4770
rect 22906 4737 22922 4754
rect 22460 4720 22662 4737
rect 21702 4682 22662 4720
rect 22720 4720 22922 4737
rect 23478 4737 23494 4754
rect 23924 4754 24512 4770
rect 23924 4737 23940 4754
rect 23478 4720 23680 4737
rect 22720 4682 23680 4720
rect 23738 4720 23940 4737
rect 24496 4737 24512 4754
rect 24942 4754 25530 4770
rect 24942 4737 24958 4754
rect 24496 4720 24698 4737
rect 23738 4682 24698 4720
rect 24756 4720 24958 4737
rect 25514 4737 25530 4754
rect 25960 4754 26548 4770
rect 25960 4737 25976 4754
rect 25514 4720 25716 4737
rect 24756 4682 25716 4720
rect 25774 4720 25976 4737
rect 26532 4737 26548 4754
rect 26978 4754 27566 4770
rect 26978 4737 26994 4754
rect 26532 4720 26734 4737
rect 25774 4682 26734 4720
rect 26792 4720 26994 4737
rect 27550 4737 27566 4754
rect 27996 4754 28584 4770
rect 27996 4737 28012 4754
rect 27550 4720 27752 4737
rect 26792 4682 27752 4720
rect 27810 4720 28012 4737
rect 28568 4737 28584 4754
rect 29014 4754 29602 4770
rect 29014 4737 29030 4754
rect 28568 4720 28770 4737
rect 27810 4682 28770 4720
rect 28828 4720 29030 4737
rect 29586 4737 29602 4754
rect 30032 4754 30620 4770
rect 30032 4737 30048 4754
rect 29586 4720 29788 4737
rect 28828 4682 29788 4720
rect 29846 4720 30048 4737
rect 30604 4737 30620 4754
rect 31050 4754 31638 4770
rect 31050 4737 31066 4754
rect 30604 4720 30806 4737
rect 29846 4682 30806 4720
rect 30864 4720 31066 4737
rect 31622 4737 31638 4754
rect 32068 4754 32656 4770
rect 32068 4737 32084 4754
rect 31622 4720 31824 4737
rect 30864 4682 31824 4720
rect 31882 4720 32084 4737
rect 32640 4737 32656 4754
rect 33086 4754 33674 4770
rect 33086 4737 33102 4754
rect 32640 4720 32842 4737
rect 31882 4682 32842 4720
rect 32900 4720 33102 4737
rect 33658 4737 33674 4754
rect 34104 4754 34692 4770
rect 34104 4737 34120 4754
rect 33658 4720 33860 4737
rect 32900 4682 33860 4720
rect 33918 4720 34120 4737
rect 34676 4737 34692 4754
rect 35122 4754 35710 4770
rect 35122 4737 35138 4754
rect 34676 4720 34878 4737
rect 33918 4682 34878 4720
rect 34936 4720 35138 4737
rect 35694 4737 35710 4754
rect 36140 4754 36728 4770
rect 36140 4737 36156 4754
rect 35694 4720 35896 4737
rect 34936 4682 35896 4720
rect 35954 4720 36156 4737
rect 36712 4737 36728 4754
rect 37158 4754 37746 4770
rect 37158 4737 37174 4754
rect 36712 4720 36914 4737
rect 35954 4682 36914 4720
rect 36972 4720 37174 4737
rect 37730 4737 37746 4754
rect 38176 4754 38764 4770
rect 38176 4737 38192 4754
rect 37730 4720 37932 4737
rect 36972 4682 37932 4720
rect 37990 4720 38192 4737
rect 38748 4737 38764 4754
rect 39194 4754 39782 4770
rect 39194 4737 39210 4754
rect 38748 4720 38950 4737
rect 37990 4682 38950 4720
rect 39008 4720 39210 4737
rect 39766 4737 39782 4754
rect 39766 4720 39968 4737
rect 39008 4682 39968 4720
rect 6578 4180 7538 4218
rect 6578 4163 6780 4180
rect 6764 4146 6780 4163
rect 7336 4163 7538 4180
rect 7596 4180 8556 4218
rect 7596 4163 7798 4180
rect 7336 4146 7352 4163
rect 6764 4130 7352 4146
rect 7782 4146 7798 4163
rect 8354 4163 8556 4180
rect 8614 4180 9574 4218
rect 8614 4163 8816 4180
rect 8354 4146 8370 4163
rect 7782 4130 8370 4146
rect 8800 4146 8816 4163
rect 9372 4163 9574 4180
rect 9632 4180 10592 4218
rect 9632 4163 9834 4180
rect 9372 4146 9388 4163
rect 8800 4130 9388 4146
rect 9818 4146 9834 4163
rect 10390 4163 10592 4180
rect 10650 4180 11610 4218
rect 10650 4163 10852 4180
rect 10390 4146 10406 4163
rect 9818 4130 10406 4146
rect 10836 4146 10852 4163
rect 11408 4163 11610 4180
rect 11668 4180 12628 4218
rect 11668 4163 11870 4180
rect 11408 4146 11424 4163
rect 10836 4130 11424 4146
rect 11854 4146 11870 4163
rect 12426 4163 12628 4180
rect 12686 4180 13646 4218
rect 12686 4163 12888 4180
rect 12426 4146 12442 4163
rect 11854 4130 12442 4146
rect 12872 4146 12888 4163
rect 13444 4163 13646 4180
rect 13704 4180 14664 4218
rect 13704 4163 13906 4180
rect 13444 4146 13460 4163
rect 12872 4130 13460 4146
rect 13890 4146 13906 4163
rect 14462 4163 14664 4180
rect 14722 4180 15682 4218
rect 14722 4163 14924 4180
rect 14462 4146 14478 4163
rect 13890 4130 14478 4146
rect 14908 4146 14924 4163
rect 15480 4163 15682 4180
rect 15740 4180 16700 4218
rect 15740 4163 15942 4180
rect 15480 4146 15496 4163
rect 14908 4130 15496 4146
rect 15926 4146 15942 4163
rect 16498 4163 16700 4180
rect 16758 4180 17718 4218
rect 16758 4163 16960 4180
rect 16498 4146 16514 4163
rect 15926 4130 16514 4146
rect 16944 4146 16960 4163
rect 17516 4163 17718 4180
rect 17516 4146 17532 4163
rect 16944 4130 17532 4146
rect 19666 4044 20626 4082
rect 19666 4027 19868 4044
rect 19852 4010 19868 4027
rect 20424 4027 20626 4044
rect 20684 4044 21644 4082
rect 20684 4027 20886 4044
rect 20424 4010 20440 4027
rect 19852 3994 20440 4010
rect 20870 4010 20886 4027
rect 21442 4027 21644 4044
rect 21702 4044 22662 4082
rect 21702 4027 21904 4044
rect 21442 4010 21458 4027
rect 20870 3994 21458 4010
rect 21888 4010 21904 4027
rect 22460 4027 22662 4044
rect 22720 4044 23680 4082
rect 22720 4027 22922 4044
rect 22460 4010 22476 4027
rect 21888 3994 22476 4010
rect 22906 4010 22922 4027
rect 23478 4027 23680 4044
rect 23738 4044 24698 4082
rect 23738 4027 23940 4044
rect 23478 4010 23494 4027
rect 22906 3994 23494 4010
rect 23924 4010 23940 4027
rect 24496 4027 24698 4044
rect 24756 4044 25716 4082
rect 24756 4027 24958 4044
rect 24496 4010 24512 4027
rect 23924 3994 24512 4010
rect 24942 4010 24958 4027
rect 25514 4027 25716 4044
rect 25774 4044 26734 4082
rect 25774 4027 25976 4044
rect 25514 4010 25530 4027
rect 24942 3994 25530 4010
rect 25960 4010 25976 4027
rect 26532 4027 26734 4044
rect 26792 4044 27752 4082
rect 26792 4027 26994 4044
rect 26532 4010 26548 4027
rect 25960 3994 26548 4010
rect 26978 4010 26994 4027
rect 27550 4027 27752 4044
rect 27810 4044 28770 4082
rect 27810 4027 28012 4044
rect 27550 4010 27566 4027
rect 26978 3994 27566 4010
rect 27996 4010 28012 4027
rect 28568 4027 28770 4044
rect 28828 4044 29788 4082
rect 28828 4027 29030 4044
rect 28568 4010 28584 4027
rect 27996 3994 28584 4010
rect 29014 4010 29030 4027
rect 29586 4027 29788 4044
rect 29846 4044 30806 4082
rect 29846 4027 30048 4044
rect 29586 4010 29602 4027
rect 29014 3994 29602 4010
rect 30032 4010 30048 4027
rect 30604 4027 30806 4044
rect 30864 4044 31824 4082
rect 30864 4027 31066 4044
rect 30604 4010 30620 4027
rect 30032 3994 30620 4010
rect 31050 4010 31066 4027
rect 31622 4027 31824 4044
rect 31882 4044 32842 4082
rect 31882 4027 32084 4044
rect 31622 4010 31638 4027
rect 31050 3994 31638 4010
rect 32068 4010 32084 4027
rect 32640 4027 32842 4044
rect 32900 4044 33860 4082
rect 32900 4027 33102 4044
rect 32640 4010 32656 4027
rect 32068 3994 32656 4010
rect 33086 4010 33102 4027
rect 33658 4027 33860 4044
rect 33918 4044 34878 4082
rect 33918 4027 34120 4044
rect 33658 4010 33674 4027
rect 33086 3994 33674 4010
rect 34104 4010 34120 4027
rect 34676 4027 34878 4044
rect 34936 4044 35896 4082
rect 34936 4027 35138 4044
rect 34676 4010 34692 4027
rect 34104 3994 34692 4010
rect 35122 4010 35138 4027
rect 35694 4027 35896 4044
rect 35954 4044 36914 4082
rect 35954 4027 36156 4044
rect 35694 4010 35710 4027
rect 35122 3994 35710 4010
rect 36140 4010 36156 4027
rect 36712 4027 36914 4044
rect 36972 4044 37932 4082
rect 36972 4027 37174 4044
rect 36712 4010 36728 4027
rect 36140 3994 36728 4010
rect 37158 4010 37174 4027
rect 37730 4027 37932 4044
rect 37990 4044 38950 4082
rect 37990 4027 38192 4044
rect 37730 4010 37746 4027
rect 37158 3994 37746 4010
rect 38176 4010 38192 4027
rect 38748 4027 38950 4044
rect 39008 4044 39968 4082
rect 39008 4027 39210 4044
rect 38748 4010 38764 4027
rect 38176 3994 38764 4010
rect 39194 4010 39210 4027
rect 39766 4027 39968 4044
rect 39766 4010 39782 4027
rect 39194 3994 39782 4010
rect 6764 3778 7352 3794
rect 6764 3761 6780 3778
rect 6578 3744 6780 3761
rect 7336 3761 7352 3778
rect 7782 3778 8370 3794
rect 7782 3761 7798 3778
rect 7336 3744 7538 3761
rect 6578 3706 7538 3744
rect 7596 3744 7798 3761
rect 8354 3761 8370 3778
rect 8800 3778 9388 3794
rect 8800 3761 8816 3778
rect 8354 3744 8556 3761
rect 7596 3706 8556 3744
rect 8614 3744 8816 3761
rect 9372 3761 9388 3778
rect 9818 3778 10406 3794
rect 9818 3761 9834 3778
rect 9372 3744 9574 3761
rect 8614 3706 9574 3744
rect 9632 3744 9834 3761
rect 10390 3761 10406 3778
rect 10836 3778 11424 3794
rect 10836 3761 10852 3778
rect 10390 3744 10592 3761
rect 9632 3706 10592 3744
rect 10650 3744 10852 3761
rect 11408 3761 11424 3778
rect 11854 3778 12442 3794
rect 11854 3761 11870 3778
rect 11408 3744 11610 3761
rect 10650 3706 11610 3744
rect 11668 3744 11870 3761
rect 12426 3761 12442 3778
rect 12872 3778 13460 3794
rect 12872 3761 12888 3778
rect 12426 3744 12628 3761
rect 11668 3706 12628 3744
rect 12686 3744 12888 3761
rect 13444 3761 13460 3778
rect 13890 3778 14478 3794
rect 13890 3761 13906 3778
rect 13444 3744 13646 3761
rect 12686 3706 13646 3744
rect 13704 3744 13906 3761
rect 14462 3761 14478 3778
rect 14908 3778 15496 3794
rect 14908 3761 14924 3778
rect 14462 3744 14664 3761
rect 13704 3706 14664 3744
rect 14722 3744 14924 3761
rect 15480 3761 15496 3778
rect 15926 3778 16514 3794
rect 15926 3761 15942 3778
rect 15480 3744 15682 3761
rect 14722 3706 15682 3744
rect 15740 3744 15942 3761
rect 16498 3761 16514 3778
rect 16944 3778 17532 3794
rect 16944 3761 16960 3778
rect 16498 3744 16700 3761
rect 15740 3706 16700 3744
rect 16758 3744 16960 3761
rect 17516 3761 17532 3778
rect 17516 3744 17718 3761
rect 16758 3706 17718 3744
rect 19852 3520 20440 3536
rect 19852 3503 19868 3520
rect 19666 3486 19868 3503
rect 20424 3503 20440 3520
rect 20870 3520 21458 3536
rect 20870 3503 20886 3520
rect 20424 3486 20626 3503
rect 19666 3448 20626 3486
rect 20684 3486 20886 3503
rect 21442 3503 21458 3520
rect 21888 3520 22476 3536
rect 21888 3503 21904 3520
rect 21442 3486 21644 3503
rect 20684 3448 21644 3486
rect 21702 3486 21904 3503
rect 22460 3503 22476 3520
rect 22906 3520 23494 3536
rect 22906 3503 22922 3520
rect 22460 3486 22662 3503
rect 21702 3448 22662 3486
rect 22720 3486 22922 3503
rect 23478 3503 23494 3520
rect 23924 3520 24512 3536
rect 23924 3503 23940 3520
rect 23478 3486 23680 3503
rect 22720 3448 23680 3486
rect 23738 3486 23940 3503
rect 24496 3503 24512 3520
rect 24942 3520 25530 3536
rect 24942 3503 24958 3520
rect 24496 3486 24698 3503
rect 23738 3448 24698 3486
rect 24756 3486 24958 3503
rect 25514 3503 25530 3520
rect 25960 3520 26548 3536
rect 25960 3503 25976 3520
rect 25514 3486 25716 3503
rect 24756 3448 25716 3486
rect 25774 3486 25976 3503
rect 26532 3503 26548 3520
rect 26978 3520 27566 3536
rect 26978 3503 26994 3520
rect 26532 3486 26734 3503
rect 25774 3448 26734 3486
rect 26792 3486 26994 3503
rect 27550 3503 27566 3520
rect 27996 3520 28584 3536
rect 27996 3503 28012 3520
rect 27550 3486 27752 3503
rect 26792 3448 27752 3486
rect 27810 3486 28012 3503
rect 28568 3503 28584 3520
rect 29014 3520 29602 3536
rect 29014 3503 29030 3520
rect 28568 3486 28770 3503
rect 27810 3448 28770 3486
rect 28828 3486 29030 3503
rect 29586 3503 29602 3520
rect 30032 3520 30620 3536
rect 30032 3503 30048 3520
rect 29586 3486 29788 3503
rect 28828 3448 29788 3486
rect 29846 3486 30048 3503
rect 30604 3503 30620 3520
rect 31050 3520 31638 3536
rect 31050 3503 31066 3520
rect 30604 3486 30806 3503
rect 29846 3448 30806 3486
rect 30864 3486 31066 3503
rect 31622 3503 31638 3520
rect 32068 3520 32656 3536
rect 32068 3503 32084 3520
rect 31622 3486 31824 3503
rect 30864 3448 31824 3486
rect 31882 3486 32084 3503
rect 32640 3503 32656 3520
rect 33086 3520 33674 3536
rect 33086 3503 33102 3520
rect 32640 3486 32842 3503
rect 31882 3448 32842 3486
rect 32900 3486 33102 3503
rect 33658 3503 33674 3520
rect 34104 3520 34692 3536
rect 34104 3503 34120 3520
rect 33658 3486 33860 3503
rect 32900 3448 33860 3486
rect 33918 3486 34120 3503
rect 34676 3503 34692 3520
rect 35122 3520 35710 3536
rect 35122 3503 35138 3520
rect 34676 3486 34878 3503
rect 33918 3448 34878 3486
rect 34936 3486 35138 3503
rect 35694 3503 35710 3520
rect 36140 3520 36728 3536
rect 36140 3503 36156 3520
rect 35694 3486 35896 3503
rect 34936 3448 35896 3486
rect 35954 3486 36156 3503
rect 36712 3503 36728 3520
rect 37158 3520 37746 3536
rect 37158 3503 37174 3520
rect 36712 3486 36914 3503
rect 35954 3448 36914 3486
rect 36972 3486 37174 3503
rect 37730 3503 37746 3520
rect 38176 3520 38764 3536
rect 38176 3503 38192 3520
rect 37730 3486 37932 3503
rect 36972 3448 37932 3486
rect 37990 3486 38192 3503
rect 38748 3503 38764 3520
rect 39194 3520 39782 3536
rect 39194 3503 39210 3520
rect 38748 3486 38950 3503
rect 37990 3448 38950 3486
rect 39008 3486 39210 3503
rect 39766 3503 39782 3520
rect 39766 3486 39968 3503
rect 39008 3448 39968 3486
rect 6578 3068 7538 3106
rect 6578 3051 6780 3068
rect 6764 3034 6780 3051
rect 7336 3051 7538 3068
rect 7596 3068 8556 3106
rect 7596 3051 7798 3068
rect 7336 3034 7352 3051
rect 6764 3018 7352 3034
rect 7782 3034 7798 3051
rect 8354 3051 8556 3068
rect 8614 3068 9574 3106
rect 8614 3051 8816 3068
rect 8354 3034 8370 3051
rect 7782 3018 8370 3034
rect 8800 3034 8816 3051
rect 9372 3051 9574 3068
rect 9632 3068 10592 3106
rect 9632 3051 9834 3068
rect 9372 3034 9388 3051
rect 8800 3018 9388 3034
rect 9818 3034 9834 3051
rect 10390 3051 10592 3068
rect 10650 3068 11610 3106
rect 10650 3051 10852 3068
rect 10390 3034 10406 3051
rect 9818 3018 10406 3034
rect 10836 3034 10852 3051
rect 11408 3051 11610 3068
rect 11668 3068 12628 3106
rect 11668 3051 11870 3068
rect 11408 3034 11424 3051
rect 10836 3018 11424 3034
rect 11854 3034 11870 3051
rect 12426 3051 12628 3068
rect 12686 3068 13646 3106
rect 12686 3051 12888 3068
rect 12426 3034 12442 3051
rect 11854 3018 12442 3034
rect 12872 3034 12888 3051
rect 13444 3051 13646 3068
rect 13704 3068 14664 3106
rect 13704 3051 13906 3068
rect 13444 3034 13460 3051
rect 12872 3018 13460 3034
rect 13890 3034 13906 3051
rect 14462 3051 14664 3068
rect 14722 3068 15682 3106
rect 14722 3051 14924 3068
rect 14462 3034 14478 3051
rect 13890 3018 14478 3034
rect 14908 3034 14924 3051
rect 15480 3051 15682 3068
rect 15740 3068 16700 3106
rect 15740 3051 15942 3068
rect 15480 3034 15496 3051
rect 14908 3018 15496 3034
rect 15926 3034 15942 3051
rect 16498 3051 16700 3068
rect 16758 3068 17718 3106
rect 16758 3051 16960 3068
rect 16498 3034 16514 3051
rect 15926 3018 16514 3034
rect 16944 3034 16960 3051
rect 17516 3051 17718 3068
rect 17516 3034 17532 3051
rect 16944 3018 17532 3034
rect 19666 2810 20626 2848
rect 19666 2793 19868 2810
rect 19852 2776 19868 2793
rect 20424 2793 20626 2810
rect 20684 2810 21644 2848
rect 20684 2793 20886 2810
rect 20424 2776 20440 2793
rect 19852 2760 20440 2776
rect 20870 2776 20886 2793
rect 21442 2793 21644 2810
rect 21702 2810 22662 2848
rect 21702 2793 21904 2810
rect 21442 2776 21458 2793
rect 20870 2760 21458 2776
rect 21888 2776 21904 2793
rect 22460 2793 22662 2810
rect 22720 2810 23680 2848
rect 22720 2793 22922 2810
rect 22460 2776 22476 2793
rect 21888 2760 22476 2776
rect 22906 2776 22922 2793
rect 23478 2793 23680 2810
rect 23738 2810 24698 2848
rect 23738 2793 23940 2810
rect 23478 2776 23494 2793
rect 22906 2760 23494 2776
rect 23924 2776 23940 2793
rect 24496 2793 24698 2810
rect 24756 2810 25716 2848
rect 24756 2793 24958 2810
rect 24496 2776 24512 2793
rect 23924 2760 24512 2776
rect 24942 2776 24958 2793
rect 25514 2793 25716 2810
rect 25774 2810 26734 2848
rect 25774 2793 25976 2810
rect 25514 2776 25530 2793
rect 24942 2760 25530 2776
rect 25960 2776 25976 2793
rect 26532 2793 26734 2810
rect 26792 2810 27752 2848
rect 26792 2793 26994 2810
rect 26532 2776 26548 2793
rect 25960 2760 26548 2776
rect 26978 2776 26994 2793
rect 27550 2793 27752 2810
rect 27810 2810 28770 2848
rect 27810 2793 28012 2810
rect 27550 2776 27566 2793
rect 26978 2760 27566 2776
rect 27996 2776 28012 2793
rect 28568 2793 28770 2810
rect 28828 2810 29788 2848
rect 28828 2793 29030 2810
rect 28568 2776 28584 2793
rect 27996 2760 28584 2776
rect 29014 2776 29030 2793
rect 29586 2793 29788 2810
rect 29846 2810 30806 2848
rect 29846 2793 30048 2810
rect 29586 2776 29602 2793
rect 29014 2760 29602 2776
rect 30032 2776 30048 2793
rect 30604 2793 30806 2810
rect 30864 2810 31824 2848
rect 30864 2793 31066 2810
rect 30604 2776 30620 2793
rect 30032 2760 30620 2776
rect 31050 2776 31066 2793
rect 31622 2793 31824 2810
rect 31882 2810 32842 2848
rect 31882 2793 32084 2810
rect 31622 2776 31638 2793
rect 31050 2760 31638 2776
rect 32068 2776 32084 2793
rect 32640 2793 32842 2810
rect 32900 2810 33860 2848
rect 32900 2793 33102 2810
rect 32640 2776 32656 2793
rect 32068 2760 32656 2776
rect 33086 2776 33102 2793
rect 33658 2793 33860 2810
rect 33918 2810 34878 2848
rect 33918 2793 34120 2810
rect 33658 2776 33674 2793
rect 33086 2760 33674 2776
rect 34104 2776 34120 2793
rect 34676 2793 34878 2810
rect 34936 2810 35896 2848
rect 34936 2793 35138 2810
rect 34676 2776 34692 2793
rect 34104 2760 34692 2776
rect 35122 2776 35138 2793
rect 35694 2793 35896 2810
rect 35954 2810 36914 2848
rect 35954 2793 36156 2810
rect 35694 2776 35710 2793
rect 35122 2760 35710 2776
rect 36140 2776 36156 2793
rect 36712 2793 36914 2810
rect 36972 2810 37932 2848
rect 36972 2793 37174 2810
rect 36712 2776 36728 2793
rect 36140 2760 36728 2776
rect 37158 2776 37174 2793
rect 37730 2793 37932 2810
rect 37990 2810 38950 2848
rect 37990 2793 38192 2810
rect 37730 2776 37746 2793
rect 37158 2760 37746 2776
rect 38176 2776 38192 2793
rect 38748 2793 38950 2810
rect 39008 2810 39968 2848
rect 39008 2793 39210 2810
rect 38748 2776 38764 2793
rect 38176 2760 38764 2776
rect 39194 2776 39210 2793
rect 39766 2793 39968 2810
rect 39766 2776 39782 2793
rect 39194 2760 39782 2776
rect 6764 2666 7352 2682
rect 6764 2649 6780 2666
rect 6578 2632 6780 2649
rect 7336 2649 7352 2666
rect 7782 2666 8370 2682
rect 7782 2649 7798 2666
rect 7336 2632 7538 2649
rect 6578 2594 7538 2632
rect 7596 2632 7798 2649
rect 8354 2649 8370 2666
rect 8800 2666 9388 2682
rect 8800 2649 8816 2666
rect 8354 2632 8556 2649
rect 7596 2594 8556 2632
rect 8614 2632 8816 2649
rect 9372 2649 9388 2666
rect 9818 2666 10406 2682
rect 9818 2649 9834 2666
rect 9372 2632 9574 2649
rect 8614 2594 9574 2632
rect 9632 2632 9834 2649
rect 10390 2649 10406 2666
rect 10836 2666 11424 2682
rect 10836 2649 10852 2666
rect 10390 2632 10592 2649
rect 9632 2594 10592 2632
rect 10650 2632 10852 2649
rect 11408 2649 11424 2666
rect 11854 2666 12442 2682
rect 11854 2649 11870 2666
rect 11408 2632 11610 2649
rect 10650 2594 11610 2632
rect 11668 2632 11870 2649
rect 12426 2649 12442 2666
rect 12872 2666 13460 2682
rect 12872 2649 12888 2666
rect 12426 2632 12628 2649
rect 11668 2594 12628 2632
rect 12686 2632 12888 2649
rect 13444 2649 13460 2666
rect 13890 2666 14478 2682
rect 13890 2649 13906 2666
rect 13444 2632 13646 2649
rect 12686 2594 13646 2632
rect 13704 2632 13906 2649
rect 14462 2649 14478 2666
rect 14908 2666 15496 2682
rect 14908 2649 14924 2666
rect 14462 2632 14664 2649
rect 13704 2594 14664 2632
rect 14722 2632 14924 2649
rect 15480 2649 15496 2666
rect 15926 2666 16514 2682
rect 15926 2649 15942 2666
rect 15480 2632 15682 2649
rect 14722 2594 15682 2632
rect 15740 2632 15942 2649
rect 16498 2649 16514 2666
rect 16944 2666 17532 2682
rect 16944 2649 16960 2666
rect 16498 2632 16700 2649
rect 15740 2594 16700 2632
rect 16758 2632 16960 2649
rect 17516 2649 17532 2666
rect 17516 2632 17718 2649
rect 16758 2594 17718 2632
rect 19852 2288 20440 2304
rect 19852 2271 19868 2288
rect 19666 2254 19868 2271
rect 20424 2271 20440 2288
rect 20870 2288 21458 2304
rect 20870 2271 20886 2288
rect 20424 2254 20626 2271
rect 19666 2216 20626 2254
rect 20684 2254 20886 2271
rect 21442 2271 21458 2288
rect 21888 2288 22476 2304
rect 21888 2271 21904 2288
rect 21442 2254 21644 2271
rect 20684 2216 21644 2254
rect 21702 2254 21904 2271
rect 22460 2271 22476 2288
rect 22906 2288 23494 2304
rect 22906 2271 22922 2288
rect 22460 2254 22662 2271
rect 21702 2216 22662 2254
rect 22720 2254 22922 2271
rect 23478 2271 23494 2288
rect 23924 2288 24512 2304
rect 23924 2271 23940 2288
rect 23478 2254 23680 2271
rect 22720 2216 23680 2254
rect 23738 2254 23940 2271
rect 24496 2271 24512 2288
rect 24942 2288 25530 2304
rect 24942 2271 24958 2288
rect 24496 2254 24698 2271
rect 23738 2216 24698 2254
rect 24756 2254 24958 2271
rect 25514 2271 25530 2288
rect 25960 2288 26548 2304
rect 25960 2271 25976 2288
rect 25514 2254 25716 2271
rect 24756 2216 25716 2254
rect 25774 2254 25976 2271
rect 26532 2271 26548 2288
rect 26978 2288 27566 2304
rect 26978 2271 26994 2288
rect 26532 2254 26734 2271
rect 25774 2216 26734 2254
rect 26792 2254 26994 2271
rect 27550 2271 27566 2288
rect 27996 2288 28584 2304
rect 27996 2271 28012 2288
rect 27550 2254 27752 2271
rect 26792 2216 27752 2254
rect 27810 2254 28012 2271
rect 28568 2271 28584 2288
rect 29014 2288 29602 2304
rect 29014 2271 29030 2288
rect 28568 2254 28770 2271
rect 27810 2216 28770 2254
rect 28828 2254 29030 2271
rect 29586 2271 29602 2288
rect 30032 2288 30620 2304
rect 30032 2271 30048 2288
rect 29586 2254 29788 2271
rect 28828 2216 29788 2254
rect 29846 2254 30048 2271
rect 30604 2271 30620 2288
rect 31050 2288 31638 2304
rect 31050 2271 31066 2288
rect 30604 2254 30806 2271
rect 29846 2216 30806 2254
rect 30864 2254 31066 2271
rect 31622 2271 31638 2288
rect 32068 2288 32656 2304
rect 32068 2271 32084 2288
rect 31622 2254 31824 2271
rect 30864 2216 31824 2254
rect 31882 2254 32084 2271
rect 32640 2271 32656 2288
rect 33086 2288 33674 2304
rect 33086 2271 33102 2288
rect 32640 2254 32842 2271
rect 31882 2216 32842 2254
rect 32900 2254 33102 2271
rect 33658 2271 33674 2288
rect 34104 2288 34692 2304
rect 34104 2271 34120 2288
rect 33658 2254 33860 2271
rect 32900 2216 33860 2254
rect 33918 2254 34120 2271
rect 34676 2271 34692 2288
rect 35122 2288 35710 2304
rect 35122 2271 35138 2288
rect 34676 2254 34878 2271
rect 33918 2216 34878 2254
rect 34936 2254 35138 2271
rect 35694 2271 35710 2288
rect 36140 2288 36728 2304
rect 36140 2271 36156 2288
rect 35694 2254 35896 2271
rect 34936 2216 35896 2254
rect 35954 2254 36156 2271
rect 36712 2271 36728 2288
rect 37158 2288 37746 2304
rect 37158 2271 37174 2288
rect 36712 2254 36914 2271
rect 35954 2216 36914 2254
rect 36972 2254 37174 2271
rect 37730 2271 37746 2288
rect 38176 2288 38764 2304
rect 38176 2271 38192 2288
rect 37730 2254 37932 2271
rect 36972 2216 37932 2254
rect 37990 2254 38192 2271
rect 38748 2271 38764 2288
rect 39194 2288 39782 2304
rect 39194 2271 39210 2288
rect 38748 2254 38950 2271
rect 37990 2216 38950 2254
rect 39008 2254 39210 2271
rect 39766 2271 39782 2288
rect 39766 2254 39968 2271
rect 39008 2216 39968 2254
rect 6578 1956 7538 1994
rect 6578 1939 6780 1956
rect 6764 1922 6780 1939
rect 7336 1939 7538 1956
rect 7596 1956 8556 1994
rect 7596 1939 7798 1956
rect 7336 1922 7352 1939
rect 6764 1906 7352 1922
rect 7782 1922 7798 1939
rect 8354 1939 8556 1956
rect 8614 1956 9574 1994
rect 8614 1939 8816 1956
rect 8354 1922 8370 1939
rect 7782 1906 8370 1922
rect 8800 1922 8816 1939
rect 9372 1939 9574 1956
rect 9632 1956 10592 1994
rect 9632 1939 9834 1956
rect 9372 1922 9388 1939
rect 8800 1906 9388 1922
rect 9818 1922 9834 1939
rect 10390 1939 10592 1956
rect 10650 1956 11610 1994
rect 10650 1939 10852 1956
rect 10390 1922 10406 1939
rect 9818 1906 10406 1922
rect 10836 1922 10852 1939
rect 11408 1939 11610 1956
rect 11668 1956 12628 1994
rect 11668 1939 11870 1956
rect 11408 1922 11424 1939
rect 10836 1906 11424 1922
rect 11854 1922 11870 1939
rect 12426 1939 12628 1956
rect 12686 1956 13646 1994
rect 12686 1939 12888 1956
rect 12426 1922 12442 1939
rect 11854 1906 12442 1922
rect 12872 1922 12888 1939
rect 13444 1939 13646 1956
rect 13704 1956 14664 1994
rect 13704 1939 13906 1956
rect 13444 1922 13460 1939
rect 12872 1906 13460 1922
rect 13890 1922 13906 1939
rect 14462 1939 14664 1956
rect 14722 1956 15682 1994
rect 14722 1939 14924 1956
rect 14462 1922 14478 1939
rect 13890 1906 14478 1922
rect 14908 1922 14924 1939
rect 15480 1939 15682 1956
rect 15740 1956 16700 1994
rect 15740 1939 15942 1956
rect 15480 1922 15496 1939
rect 14908 1906 15496 1922
rect 15926 1922 15942 1939
rect 16498 1939 16700 1956
rect 16758 1956 17718 1994
rect 16758 1939 16960 1956
rect 16498 1922 16514 1939
rect 15926 1906 16514 1922
rect 16944 1922 16960 1939
rect 17516 1939 17718 1956
rect 17516 1922 17532 1939
rect 16944 1906 17532 1922
rect 19666 1578 20626 1616
rect 6764 1554 7352 1570
rect 6764 1537 6780 1554
rect 6578 1520 6780 1537
rect 7336 1537 7352 1554
rect 7782 1554 8370 1570
rect 7782 1537 7798 1554
rect 7336 1520 7538 1537
rect 6578 1482 7538 1520
rect 7596 1520 7798 1537
rect 8354 1537 8370 1554
rect 8800 1554 9388 1570
rect 8800 1537 8816 1554
rect 8354 1520 8556 1537
rect 7596 1482 8556 1520
rect 8614 1520 8816 1537
rect 9372 1537 9388 1554
rect 9818 1554 10406 1570
rect 9818 1537 9834 1554
rect 9372 1520 9574 1537
rect 8614 1482 9574 1520
rect 9632 1520 9834 1537
rect 10390 1537 10406 1554
rect 10836 1554 11424 1570
rect 10836 1537 10852 1554
rect 10390 1520 10592 1537
rect 9632 1482 10592 1520
rect 10650 1520 10852 1537
rect 11408 1537 11424 1554
rect 11854 1554 12442 1570
rect 11854 1537 11870 1554
rect 11408 1520 11610 1537
rect 10650 1482 11610 1520
rect 11668 1520 11870 1537
rect 12426 1537 12442 1554
rect 12872 1554 13460 1570
rect 12872 1537 12888 1554
rect 12426 1520 12628 1537
rect 11668 1482 12628 1520
rect 12686 1520 12888 1537
rect 13444 1537 13460 1554
rect 13890 1554 14478 1570
rect 13890 1537 13906 1554
rect 13444 1520 13646 1537
rect 12686 1482 13646 1520
rect 13704 1520 13906 1537
rect 14462 1537 14478 1554
rect 14908 1554 15496 1570
rect 14908 1537 14924 1554
rect 14462 1520 14664 1537
rect 13704 1482 14664 1520
rect 14722 1520 14924 1537
rect 15480 1537 15496 1554
rect 15926 1554 16514 1570
rect 15926 1537 15942 1554
rect 15480 1520 15682 1537
rect 14722 1482 15682 1520
rect 15740 1520 15942 1537
rect 16498 1537 16514 1554
rect 16944 1554 17532 1570
rect 19666 1561 19868 1578
rect 16944 1537 16960 1554
rect 16498 1520 16700 1537
rect 15740 1482 16700 1520
rect 16758 1520 16960 1537
rect 17516 1537 17532 1554
rect 19852 1544 19868 1561
rect 20424 1561 20626 1578
rect 20684 1578 21644 1616
rect 20684 1561 20886 1578
rect 20424 1544 20440 1561
rect 17516 1520 17718 1537
rect 19852 1528 20440 1544
rect 20870 1544 20886 1561
rect 21442 1561 21644 1578
rect 21702 1578 22662 1616
rect 21702 1561 21904 1578
rect 21442 1544 21458 1561
rect 20870 1528 21458 1544
rect 21888 1544 21904 1561
rect 22460 1561 22662 1578
rect 22720 1578 23680 1616
rect 22720 1561 22922 1578
rect 22460 1544 22476 1561
rect 21888 1528 22476 1544
rect 22906 1544 22922 1561
rect 23478 1561 23680 1578
rect 23738 1578 24698 1616
rect 23738 1561 23940 1578
rect 23478 1544 23494 1561
rect 22906 1528 23494 1544
rect 23924 1544 23940 1561
rect 24496 1561 24698 1578
rect 24756 1578 25716 1616
rect 24756 1561 24958 1578
rect 24496 1544 24512 1561
rect 23924 1528 24512 1544
rect 24942 1544 24958 1561
rect 25514 1561 25716 1578
rect 25774 1578 26734 1616
rect 25774 1561 25976 1578
rect 25514 1544 25530 1561
rect 24942 1528 25530 1544
rect 25960 1544 25976 1561
rect 26532 1561 26734 1578
rect 26792 1578 27752 1616
rect 26792 1561 26994 1578
rect 26532 1544 26548 1561
rect 25960 1528 26548 1544
rect 26978 1544 26994 1561
rect 27550 1561 27752 1578
rect 27810 1578 28770 1616
rect 27810 1561 28012 1578
rect 27550 1544 27566 1561
rect 26978 1528 27566 1544
rect 27996 1544 28012 1561
rect 28568 1561 28770 1578
rect 28828 1578 29788 1616
rect 28828 1561 29030 1578
rect 28568 1544 28584 1561
rect 27996 1528 28584 1544
rect 29014 1544 29030 1561
rect 29586 1561 29788 1578
rect 29846 1578 30806 1616
rect 29846 1561 30048 1578
rect 29586 1544 29602 1561
rect 29014 1528 29602 1544
rect 30032 1544 30048 1561
rect 30604 1561 30806 1578
rect 30864 1578 31824 1616
rect 30864 1561 31066 1578
rect 30604 1544 30620 1561
rect 30032 1528 30620 1544
rect 31050 1544 31066 1561
rect 31622 1561 31824 1578
rect 31882 1578 32842 1616
rect 31882 1561 32084 1578
rect 31622 1544 31638 1561
rect 31050 1528 31638 1544
rect 32068 1544 32084 1561
rect 32640 1561 32842 1578
rect 32900 1578 33860 1616
rect 32900 1561 33102 1578
rect 32640 1544 32656 1561
rect 32068 1528 32656 1544
rect 33086 1544 33102 1561
rect 33658 1561 33860 1578
rect 33918 1578 34878 1616
rect 33918 1561 34120 1578
rect 33658 1544 33674 1561
rect 33086 1528 33674 1544
rect 34104 1544 34120 1561
rect 34676 1561 34878 1578
rect 34936 1578 35896 1616
rect 34936 1561 35138 1578
rect 34676 1544 34692 1561
rect 34104 1528 34692 1544
rect 35122 1544 35138 1561
rect 35694 1561 35896 1578
rect 35954 1578 36914 1616
rect 35954 1561 36156 1578
rect 35694 1544 35710 1561
rect 35122 1528 35710 1544
rect 36140 1544 36156 1561
rect 36712 1561 36914 1578
rect 36972 1578 37932 1616
rect 36972 1561 37174 1578
rect 36712 1544 36728 1561
rect 36140 1528 36728 1544
rect 37158 1544 37174 1561
rect 37730 1561 37932 1578
rect 37990 1578 38950 1616
rect 37990 1561 38192 1578
rect 37730 1544 37746 1561
rect 37158 1528 37746 1544
rect 38176 1544 38192 1561
rect 38748 1561 38950 1578
rect 39008 1578 39968 1616
rect 39008 1561 39210 1578
rect 38748 1544 38764 1561
rect 38176 1528 38764 1544
rect 39194 1544 39210 1561
rect 39766 1561 39968 1578
rect 39766 1544 39782 1561
rect 39194 1528 39782 1544
rect 16758 1482 17718 1520
rect 19852 1054 20440 1070
rect 19852 1037 19868 1054
rect 19666 1020 19868 1037
rect 20424 1037 20440 1054
rect 20870 1054 21458 1070
rect 20870 1037 20886 1054
rect 20424 1020 20626 1037
rect 19666 982 20626 1020
rect 20684 1020 20886 1037
rect 21442 1037 21458 1054
rect 21888 1054 22476 1070
rect 21888 1037 21904 1054
rect 21442 1020 21644 1037
rect 20684 982 21644 1020
rect 21702 1020 21904 1037
rect 22460 1037 22476 1054
rect 22906 1054 23494 1070
rect 22906 1037 22922 1054
rect 22460 1020 22662 1037
rect 21702 982 22662 1020
rect 22720 1020 22922 1037
rect 23478 1037 23494 1054
rect 23924 1054 24512 1070
rect 23924 1037 23940 1054
rect 23478 1020 23680 1037
rect 22720 982 23680 1020
rect 23738 1020 23940 1037
rect 24496 1037 24512 1054
rect 24942 1054 25530 1070
rect 24942 1037 24958 1054
rect 24496 1020 24698 1037
rect 23738 982 24698 1020
rect 24756 1020 24958 1037
rect 25514 1037 25530 1054
rect 25960 1054 26548 1070
rect 25960 1037 25976 1054
rect 25514 1020 25716 1037
rect 24756 982 25716 1020
rect 25774 1020 25976 1037
rect 26532 1037 26548 1054
rect 26978 1054 27566 1070
rect 26978 1037 26994 1054
rect 26532 1020 26734 1037
rect 25774 982 26734 1020
rect 26792 1020 26994 1037
rect 27550 1037 27566 1054
rect 27996 1054 28584 1070
rect 27996 1037 28012 1054
rect 27550 1020 27752 1037
rect 26792 982 27752 1020
rect 27810 1020 28012 1037
rect 28568 1037 28584 1054
rect 29014 1054 29602 1070
rect 29014 1037 29030 1054
rect 28568 1020 28770 1037
rect 27810 982 28770 1020
rect 28828 1020 29030 1037
rect 29586 1037 29602 1054
rect 30032 1054 30620 1070
rect 30032 1037 30048 1054
rect 29586 1020 29788 1037
rect 28828 982 29788 1020
rect 29846 1020 30048 1037
rect 30604 1037 30620 1054
rect 31050 1054 31638 1070
rect 31050 1037 31066 1054
rect 30604 1020 30806 1037
rect 29846 982 30806 1020
rect 30864 1020 31066 1037
rect 31622 1037 31638 1054
rect 32068 1054 32656 1070
rect 32068 1037 32084 1054
rect 31622 1020 31824 1037
rect 30864 982 31824 1020
rect 31882 1020 32084 1037
rect 32640 1037 32656 1054
rect 33086 1054 33674 1070
rect 33086 1037 33102 1054
rect 32640 1020 32842 1037
rect 31882 982 32842 1020
rect 32900 1020 33102 1037
rect 33658 1037 33674 1054
rect 34104 1054 34692 1070
rect 34104 1037 34120 1054
rect 33658 1020 33860 1037
rect 32900 982 33860 1020
rect 33918 1020 34120 1037
rect 34676 1037 34692 1054
rect 35122 1054 35710 1070
rect 35122 1037 35138 1054
rect 34676 1020 34878 1037
rect 33918 982 34878 1020
rect 34936 1020 35138 1037
rect 35694 1037 35710 1054
rect 36140 1054 36728 1070
rect 36140 1037 36156 1054
rect 35694 1020 35896 1037
rect 34936 982 35896 1020
rect 35954 1020 36156 1037
rect 36712 1037 36728 1054
rect 37158 1054 37746 1070
rect 37158 1037 37174 1054
rect 36712 1020 36914 1037
rect 35954 982 36914 1020
rect 36972 1020 37174 1037
rect 37730 1037 37746 1054
rect 38176 1054 38764 1070
rect 38176 1037 38192 1054
rect 37730 1020 37932 1037
rect 36972 982 37932 1020
rect 37990 1020 38192 1037
rect 38748 1037 38764 1054
rect 39194 1054 39782 1070
rect 39194 1037 39210 1054
rect 38748 1020 38950 1037
rect 37990 982 38950 1020
rect 39008 1020 39210 1037
rect 39766 1037 39782 1054
rect 39766 1020 39968 1037
rect 39008 982 39968 1020
rect 6578 844 7538 882
rect 6578 827 6780 844
rect 6764 810 6780 827
rect 7336 827 7538 844
rect 7596 844 8556 882
rect 7596 827 7798 844
rect 7336 810 7352 827
rect 6764 794 7352 810
rect 7782 810 7798 827
rect 8354 827 8556 844
rect 8614 844 9574 882
rect 8614 827 8816 844
rect 8354 810 8370 827
rect 7782 794 8370 810
rect 8800 810 8816 827
rect 9372 827 9574 844
rect 9632 844 10592 882
rect 9632 827 9834 844
rect 9372 810 9388 827
rect 8800 794 9388 810
rect 9818 810 9834 827
rect 10390 827 10592 844
rect 10650 844 11610 882
rect 10650 827 10852 844
rect 10390 810 10406 827
rect 9818 794 10406 810
rect 10836 810 10852 827
rect 11408 827 11610 844
rect 11668 844 12628 882
rect 11668 827 11870 844
rect 11408 810 11424 827
rect 10836 794 11424 810
rect 11854 810 11870 827
rect 12426 827 12628 844
rect 12686 844 13646 882
rect 12686 827 12888 844
rect 12426 810 12442 827
rect 11854 794 12442 810
rect 12872 810 12888 827
rect 13444 827 13646 844
rect 13704 844 14664 882
rect 13704 827 13906 844
rect 13444 810 13460 827
rect 12872 794 13460 810
rect 13890 810 13906 827
rect 14462 827 14664 844
rect 14722 844 15682 882
rect 14722 827 14924 844
rect 14462 810 14478 827
rect 13890 794 14478 810
rect 14908 810 14924 827
rect 15480 827 15682 844
rect 15740 844 16700 882
rect 15740 827 15942 844
rect 15480 810 15496 827
rect 14908 794 15496 810
rect 15926 810 15942 827
rect 16498 827 16700 844
rect 16758 844 17718 882
rect 16758 827 16960 844
rect 16498 810 16514 827
rect 15926 794 16514 810
rect 16944 810 16960 827
rect 17516 827 17718 844
rect 17516 810 17532 827
rect 16944 794 17532 810
rect 19666 344 20626 382
rect 19666 327 19868 344
rect 19852 310 19868 327
rect 20424 327 20626 344
rect 20684 344 21644 382
rect 20684 327 20886 344
rect 20424 310 20440 327
rect 19852 294 20440 310
rect 20870 310 20886 327
rect 21442 327 21644 344
rect 21702 344 22662 382
rect 21702 327 21904 344
rect 21442 310 21458 327
rect 20870 294 21458 310
rect 21888 310 21904 327
rect 22460 327 22662 344
rect 22720 344 23680 382
rect 22720 327 22922 344
rect 22460 310 22476 327
rect 21888 294 22476 310
rect 22906 310 22922 327
rect 23478 327 23680 344
rect 23738 344 24698 382
rect 23738 327 23940 344
rect 23478 310 23494 327
rect 22906 294 23494 310
rect 23924 310 23940 327
rect 24496 327 24698 344
rect 24756 344 25716 382
rect 24756 327 24958 344
rect 24496 310 24512 327
rect 23924 294 24512 310
rect 24942 310 24958 327
rect 25514 327 25716 344
rect 25774 344 26734 382
rect 25774 327 25976 344
rect 25514 310 25530 327
rect 24942 294 25530 310
rect 25960 310 25976 327
rect 26532 327 26734 344
rect 26792 344 27752 382
rect 26792 327 26994 344
rect 26532 310 26548 327
rect 25960 294 26548 310
rect 26978 310 26994 327
rect 27550 327 27752 344
rect 27810 344 28770 382
rect 27810 327 28012 344
rect 27550 310 27566 327
rect 26978 294 27566 310
rect 27996 310 28012 327
rect 28568 327 28770 344
rect 28828 344 29788 382
rect 28828 327 29030 344
rect 28568 310 28584 327
rect 27996 294 28584 310
rect 29014 310 29030 327
rect 29586 327 29788 344
rect 29846 344 30806 382
rect 29846 327 30048 344
rect 29586 310 29602 327
rect 29014 294 29602 310
rect 30032 310 30048 327
rect 30604 327 30806 344
rect 30864 344 31824 382
rect 30864 327 31066 344
rect 30604 310 30620 327
rect 30032 294 30620 310
rect 31050 310 31066 327
rect 31622 327 31824 344
rect 31882 344 32842 382
rect 31882 327 32084 344
rect 31622 310 31638 327
rect 31050 294 31638 310
rect 32068 310 32084 327
rect 32640 327 32842 344
rect 32900 344 33860 382
rect 32900 327 33102 344
rect 32640 310 32656 327
rect 32068 294 32656 310
rect 33086 310 33102 327
rect 33658 327 33860 344
rect 33918 344 34878 382
rect 33918 327 34120 344
rect 33658 310 33674 327
rect 33086 294 33674 310
rect 34104 310 34120 327
rect 34676 327 34878 344
rect 34936 344 35896 382
rect 34936 327 35138 344
rect 34676 310 34692 327
rect 34104 294 34692 310
rect 35122 310 35138 327
rect 35694 327 35896 344
rect 35954 344 36914 382
rect 35954 327 36156 344
rect 35694 310 35710 327
rect 35122 294 35710 310
rect 36140 310 36156 327
rect 36712 327 36914 344
rect 36972 344 37932 382
rect 36972 327 37174 344
rect 36712 310 36728 327
rect 36140 294 36728 310
rect 37158 310 37174 327
rect 37730 327 37932 344
rect 37990 344 38950 382
rect 37990 327 38192 344
rect 37730 310 37746 327
rect 37158 294 37746 310
rect 38176 310 38192 327
rect 38748 327 38950 344
rect 39008 344 39968 382
rect 39008 327 39210 344
rect 38748 310 38764 327
rect 38176 294 38764 310
rect 39194 310 39210 327
rect 39766 327 39968 344
rect 39766 310 39782 327
rect 39194 294 39782 310
rect 7222 12 7810 28
rect 7222 -5 7238 12
rect 7036 -22 7238 -5
rect 7794 -5 7810 12
rect 8240 12 8828 28
rect 8240 -5 8256 12
rect 7794 -22 7996 -5
rect 7036 -60 7996 -22
rect 8054 -22 8256 -5
rect 8812 -5 8828 12
rect 9258 12 9846 28
rect 9258 -5 9274 12
rect 8812 -22 9014 -5
rect 8054 -60 9014 -22
rect 9072 -22 9274 -5
rect 9830 -5 9846 12
rect 10276 12 10864 28
rect 10276 -5 10292 12
rect 9830 -22 10032 -5
rect 9072 -60 10032 -22
rect 10090 -22 10292 -5
rect 10848 -5 10864 12
rect 11294 12 11882 28
rect 11294 -5 11310 12
rect 10848 -22 11050 -5
rect 10090 -60 11050 -22
rect 11108 -22 11310 -5
rect 11866 -5 11882 12
rect 12312 12 12900 28
rect 12312 -5 12328 12
rect 11866 -22 12068 -5
rect 11108 -60 12068 -22
rect 12126 -22 12328 -5
rect 12884 -5 12900 12
rect 13330 12 13918 28
rect 13330 -5 13346 12
rect 12884 -22 13086 -5
rect 12126 -60 13086 -22
rect 13144 -22 13346 -5
rect 13902 -5 13918 12
rect 14348 12 14936 28
rect 14348 -5 14364 12
rect 13902 -22 14104 -5
rect 13144 -60 14104 -22
rect 14162 -22 14364 -5
rect 14920 -5 14936 12
rect 15366 12 15954 28
rect 15366 -5 15382 12
rect 14920 -22 15122 -5
rect 14162 -60 15122 -22
rect 15180 -22 15382 -5
rect 15938 -5 15954 12
rect 16384 12 16972 28
rect 16384 -5 16400 12
rect 15938 -22 16140 -5
rect 15180 -60 16140 -22
rect 16198 -22 16400 -5
rect 16956 -5 16972 12
rect 16956 -22 17158 -5
rect 16198 -60 17158 -22
rect 19852 -178 20440 -162
rect 19852 -195 19868 -178
rect 19666 -212 19868 -195
rect 20424 -195 20440 -178
rect 20870 -178 21458 -162
rect 20870 -195 20886 -178
rect 20424 -212 20626 -195
rect 19666 -250 20626 -212
rect 20684 -212 20886 -195
rect 21442 -195 21458 -178
rect 21888 -178 22476 -162
rect 21888 -195 21904 -178
rect 21442 -212 21644 -195
rect 20684 -250 21644 -212
rect 21702 -212 21904 -195
rect 22460 -195 22476 -178
rect 22906 -178 23494 -162
rect 22906 -195 22922 -178
rect 22460 -212 22662 -195
rect 21702 -250 22662 -212
rect 22720 -212 22922 -195
rect 23478 -195 23494 -178
rect 23924 -178 24512 -162
rect 23924 -195 23940 -178
rect 23478 -212 23680 -195
rect 22720 -250 23680 -212
rect 23738 -212 23940 -195
rect 24496 -195 24512 -178
rect 24942 -178 25530 -162
rect 24942 -195 24958 -178
rect 24496 -212 24698 -195
rect 23738 -250 24698 -212
rect 24756 -212 24958 -195
rect 25514 -195 25530 -178
rect 25960 -178 26548 -162
rect 25960 -195 25976 -178
rect 25514 -212 25716 -195
rect 24756 -250 25716 -212
rect 25774 -212 25976 -195
rect 26532 -195 26548 -178
rect 26978 -178 27566 -162
rect 26978 -195 26994 -178
rect 26532 -212 26734 -195
rect 25774 -250 26734 -212
rect 26792 -212 26994 -195
rect 27550 -195 27566 -178
rect 27996 -178 28584 -162
rect 27996 -195 28012 -178
rect 27550 -212 27752 -195
rect 26792 -250 27752 -212
rect 27810 -212 28012 -195
rect 28568 -195 28584 -178
rect 29014 -178 29602 -162
rect 29014 -195 29030 -178
rect 28568 -212 28770 -195
rect 27810 -250 28770 -212
rect 28828 -212 29030 -195
rect 29586 -195 29602 -178
rect 30032 -178 30620 -162
rect 30032 -195 30048 -178
rect 29586 -212 29788 -195
rect 28828 -250 29788 -212
rect 29846 -212 30048 -195
rect 30604 -195 30620 -178
rect 31050 -178 31638 -162
rect 31050 -195 31066 -178
rect 30604 -212 30806 -195
rect 29846 -250 30806 -212
rect 30864 -212 31066 -195
rect 31622 -195 31638 -178
rect 32068 -178 32656 -162
rect 32068 -195 32084 -178
rect 31622 -212 31824 -195
rect 30864 -250 31824 -212
rect 31882 -212 32084 -195
rect 32640 -195 32656 -178
rect 33086 -178 33674 -162
rect 33086 -195 33102 -178
rect 32640 -212 32842 -195
rect 31882 -250 32842 -212
rect 32900 -212 33102 -195
rect 33658 -195 33674 -178
rect 34104 -178 34692 -162
rect 34104 -195 34120 -178
rect 33658 -212 33860 -195
rect 32900 -250 33860 -212
rect 33918 -212 34120 -195
rect 34676 -195 34692 -178
rect 35122 -178 35710 -162
rect 35122 -195 35138 -178
rect 34676 -212 34878 -195
rect 33918 -250 34878 -212
rect 34936 -212 35138 -195
rect 35694 -195 35710 -178
rect 36140 -178 36728 -162
rect 36140 -195 36156 -178
rect 35694 -212 35896 -195
rect 34936 -250 35896 -212
rect 35954 -212 36156 -195
rect 36712 -195 36728 -178
rect 37158 -178 37746 -162
rect 37158 -195 37174 -178
rect 36712 -212 36914 -195
rect 35954 -250 36914 -212
rect 36972 -212 37174 -195
rect 37730 -195 37746 -178
rect 38176 -178 38764 -162
rect 38176 -195 38192 -178
rect 37730 -212 37932 -195
rect 36972 -250 37932 -212
rect 37990 -212 38192 -195
rect 38748 -195 38764 -178
rect 39194 -178 39782 -162
rect 39194 -195 39210 -178
rect 38748 -212 38950 -195
rect 37990 -250 38950 -212
rect 39008 -212 39210 -195
rect 39766 -195 39782 -178
rect 39766 -212 39968 -195
rect 39008 -250 39968 -212
rect 7036 -698 7996 -660
rect 7036 -715 7238 -698
rect 7222 -732 7238 -715
rect 7794 -715 7996 -698
rect 8054 -698 9014 -660
rect 8054 -715 8256 -698
rect 7794 -732 7810 -715
rect 7222 -748 7810 -732
rect 8240 -732 8256 -715
rect 8812 -715 9014 -698
rect 9072 -698 10032 -660
rect 9072 -715 9274 -698
rect 8812 -732 8828 -715
rect 8240 -748 8828 -732
rect 9258 -732 9274 -715
rect 9830 -715 10032 -698
rect 10090 -698 11050 -660
rect 10090 -715 10292 -698
rect 9830 -732 9846 -715
rect 9258 -748 9846 -732
rect 10276 -732 10292 -715
rect 10848 -715 11050 -698
rect 11108 -698 12068 -660
rect 11108 -715 11310 -698
rect 10848 -732 10864 -715
rect 10276 -748 10864 -732
rect 11294 -732 11310 -715
rect 11866 -715 12068 -698
rect 12126 -698 13086 -660
rect 12126 -715 12328 -698
rect 11866 -732 11882 -715
rect 11294 -748 11882 -732
rect 12312 -732 12328 -715
rect 12884 -715 13086 -698
rect 13144 -698 14104 -660
rect 13144 -715 13346 -698
rect 12884 -732 12900 -715
rect 12312 -748 12900 -732
rect 13330 -732 13346 -715
rect 13902 -715 14104 -698
rect 14162 -698 15122 -660
rect 14162 -715 14364 -698
rect 13902 -732 13918 -715
rect 13330 -748 13918 -732
rect 14348 -732 14364 -715
rect 14920 -715 15122 -698
rect 15180 -698 16140 -660
rect 15180 -715 15382 -698
rect 14920 -732 14936 -715
rect 14348 -748 14936 -732
rect 15366 -732 15382 -715
rect 15938 -715 16140 -698
rect 16198 -698 17158 -660
rect 16198 -715 16400 -698
rect 15938 -732 15954 -715
rect 15366 -748 15954 -732
rect 16384 -732 16400 -715
rect 16956 -715 17158 -698
rect 16956 -732 16972 -715
rect 16384 -748 16972 -732
rect 19666 -888 20626 -850
rect 19666 -905 19868 -888
rect 19852 -922 19868 -905
rect 20424 -905 20626 -888
rect 20684 -888 21644 -850
rect 20684 -905 20886 -888
rect 20424 -922 20440 -905
rect 19852 -938 20440 -922
rect 20870 -922 20886 -905
rect 21442 -905 21644 -888
rect 21702 -888 22662 -850
rect 21702 -905 21904 -888
rect 21442 -922 21458 -905
rect 20870 -938 21458 -922
rect 21888 -922 21904 -905
rect 22460 -905 22662 -888
rect 22720 -888 23680 -850
rect 22720 -905 22922 -888
rect 22460 -922 22476 -905
rect 21888 -938 22476 -922
rect 22906 -922 22922 -905
rect 23478 -905 23680 -888
rect 23738 -888 24698 -850
rect 23738 -905 23940 -888
rect 23478 -922 23494 -905
rect 22906 -938 23494 -922
rect 23924 -922 23940 -905
rect 24496 -905 24698 -888
rect 24756 -888 25716 -850
rect 24756 -905 24958 -888
rect 24496 -922 24512 -905
rect 23924 -938 24512 -922
rect 24942 -922 24958 -905
rect 25514 -905 25716 -888
rect 25774 -888 26734 -850
rect 25774 -905 25976 -888
rect 25514 -922 25530 -905
rect 24942 -938 25530 -922
rect 25960 -922 25976 -905
rect 26532 -905 26734 -888
rect 26792 -888 27752 -850
rect 26792 -905 26994 -888
rect 26532 -922 26548 -905
rect 25960 -938 26548 -922
rect 26978 -922 26994 -905
rect 27550 -905 27752 -888
rect 27810 -888 28770 -850
rect 27810 -905 28012 -888
rect 27550 -922 27566 -905
rect 26978 -938 27566 -922
rect 27996 -922 28012 -905
rect 28568 -905 28770 -888
rect 28828 -888 29788 -850
rect 28828 -905 29030 -888
rect 28568 -922 28584 -905
rect 27996 -938 28584 -922
rect 29014 -922 29030 -905
rect 29586 -905 29788 -888
rect 29846 -888 30806 -850
rect 29846 -905 30048 -888
rect 29586 -922 29602 -905
rect 29014 -938 29602 -922
rect 30032 -922 30048 -905
rect 30604 -905 30806 -888
rect 30864 -888 31824 -850
rect 30864 -905 31066 -888
rect 30604 -922 30620 -905
rect 30032 -938 30620 -922
rect 31050 -922 31066 -905
rect 31622 -905 31824 -888
rect 31882 -888 32842 -850
rect 31882 -905 32084 -888
rect 31622 -922 31638 -905
rect 31050 -938 31638 -922
rect 32068 -922 32084 -905
rect 32640 -905 32842 -888
rect 32900 -888 33860 -850
rect 32900 -905 33102 -888
rect 32640 -922 32656 -905
rect 32068 -938 32656 -922
rect 33086 -922 33102 -905
rect 33658 -905 33860 -888
rect 33918 -888 34878 -850
rect 33918 -905 34120 -888
rect 33658 -922 33674 -905
rect 33086 -938 33674 -922
rect 34104 -922 34120 -905
rect 34676 -905 34878 -888
rect 34936 -888 35896 -850
rect 34936 -905 35138 -888
rect 34676 -922 34692 -905
rect 34104 -938 34692 -922
rect 35122 -922 35138 -905
rect 35694 -905 35896 -888
rect 35954 -888 36914 -850
rect 35954 -905 36156 -888
rect 35694 -922 35710 -905
rect 35122 -938 35710 -922
rect 36140 -922 36156 -905
rect 36712 -905 36914 -888
rect 36972 -888 37932 -850
rect 36972 -905 37174 -888
rect 36712 -922 36728 -905
rect 36140 -938 36728 -922
rect 37158 -922 37174 -905
rect 37730 -905 37932 -888
rect 37990 -888 38950 -850
rect 37990 -905 38192 -888
rect 37730 -922 37746 -905
rect 37158 -938 37746 -922
rect 38176 -922 38192 -905
rect 38748 -905 38950 -888
rect 39008 -888 39968 -850
rect 39008 -905 39210 -888
rect 38748 -922 38764 -905
rect 38176 -938 38764 -922
rect 39194 -922 39210 -905
rect 39766 -905 39968 -888
rect 39766 -922 39782 -905
rect 39194 -938 39782 -922
<< polycont >>
rect 23776 26601 24332 26635
rect 24794 26601 25350 26635
rect 25812 26601 26368 26635
rect 26830 26601 27386 26635
rect 27848 26601 28404 26635
rect 28866 26601 29422 26635
rect 29884 26601 30440 26635
rect 30902 26601 31458 26635
rect 31920 26601 32476 26635
rect 32938 26601 33494 26635
rect 33956 26601 34512 26635
rect 34974 26601 35530 26635
rect 35992 26601 36548 26635
rect 37010 26601 37566 26635
rect 38028 26601 38584 26635
rect 39046 26601 39602 26635
rect 23776 25873 24332 25907
rect 24794 25873 25350 25907
rect 25812 25873 26368 25907
rect 26830 25873 27386 25907
rect 27848 25873 28404 25907
rect 28866 25873 29422 25907
rect 29884 25873 30440 25907
rect 30902 25873 31458 25907
rect 31920 25873 32476 25907
rect 32938 25873 33494 25907
rect 33956 25873 34512 25907
rect 34974 25873 35530 25907
rect 35992 25873 36548 25907
rect 37010 25873 37566 25907
rect 38028 25873 38584 25907
rect 39046 25873 39602 25907
rect 23776 25465 24332 25499
rect 24794 25465 25350 25499
rect 25812 25465 26368 25499
rect 26830 25465 27386 25499
rect 27848 25465 28404 25499
rect 28866 25465 29422 25499
rect 29884 25465 30440 25499
rect 30902 25465 31458 25499
rect 31920 25465 32476 25499
rect 32938 25465 33494 25499
rect 33956 25465 34512 25499
rect 34974 25465 35530 25499
rect 35992 25465 36548 25499
rect 37010 25465 37566 25499
rect 38028 25465 38584 25499
rect 39046 25465 39602 25499
rect 23776 24737 24332 24771
rect 24794 24737 25350 24771
rect 25812 24737 26368 24771
rect 26830 24737 27386 24771
rect 27848 24737 28404 24771
rect 28866 24737 29422 24771
rect 29884 24737 30440 24771
rect 30902 24737 31458 24771
rect 31920 24737 32476 24771
rect 32938 24737 33494 24771
rect 33956 24737 34512 24771
rect 34974 24737 35530 24771
rect 35992 24737 36548 24771
rect 37010 24737 37566 24771
rect 38028 24737 38584 24771
rect 39046 24737 39602 24771
rect 23776 24329 24332 24363
rect 24794 24329 25350 24363
rect 25812 24329 26368 24363
rect 26830 24329 27386 24363
rect 27848 24329 28404 24363
rect 28866 24329 29422 24363
rect 29884 24329 30440 24363
rect 30902 24329 31458 24363
rect 31920 24329 32476 24363
rect 32938 24329 33494 24363
rect 33956 24329 34512 24363
rect 34974 24329 35530 24363
rect 35992 24329 36548 24363
rect 37010 24329 37566 24363
rect 38028 24329 38584 24363
rect 39046 24329 39602 24363
rect 23776 23601 24332 23635
rect 24794 23601 25350 23635
rect 25812 23601 26368 23635
rect 26830 23601 27386 23635
rect 27848 23601 28404 23635
rect 28866 23601 29422 23635
rect 29884 23601 30440 23635
rect 30902 23601 31458 23635
rect 31920 23601 32476 23635
rect 32938 23601 33494 23635
rect 33956 23601 34512 23635
rect 34974 23601 35530 23635
rect 35992 23601 36548 23635
rect 37010 23601 37566 23635
rect 38028 23601 38584 23635
rect 39046 23601 39602 23635
rect 24970 22691 25526 22725
rect 25988 22691 26544 22725
rect 27006 22691 27562 22725
rect 28024 22691 28580 22725
rect 29042 22691 29598 22725
rect 30060 22691 30616 22725
rect 31078 22691 31634 22725
rect 32096 22691 32652 22725
rect 33114 22691 33670 22725
rect 34132 22691 34688 22725
rect 35150 22691 35706 22725
rect 36168 22691 36724 22725
rect 37186 22691 37742 22725
rect 38204 22691 38760 22725
rect 24970 21963 25526 21997
rect 25988 21963 26544 21997
rect 27006 21963 27562 21997
rect 28024 21963 28580 21997
rect 29042 21963 29598 21997
rect 30060 21963 30616 21997
rect 31078 21963 31634 21997
rect 32096 21963 32652 21997
rect 33114 21963 33670 21997
rect 34132 21963 34688 21997
rect 35150 21963 35706 21997
rect 36168 21963 36724 21997
rect 37186 21963 37742 21997
rect 38204 21963 38760 21997
rect 24970 21659 25526 21693
rect 25988 21659 26544 21693
rect 27006 21659 27562 21693
rect 28024 21659 28580 21693
rect 29042 21659 29598 21693
rect 30060 21659 30616 21693
rect 31078 21659 31634 21693
rect 32096 21659 32652 21693
rect 33114 21659 33670 21693
rect 34132 21659 34688 21693
rect 35150 21659 35706 21693
rect 36168 21659 36724 21693
rect 37186 21659 37742 21693
rect 38204 21659 38760 21693
rect 24970 20931 25526 20965
rect 25988 20931 26544 20965
rect 27006 20931 27562 20965
rect 28024 20931 28580 20965
rect 29042 20931 29598 20965
rect 30060 20931 30616 20965
rect 31078 20931 31634 20965
rect 32096 20931 32652 20965
rect 33114 20931 33670 20965
rect 34132 20931 34688 20965
rect 35150 20931 35706 20965
rect 36168 20931 36724 20965
rect 37186 20931 37742 20965
rect 38204 20931 38760 20965
rect 24762 20055 25318 20089
rect 25780 20055 26336 20089
rect 26798 20055 27354 20089
rect 27816 20055 28372 20089
rect 28834 20055 29390 20089
rect 29852 20055 30408 20089
rect 30870 20055 31426 20089
rect 31888 20055 32444 20089
rect 32906 20055 33462 20089
rect 33924 20055 34480 20089
rect 34942 20055 35498 20089
rect 35960 20055 36516 20089
rect 36978 20055 37534 20089
rect 37996 20055 38552 20089
rect 39014 20055 39570 20089
rect 19458 19951 20014 19985
rect 20476 19951 21032 19985
rect 21494 19951 22050 19985
rect 22512 19951 23068 19985
rect 24762 19327 25318 19361
rect 25780 19327 26336 19361
rect 26798 19327 27354 19361
rect 27816 19327 28372 19361
rect 28834 19327 29390 19361
rect 29852 19327 30408 19361
rect 30870 19327 31426 19361
rect 31888 19327 32444 19361
rect 32906 19327 33462 19361
rect 33924 19327 34480 19361
rect 34942 19327 35498 19361
rect 35960 19327 36516 19361
rect 36978 19327 37534 19361
rect 37996 19327 38552 19361
rect 39014 19327 39570 19361
rect 19458 19223 20014 19257
rect 20476 19223 21032 19257
rect 21494 19223 22050 19257
rect 22512 19223 23068 19257
rect 19458 18919 20014 18953
rect 20476 18919 21032 18953
rect 21494 18919 22050 18953
rect 22512 18919 23068 18953
rect 24762 18799 25318 18833
rect 25780 18799 26336 18833
rect 26798 18799 27354 18833
rect 27816 18799 28372 18833
rect 28834 18799 29390 18833
rect 29852 18799 30408 18833
rect 30870 18799 31426 18833
rect 31888 18799 32444 18833
rect 32906 18799 33462 18833
rect 33924 18799 34480 18833
rect 34942 18799 35498 18833
rect 35960 18799 36516 18833
rect 36978 18799 37534 18833
rect 37996 18799 38552 18833
rect 39014 18799 39570 18833
rect 19458 18191 20014 18225
rect 20476 18191 21032 18225
rect 21494 18191 22050 18225
rect 22512 18191 23068 18225
rect 24762 18071 25318 18105
rect 25780 18071 26336 18105
rect 26798 18071 27354 18105
rect 27816 18071 28372 18105
rect 28834 18071 29390 18105
rect 29852 18071 30408 18105
rect 30870 18071 31426 18105
rect 31888 18071 32444 18105
rect 32906 18071 33462 18105
rect 33924 18071 34480 18105
rect 34942 18071 35498 18105
rect 35960 18071 36516 18105
rect 36978 18071 37534 18105
rect 37996 18071 38552 18105
rect 39014 18071 39570 18105
rect 19458 17887 20014 17921
rect 20476 17887 21032 17921
rect 21494 17887 22050 17921
rect 22512 17887 23068 17921
rect 24762 17543 25318 17577
rect 25780 17543 26336 17577
rect 26798 17543 27354 17577
rect 27816 17543 28372 17577
rect 28834 17543 29390 17577
rect 29852 17543 30408 17577
rect 30870 17543 31426 17577
rect 31888 17543 32444 17577
rect 32906 17543 33462 17577
rect 33924 17543 34480 17577
rect 34942 17543 35498 17577
rect 35960 17543 36516 17577
rect 36978 17543 37534 17577
rect 37996 17543 38552 17577
rect 39014 17543 39570 17577
rect 19458 17159 20014 17193
rect 20476 17159 21032 17193
rect 21494 17159 22050 17193
rect 22512 17159 23068 17193
rect 19458 16855 20014 16889
rect 20476 16855 21032 16889
rect 21494 16855 22050 16889
rect 22512 16855 23068 16889
rect 24762 16815 25318 16849
rect 25780 16815 26336 16849
rect 26798 16815 27354 16849
rect 27816 16815 28372 16849
rect 28834 16815 29390 16849
rect 29852 16815 30408 16849
rect 30870 16815 31426 16849
rect 31888 16815 32444 16849
rect 32906 16815 33462 16849
rect 33924 16815 34480 16849
rect 34942 16815 35498 16849
rect 35960 16815 36516 16849
rect 36978 16815 37534 16849
rect 37996 16815 38552 16849
rect 39014 16815 39570 16849
rect 24762 16287 25318 16321
rect 25780 16287 26336 16321
rect 26798 16287 27354 16321
rect 27816 16287 28372 16321
rect 28834 16287 29390 16321
rect 29852 16287 30408 16321
rect 30870 16287 31426 16321
rect 31888 16287 32444 16321
rect 32906 16287 33462 16321
rect 33924 16287 34480 16321
rect 34942 16287 35498 16321
rect 35960 16287 36516 16321
rect 36978 16287 37534 16321
rect 37996 16287 38552 16321
rect 39014 16287 39570 16321
rect 19458 16127 20014 16161
rect 20476 16127 21032 16161
rect 21494 16127 22050 16161
rect 22512 16127 23068 16161
rect 24762 15559 25318 15593
rect 25780 15559 26336 15593
rect 26798 15559 27354 15593
rect 27816 15559 28372 15593
rect 28834 15559 29390 15593
rect 29852 15559 30408 15593
rect 30870 15559 31426 15593
rect 31888 15559 32444 15593
rect 32906 15559 33462 15593
rect 33924 15559 34480 15593
rect 34942 15559 35498 15593
rect 35960 15559 36516 15593
rect 36978 15559 37534 15593
rect 37996 15559 38552 15593
rect 39014 15559 39570 15593
rect 382 480 482 514
rect 640 480 740 514
rect 898 480 998 514
rect 1156 480 1256 514
rect 1414 480 1514 514
rect 1672 480 1772 514
rect 1930 480 2030 514
rect 2188 480 2288 514
rect 2446 480 2546 514
rect 2704 480 2804 514
rect 2962 480 3062 514
rect 3220 480 3320 514
rect 3478 480 3578 514
rect 3736 480 3836 514
rect 382 -30 482 4
rect 640 -30 740 4
rect 898 -30 998 4
rect 1156 -30 1256 4
rect 1414 -30 1514 4
rect 1672 -30 1772 4
rect 1930 -30 2030 4
rect 2188 -30 2288 4
rect 2446 -30 2546 4
rect 2704 -30 2804 4
rect 2962 -30 3062 4
rect 3220 -30 3320 4
rect 3478 -30 3578 4
rect 3736 -30 3836 4
rect 382 -520 482 -486
rect 640 -520 740 -486
rect 898 -520 998 -486
rect 1156 -520 1256 -486
rect 1414 -520 1514 -486
rect 1672 -520 1772 -486
rect 1930 -520 2030 -486
rect 2188 -520 2288 -486
rect 2446 -520 2546 -486
rect 2704 -520 2804 -486
rect 2962 -520 3062 -486
rect 3220 -520 3320 -486
rect 3478 -520 3578 -486
rect 3736 -520 3836 -486
rect 382 -1030 482 -996
rect 640 -1030 740 -996
rect 898 -1030 998 -996
rect 1156 -1030 1256 -996
rect 1414 -1030 1514 -996
rect 1672 -1030 1772 -996
rect 1930 -1030 2030 -996
rect 2188 -1030 2288 -996
rect 2446 -1030 2546 -996
rect 2704 -1030 2804 -996
rect 2962 -1030 3062 -996
rect 3220 -1030 3320 -996
rect 3478 -1030 3578 -996
rect 3736 -1030 3836 -996
rect 19870 13082 20426 13116
rect 20888 13082 21444 13116
rect 21906 13082 22462 13116
rect 22924 13082 23480 13116
rect 23942 13082 24498 13116
rect 24960 13082 25516 13116
rect 25978 13082 26534 13116
rect 26996 13082 27552 13116
rect 28014 13082 28570 13116
rect 29032 13082 29588 13116
rect 30050 13082 30606 13116
rect 31068 13082 31624 13116
rect 32086 13082 32642 13116
rect 33104 13082 33660 13116
rect 34122 13082 34678 13116
rect 35140 13082 35696 13116
rect 36158 13082 36714 13116
rect 37176 13082 37732 13116
rect 38194 13082 38750 13116
rect 39212 13082 39768 13116
rect 8104 12606 8660 12640
rect 9122 12606 9678 12640
rect 10140 12606 10696 12640
rect 11158 12606 11714 12640
rect 12176 12606 12732 12640
rect 13194 12606 13750 12640
rect 14212 12606 14768 12640
rect 15230 12606 15786 12640
rect 16248 12606 16804 12640
rect 19870 12372 20426 12406
rect 20888 12372 21444 12406
rect 21906 12372 22462 12406
rect 22924 12372 23480 12406
rect 23942 12372 24498 12406
rect 24960 12372 25516 12406
rect 25978 12372 26534 12406
rect 26996 12372 27552 12406
rect 28014 12372 28570 12406
rect 29032 12372 29588 12406
rect 30050 12372 30606 12406
rect 31068 12372 31624 12406
rect 32086 12372 32642 12406
rect 33104 12372 33660 12406
rect 34122 12372 34678 12406
rect 35140 12372 35696 12406
rect 36158 12372 36714 12406
rect 37176 12372 37732 12406
rect 38194 12372 38750 12406
rect 39212 12372 39768 12406
rect 19870 12264 20426 12298
rect 20888 12264 21444 12298
rect 21906 12264 22462 12298
rect 22924 12264 23480 12298
rect 23942 12264 24498 12298
rect 24960 12264 25516 12298
rect 25978 12264 26534 12298
rect 26996 12264 27552 12298
rect 28014 12264 28570 12298
rect 29032 12264 29588 12298
rect 30050 12264 30606 12298
rect 31068 12264 31624 12298
rect 32086 12264 32642 12298
rect 33104 12264 33660 12298
rect 34122 12264 34678 12298
rect 35140 12264 35696 12298
rect 36158 12264 36714 12298
rect 37176 12264 37732 12298
rect 38194 12264 38750 12298
rect 39212 12264 39768 12298
rect 8104 11896 8660 11930
rect 9122 11896 9678 11930
rect 8104 11788 8660 11822
rect 10140 11896 10696 11930
rect 9122 11788 9678 11822
rect 11158 11896 11714 11930
rect 10140 11788 10696 11822
rect 12176 11896 12732 11930
rect 11158 11788 11714 11822
rect 13194 11896 13750 11930
rect 12176 11788 12732 11822
rect 14212 11896 14768 11930
rect 13194 11788 13750 11822
rect 15230 11896 15786 11930
rect 14212 11788 14768 11822
rect 16248 11896 16804 11930
rect 15230 11788 15786 11822
rect 16248 11788 16804 11822
rect 19870 11554 20426 11588
rect 20888 11554 21444 11588
rect 21906 11554 22462 11588
rect 22924 11554 23480 11588
rect 23942 11554 24498 11588
rect 24960 11554 25516 11588
rect 25978 11554 26534 11588
rect 26996 11554 27552 11588
rect 28014 11554 28570 11588
rect 29032 11554 29588 11588
rect 30050 11554 30606 11588
rect 31068 11554 31624 11588
rect 32086 11554 32642 11588
rect 33104 11554 33660 11588
rect 34122 11554 34678 11588
rect 35140 11554 35696 11588
rect 36158 11554 36714 11588
rect 37176 11554 37732 11588
rect 38194 11554 38750 11588
rect 39212 11554 39768 11588
rect 8104 11078 8660 11112
rect 9122 11078 9678 11112
rect 8104 10970 8660 11004
rect 10140 11078 10696 11112
rect 9122 10970 9678 11004
rect 11158 11078 11714 11112
rect 10140 10970 10696 11004
rect 12176 11078 12732 11112
rect 11158 10970 11714 11004
rect 13194 11078 13750 11112
rect 12176 10970 12732 11004
rect 14212 11078 14768 11112
rect 13194 10970 13750 11004
rect 15230 11078 15786 11112
rect 14212 10970 14768 11004
rect 16248 11078 16804 11112
rect 15230 10970 15786 11004
rect 16248 10970 16804 11004
rect 19870 10886 20426 10920
rect 20888 10886 21444 10920
rect 21906 10886 22462 10920
rect 22924 10886 23480 10920
rect 23942 10886 24498 10920
rect 24960 10886 25516 10920
rect 25978 10886 26534 10920
rect 26996 10886 27552 10920
rect 28014 10886 28570 10920
rect 29032 10886 29588 10920
rect 30050 10886 30606 10920
rect 31068 10886 31624 10920
rect 32086 10886 32642 10920
rect 33104 10886 33660 10920
rect 34122 10886 34678 10920
rect 35140 10886 35696 10920
rect 36158 10886 36714 10920
rect 37176 10886 37732 10920
rect 38194 10886 38750 10920
rect 39212 10886 39768 10920
rect 8104 10260 8660 10294
rect 9122 10260 9678 10294
rect 8104 10152 8660 10186
rect 10140 10260 10696 10294
rect 9122 10152 9678 10186
rect 11158 10260 11714 10294
rect 10140 10152 10696 10186
rect 12176 10260 12732 10294
rect 11158 10152 11714 10186
rect 13194 10260 13750 10294
rect 12176 10152 12732 10186
rect 14212 10260 14768 10294
rect 13194 10152 13750 10186
rect 15230 10260 15786 10294
rect 14212 10152 14768 10186
rect 16248 10260 16804 10294
rect 15230 10152 15786 10186
rect 16248 10152 16804 10186
rect 19870 10176 20426 10210
rect 20888 10176 21444 10210
rect 21906 10176 22462 10210
rect 22924 10176 23480 10210
rect 23942 10176 24498 10210
rect 24960 10176 25516 10210
rect 25978 10176 26534 10210
rect 26996 10176 27552 10210
rect 28014 10176 28570 10210
rect 29032 10176 29588 10210
rect 30050 10176 30606 10210
rect 31068 10176 31624 10210
rect 32086 10176 32642 10210
rect 33104 10176 33660 10210
rect 34122 10176 34678 10210
rect 35140 10176 35696 10210
rect 36158 10176 36714 10210
rect 37176 10176 37732 10210
rect 38194 10176 38750 10210
rect 39212 10176 39768 10210
rect 19870 9654 20426 9688
rect 20888 9654 21444 9688
rect 21906 9654 22462 9688
rect 22924 9654 23480 9688
rect 23942 9654 24498 9688
rect 24960 9654 25516 9688
rect 25978 9654 26534 9688
rect 26996 9654 27552 9688
rect 28014 9654 28570 9688
rect 29032 9654 29588 9688
rect 30050 9654 30606 9688
rect 31068 9654 31624 9688
rect 32086 9654 32642 9688
rect 33104 9654 33660 9688
rect 34122 9654 34678 9688
rect 35140 9654 35696 9688
rect 36158 9654 36714 9688
rect 37176 9654 37732 9688
rect 38194 9654 38750 9688
rect 39212 9654 39768 9688
rect 8104 9442 8660 9476
rect 9122 9442 9678 9476
rect 8104 9334 8660 9368
rect 10140 9442 10696 9476
rect 9122 9334 9678 9368
rect 11158 9442 11714 9476
rect 10140 9334 10696 9368
rect 12176 9442 12732 9476
rect 11158 9334 11714 9368
rect 13194 9442 13750 9476
rect 12176 9334 12732 9368
rect 14212 9442 14768 9476
rect 13194 9334 13750 9368
rect 15230 9442 15786 9476
rect 14212 9334 14768 9368
rect 16248 9442 16804 9476
rect 15230 9334 15786 9368
rect 16248 9334 16804 9368
rect 19870 8944 20426 8978
rect 20888 8944 21444 8978
rect 21906 8944 22462 8978
rect 22924 8944 23480 8978
rect 23942 8944 24498 8978
rect 24960 8944 25516 8978
rect 25978 8944 26534 8978
rect 26996 8944 27552 8978
rect 28014 8944 28570 8978
rect 29032 8944 29588 8978
rect 30050 8944 30606 8978
rect 31068 8944 31624 8978
rect 32086 8944 32642 8978
rect 33104 8944 33660 8978
rect 34122 8944 34678 8978
rect 35140 8944 35696 8978
rect 36158 8944 36714 8978
rect 37176 8944 37732 8978
rect 38194 8944 38750 8978
rect 39212 8944 39768 8978
rect 8104 8624 8660 8658
rect 9122 8624 9678 8658
rect 8104 8516 8660 8550
rect 10140 8624 10696 8658
rect 9122 8516 9678 8550
rect 11158 8624 11714 8658
rect 10140 8516 10696 8550
rect 12176 8624 12732 8658
rect 11158 8516 11714 8550
rect 13194 8624 13750 8658
rect 12176 8516 12732 8550
rect 14212 8624 14768 8658
rect 13194 8516 13750 8550
rect 15230 8624 15786 8658
rect 14212 8516 14768 8550
rect 16248 8624 16804 8658
rect 15230 8516 15786 8550
rect 16248 8516 16804 8550
rect 19868 8420 20424 8454
rect 20886 8420 21442 8454
rect 21904 8420 22460 8454
rect 22922 8420 23478 8454
rect 23940 8420 24496 8454
rect 24958 8420 25514 8454
rect 25976 8420 26532 8454
rect 26994 8420 27550 8454
rect 28012 8420 28568 8454
rect 29030 8420 29586 8454
rect 30048 8420 30604 8454
rect 31066 8420 31622 8454
rect 32084 8420 32640 8454
rect 33102 8420 33658 8454
rect 34120 8420 34676 8454
rect 35138 8420 35694 8454
rect 36156 8420 36712 8454
rect 37174 8420 37730 8454
rect 38192 8420 38748 8454
rect 39210 8420 39766 8454
rect 8104 7806 8660 7840
rect 9122 7806 9678 7840
rect 8104 7698 8660 7732
rect 10140 7806 10696 7840
rect 9122 7698 9678 7732
rect 11158 7806 11714 7840
rect 10140 7698 10696 7732
rect 12176 7806 12732 7840
rect 11158 7698 11714 7732
rect 13194 7806 13750 7840
rect 12176 7698 12732 7732
rect 14212 7806 14768 7840
rect 13194 7698 13750 7732
rect 15230 7806 15786 7840
rect 14212 7698 14768 7732
rect 16248 7806 16804 7840
rect 15230 7698 15786 7732
rect 16248 7698 16804 7732
rect 19868 7710 20424 7744
rect 20886 7710 21442 7744
rect 21904 7710 22460 7744
rect 22922 7710 23478 7744
rect 23940 7710 24496 7744
rect 24958 7710 25514 7744
rect 25976 7710 26532 7744
rect 26994 7710 27550 7744
rect 28012 7710 28568 7744
rect 29030 7710 29586 7744
rect 30048 7710 30604 7744
rect 31066 7710 31622 7744
rect 32084 7710 32640 7744
rect 33102 7710 33658 7744
rect 34120 7710 34676 7744
rect 35138 7710 35694 7744
rect 36156 7710 36712 7744
rect 37174 7710 37730 7744
rect 38192 7710 38748 7744
rect 39210 7710 39766 7744
rect 19868 7186 20424 7220
rect 20886 7186 21442 7220
rect 21904 7186 22460 7220
rect 22922 7186 23478 7220
rect 23940 7186 24496 7220
rect 24958 7186 25514 7220
rect 25976 7186 26532 7220
rect 26994 7186 27550 7220
rect 28012 7186 28568 7220
rect 29030 7186 29586 7220
rect 30048 7186 30604 7220
rect 31066 7186 31622 7220
rect 32084 7186 32640 7220
rect 33102 7186 33658 7220
rect 34120 7186 34676 7220
rect 35138 7186 35694 7220
rect 36156 7186 36712 7220
rect 37174 7186 37730 7220
rect 38192 7186 38748 7220
rect 39210 7186 39766 7220
rect 8104 6988 8660 7022
rect 9122 6988 9678 7022
rect 8104 6880 8660 6914
rect 10140 6988 10696 7022
rect 9122 6880 9678 6914
rect 11158 6988 11714 7022
rect 10140 6880 10696 6914
rect 12176 6988 12732 7022
rect 11158 6880 11714 6914
rect 13194 6988 13750 7022
rect 12176 6880 12732 6914
rect 14212 6988 14768 7022
rect 13194 6880 13750 6914
rect 15230 6988 15786 7022
rect 14212 6880 14768 6914
rect 16248 6988 16804 7022
rect 15230 6880 15786 6914
rect 16248 6880 16804 6914
rect 19868 6476 20424 6510
rect 20886 6476 21442 6510
rect 21904 6476 22460 6510
rect 22922 6476 23478 6510
rect 23940 6476 24496 6510
rect 24958 6476 25514 6510
rect 25976 6476 26532 6510
rect 26994 6476 27550 6510
rect 28012 6476 28568 6510
rect 29030 6476 29586 6510
rect 30048 6476 30604 6510
rect 31066 6476 31622 6510
rect 32084 6476 32640 6510
rect 33102 6476 33658 6510
rect 34120 6476 34676 6510
rect 35138 6476 35694 6510
rect 36156 6476 36712 6510
rect 37174 6476 37730 6510
rect 38192 6476 38748 6510
rect 39210 6476 39766 6510
rect 8104 6170 8660 6204
rect 9122 6170 9678 6204
rect 10140 6170 10696 6204
rect 11158 6170 11714 6204
rect 12176 6170 12732 6204
rect 13194 6170 13750 6204
rect 14212 6170 14768 6204
rect 15230 6170 15786 6204
rect 16248 6170 16804 6204
rect 19868 5954 20424 5988
rect 20886 5954 21442 5988
rect 21904 5954 22460 5988
rect 22922 5954 23478 5988
rect 23940 5954 24496 5988
rect 24958 5954 25514 5988
rect 25976 5954 26532 5988
rect 26994 5954 27550 5988
rect 28012 5954 28568 5988
rect 29030 5954 29586 5988
rect 30048 5954 30604 5988
rect 31066 5954 31622 5988
rect 32084 5954 32640 5988
rect 33102 5954 33658 5988
rect 34120 5954 34676 5988
rect 35138 5954 35694 5988
rect 36156 5954 36712 5988
rect 37174 5954 37730 5988
rect 38192 5954 38748 5988
rect 39210 5954 39766 5988
rect 19868 5244 20424 5278
rect 20886 5244 21442 5278
rect 21904 5244 22460 5278
rect 22922 5244 23478 5278
rect 23940 5244 24496 5278
rect 24958 5244 25514 5278
rect 25976 5244 26532 5278
rect 26994 5244 27550 5278
rect 28012 5244 28568 5278
rect 29030 5244 29586 5278
rect 30048 5244 30604 5278
rect 31066 5244 31622 5278
rect 32084 5244 32640 5278
rect 33102 5244 33658 5278
rect 34120 5244 34676 5278
rect 35138 5244 35694 5278
rect 36156 5244 36712 5278
rect 37174 5244 37730 5278
rect 38192 5244 38748 5278
rect 39210 5244 39766 5278
rect 6780 4856 7336 4890
rect 7798 4856 8354 4890
rect 8816 4856 9372 4890
rect 9834 4856 10390 4890
rect 10852 4856 11408 4890
rect 11870 4856 12426 4890
rect 12888 4856 13444 4890
rect 13906 4856 14462 4890
rect 14924 4856 15480 4890
rect 15942 4856 16498 4890
rect 16960 4856 17516 4890
rect 19868 4720 20424 4754
rect 20886 4720 21442 4754
rect 21904 4720 22460 4754
rect 22922 4720 23478 4754
rect 23940 4720 24496 4754
rect 24958 4720 25514 4754
rect 25976 4720 26532 4754
rect 26994 4720 27550 4754
rect 28012 4720 28568 4754
rect 29030 4720 29586 4754
rect 30048 4720 30604 4754
rect 31066 4720 31622 4754
rect 32084 4720 32640 4754
rect 33102 4720 33658 4754
rect 34120 4720 34676 4754
rect 35138 4720 35694 4754
rect 36156 4720 36712 4754
rect 37174 4720 37730 4754
rect 38192 4720 38748 4754
rect 39210 4720 39766 4754
rect 6780 4146 7336 4180
rect 7798 4146 8354 4180
rect 8816 4146 9372 4180
rect 9834 4146 10390 4180
rect 10852 4146 11408 4180
rect 11870 4146 12426 4180
rect 12888 4146 13444 4180
rect 13906 4146 14462 4180
rect 14924 4146 15480 4180
rect 15942 4146 16498 4180
rect 16960 4146 17516 4180
rect 19868 4010 20424 4044
rect 20886 4010 21442 4044
rect 21904 4010 22460 4044
rect 22922 4010 23478 4044
rect 23940 4010 24496 4044
rect 24958 4010 25514 4044
rect 25976 4010 26532 4044
rect 26994 4010 27550 4044
rect 28012 4010 28568 4044
rect 29030 4010 29586 4044
rect 30048 4010 30604 4044
rect 31066 4010 31622 4044
rect 32084 4010 32640 4044
rect 33102 4010 33658 4044
rect 34120 4010 34676 4044
rect 35138 4010 35694 4044
rect 36156 4010 36712 4044
rect 37174 4010 37730 4044
rect 38192 4010 38748 4044
rect 39210 4010 39766 4044
rect 6780 3744 7336 3778
rect 7798 3744 8354 3778
rect 8816 3744 9372 3778
rect 9834 3744 10390 3778
rect 10852 3744 11408 3778
rect 11870 3744 12426 3778
rect 12888 3744 13444 3778
rect 13906 3744 14462 3778
rect 14924 3744 15480 3778
rect 15942 3744 16498 3778
rect 16960 3744 17516 3778
rect 19868 3486 20424 3520
rect 20886 3486 21442 3520
rect 21904 3486 22460 3520
rect 22922 3486 23478 3520
rect 23940 3486 24496 3520
rect 24958 3486 25514 3520
rect 25976 3486 26532 3520
rect 26994 3486 27550 3520
rect 28012 3486 28568 3520
rect 29030 3486 29586 3520
rect 30048 3486 30604 3520
rect 31066 3486 31622 3520
rect 32084 3486 32640 3520
rect 33102 3486 33658 3520
rect 34120 3486 34676 3520
rect 35138 3486 35694 3520
rect 36156 3486 36712 3520
rect 37174 3486 37730 3520
rect 38192 3486 38748 3520
rect 39210 3486 39766 3520
rect 6780 3034 7336 3068
rect 7798 3034 8354 3068
rect 8816 3034 9372 3068
rect 9834 3034 10390 3068
rect 10852 3034 11408 3068
rect 11870 3034 12426 3068
rect 12888 3034 13444 3068
rect 13906 3034 14462 3068
rect 14924 3034 15480 3068
rect 15942 3034 16498 3068
rect 16960 3034 17516 3068
rect 19868 2776 20424 2810
rect 20886 2776 21442 2810
rect 21904 2776 22460 2810
rect 22922 2776 23478 2810
rect 23940 2776 24496 2810
rect 24958 2776 25514 2810
rect 25976 2776 26532 2810
rect 26994 2776 27550 2810
rect 28012 2776 28568 2810
rect 29030 2776 29586 2810
rect 30048 2776 30604 2810
rect 31066 2776 31622 2810
rect 32084 2776 32640 2810
rect 33102 2776 33658 2810
rect 34120 2776 34676 2810
rect 35138 2776 35694 2810
rect 36156 2776 36712 2810
rect 37174 2776 37730 2810
rect 38192 2776 38748 2810
rect 39210 2776 39766 2810
rect 6780 2632 7336 2666
rect 7798 2632 8354 2666
rect 8816 2632 9372 2666
rect 9834 2632 10390 2666
rect 10852 2632 11408 2666
rect 11870 2632 12426 2666
rect 12888 2632 13444 2666
rect 13906 2632 14462 2666
rect 14924 2632 15480 2666
rect 15942 2632 16498 2666
rect 16960 2632 17516 2666
rect 19868 2254 20424 2288
rect 20886 2254 21442 2288
rect 21904 2254 22460 2288
rect 22922 2254 23478 2288
rect 23940 2254 24496 2288
rect 24958 2254 25514 2288
rect 25976 2254 26532 2288
rect 26994 2254 27550 2288
rect 28012 2254 28568 2288
rect 29030 2254 29586 2288
rect 30048 2254 30604 2288
rect 31066 2254 31622 2288
rect 32084 2254 32640 2288
rect 33102 2254 33658 2288
rect 34120 2254 34676 2288
rect 35138 2254 35694 2288
rect 36156 2254 36712 2288
rect 37174 2254 37730 2288
rect 38192 2254 38748 2288
rect 39210 2254 39766 2288
rect 6780 1922 7336 1956
rect 7798 1922 8354 1956
rect 8816 1922 9372 1956
rect 9834 1922 10390 1956
rect 10852 1922 11408 1956
rect 11870 1922 12426 1956
rect 12888 1922 13444 1956
rect 13906 1922 14462 1956
rect 14924 1922 15480 1956
rect 15942 1922 16498 1956
rect 16960 1922 17516 1956
rect 6780 1520 7336 1554
rect 7798 1520 8354 1554
rect 8816 1520 9372 1554
rect 9834 1520 10390 1554
rect 10852 1520 11408 1554
rect 11870 1520 12426 1554
rect 12888 1520 13444 1554
rect 13906 1520 14462 1554
rect 14924 1520 15480 1554
rect 15942 1520 16498 1554
rect 16960 1520 17516 1554
rect 19868 1544 20424 1578
rect 20886 1544 21442 1578
rect 21904 1544 22460 1578
rect 22922 1544 23478 1578
rect 23940 1544 24496 1578
rect 24958 1544 25514 1578
rect 25976 1544 26532 1578
rect 26994 1544 27550 1578
rect 28012 1544 28568 1578
rect 29030 1544 29586 1578
rect 30048 1544 30604 1578
rect 31066 1544 31622 1578
rect 32084 1544 32640 1578
rect 33102 1544 33658 1578
rect 34120 1544 34676 1578
rect 35138 1544 35694 1578
rect 36156 1544 36712 1578
rect 37174 1544 37730 1578
rect 38192 1544 38748 1578
rect 39210 1544 39766 1578
rect 19868 1020 20424 1054
rect 20886 1020 21442 1054
rect 21904 1020 22460 1054
rect 22922 1020 23478 1054
rect 23940 1020 24496 1054
rect 24958 1020 25514 1054
rect 25976 1020 26532 1054
rect 26994 1020 27550 1054
rect 28012 1020 28568 1054
rect 29030 1020 29586 1054
rect 30048 1020 30604 1054
rect 31066 1020 31622 1054
rect 32084 1020 32640 1054
rect 33102 1020 33658 1054
rect 34120 1020 34676 1054
rect 35138 1020 35694 1054
rect 36156 1020 36712 1054
rect 37174 1020 37730 1054
rect 38192 1020 38748 1054
rect 39210 1020 39766 1054
rect 6780 810 7336 844
rect 7798 810 8354 844
rect 8816 810 9372 844
rect 9834 810 10390 844
rect 10852 810 11408 844
rect 11870 810 12426 844
rect 12888 810 13444 844
rect 13906 810 14462 844
rect 14924 810 15480 844
rect 15942 810 16498 844
rect 16960 810 17516 844
rect 19868 310 20424 344
rect 20886 310 21442 344
rect 21904 310 22460 344
rect 22922 310 23478 344
rect 23940 310 24496 344
rect 24958 310 25514 344
rect 25976 310 26532 344
rect 26994 310 27550 344
rect 28012 310 28568 344
rect 29030 310 29586 344
rect 30048 310 30604 344
rect 31066 310 31622 344
rect 32084 310 32640 344
rect 33102 310 33658 344
rect 34120 310 34676 344
rect 35138 310 35694 344
rect 36156 310 36712 344
rect 37174 310 37730 344
rect 38192 310 38748 344
rect 39210 310 39766 344
rect 7238 -22 7794 12
rect 8256 -22 8812 12
rect 9274 -22 9830 12
rect 10292 -22 10848 12
rect 11310 -22 11866 12
rect 12328 -22 12884 12
rect 13346 -22 13902 12
rect 14364 -22 14920 12
rect 15382 -22 15938 12
rect 16400 -22 16956 12
rect 19868 -212 20424 -178
rect 20886 -212 21442 -178
rect 21904 -212 22460 -178
rect 22922 -212 23478 -178
rect 23940 -212 24496 -178
rect 24958 -212 25514 -178
rect 25976 -212 26532 -178
rect 26994 -212 27550 -178
rect 28012 -212 28568 -178
rect 29030 -212 29586 -178
rect 30048 -212 30604 -178
rect 31066 -212 31622 -178
rect 32084 -212 32640 -178
rect 33102 -212 33658 -178
rect 34120 -212 34676 -178
rect 35138 -212 35694 -178
rect 36156 -212 36712 -178
rect 37174 -212 37730 -178
rect 38192 -212 38748 -178
rect 39210 -212 39766 -178
rect 7238 -732 7794 -698
rect 8256 -732 8812 -698
rect 9274 -732 9830 -698
rect 10292 -732 10848 -698
rect 11310 -732 11866 -698
rect 12328 -732 12884 -698
rect 13346 -732 13902 -698
rect 14364 -732 14920 -698
rect 15382 -732 15938 -698
rect 16400 -732 16956 -698
rect 19868 -922 20424 -888
rect 20886 -922 21442 -888
rect 21904 -922 22460 -888
rect 22922 -922 23478 -888
rect 23940 -922 24496 -888
rect 24958 -922 25514 -888
rect 25976 -922 26532 -888
rect 26994 -922 27550 -888
rect 28012 -922 28568 -888
rect 29030 -922 29586 -888
rect 30048 -922 30604 -888
rect 31066 -922 31622 -888
rect 32084 -922 32640 -888
rect 33102 -922 33658 -888
rect 34120 -922 34676 -888
rect 35138 -922 35694 -888
rect 36156 -922 36712 -888
rect 37174 -922 37730 -888
rect 38192 -922 38748 -888
rect 39210 -922 39766 -888
<< locali >>
rect 17418 29240 17518 29402
rect 41762 29240 41862 29402
rect 24008 26858 24098 26888
rect 24008 26824 24036 26858
rect 24070 26824 24098 26858
rect 24008 26796 24098 26824
rect 25026 26858 25116 26888
rect 25026 26824 25054 26858
rect 25088 26824 25116 26858
rect 25026 26796 25116 26824
rect 26044 26858 26134 26888
rect 26044 26824 26072 26858
rect 26106 26824 26134 26858
rect 26044 26796 26134 26824
rect 27062 26858 27152 26888
rect 27062 26824 27090 26858
rect 27124 26824 27152 26858
rect 27062 26796 27152 26824
rect 28080 26858 28170 26888
rect 28080 26824 28108 26858
rect 28142 26824 28170 26858
rect 28080 26796 28170 26824
rect 29098 26858 29188 26888
rect 29098 26824 29126 26858
rect 29160 26824 29188 26858
rect 29098 26796 29188 26824
rect 30116 26858 30206 26888
rect 30116 26824 30144 26858
rect 30178 26824 30206 26858
rect 30116 26796 30206 26824
rect 31134 26858 31224 26888
rect 31134 26824 31162 26858
rect 31196 26824 31224 26858
rect 31134 26796 31224 26824
rect 32152 26858 32242 26888
rect 32152 26824 32180 26858
rect 32214 26824 32242 26858
rect 32152 26796 32242 26824
rect 33170 26858 33260 26888
rect 33170 26824 33198 26858
rect 33232 26824 33260 26858
rect 33170 26796 33260 26824
rect 34188 26858 34278 26888
rect 34188 26824 34216 26858
rect 34250 26824 34278 26858
rect 34188 26796 34278 26824
rect 35206 26858 35296 26888
rect 35206 26824 35234 26858
rect 35268 26824 35296 26858
rect 35206 26796 35296 26824
rect 36224 26858 36314 26888
rect 36224 26824 36252 26858
rect 36286 26824 36314 26858
rect 36224 26796 36314 26824
rect 37242 26858 37332 26888
rect 37242 26824 37270 26858
rect 37304 26824 37332 26858
rect 37242 26796 37332 26824
rect 38260 26858 38350 26888
rect 38260 26824 38288 26858
rect 38322 26824 38350 26858
rect 38260 26796 38350 26824
rect 39278 26858 39368 26888
rect 39278 26824 39306 26858
rect 39340 26824 39368 26858
rect 39278 26796 39368 26824
rect 23760 26601 23776 26635
rect 24332 26601 24348 26635
rect 24778 26601 24794 26635
rect 25350 26601 25366 26635
rect 25796 26601 25812 26635
rect 26368 26601 26384 26635
rect 26814 26601 26830 26635
rect 27386 26601 27402 26635
rect 27832 26601 27848 26635
rect 28404 26601 28420 26635
rect 28850 26601 28866 26635
rect 29422 26601 29438 26635
rect 29868 26601 29884 26635
rect 30440 26601 30456 26635
rect 30886 26601 30902 26635
rect 31458 26601 31474 26635
rect 31904 26601 31920 26635
rect 32476 26601 32492 26635
rect 32922 26601 32938 26635
rect 33494 26601 33510 26635
rect 33940 26601 33956 26635
rect 34512 26601 34528 26635
rect 34958 26601 34974 26635
rect 35530 26601 35546 26635
rect 35976 26601 35992 26635
rect 36548 26601 36564 26635
rect 36994 26601 37010 26635
rect 37566 26601 37582 26635
rect 38012 26601 38028 26635
rect 38584 26601 38600 26635
rect 39030 26601 39046 26635
rect 39602 26601 39618 26635
rect 23528 26542 23562 26558
rect 23528 25950 23562 25966
rect 24546 26542 24580 26558
rect 24546 25950 24580 25966
rect 25564 26542 25598 26558
rect 25564 25950 25598 25966
rect 26582 26542 26616 26558
rect 26582 25950 26616 25966
rect 27600 26542 27634 26558
rect 27600 25950 27634 25966
rect 28618 26542 28652 26558
rect 28618 25950 28652 25966
rect 29636 26542 29670 26558
rect 29636 25950 29670 25966
rect 30654 26542 30688 26558
rect 30654 25950 30688 25966
rect 31672 26542 31706 26558
rect 31672 25950 31706 25966
rect 32690 26542 32724 26558
rect 32690 25950 32724 25966
rect 33708 26542 33742 26558
rect 33708 25950 33742 25966
rect 34726 26542 34760 26558
rect 34726 25950 34760 25966
rect 35744 26542 35778 26558
rect 35744 25950 35778 25966
rect 36762 26542 36796 26558
rect 36762 25950 36796 25966
rect 37780 26542 37814 26558
rect 37780 25950 37814 25966
rect 38798 26542 38832 26558
rect 38798 25950 38832 25966
rect 39816 26542 39850 26558
rect 39816 25950 39850 25966
rect 23760 25873 23776 25907
rect 24332 25873 24348 25907
rect 24778 25873 24794 25907
rect 25350 25873 25366 25907
rect 25796 25873 25812 25907
rect 26368 25873 26384 25907
rect 26814 25873 26830 25907
rect 27386 25873 27402 25907
rect 27832 25873 27848 25907
rect 28404 25873 28420 25907
rect 28850 25873 28866 25907
rect 29422 25873 29438 25907
rect 29868 25873 29884 25907
rect 30440 25873 30456 25907
rect 30886 25873 30902 25907
rect 31458 25873 31474 25907
rect 31904 25873 31920 25907
rect 32476 25873 32492 25907
rect 32922 25873 32938 25907
rect 33494 25873 33510 25907
rect 33940 25873 33956 25907
rect 34512 25873 34528 25907
rect 34958 25873 34974 25907
rect 35530 25873 35546 25907
rect 35976 25873 35992 25907
rect 36548 25873 36564 25907
rect 36994 25873 37010 25907
rect 37566 25873 37582 25907
rect 38012 25873 38028 25907
rect 38584 25873 38600 25907
rect 39030 25873 39046 25907
rect 39602 25873 39618 25907
rect 24030 25704 24120 25734
rect 24030 25670 24058 25704
rect 24092 25670 24120 25704
rect 24030 25642 24120 25670
rect 25048 25704 25138 25734
rect 25048 25670 25076 25704
rect 25110 25670 25138 25704
rect 25048 25642 25138 25670
rect 26066 25704 26156 25734
rect 26066 25670 26094 25704
rect 26128 25670 26156 25704
rect 26066 25642 26156 25670
rect 27084 25704 27174 25734
rect 27084 25670 27112 25704
rect 27146 25670 27174 25704
rect 27084 25642 27174 25670
rect 28102 25704 28192 25734
rect 28102 25670 28130 25704
rect 28164 25670 28192 25704
rect 28102 25642 28192 25670
rect 29120 25704 29210 25734
rect 29120 25670 29148 25704
rect 29182 25670 29210 25704
rect 29120 25642 29210 25670
rect 30138 25704 30228 25734
rect 30138 25670 30166 25704
rect 30200 25670 30228 25704
rect 30138 25642 30228 25670
rect 31156 25704 31246 25734
rect 31156 25670 31184 25704
rect 31218 25670 31246 25704
rect 31156 25642 31246 25670
rect 32174 25704 32264 25734
rect 32174 25670 32202 25704
rect 32236 25670 32264 25704
rect 32174 25642 32264 25670
rect 33192 25704 33282 25734
rect 33192 25670 33220 25704
rect 33254 25670 33282 25704
rect 33192 25642 33282 25670
rect 34210 25704 34300 25734
rect 34210 25670 34238 25704
rect 34272 25670 34300 25704
rect 34210 25642 34300 25670
rect 35228 25704 35318 25734
rect 35228 25670 35256 25704
rect 35290 25670 35318 25704
rect 35228 25642 35318 25670
rect 36246 25704 36336 25734
rect 36246 25670 36274 25704
rect 36308 25670 36336 25704
rect 36246 25642 36336 25670
rect 37264 25704 37354 25734
rect 37264 25670 37292 25704
rect 37326 25670 37354 25704
rect 37264 25642 37354 25670
rect 38282 25704 38372 25734
rect 38282 25670 38310 25704
rect 38344 25670 38372 25704
rect 38282 25642 38372 25670
rect 39300 25704 39390 25734
rect 39300 25670 39328 25704
rect 39362 25670 39390 25704
rect 39300 25642 39390 25670
rect 23760 25465 23776 25499
rect 24332 25465 24348 25499
rect 24778 25465 24794 25499
rect 25350 25465 25366 25499
rect 25796 25465 25812 25499
rect 26368 25465 26384 25499
rect 26814 25465 26830 25499
rect 27386 25465 27402 25499
rect 27832 25465 27848 25499
rect 28404 25465 28420 25499
rect 28850 25465 28866 25499
rect 29422 25465 29438 25499
rect 29868 25465 29884 25499
rect 30440 25465 30456 25499
rect 30886 25465 30902 25499
rect 31458 25465 31474 25499
rect 31904 25465 31920 25499
rect 32476 25465 32492 25499
rect 32922 25465 32938 25499
rect 33494 25465 33510 25499
rect 33940 25465 33956 25499
rect 34512 25465 34528 25499
rect 34958 25465 34974 25499
rect 35530 25465 35546 25499
rect 35976 25465 35992 25499
rect 36548 25465 36564 25499
rect 36994 25465 37010 25499
rect 37566 25465 37582 25499
rect 38012 25465 38028 25499
rect 38584 25465 38600 25499
rect 39030 25465 39046 25499
rect 39602 25465 39618 25499
rect 23528 25406 23562 25422
rect 23528 24814 23562 24830
rect 24546 25406 24580 25422
rect 24546 24814 24580 24830
rect 25564 25406 25598 25422
rect 25564 24814 25598 24830
rect 26582 25406 26616 25422
rect 26582 24814 26616 24830
rect 27600 25406 27634 25422
rect 27600 24814 27634 24830
rect 28618 25406 28652 25422
rect 28618 24814 28652 24830
rect 29636 25406 29670 25422
rect 29636 24814 29670 24830
rect 30654 25406 30688 25422
rect 30654 24814 30688 24830
rect 31672 25406 31706 25422
rect 31672 24814 31706 24830
rect 32690 25406 32724 25422
rect 32690 24814 32724 24830
rect 33708 25406 33742 25422
rect 33708 24814 33742 24830
rect 34726 25406 34760 25422
rect 34726 24814 34760 24830
rect 35744 25406 35778 25422
rect 35744 24814 35778 24830
rect 36762 25406 36796 25422
rect 36762 24814 36796 24830
rect 37780 25406 37814 25422
rect 37780 24814 37814 24830
rect 38798 25406 38832 25422
rect 38798 24814 38832 24830
rect 39816 25406 39850 25422
rect 39816 24814 39850 24830
rect 23760 24737 23776 24771
rect 24332 24737 24348 24771
rect 24778 24737 24794 24771
rect 25350 24737 25366 24771
rect 25796 24737 25812 24771
rect 26368 24737 26384 24771
rect 26814 24737 26830 24771
rect 27386 24737 27402 24771
rect 27832 24737 27848 24771
rect 28404 24737 28420 24771
rect 28850 24737 28866 24771
rect 29422 24737 29438 24771
rect 29868 24737 29884 24771
rect 30440 24737 30456 24771
rect 30886 24737 30902 24771
rect 31458 24737 31474 24771
rect 31904 24737 31920 24771
rect 32476 24737 32492 24771
rect 32922 24737 32938 24771
rect 33494 24737 33510 24771
rect 33940 24737 33956 24771
rect 34512 24737 34528 24771
rect 34958 24737 34974 24771
rect 35530 24737 35546 24771
rect 35976 24737 35992 24771
rect 36548 24737 36564 24771
rect 36994 24737 37010 24771
rect 37566 24737 37582 24771
rect 38012 24737 38028 24771
rect 38584 24737 38600 24771
rect 39030 24737 39046 24771
rect 39602 24737 39618 24771
rect 24008 24572 24098 24602
rect 24008 24538 24036 24572
rect 24070 24538 24098 24572
rect 24008 24510 24098 24538
rect 25026 24572 25116 24602
rect 25026 24538 25054 24572
rect 25088 24538 25116 24572
rect 25026 24510 25116 24538
rect 26044 24572 26134 24602
rect 26044 24538 26072 24572
rect 26106 24538 26134 24572
rect 26044 24510 26134 24538
rect 27062 24572 27152 24602
rect 27062 24538 27090 24572
rect 27124 24538 27152 24572
rect 27062 24510 27152 24538
rect 28080 24572 28170 24602
rect 28080 24538 28108 24572
rect 28142 24538 28170 24572
rect 28080 24510 28170 24538
rect 29098 24572 29188 24602
rect 29098 24538 29126 24572
rect 29160 24538 29188 24572
rect 29098 24510 29188 24538
rect 30116 24572 30206 24602
rect 30116 24538 30144 24572
rect 30178 24538 30206 24572
rect 30116 24510 30206 24538
rect 31134 24572 31224 24602
rect 31134 24538 31162 24572
rect 31196 24538 31224 24572
rect 31134 24510 31224 24538
rect 32152 24572 32242 24602
rect 32152 24538 32180 24572
rect 32214 24538 32242 24572
rect 32152 24510 32242 24538
rect 33170 24572 33260 24602
rect 33170 24538 33198 24572
rect 33232 24538 33260 24572
rect 33170 24510 33260 24538
rect 34188 24572 34278 24602
rect 34188 24538 34216 24572
rect 34250 24538 34278 24572
rect 34188 24510 34278 24538
rect 35206 24572 35296 24602
rect 35206 24538 35234 24572
rect 35268 24538 35296 24572
rect 35206 24510 35296 24538
rect 36224 24572 36314 24602
rect 36224 24538 36252 24572
rect 36286 24538 36314 24572
rect 36224 24510 36314 24538
rect 37242 24572 37332 24602
rect 37242 24538 37270 24572
rect 37304 24538 37332 24572
rect 37242 24510 37332 24538
rect 38260 24572 38350 24602
rect 38260 24538 38288 24572
rect 38322 24538 38350 24572
rect 38260 24510 38350 24538
rect 39278 24572 39368 24602
rect 39278 24538 39306 24572
rect 39340 24538 39368 24572
rect 39278 24510 39368 24538
rect 23760 24329 23776 24363
rect 24332 24329 24348 24363
rect 24778 24329 24794 24363
rect 25350 24329 25366 24363
rect 25796 24329 25812 24363
rect 26368 24329 26384 24363
rect 26814 24329 26830 24363
rect 27386 24329 27402 24363
rect 27832 24329 27848 24363
rect 28404 24329 28420 24363
rect 28850 24329 28866 24363
rect 29422 24329 29438 24363
rect 29868 24329 29884 24363
rect 30440 24329 30456 24363
rect 30886 24329 30902 24363
rect 31458 24329 31474 24363
rect 31904 24329 31920 24363
rect 32476 24329 32492 24363
rect 32922 24329 32938 24363
rect 33494 24329 33510 24363
rect 33940 24329 33956 24363
rect 34512 24329 34528 24363
rect 34958 24329 34974 24363
rect 35530 24329 35546 24363
rect 35976 24329 35992 24363
rect 36548 24329 36564 24363
rect 36994 24329 37010 24363
rect 37566 24329 37582 24363
rect 38012 24329 38028 24363
rect 38584 24329 38600 24363
rect 39030 24329 39046 24363
rect 39602 24329 39618 24363
rect 23528 24270 23562 24286
rect 23528 23678 23562 23694
rect 24546 24270 24580 24286
rect 24546 23678 24580 23694
rect 25564 24270 25598 24286
rect 25564 23678 25598 23694
rect 26582 24270 26616 24286
rect 26582 23678 26616 23694
rect 27600 24270 27634 24286
rect 27600 23678 27634 23694
rect 28618 24270 28652 24286
rect 28618 23678 28652 23694
rect 29636 24270 29670 24286
rect 29636 23678 29670 23694
rect 30654 24270 30688 24286
rect 30654 23678 30688 23694
rect 31672 24270 31706 24286
rect 31672 23678 31706 23694
rect 32690 24270 32724 24286
rect 32690 23678 32724 23694
rect 33708 24270 33742 24286
rect 33708 23678 33742 23694
rect 34726 24270 34760 24286
rect 34726 23678 34760 23694
rect 35744 24270 35778 24286
rect 35744 23678 35778 23694
rect 36762 24270 36796 24286
rect 36762 23678 36796 23694
rect 37780 24270 37814 24286
rect 37780 23678 37814 23694
rect 38798 24270 38832 24286
rect 38798 23678 38832 23694
rect 39816 24270 39850 24286
rect 39816 23678 39850 23694
rect 23760 23601 23776 23635
rect 24332 23601 24348 23635
rect 24778 23601 24794 23635
rect 25350 23601 25366 23635
rect 25796 23601 25812 23635
rect 26368 23601 26384 23635
rect 26814 23601 26830 23635
rect 27386 23601 27402 23635
rect 27832 23601 27848 23635
rect 28404 23601 28420 23635
rect 28850 23601 28866 23635
rect 29422 23601 29438 23635
rect 29868 23601 29884 23635
rect 30440 23601 30456 23635
rect 30886 23601 30902 23635
rect 31458 23601 31474 23635
rect 31904 23601 31920 23635
rect 32476 23601 32492 23635
rect 32922 23601 32938 23635
rect 33494 23601 33510 23635
rect 33940 23601 33956 23635
rect 34512 23601 34528 23635
rect 34958 23601 34974 23635
rect 35530 23601 35546 23635
rect 35976 23601 35992 23635
rect 36548 23601 36564 23635
rect 36994 23601 37010 23635
rect 37566 23601 37582 23635
rect 38012 23601 38028 23635
rect 38584 23601 38600 23635
rect 39030 23601 39046 23635
rect 39602 23601 39618 23635
rect 24008 23190 24098 23220
rect 24008 23156 24036 23190
rect 24070 23156 24098 23190
rect 24008 23128 24098 23156
rect 25026 23190 25116 23220
rect 25026 23156 25054 23190
rect 25088 23156 25116 23190
rect 25026 23128 25116 23156
rect 26044 23190 26134 23220
rect 26044 23156 26072 23190
rect 26106 23156 26134 23190
rect 26044 23128 26134 23156
rect 27062 23190 27152 23220
rect 27062 23156 27090 23190
rect 27124 23156 27152 23190
rect 27062 23128 27152 23156
rect 28080 23190 28170 23220
rect 28080 23156 28108 23190
rect 28142 23156 28170 23190
rect 28080 23128 28170 23156
rect 29098 23190 29188 23220
rect 29098 23156 29126 23190
rect 29160 23156 29188 23190
rect 29098 23128 29188 23156
rect 30116 23190 30206 23220
rect 30116 23156 30144 23190
rect 30178 23156 30206 23190
rect 30116 23128 30206 23156
rect 31134 23190 31224 23220
rect 31134 23156 31162 23190
rect 31196 23156 31224 23190
rect 31134 23128 31224 23156
rect 32152 23190 32242 23220
rect 32152 23156 32180 23190
rect 32214 23156 32242 23190
rect 32152 23128 32242 23156
rect 33170 23190 33260 23220
rect 33170 23156 33198 23190
rect 33232 23156 33260 23190
rect 33170 23128 33260 23156
rect 34188 23190 34278 23220
rect 34188 23156 34216 23190
rect 34250 23156 34278 23190
rect 34188 23128 34278 23156
rect 35206 23190 35296 23220
rect 35206 23156 35234 23190
rect 35268 23156 35296 23190
rect 35206 23128 35296 23156
rect 36224 23190 36314 23220
rect 36224 23156 36252 23190
rect 36286 23156 36314 23190
rect 36224 23128 36314 23156
rect 37242 23190 37332 23220
rect 37242 23156 37270 23190
rect 37304 23156 37332 23190
rect 37242 23128 37332 23156
rect 38260 23190 38350 23220
rect 38260 23156 38288 23190
rect 38322 23156 38350 23190
rect 38260 23128 38350 23156
rect 39278 23190 39368 23220
rect 39278 23156 39306 23190
rect 39340 23156 39368 23190
rect 39278 23128 39368 23156
rect 24954 22691 24970 22725
rect 25526 22691 25542 22725
rect 25972 22691 25988 22725
rect 26544 22691 26560 22725
rect 26990 22691 27006 22725
rect 27562 22691 27578 22725
rect 28008 22691 28024 22725
rect 28580 22691 28596 22725
rect 29026 22691 29042 22725
rect 29598 22691 29614 22725
rect 30044 22691 30060 22725
rect 30616 22691 30632 22725
rect 31062 22691 31078 22725
rect 31634 22691 31650 22725
rect 32080 22691 32096 22725
rect 32652 22691 32668 22725
rect 33098 22691 33114 22725
rect 33670 22691 33686 22725
rect 34116 22691 34132 22725
rect 34688 22691 34704 22725
rect 35134 22691 35150 22725
rect 35706 22691 35722 22725
rect 36152 22691 36168 22725
rect 36724 22691 36740 22725
rect 37170 22691 37186 22725
rect 37742 22691 37758 22725
rect 38188 22691 38204 22725
rect 38760 22691 38776 22725
rect 24722 22632 24756 22648
rect 24722 22040 24756 22056
rect 25740 22632 25774 22648
rect 25740 22040 25774 22056
rect 26758 22632 26792 22648
rect 26758 22040 26792 22056
rect 27776 22632 27810 22648
rect 27776 22040 27810 22056
rect 28794 22632 28828 22648
rect 28794 22040 28828 22056
rect 29812 22632 29846 22648
rect 29812 22040 29846 22056
rect 30830 22632 30864 22648
rect 30830 22040 30864 22056
rect 31848 22632 31882 22648
rect 31848 22040 31882 22056
rect 32866 22632 32900 22648
rect 32866 22040 32900 22056
rect 33884 22632 33918 22648
rect 33884 22040 33918 22056
rect 34902 22632 34936 22648
rect 34902 22040 34936 22056
rect 35920 22632 35954 22648
rect 35920 22040 35954 22056
rect 36938 22632 36972 22648
rect 36938 22040 36972 22056
rect 37956 22632 37990 22648
rect 37956 22040 37990 22056
rect 38974 22632 39008 22648
rect 38974 22040 39008 22056
rect 24954 21963 24970 21997
rect 25526 21963 25542 21997
rect 25972 21963 25988 21997
rect 26544 21963 26560 21997
rect 26990 21963 27006 21997
rect 27562 21963 27578 21997
rect 28008 21963 28024 21997
rect 28580 21963 28596 21997
rect 29026 21963 29042 21997
rect 29598 21963 29614 21997
rect 30044 21963 30060 21997
rect 30616 21963 30632 21997
rect 31062 21963 31078 21997
rect 31634 21963 31650 21997
rect 32080 21963 32096 21997
rect 32652 21963 32668 21997
rect 33098 21963 33114 21997
rect 33670 21963 33686 21997
rect 34116 21963 34132 21997
rect 34688 21963 34704 21997
rect 35134 21963 35150 21997
rect 35706 21963 35722 21997
rect 36152 21963 36168 21997
rect 36724 21963 36740 21997
rect 37170 21963 37186 21997
rect 37742 21963 37758 21997
rect 38188 21963 38204 21997
rect 38760 21963 38776 21997
rect 24696 21842 24786 21872
rect 24696 21808 24724 21842
rect 24758 21808 24786 21842
rect 24696 21780 24786 21808
rect 25714 21842 25804 21872
rect 25714 21808 25742 21842
rect 25776 21808 25804 21842
rect 25714 21780 25804 21808
rect 26732 21842 26822 21872
rect 26732 21808 26760 21842
rect 26794 21808 26822 21842
rect 26732 21780 26822 21808
rect 27750 21842 27840 21872
rect 27750 21808 27778 21842
rect 27812 21808 27840 21842
rect 27750 21780 27840 21808
rect 28768 21842 28858 21872
rect 28768 21808 28796 21842
rect 28830 21808 28858 21842
rect 28768 21780 28858 21808
rect 29786 21842 29876 21872
rect 29786 21808 29814 21842
rect 29848 21808 29876 21842
rect 29786 21780 29876 21808
rect 30804 21842 30894 21872
rect 30804 21808 30832 21842
rect 30866 21808 30894 21842
rect 30804 21780 30894 21808
rect 31822 21842 31912 21872
rect 31822 21808 31850 21842
rect 31884 21808 31912 21842
rect 31822 21780 31912 21808
rect 32840 21842 32930 21872
rect 32840 21808 32868 21842
rect 32902 21808 32930 21842
rect 32840 21780 32930 21808
rect 33858 21842 33948 21872
rect 33858 21808 33886 21842
rect 33920 21808 33948 21842
rect 33858 21780 33948 21808
rect 34876 21842 34966 21872
rect 34876 21808 34904 21842
rect 34938 21808 34966 21842
rect 34876 21780 34966 21808
rect 35894 21842 35984 21872
rect 35894 21808 35922 21842
rect 35956 21808 35984 21842
rect 35894 21780 35984 21808
rect 36912 21842 37002 21872
rect 36912 21808 36940 21842
rect 36974 21808 37002 21842
rect 36912 21780 37002 21808
rect 37930 21842 38020 21872
rect 37930 21808 37958 21842
rect 37992 21808 38020 21842
rect 37930 21780 38020 21808
rect 38948 21842 39038 21872
rect 38948 21808 38976 21842
rect 39010 21808 39038 21842
rect 38948 21780 39038 21808
rect 24954 21659 24970 21693
rect 25526 21659 25542 21693
rect 25972 21659 25988 21693
rect 26544 21659 26560 21693
rect 26990 21659 27006 21693
rect 27562 21659 27578 21693
rect 28008 21659 28024 21693
rect 28580 21659 28596 21693
rect 29026 21659 29042 21693
rect 29598 21659 29614 21693
rect 30044 21659 30060 21693
rect 30616 21659 30632 21693
rect 31062 21659 31078 21693
rect 31634 21659 31650 21693
rect 32080 21659 32096 21693
rect 32652 21659 32668 21693
rect 33098 21659 33114 21693
rect 33670 21659 33686 21693
rect 34116 21659 34132 21693
rect 34688 21659 34704 21693
rect 35134 21659 35150 21693
rect 35706 21659 35722 21693
rect 36152 21659 36168 21693
rect 36724 21659 36740 21693
rect 37170 21659 37186 21693
rect 37742 21659 37758 21693
rect 38188 21659 38204 21693
rect 38760 21659 38776 21693
rect 24722 21600 24756 21616
rect 24722 21008 24756 21024
rect 25740 21600 25774 21616
rect 25740 21008 25774 21024
rect 26758 21600 26792 21616
rect 26758 21008 26792 21024
rect 27776 21600 27810 21616
rect 27776 21008 27810 21024
rect 28794 21600 28828 21616
rect 28794 21008 28828 21024
rect 29812 21600 29846 21616
rect 29812 21008 29846 21024
rect 30830 21600 30864 21616
rect 30830 21008 30864 21024
rect 31848 21600 31882 21616
rect 31848 21008 31882 21024
rect 32866 21600 32900 21616
rect 32866 21008 32900 21024
rect 33884 21600 33918 21616
rect 33884 21008 33918 21024
rect 34902 21600 34936 21616
rect 34902 21008 34936 21024
rect 35920 21600 35954 21616
rect 35920 21008 35954 21024
rect 36938 21600 36972 21616
rect 36938 21008 36972 21024
rect 37956 21600 37990 21616
rect 37956 21008 37990 21024
rect 38974 21600 39008 21616
rect 38974 21008 39008 21024
rect 24954 20931 24970 20965
rect 25526 20931 25542 20965
rect 25972 20931 25988 20965
rect 26544 20931 26560 20965
rect 26990 20931 27006 20965
rect 27562 20931 27578 20965
rect 28008 20931 28024 20965
rect 28580 20931 28596 20965
rect 29026 20931 29042 20965
rect 29598 20931 29614 20965
rect 30044 20931 30060 20965
rect 30616 20931 30632 20965
rect 31062 20931 31078 20965
rect 31634 20931 31650 20965
rect 32080 20931 32096 20965
rect 32652 20931 32668 20965
rect 33098 20931 33114 20965
rect 33670 20931 33686 20965
rect 34116 20931 34132 20965
rect 34688 20931 34704 20965
rect 35134 20931 35150 20965
rect 35706 20931 35722 20965
rect 36152 20931 36168 20965
rect 36724 20931 36740 20965
rect 37170 20931 37186 20965
rect 37742 20931 37758 20965
rect 38188 20931 38204 20965
rect 38760 20931 38776 20965
rect 24302 20564 24392 20594
rect 24302 20530 24330 20564
rect 24364 20530 24392 20564
rect 24302 20502 24392 20530
rect 25320 20564 25410 20594
rect 25320 20530 25348 20564
rect 25382 20530 25410 20564
rect 25320 20502 25410 20530
rect 26338 20564 26428 20594
rect 26338 20530 26366 20564
rect 26400 20530 26428 20564
rect 26338 20502 26428 20530
rect 27356 20564 27446 20594
rect 27356 20530 27384 20564
rect 27418 20530 27446 20564
rect 27356 20502 27446 20530
rect 28374 20564 28464 20594
rect 28374 20530 28402 20564
rect 28436 20530 28464 20564
rect 28374 20502 28464 20530
rect 29392 20564 29482 20594
rect 29392 20530 29420 20564
rect 29454 20530 29482 20564
rect 29392 20502 29482 20530
rect 30410 20564 30500 20594
rect 30410 20530 30438 20564
rect 30472 20530 30500 20564
rect 30410 20502 30500 20530
rect 31428 20564 31518 20594
rect 31428 20530 31456 20564
rect 31490 20530 31518 20564
rect 31428 20502 31518 20530
rect 32446 20564 32536 20594
rect 32446 20530 32474 20564
rect 32508 20530 32536 20564
rect 32446 20502 32536 20530
rect 33464 20564 33554 20594
rect 33464 20530 33492 20564
rect 33526 20530 33554 20564
rect 33464 20502 33554 20530
rect 34482 20564 34572 20594
rect 34482 20530 34510 20564
rect 34544 20530 34572 20564
rect 34482 20502 34572 20530
rect 35500 20564 35590 20594
rect 35500 20530 35528 20564
rect 35562 20530 35590 20564
rect 35500 20502 35590 20530
rect 36518 20564 36608 20594
rect 36518 20530 36546 20564
rect 36580 20530 36608 20564
rect 36518 20502 36608 20530
rect 37536 20564 37626 20594
rect 37536 20530 37564 20564
rect 37598 20530 37626 20564
rect 37536 20502 37626 20530
rect 38554 20564 38644 20594
rect 38554 20530 38582 20564
rect 38616 20530 38644 20564
rect 38554 20502 38644 20530
rect 39572 20564 39662 20594
rect 39572 20530 39600 20564
rect 39634 20530 39662 20564
rect 39572 20502 39662 20530
rect 19704 20254 19794 20284
rect 19704 20220 19732 20254
rect 19766 20220 19794 20254
rect 19704 20192 19794 20220
rect 20722 20254 20812 20284
rect 20722 20220 20750 20254
rect 20784 20220 20812 20254
rect 20722 20192 20812 20220
rect 21740 20254 21830 20284
rect 21740 20220 21768 20254
rect 21802 20220 21830 20254
rect 21740 20192 21830 20220
rect 22758 20254 22848 20284
rect 22758 20220 22786 20254
rect 22820 20220 22848 20254
rect 22758 20192 22848 20220
rect 24746 20055 24762 20089
rect 25318 20055 25334 20089
rect 25764 20055 25780 20089
rect 26336 20055 26352 20089
rect 26782 20055 26798 20089
rect 27354 20055 27370 20089
rect 27800 20055 27816 20089
rect 28372 20055 28388 20089
rect 28818 20055 28834 20089
rect 29390 20055 29406 20089
rect 29836 20055 29852 20089
rect 30408 20055 30424 20089
rect 30854 20055 30870 20089
rect 31426 20055 31442 20089
rect 31872 20055 31888 20089
rect 32444 20055 32460 20089
rect 32890 20055 32906 20089
rect 33462 20055 33478 20089
rect 33908 20055 33924 20089
rect 34480 20055 34496 20089
rect 34926 20055 34942 20089
rect 35498 20055 35514 20089
rect 35944 20055 35960 20089
rect 36516 20055 36532 20089
rect 36962 20055 36978 20089
rect 37534 20055 37550 20089
rect 37980 20055 37996 20089
rect 38552 20055 38568 20089
rect 38998 20055 39014 20089
rect 39570 20055 39586 20089
rect 24514 19996 24548 20012
rect 19442 19951 19458 19985
rect 20014 19951 20030 19985
rect 20460 19951 20476 19985
rect 21032 19951 21048 19985
rect 21478 19951 21494 19985
rect 22050 19951 22066 19985
rect 22496 19951 22512 19985
rect 23068 19951 23084 19985
rect 19210 19892 19244 19908
rect 19210 19300 19244 19316
rect 20228 19892 20262 19908
rect 20228 19300 20262 19316
rect 21246 19892 21280 19908
rect 21246 19300 21280 19316
rect 22264 19892 22298 19908
rect 22264 19300 22298 19316
rect 23282 19892 23316 19908
rect 24514 19404 24548 19420
rect 25532 19996 25566 20012
rect 25532 19404 25566 19420
rect 26550 19996 26584 20012
rect 26550 19404 26584 19420
rect 27568 19996 27602 20012
rect 27568 19404 27602 19420
rect 28586 19996 28620 20012
rect 28586 19404 28620 19420
rect 29604 19996 29638 20012
rect 29604 19404 29638 19420
rect 30622 19996 30656 20012
rect 30622 19404 30656 19420
rect 31640 19996 31674 20012
rect 31640 19404 31674 19420
rect 32658 19996 32692 20012
rect 32658 19404 32692 19420
rect 33676 19996 33710 20012
rect 33676 19404 33710 19420
rect 34694 19996 34728 20012
rect 34694 19404 34728 19420
rect 35712 19996 35746 20012
rect 35712 19404 35746 19420
rect 36730 19996 36764 20012
rect 36730 19404 36764 19420
rect 37748 19996 37782 20012
rect 37748 19404 37782 19420
rect 38766 19996 38800 20012
rect 38766 19404 38800 19420
rect 39784 19996 39818 20012
rect 39784 19404 39818 19420
rect 24746 19327 24762 19361
rect 25318 19327 25334 19361
rect 25764 19327 25780 19361
rect 26336 19327 26352 19361
rect 26782 19327 26798 19361
rect 27354 19327 27370 19361
rect 27800 19327 27816 19361
rect 28372 19327 28388 19361
rect 28818 19327 28834 19361
rect 29390 19327 29406 19361
rect 29836 19327 29852 19361
rect 30408 19327 30424 19361
rect 30854 19327 30870 19361
rect 31426 19327 31442 19361
rect 31872 19327 31888 19361
rect 32444 19327 32460 19361
rect 32890 19327 32906 19361
rect 33462 19327 33478 19361
rect 33908 19327 33924 19361
rect 34480 19327 34496 19361
rect 34926 19327 34942 19361
rect 35498 19327 35514 19361
rect 35944 19327 35960 19361
rect 36516 19327 36532 19361
rect 36962 19327 36978 19361
rect 37534 19327 37550 19361
rect 37980 19327 37996 19361
rect 38552 19327 38568 19361
rect 38998 19327 39014 19361
rect 39570 19327 39586 19361
rect 23282 19300 23316 19316
rect 19442 19223 19458 19257
rect 20014 19223 20030 19257
rect 20460 19223 20476 19257
rect 21032 19223 21048 19257
rect 21478 19223 21494 19257
rect 22050 19223 22066 19257
rect 22496 19223 22512 19257
rect 23068 19223 23084 19257
rect 19180 19100 19270 19130
rect 19180 19066 19208 19100
rect 19242 19066 19270 19100
rect 19180 19038 19270 19066
rect 20198 19100 20288 19130
rect 20198 19066 20226 19100
rect 20260 19066 20288 19100
rect 20198 19038 20288 19066
rect 21216 19100 21306 19130
rect 21216 19066 21244 19100
rect 21278 19066 21306 19100
rect 21216 19038 21306 19066
rect 22234 19100 22324 19130
rect 22234 19066 22262 19100
rect 22296 19066 22324 19100
rect 22234 19038 22324 19066
rect 24392 19116 24482 19146
rect 24392 19082 24420 19116
rect 24454 19082 24482 19116
rect 24392 19054 24482 19082
rect 25410 19116 25500 19146
rect 25410 19082 25438 19116
rect 25472 19082 25500 19116
rect 25410 19054 25500 19082
rect 26428 19116 26518 19146
rect 26428 19082 26456 19116
rect 26490 19082 26518 19116
rect 26428 19054 26518 19082
rect 27446 19116 27536 19146
rect 27446 19082 27474 19116
rect 27508 19082 27536 19116
rect 27446 19054 27536 19082
rect 28464 19116 28554 19146
rect 28464 19082 28492 19116
rect 28526 19082 28554 19116
rect 28464 19054 28554 19082
rect 29482 19116 29572 19146
rect 29482 19082 29510 19116
rect 29544 19082 29572 19116
rect 29482 19054 29572 19082
rect 30500 19116 30590 19146
rect 30500 19082 30528 19116
rect 30562 19082 30590 19116
rect 30500 19054 30590 19082
rect 31518 19116 31608 19146
rect 31518 19082 31546 19116
rect 31580 19082 31608 19116
rect 31518 19054 31608 19082
rect 32536 19116 32626 19146
rect 32536 19082 32564 19116
rect 32598 19082 32626 19116
rect 32536 19054 32626 19082
rect 33554 19116 33644 19146
rect 33554 19082 33582 19116
rect 33616 19082 33644 19116
rect 33554 19054 33644 19082
rect 34572 19116 34662 19146
rect 34572 19082 34600 19116
rect 34634 19082 34662 19116
rect 34572 19054 34662 19082
rect 35590 19116 35680 19146
rect 35590 19082 35618 19116
rect 35652 19082 35680 19116
rect 35590 19054 35680 19082
rect 36608 19116 36698 19146
rect 36608 19082 36636 19116
rect 36670 19082 36698 19116
rect 36608 19054 36698 19082
rect 37626 19116 37716 19146
rect 37626 19082 37654 19116
rect 37688 19082 37716 19116
rect 37626 19054 37716 19082
rect 38644 19116 38734 19146
rect 38644 19082 38672 19116
rect 38706 19082 38734 19116
rect 38644 19054 38734 19082
rect 39662 19116 39752 19146
rect 39662 19082 39690 19116
rect 39724 19082 39752 19116
rect 39662 19054 39752 19082
rect 19442 18919 19458 18953
rect 20014 18919 20030 18953
rect 20460 18919 20476 18953
rect 21032 18919 21048 18953
rect 21478 18919 21494 18953
rect 22050 18919 22066 18953
rect 22496 18919 22512 18953
rect 23068 18919 23084 18953
rect 19210 18860 19244 18876
rect 19210 18268 19244 18284
rect 20228 18860 20262 18876
rect 20228 18268 20262 18284
rect 21246 18860 21280 18876
rect 21246 18268 21280 18284
rect 22264 18860 22298 18876
rect 22264 18268 22298 18284
rect 23282 18860 23316 18876
rect 24746 18799 24762 18833
rect 25318 18799 25334 18833
rect 25764 18799 25780 18833
rect 26336 18799 26352 18833
rect 26782 18799 26798 18833
rect 27354 18799 27370 18833
rect 27800 18799 27816 18833
rect 28372 18799 28388 18833
rect 28818 18799 28834 18833
rect 29390 18799 29406 18833
rect 29836 18799 29852 18833
rect 30408 18799 30424 18833
rect 30854 18799 30870 18833
rect 31426 18799 31442 18833
rect 31872 18799 31888 18833
rect 32444 18799 32460 18833
rect 32890 18799 32906 18833
rect 33462 18799 33478 18833
rect 33908 18799 33924 18833
rect 34480 18799 34496 18833
rect 34926 18799 34942 18833
rect 35498 18799 35514 18833
rect 35944 18799 35960 18833
rect 36516 18799 36532 18833
rect 36962 18799 36978 18833
rect 37534 18799 37550 18833
rect 37980 18799 37996 18833
rect 38552 18799 38568 18833
rect 38998 18799 39014 18833
rect 39570 18799 39586 18833
rect 23282 18268 23316 18284
rect 24514 18740 24548 18756
rect 19442 18191 19458 18225
rect 20014 18191 20030 18225
rect 20460 18191 20476 18225
rect 21032 18191 21048 18225
rect 21478 18191 21494 18225
rect 22050 18191 22066 18225
rect 22496 18191 22512 18225
rect 23068 18191 23084 18225
rect 24514 18148 24548 18164
rect 25532 18740 25566 18756
rect 25532 18148 25566 18164
rect 26550 18740 26584 18756
rect 26550 18148 26584 18164
rect 27568 18740 27602 18756
rect 27568 18148 27602 18164
rect 28586 18740 28620 18756
rect 28586 18148 28620 18164
rect 29604 18740 29638 18756
rect 29604 18148 29638 18164
rect 30622 18740 30656 18756
rect 30622 18148 30656 18164
rect 31640 18740 31674 18756
rect 31640 18148 31674 18164
rect 32658 18740 32692 18756
rect 32658 18148 32692 18164
rect 33676 18740 33710 18756
rect 33676 18148 33710 18164
rect 34694 18740 34728 18756
rect 34694 18148 34728 18164
rect 35712 18740 35746 18756
rect 35712 18148 35746 18164
rect 36730 18740 36764 18756
rect 36730 18148 36764 18164
rect 37748 18740 37782 18756
rect 37748 18148 37782 18164
rect 38766 18740 38800 18756
rect 38766 18148 38800 18164
rect 39784 18740 39818 18756
rect 39784 18148 39818 18164
rect 19190 18072 19280 18102
rect 19190 18038 19218 18072
rect 19252 18038 19280 18072
rect 19190 18010 19280 18038
rect 20208 18072 20298 18102
rect 20208 18038 20236 18072
rect 20270 18038 20298 18072
rect 20208 18010 20298 18038
rect 21226 18072 21316 18102
rect 21226 18038 21254 18072
rect 21288 18038 21316 18072
rect 21226 18010 21316 18038
rect 22244 18072 22334 18102
rect 22244 18038 22272 18072
rect 22306 18038 22334 18072
rect 24746 18071 24762 18105
rect 25318 18071 25334 18105
rect 25764 18071 25780 18105
rect 26336 18071 26352 18105
rect 26782 18071 26798 18105
rect 27354 18071 27370 18105
rect 27800 18071 27816 18105
rect 28372 18071 28388 18105
rect 28818 18071 28834 18105
rect 29390 18071 29406 18105
rect 29836 18071 29852 18105
rect 30408 18071 30424 18105
rect 30854 18071 30870 18105
rect 31426 18071 31442 18105
rect 31872 18071 31888 18105
rect 32444 18071 32460 18105
rect 32890 18071 32906 18105
rect 33462 18071 33478 18105
rect 33908 18071 33924 18105
rect 34480 18071 34496 18105
rect 34926 18071 34942 18105
rect 35498 18071 35514 18105
rect 35944 18071 35960 18105
rect 36516 18071 36532 18105
rect 36962 18071 36978 18105
rect 37534 18071 37550 18105
rect 37980 18071 37996 18105
rect 38552 18071 38568 18105
rect 38998 18071 39014 18105
rect 39570 18071 39586 18105
rect 22244 18010 22334 18038
rect 19442 17887 19458 17921
rect 20014 17887 20030 17921
rect 20460 17887 20476 17921
rect 21032 17887 21048 17921
rect 21478 17887 21494 17921
rect 22050 17887 22066 17921
rect 22496 17887 22512 17921
rect 23068 17887 23084 17921
rect 24416 17848 24506 17878
rect 19210 17828 19244 17844
rect 19210 17236 19244 17252
rect 20228 17828 20262 17844
rect 20228 17236 20262 17252
rect 21246 17828 21280 17844
rect 21246 17236 21280 17252
rect 22264 17828 22298 17844
rect 22264 17236 22298 17252
rect 23282 17828 23316 17844
rect 24416 17814 24444 17848
rect 24478 17814 24506 17848
rect 24416 17786 24506 17814
rect 25434 17848 25524 17878
rect 25434 17814 25462 17848
rect 25496 17814 25524 17848
rect 25434 17786 25524 17814
rect 26452 17848 26542 17878
rect 26452 17814 26480 17848
rect 26514 17814 26542 17848
rect 26452 17786 26542 17814
rect 27470 17848 27560 17878
rect 27470 17814 27498 17848
rect 27532 17814 27560 17848
rect 27470 17786 27560 17814
rect 28488 17848 28578 17878
rect 28488 17814 28516 17848
rect 28550 17814 28578 17848
rect 28488 17786 28578 17814
rect 29506 17848 29596 17878
rect 29506 17814 29534 17848
rect 29568 17814 29596 17848
rect 29506 17786 29596 17814
rect 30524 17848 30614 17878
rect 30524 17814 30552 17848
rect 30586 17814 30614 17848
rect 30524 17786 30614 17814
rect 31542 17848 31632 17878
rect 31542 17814 31570 17848
rect 31604 17814 31632 17848
rect 31542 17786 31632 17814
rect 32560 17848 32650 17878
rect 32560 17814 32588 17848
rect 32622 17814 32650 17848
rect 32560 17786 32650 17814
rect 33578 17848 33668 17878
rect 33578 17814 33606 17848
rect 33640 17814 33668 17848
rect 33578 17786 33668 17814
rect 34596 17848 34686 17878
rect 34596 17814 34624 17848
rect 34658 17814 34686 17848
rect 34596 17786 34686 17814
rect 35614 17848 35704 17878
rect 35614 17814 35642 17848
rect 35676 17814 35704 17848
rect 35614 17786 35704 17814
rect 36632 17848 36722 17878
rect 36632 17814 36660 17848
rect 36694 17814 36722 17848
rect 36632 17786 36722 17814
rect 37650 17848 37740 17878
rect 37650 17814 37678 17848
rect 37712 17814 37740 17848
rect 37650 17786 37740 17814
rect 38668 17848 38758 17878
rect 38668 17814 38696 17848
rect 38730 17814 38758 17848
rect 38668 17786 38758 17814
rect 39686 17848 39776 17878
rect 39686 17814 39714 17848
rect 39748 17814 39776 17848
rect 39686 17786 39776 17814
rect 24746 17543 24762 17577
rect 25318 17543 25334 17577
rect 25764 17543 25780 17577
rect 26336 17543 26352 17577
rect 26782 17543 26798 17577
rect 27354 17543 27370 17577
rect 27800 17543 27816 17577
rect 28372 17543 28388 17577
rect 28818 17543 28834 17577
rect 29390 17543 29406 17577
rect 29836 17543 29852 17577
rect 30408 17543 30424 17577
rect 30854 17543 30870 17577
rect 31426 17543 31442 17577
rect 31872 17543 31888 17577
rect 32444 17543 32460 17577
rect 32890 17543 32906 17577
rect 33462 17543 33478 17577
rect 33908 17543 33924 17577
rect 34480 17543 34496 17577
rect 34926 17543 34942 17577
rect 35498 17543 35514 17577
rect 35944 17543 35960 17577
rect 36516 17543 36532 17577
rect 36962 17543 36978 17577
rect 37534 17543 37550 17577
rect 37980 17543 37996 17577
rect 38552 17543 38568 17577
rect 38998 17543 39014 17577
rect 39570 17543 39586 17577
rect 23282 17236 23316 17252
rect 24514 17484 24548 17500
rect 19442 17159 19458 17193
rect 20014 17159 20030 17193
rect 20460 17159 20476 17193
rect 21032 17159 21048 17193
rect 21478 17159 21494 17193
rect 22050 17159 22066 17193
rect 22496 17159 22512 17193
rect 23068 17159 23084 17193
rect 19180 17044 19270 17074
rect 19180 17010 19208 17044
rect 19242 17010 19270 17044
rect 19180 16982 19270 17010
rect 20198 17044 20288 17074
rect 20198 17010 20226 17044
rect 20260 17010 20288 17044
rect 20198 16982 20288 17010
rect 21216 17044 21306 17074
rect 21216 17010 21244 17044
rect 21278 17010 21306 17044
rect 21216 16982 21306 17010
rect 22234 17044 22324 17074
rect 22234 17010 22262 17044
rect 22296 17010 22324 17044
rect 22234 16982 22324 17010
rect 24514 16892 24548 16908
rect 25532 17484 25566 17500
rect 25532 16892 25566 16908
rect 26550 17484 26584 17500
rect 26550 16892 26584 16908
rect 27568 17484 27602 17500
rect 27568 16892 27602 16908
rect 28586 17484 28620 17500
rect 28586 16892 28620 16908
rect 29604 17484 29638 17500
rect 29604 16892 29638 16908
rect 30622 17484 30656 17500
rect 30622 16892 30656 16908
rect 31640 17484 31674 17500
rect 31640 16892 31674 16908
rect 32658 17484 32692 17500
rect 32658 16892 32692 16908
rect 33676 17484 33710 17500
rect 33676 16892 33710 16908
rect 34694 17484 34728 17500
rect 34694 16892 34728 16908
rect 35712 17484 35746 17500
rect 35712 16892 35746 16908
rect 36730 17484 36764 17500
rect 36730 16892 36764 16908
rect 37748 17484 37782 17500
rect 37748 16892 37782 16908
rect 38766 17484 38800 17500
rect 38766 16892 38800 16908
rect 39784 17484 39818 17500
rect 39784 16892 39818 16908
rect 19442 16855 19458 16889
rect 20014 16855 20030 16889
rect 20460 16855 20476 16889
rect 21032 16855 21048 16889
rect 21478 16855 21494 16889
rect 22050 16855 22066 16889
rect 22496 16855 22512 16889
rect 23068 16855 23084 16889
rect 24746 16815 24762 16849
rect 25318 16815 25334 16849
rect 25764 16815 25780 16849
rect 26336 16815 26352 16849
rect 26782 16815 26798 16849
rect 27354 16815 27370 16849
rect 27800 16815 27816 16849
rect 28372 16815 28388 16849
rect 28818 16815 28834 16849
rect 29390 16815 29406 16849
rect 29836 16815 29852 16849
rect 30408 16815 30424 16849
rect 30854 16815 30870 16849
rect 31426 16815 31442 16849
rect 31872 16815 31888 16849
rect 32444 16815 32460 16849
rect 32890 16815 32906 16849
rect 33462 16815 33478 16849
rect 33908 16815 33924 16849
rect 34480 16815 34496 16849
rect 34926 16815 34942 16849
rect 35498 16815 35514 16849
rect 35944 16815 35960 16849
rect 36516 16815 36532 16849
rect 36962 16815 36978 16849
rect 37534 16815 37550 16849
rect 37980 16815 37996 16849
rect 38552 16815 38568 16849
rect 38998 16815 39014 16849
rect 39570 16815 39586 16849
rect 19210 16796 19244 16812
rect 19210 16204 19244 16220
rect 20228 16796 20262 16812
rect 20228 16204 20262 16220
rect 21246 16796 21280 16812
rect 21246 16204 21280 16220
rect 22264 16796 22298 16812
rect 22264 16204 22298 16220
rect 23282 16796 23316 16812
rect 24280 16604 24370 16634
rect 24280 16570 24308 16604
rect 24342 16570 24370 16604
rect 24280 16542 24370 16570
rect 25298 16604 25388 16634
rect 25298 16570 25326 16604
rect 25360 16570 25388 16604
rect 25298 16542 25388 16570
rect 26316 16604 26406 16634
rect 26316 16570 26344 16604
rect 26378 16570 26406 16604
rect 26316 16542 26406 16570
rect 27334 16604 27424 16634
rect 27334 16570 27362 16604
rect 27396 16570 27424 16604
rect 27334 16542 27424 16570
rect 28352 16604 28442 16634
rect 28352 16570 28380 16604
rect 28414 16570 28442 16604
rect 28352 16542 28442 16570
rect 29370 16604 29460 16634
rect 29370 16570 29398 16604
rect 29432 16570 29460 16604
rect 29370 16542 29460 16570
rect 30388 16604 30478 16634
rect 30388 16570 30416 16604
rect 30450 16570 30478 16604
rect 30388 16542 30478 16570
rect 31406 16604 31496 16634
rect 31406 16570 31434 16604
rect 31468 16570 31496 16604
rect 31406 16542 31496 16570
rect 32424 16604 32514 16634
rect 32424 16570 32452 16604
rect 32486 16570 32514 16604
rect 32424 16542 32514 16570
rect 33442 16604 33532 16634
rect 33442 16570 33470 16604
rect 33504 16570 33532 16604
rect 33442 16542 33532 16570
rect 34460 16604 34550 16634
rect 34460 16570 34488 16604
rect 34522 16570 34550 16604
rect 34460 16542 34550 16570
rect 35478 16604 35568 16634
rect 35478 16570 35506 16604
rect 35540 16570 35568 16604
rect 35478 16542 35568 16570
rect 36496 16604 36586 16634
rect 36496 16570 36524 16604
rect 36558 16570 36586 16604
rect 36496 16542 36586 16570
rect 37514 16604 37604 16634
rect 37514 16570 37542 16604
rect 37576 16570 37604 16604
rect 37514 16542 37604 16570
rect 38532 16604 38622 16634
rect 38532 16570 38560 16604
rect 38594 16570 38622 16604
rect 38532 16542 38622 16570
rect 39550 16604 39640 16634
rect 39550 16570 39578 16604
rect 39612 16570 39640 16604
rect 39550 16542 39640 16570
rect 24746 16287 24762 16321
rect 25318 16287 25334 16321
rect 25764 16287 25780 16321
rect 26336 16287 26352 16321
rect 26782 16287 26798 16321
rect 27354 16287 27370 16321
rect 27800 16287 27816 16321
rect 28372 16287 28388 16321
rect 28818 16287 28834 16321
rect 29390 16287 29406 16321
rect 29836 16287 29852 16321
rect 30408 16287 30424 16321
rect 30854 16287 30870 16321
rect 31426 16287 31442 16321
rect 31872 16287 31888 16321
rect 32444 16287 32460 16321
rect 32890 16287 32906 16321
rect 33462 16287 33478 16321
rect 33908 16287 33924 16321
rect 34480 16287 34496 16321
rect 34926 16287 34942 16321
rect 35498 16287 35514 16321
rect 35944 16287 35960 16321
rect 36516 16287 36532 16321
rect 36962 16287 36978 16321
rect 37534 16287 37550 16321
rect 37980 16287 37996 16321
rect 38552 16287 38568 16321
rect 38998 16287 39014 16321
rect 39570 16287 39586 16321
rect 23282 16204 23316 16220
rect 24514 16228 24548 16244
rect 19442 16127 19458 16161
rect 20014 16127 20030 16161
rect 20460 16127 20476 16161
rect 21032 16127 21048 16161
rect 21478 16127 21494 16161
rect 22050 16127 22066 16161
rect 22496 16127 22512 16161
rect 23068 16127 23084 16161
rect 19704 15892 19794 15922
rect 19704 15858 19732 15892
rect 19766 15858 19794 15892
rect 19704 15830 19794 15858
rect 20722 15892 20812 15922
rect 20722 15858 20750 15892
rect 20784 15858 20812 15892
rect 20722 15830 20812 15858
rect 21740 15892 21830 15922
rect 21740 15858 21768 15892
rect 21802 15858 21830 15892
rect 21740 15830 21830 15858
rect 22758 15892 22848 15922
rect 22758 15858 22786 15892
rect 22820 15858 22848 15892
rect 22758 15830 22848 15858
rect 24514 15636 24548 15652
rect 25532 16228 25566 16244
rect 25532 15636 25566 15652
rect 26550 16228 26584 16244
rect 26550 15636 26584 15652
rect 27568 16228 27602 16244
rect 27568 15636 27602 15652
rect 28586 16228 28620 16244
rect 28586 15636 28620 15652
rect 29604 16228 29638 16244
rect 29604 15636 29638 15652
rect 30622 16228 30656 16244
rect 30622 15636 30656 15652
rect 31640 16228 31674 16244
rect 31640 15636 31674 15652
rect 32658 16228 32692 16244
rect 32658 15636 32692 15652
rect 33676 16228 33710 16244
rect 33676 15636 33710 15652
rect 34694 16228 34728 16244
rect 34694 15636 34728 15652
rect 35712 16228 35746 16244
rect 35712 15636 35746 15652
rect 36730 16228 36764 16244
rect 36730 15636 36764 15652
rect 37748 16228 37782 16244
rect 37748 15636 37782 15652
rect 38766 16228 38800 16244
rect 38766 15636 38800 15652
rect 39784 16228 39818 16244
rect 39784 15636 39818 15652
rect 24746 15559 24762 15593
rect 25318 15559 25334 15593
rect 25764 15559 25780 15593
rect 26336 15559 26352 15593
rect 26782 15559 26798 15593
rect 27354 15559 27370 15593
rect 27800 15559 27816 15593
rect 28372 15559 28388 15593
rect 28818 15559 28834 15593
rect 29390 15559 29406 15593
rect 29836 15559 29852 15593
rect 30408 15559 30424 15593
rect 30854 15559 30870 15593
rect 31426 15559 31442 15593
rect 31872 15559 31888 15593
rect 32444 15559 32460 15593
rect 32890 15559 32906 15593
rect 33462 15559 33478 15593
rect 33908 15559 33924 15593
rect 34480 15559 34496 15593
rect 34926 15559 34942 15593
rect 35498 15559 35514 15593
rect 35944 15559 35960 15593
rect 36516 15559 36532 15593
rect 36962 15559 36978 15593
rect 37534 15559 37550 15593
rect 37980 15559 37996 15593
rect 38552 15559 38568 15593
rect 38998 15559 39014 15593
rect 39570 15559 39586 15593
rect 17418 14732 17518 14894
rect 41762 14732 41862 14894
rect 4718 13740 4818 13902
rect 41862 13740 41962 13902
rect 20126 13296 20208 13320
rect 20126 13262 20150 13296
rect 20184 13262 20208 13296
rect 20126 13238 20208 13262
rect 21144 13296 21226 13320
rect 21144 13262 21168 13296
rect 21202 13262 21226 13296
rect 21144 13238 21226 13262
rect 22162 13296 22244 13320
rect 22162 13262 22186 13296
rect 22220 13262 22244 13296
rect 22162 13238 22244 13262
rect 23180 13296 23262 13320
rect 23180 13262 23204 13296
rect 23238 13262 23262 13296
rect 23180 13238 23262 13262
rect 24198 13296 24280 13320
rect 24198 13262 24222 13296
rect 24256 13262 24280 13296
rect 24198 13238 24280 13262
rect 25216 13296 25298 13320
rect 25216 13262 25240 13296
rect 25274 13262 25298 13296
rect 25216 13238 25298 13262
rect 26234 13296 26316 13320
rect 26234 13262 26258 13296
rect 26292 13262 26316 13296
rect 26234 13238 26316 13262
rect 27252 13296 27334 13320
rect 27252 13262 27276 13296
rect 27310 13262 27334 13296
rect 27252 13238 27334 13262
rect 28270 13296 28352 13320
rect 28270 13262 28294 13296
rect 28328 13262 28352 13296
rect 28270 13238 28352 13262
rect 29288 13296 29370 13320
rect 29288 13262 29312 13296
rect 29346 13262 29370 13296
rect 29288 13238 29370 13262
rect 30306 13296 30388 13320
rect 30306 13262 30330 13296
rect 30364 13262 30388 13296
rect 30306 13238 30388 13262
rect 31324 13296 31406 13320
rect 31324 13262 31348 13296
rect 31382 13262 31406 13296
rect 31324 13238 31406 13262
rect 32342 13296 32424 13320
rect 32342 13262 32366 13296
rect 32400 13262 32424 13296
rect 32342 13238 32424 13262
rect 33360 13296 33442 13320
rect 33360 13262 33384 13296
rect 33418 13262 33442 13296
rect 33360 13238 33442 13262
rect 34378 13296 34460 13320
rect 34378 13262 34402 13296
rect 34436 13262 34460 13296
rect 34378 13238 34460 13262
rect 35396 13296 35478 13320
rect 35396 13262 35420 13296
rect 35454 13262 35478 13296
rect 35396 13238 35478 13262
rect 36414 13296 36496 13320
rect 36414 13262 36438 13296
rect 36472 13262 36496 13296
rect 36414 13238 36496 13262
rect 37432 13296 37514 13320
rect 37432 13262 37456 13296
rect 37490 13262 37514 13296
rect 37432 13238 37514 13262
rect 38450 13296 38532 13320
rect 38450 13262 38474 13296
rect 38508 13262 38532 13296
rect 38450 13238 38532 13262
rect 39468 13296 39550 13320
rect 39468 13262 39492 13296
rect 39526 13262 39550 13296
rect 39468 13238 39550 13262
rect 19854 13082 19870 13116
rect 20426 13082 20442 13116
rect 20872 13082 20888 13116
rect 21444 13082 21460 13116
rect 21890 13082 21906 13116
rect 22462 13082 22478 13116
rect 22908 13082 22924 13116
rect 23480 13082 23496 13116
rect 23926 13082 23942 13116
rect 24498 13082 24514 13116
rect 24944 13082 24960 13116
rect 25516 13082 25532 13116
rect 25962 13082 25978 13116
rect 26534 13082 26550 13116
rect 26980 13082 26996 13116
rect 27552 13082 27568 13116
rect 27998 13082 28014 13116
rect 28570 13082 28586 13116
rect 29016 13082 29032 13116
rect 29588 13082 29604 13116
rect 30034 13082 30050 13116
rect 30606 13082 30622 13116
rect 31052 13082 31068 13116
rect 31624 13082 31640 13116
rect 32070 13082 32086 13116
rect 32642 13082 32658 13116
rect 33088 13082 33104 13116
rect 33660 13082 33676 13116
rect 34106 13082 34122 13116
rect 34678 13082 34694 13116
rect 35124 13082 35140 13116
rect 35696 13082 35712 13116
rect 36142 13082 36158 13116
rect 36714 13082 36730 13116
rect 37160 13082 37176 13116
rect 37732 13082 37748 13116
rect 38178 13082 38194 13116
rect 38750 13082 38766 13116
rect 39196 13082 39212 13116
rect 39768 13082 39784 13116
rect -202 780 -102 942
rect 4302 780 4402 942
rect 366 480 382 514
rect 482 480 498 514
rect 624 480 640 514
rect 740 480 756 514
rect 882 480 898 514
rect 998 480 1014 514
rect 1140 480 1156 514
rect 1256 480 1272 514
rect 1398 480 1414 514
rect 1514 480 1530 514
rect 1656 480 1672 514
rect 1772 480 1788 514
rect 1914 480 1930 514
rect 2030 480 2046 514
rect 2172 480 2188 514
rect 2288 480 2304 514
rect 2430 480 2446 514
rect 2546 480 2562 514
rect 2688 480 2704 514
rect 2804 480 2820 514
rect 2946 480 2962 514
rect 3062 480 3078 514
rect 3204 480 3220 514
rect 3320 480 3336 514
rect 3462 480 3478 514
rect 3578 480 3594 514
rect 3720 480 3736 514
rect 3836 480 3852 514
rect 286 430 320 446
rect 286 38 320 54
rect 544 430 578 446
rect 544 38 578 54
rect 802 430 836 446
rect 802 38 836 54
rect 1060 430 1094 446
rect 1060 38 1094 54
rect 1318 430 1352 446
rect 1318 38 1352 54
rect 1576 430 1610 446
rect 1576 38 1610 54
rect 1834 430 1868 446
rect 1834 38 1868 54
rect 2092 430 2126 446
rect 2092 38 2126 54
rect 2350 430 2384 446
rect 2350 38 2384 54
rect 2608 430 2642 446
rect 2608 38 2642 54
rect 2866 430 2900 446
rect 2866 38 2900 54
rect 3124 430 3158 446
rect 3124 38 3158 54
rect 3382 430 3416 446
rect 3382 38 3416 54
rect 3640 430 3674 446
rect 3640 38 3674 54
rect 3898 430 3932 446
rect 3898 38 3932 54
rect 366 -30 382 4
rect 482 -30 498 4
rect 624 -30 640 4
rect 740 -30 756 4
rect 882 -30 898 4
rect 998 -30 1014 4
rect 1140 -30 1156 4
rect 1256 -30 1272 4
rect 1398 -30 1414 4
rect 1514 -30 1530 4
rect 1656 -30 1672 4
rect 1772 -30 1788 4
rect 1914 -30 1930 4
rect 2030 -30 2046 4
rect 2172 -30 2188 4
rect 2288 -30 2304 4
rect 2430 -30 2446 4
rect 2546 -30 2562 4
rect 2688 -30 2704 4
rect 2804 -30 2820 4
rect 2946 -30 2962 4
rect 3062 -30 3078 4
rect 3204 -30 3220 4
rect 3320 -30 3336 4
rect 3462 -30 3478 4
rect 3578 -30 3594 4
rect 3720 -30 3736 4
rect 3836 -30 3852 4
rect 366 -520 382 -486
rect 482 -520 498 -486
rect 624 -520 640 -486
rect 740 -520 756 -486
rect 882 -520 898 -486
rect 998 -520 1014 -486
rect 1140 -520 1156 -486
rect 1256 -520 1272 -486
rect 1398 -520 1414 -486
rect 1514 -520 1530 -486
rect 1656 -520 1672 -486
rect 1772 -520 1788 -486
rect 1914 -520 1930 -486
rect 2030 -520 2046 -486
rect 2172 -520 2188 -486
rect 2288 -520 2304 -486
rect 2430 -520 2446 -486
rect 2546 -520 2562 -486
rect 2688 -520 2704 -486
rect 2804 -520 2820 -486
rect 2946 -520 2962 -486
rect 3062 -520 3078 -486
rect 3204 -520 3220 -486
rect 3320 -520 3336 -486
rect 3462 -520 3478 -486
rect 3578 -520 3594 -486
rect 3720 -520 3736 -486
rect 3836 -520 3852 -486
rect 286 -570 320 -554
rect 286 -962 320 -946
rect 544 -570 578 -554
rect 544 -962 578 -946
rect 802 -570 836 -554
rect 802 -962 836 -946
rect 1060 -570 1094 -554
rect 1060 -962 1094 -946
rect 1318 -570 1352 -554
rect 1318 -962 1352 -946
rect 1576 -570 1610 -554
rect 1576 -962 1610 -946
rect 1834 -570 1868 -554
rect 1834 -962 1868 -946
rect 2092 -570 2126 -554
rect 2092 -962 2126 -946
rect 2350 -570 2384 -554
rect 2350 -962 2384 -946
rect 2608 -570 2642 -554
rect 2608 -962 2642 -946
rect 2866 -570 2900 -554
rect 2866 -962 2900 -946
rect 3124 -570 3158 -554
rect 3124 -962 3158 -946
rect 3382 -570 3416 -554
rect 3382 -962 3416 -946
rect 3640 -570 3674 -554
rect 3640 -962 3674 -946
rect 3898 -570 3932 -554
rect 3898 -962 3932 -946
rect 366 -1030 382 -996
rect 482 -1030 498 -996
rect 624 -1030 640 -996
rect 740 -1030 756 -996
rect 882 -1030 898 -996
rect 998 -1030 1014 -996
rect 1140 -1030 1156 -996
rect 1256 -1030 1272 -996
rect 1398 -1030 1414 -996
rect 1514 -1030 1530 -996
rect 1656 -1030 1672 -996
rect 1772 -1030 1788 -996
rect 1914 -1030 1930 -996
rect 2030 -1030 2046 -996
rect 2172 -1030 2188 -996
rect 2288 -1030 2304 -996
rect 2430 -1030 2446 -996
rect 2546 -1030 2562 -996
rect 2688 -1030 2704 -996
rect 2804 -1030 2820 -996
rect 2946 -1030 2962 -996
rect 3062 -1030 3078 -996
rect 3204 -1030 3220 -996
rect 3320 -1030 3336 -996
rect 3462 -1030 3478 -996
rect 3578 -1030 3594 -996
rect 3720 -1030 3736 -996
rect 3836 -1030 3852 -996
rect -202 -2042 -102 -1880
rect 4302 -2042 4402 -1880
rect 19622 13032 19656 13048
rect 7832 12694 7914 12718
rect 7832 12660 7856 12694
rect 7890 12660 7914 12694
rect 7832 12636 7914 12660
rect 8850 12694 8932 12718
rect 8850 12660 8874 12694
rect 8908 12660 8932 12694
rect 8088 12606 8104 12640
rect 8660 12606 8676 12640
rect 8850 12636 8932 12660
rect 9868 12694 9950 12718
rect 9868 12660 9892 12694
rect 9926 12660 9950 12694
rect 9106 12606 9122 12640
rect 9678 12606 9694 12640
rect 9868 12636 9950 12660
rect 10886 12694 10968 12718
rect 10886 12660 10910 12694
rect 10944 12660 10968 12694
rect 10124 12606 10140 12640
rect 10696 12606 10712 12640
rect 10886 12636 10968 12660
rect 11904 12694 11986 12718
rect 11904 12660 11928 12694
rect 11962 12660 11986 12694
rect 11142 12606 11158 12640
rect 11714 12606 11730 12640
rect 11904 12636 11986 12660
rect 12922 12694 13004 12718
rect 12922 12660 12946 12694
rect 12980 12660 13004 12694
rect 12160 12606 12176 12640
rect 12732 12606 12748 12640
rect 12922 12636 13004 12660
rect 13940 12694 14022 12718
rect 13940 12660 13964 12694
rect 13998 12660 14022 12694
rect 13178 12606 13194 12640
rect 13750 12606 13766 12640
rect 13940 12636 14022 12660
rect 14958 12694 15040 12718
rect 14958 12660 14982 12694
rect 15016 12660 15040 12694
rect 14196 12606 14212 12640
rect 14768 12606 14784 12640
rect 14958 12636 15040 12660
rect 15976 12694 16058 12718
rect 15976 12660 16000 12694
rect 16034 12660 16058 12694
rect 15214 12606 15230 12640
rect 15786 12606 15802 12640
rect 15976 12636 16058 12660
rect 17004 12694 17086 12718
rect 17004 12660 17028 12694
rect 17062 12660 17086 12694
rect 16232 12606 16248 12640
rect 16804 12606 16820 12640
rect 17004 12636 17086 12660
rect 7856 12556 7890 12572
rect 7856 11964 7890 11980
rect 8874 12556 8908 12572
rect 8874 11964 8908 11980
rect 9892 12556 9926 12572
rect 9892 11964 9926 11980
rect 10910 12556 10944 12572
rect 10910 11964 10944 11980
rect 11928 12556 11962 12572
rect 11928 11964 11962 11980
rect 12946 12556 12980 12572
rect 12946 11964 12980 11980
rect 13964 12556 13998 12572
rect 13964 11964 13998 11980
rect 14982 12556 15016 12572
rect 14982 11964 15016 11980
rect 16000 12556 16034 12572
rect 16000 11964 16034 11980
rect 17018 12556 17052 12572
rect 19622 12440 19656 12456
rect 20640 13032 20674 13048
rect 20640 12440 20674 12456
rect 21658 13032 21692 13048
rect 21658 12440 21692 12456
rect 22676 13032 22710 13048
rect 22676 12440 22710 12456
rect 23694 13032 23728 13048
rect 23694 12440 23728 12456
rect 24712 13032 24746 13048
rect 24712 12440 24746 12456
rect 25730 13032 25764 13048
rect 25730 12440 25764 12456
rect 26748 13032 26782 13048
rect 26748 12440 26782 12456
rect 27766 13032 27800 13048
rect 27766 12440 27800 12456
rect 28784 13032 28818 13048
rect 28784 12440 28818 12456
rect 29802 13032 29836 13048
rect 29802 12440 29836 12456
rect 30820 13032 30854 13048
rect 30820 12440 30854 12456
rect 31838 13032 31872 13048
rect 31838 12440 31872 12456
rect 32856 13032 32890 13048
rect 32856 12440 32890 12456
rect 33874 13032 33908 13048
rect 33874 12440 33908 12456
rect 34892 13032 34926 13048
rect 34892 12440 34926 12456
rect 35910 13032 35944 13048
rect 35910 12440 35944 12456
rect 36928 13032 36962 13048
rect 36928 12440 36962 12456
rect 37946 13032 37980 13048
rect 37946 12440 37980 12456
rect 38964 13032 38998 13048
rect 38964 12440 38998 12456
rect 39982 13032 40016 13048
rect 39982 12440 40016 12456
rect 19854 12372 19870 12406
rect 20426 12372 20442 12406
rect 20872 12372 20888 12406
rect 21444 12372 21460 12406
rect 21890 12372 21906 12406
rect 22462 12372 22478 12406
rect 22908 12372 22924 12406
rect 23480 12372 23496 12406
rect 23926 12372 23942 12406
rect 24498 12372 24514 12406
rect 24944 12372 24960 12406
rect 25516 12372 25532 12406
rect 25962 12372 25978 12406
rect 26534 12372 26550 12406
rect 26980 12372 26996 12406
rect 27552 12372 27568 12406
rect 27998 12372 28014 12406
rect 28570 12372 28586 12406
rect 29016 12372 29032 12406
rect 29588 12372 29604 12406
rect 30034 12372 30050 12406
rect 30606 12372 30622 12406
rect 31052 12372 31068 12406
rect 31624 12372 31640 12406
rect 32070 12372 32086 12406
rect 32642 12372 32658 12406
rect 33088 12372 33104 12406
rect 33660 12372 33676 12406
rect 34106 12372 34122 12406
rect 34678 12372 34694 12406
rect 35124 12372 35140 12406
rect 35696 12372 35712 12406
rect 36142 12372 36158 12406
rect 36714 12372 36730 12406
rect 37160 12372 37176 12406
rect 37732 12372 37748 12406
rect 38178 12372 38194 12406
rect 38750 12372 38766 12406
rect 39196 12372 39212 12406
rect 39768 12372 39784 12406
rect 19854 12264 19870 12298
rect 20426 12264 20442 12298
rect 20872 12264 20888 12298
rect 21444 12264 21460 12298
rect 21890 12264 21906 12298
rect 22462 12264 22478 12298
rect 22908 12264 22924 12298
rect 23480 12264 23496 12298
rect 23926 12264 23942 12298
rect 24498 12264 24514 12298
rect 24944 12264 24960 12298
rect 25516 12264 25532 12298
rect 25962 12264 25978 12298
rect 26534 12264 26550 12298
rect 26980 12264 26996 12298
rect 27552 12264 27568 12298
rect 27998 12264 28014 12298
rect 28570 12264 28586 12298
rect 29016 12264 29032 12298
rect 29588 12264 29604 12298
rect 30034 12264 30050 12298
rect 30606 12264 30622 12298
rect 31052 12264 31068 12298
rect 31624 12264 31640 12298
rect 32070 12264 32086 12298
rect 32642 12264 32658 12298
rect 33088 12264 33104 12298
rect 33660 12264 33676 12298
rect 34106 12264 34122 12298
rect 34678 12264 34694 12298
rect 35124 12264 35140 12298
rect 35696 12264 35712 12298
rect 36142 12264 36158 12298
rect 36714 12264 36730 12298
rect 37160 12264 37176 12298
rect 37732 12264 37748 12298
rect 38178 12264 38194 12298
rect 38750 12264 38766 12298
rect 39196 12264 39212 12298
rect 39768 12264 39784 12298
rect 17018 11964 17052 11980
rect 19622 12214 19656 12230
rect 7832 11876 7914 11900
rect 8088 11896 8104 11930
rect 8660 11896 8676 11930
rect 7832 11842 7856 11876
rect 7890 11842 7914 11876
rect 7832 11818 7914 11842
rect 8850 11876 8932 11900
rect 9106 11896 9122 11930
rect 9678 11896 9694 11930
rect 8850 11842 8874 11876
rect 8908 11842 8932 11876
rect 8088 11788 8104 11822
rect 8660 11788 8676 11822
rect 8850 11818 8932 11842
rect 9868 11876 9950 11900
rect 10124 11896 10140 11930
rect 10696 11896 10712 11930
rect 9868 11842 9892 11876
rect 9926 11842 9950 11876
rect 9106 11788 9122 11822
rect 9678 11788 9694 11822
rect 9868 11818 9950 11842
rect 10886 11876 10968 11900
rect 11142 11896 11158 11930
rect 11714 11896 11730 11930
rect 10886 11842 10910 11876
rect 10944 11842 10968 11876
rect 10124 11788 10140 11822
rect 10696 11788 10712 11822
rect 10886 11818 10968 11842
rect 11904 11876 11986 11900
rect 12160 11896 12176 11930
rect 12732 11896 12748 11930
rect 11904 11842 11928 11876
rect 11962 11842 11986 11876
rect 11142 11788 11158 11822
rect 11714 11788 11730 11822
rect 11904 11818 11986 11842
rect 12922 11876 13004 11900
rect 13178 11896 13194 11930
rect 13750 11896 13766 11930
rect 12922 11842 12946 11876
rect 12980 11842 13004 11876
rect 12160 11788 12176 11822
rect 12732 11788 12748 11822
rect 12922 11818 13004 11842
rect 13940 11876 14022 11900
rect 14196 11896 14212 11930
rect 14768 11896 14784 11930
rect 13940 11842 13964 11876
rect 13998 11842 14022 11876
rect 13178 11788 13194 11822
rect 13750 11788 13766 11822
rect 13940 11818 14022 11842
rect 14958 11876 15040 11900
rect 15214 11896 15230 11930
rect 15786 11896 15802 11930
rect 14958 11842 14982 11876
rect 15016 11842 15040 11876
rect 14196 11788 14212 11822
rect 14768 11788 14784 11822
rect 14958 11818 15040 11842
rect 15976 11876 16058 11900
rect 16232 11896 16248 11930
rect 16804 11896 16820 11930
rect 15976 11842 16000 11876
rect 16034 11842 16058 11876
rect 15214 11788 15230 11822
rect 15786 11788 15802 11822
rect 15976 11818 16058 11842
rect 17004 11876 17086 11900
rect 17004 11842 17028 11876
rect 17062 11842 17086 11876
rect 16232 11788 16248 11822
rect 16804 11788 16820 11822
rect 17004 11818 17086 11842
rect 13448 11786 13508 11788
rect 7856 11738 7890 11754
rect 7856 11146 7890 11162
rect 8874 11738 8908 11754
rect 8874 11146 8908 11162
rect 9892 11738 9926 11754
rect 9892 11146 9926 11162
rect 10910 11738 10944 11754
rect 10910 11146 10944 11162
rect 11928 11738 11962 11754
rect 11928 11146 11962 11162
rect 12946 11738 12980 11754
rect 12946 11146 12980 11162
rect 13964 11738 13998 11754
rect 13964 11146 13998 11162
rect 14982 11738 15016 11754
rect 14982 11146 15016 11162
rect 16000 11738 16034 11754
rect 16000 11146 16034 11162
rect 17018 11738 17052 11754
rect 19622 11622 19656 11638
rect 20640 12214 20674 12230
rect 20640 11622 20674 11638
rect 21658 12214 21692 12230
rect 21658 11622 21692 11638
rect 22676 12214 22710 12230
rect 22676 11622 22710 11638
rect 23694 12214 23728 12230
rect 23694 11622 23728 11638
rect 24712 12214 24746 12230
rect 24712 11622 24746 11638
rect 25730 12214 25764 12230
rect 25730 11622 25764 11638
rect 26748 12214 26782 12230
rect 26748 11622 26782 11638
rect 27766 12214 27800 12230
rect 27766 11622 27800 11638
rect 28784 12214 28818 12230
rect 28784 11622 28818 11638
rect 29802 12214 29836 12230
rect 29802 11622 29836 11638
rect 30820 12214 30854 12230
rect 30820 11622 30854 11638
rect 31838 12214 31872 12230
rect 31838 11622 31872 11638
rect 32856 12214 32890 12230
rect 32856 11622 32890 11638
rect 33874 12214 33908 12230
rect 33874 11622 33908 11638
rect 34892 12214 34926 12230
rect 34892 11622 34926 11638
rect 35910 12214 35944 12230
rect 35910 11622 35944 11638
rect 36928 12214 36962 12230
rect 36928 11622 36962 11638
rect 37946 12214 37980 12230
rect 37946 11622 37980 11638
rect 38964 12214 38998 12230
rect 38964 11622 38998 11638
rect 39982 12214 40016 12230
rect 39982 11622 40016 11638
rect 19854 11554 19870 11588
rect 20426 11554 20442 11588
rect 20872 11554 20888 11588
rect 21444 11554 21460 11588
rect 21890 11554 21906 11588
rect 22462 11554 22478 11588
rect 22908 11554 22924 11588
rect 23480 11554 23496 11588
rect 23926 11554 23942 11588
rect 24498 11554 24514 11588
rect 24944 11554 24960 11588
rect 25516 11554 25532 11588
rect 25962 11554 25978 11588
rect 26534 11554 26550 11588
rect 26980 11554 26996 11588
rect 27552 11554 27568 11588
rect 27998 11554 28014 11588
rect 28570 11554 28586 11588
rect 29016 11554 29032 11588
rect 29588 11554 29604 11588
rect 30034 11554 30050 11588
rect 30606 11554 30622 11588
rect 31052 11554 31068 11588
rect 31624 11554 31640 11588
rect 32070 11554 32086 11588
rect 32642 11554 32658 11588
rect 33088 11554 33104 11588
rect 33660 11554 33676 11588
rect 34106 11554 34122 11588
rect 34678 11554 34694 11588
rect 35124 11554 35140 11588
rect 35696 11554 35712 11588
rect 36142 11554 36158 11588
rect 36714 11554 36730 11588
rect 37160 11554 37176 11588
rect 37732 11554 37748 11588
rect 38178 11554 38194 11588
rect 38750 11554 38766 11588
rect 39196 11554 39212 11588
rect 39768 11554 39784 11588
rect 20138 11270 20220 11294
rect 20138 11236 20162 11270
rect 20196 11236 20220 11270
rect 20138 11212 20220 11236
rect 21156 11270 21238 11294
rect 21156 11236 21180 11270
rect 21214 11236 21238 11270
rect 21156 11212 21238 11236
rect 22174 11270 22256 11294
rect 22174 11236 22198 11270
rect 22232 11236 22256 11270
rect 22174 11212 22256 11236
rect 23192 11270 23274 11294
rect 23192 11236 23216 11270
rect 23250 11236 23274 11270
rect 23192 11212 23274 11236
rect 24210 11270 24292 11294
rect 24210 11236 24234 11270
rect 24268 11236 24292 11270
rect 24210 11212 24292 11236
rect 25228 11270 25310 11294
rect 25228 11236 25252 11270
rect 25286 11236 25310 11270
rect 25228 11212 25310 11236
rect 26246 11270 26328 11294
rect 26246 11236 26270 11270
rect 26304 11236 26328 11270
rect 26246 11212 26328 11236
rect 27264 11270 27346 11294
rect 27264 11236 27288 11270
rect 27322 11236 27346 11270
rect 27264 11212 27346 11236
rect 28282 11270 28364 11294
rect 28282 11236 28306 11270
rect 28340 11236 28364 11270
rect 28282 11212 28364 11236
rect 29300 11270 29382 11294
rect 29300 11236 29324 11270
rect 29358 11236 29382 11270
rect 29300 11212 29382 11236
rect 30318 11270 30400 11294
rect 30318 11236 30342 11270
rect 30376 11236 30400 11270
rect 30318 11212 30400 11236
rect 31336 11270 31418 11294
rect 31336 11236 31360 11270
rect 31394 11236 31418 11270
rect 31336 11212 31418 11236
rect 32354 11270 32436 11294
rect 32354 11236 32378 11270
rect 32412 11236 32436 11270
rect 32354 11212 32436 11236
rect 33372 11270 33454 11294
rect 33372 11236 33396 11270
rect 33430 11236 33454 11270
rect 33372 11212 33454 11236
rect 34390 11270 34472 11294
rect 34390 11236 34414 11270
rect 34448 11236 34472 11270
rect 34390 11212 34472 11236
rect 35408 11270 35490 11294
rect 35408 11236 35432 11270
rect 35466 11236 35490 11270
rect 35408 11212 35490 11236
rect 36426 11270 36508 11294
rect 36426 11236 36450 11270
rect 36484 11236 36508 11270
rect 36426 11212 36508 11236
rect 37444 11270 37526 11294
rect 37444 11236 37468 11270
rect 37502 11236 37526 11270
rect 37444 11212 37526 11236
rect 38462 11270 38544 11294
rect 38462 11236 38486 11270
rect 38520 11236 38544 11270
rect 38462 11212 38544 11236
rect 39480 11270 39562 11294
rect 39480 11236 39504 11270
rect 39538 11236 39562 11270
rect 39480 11212 39562 11236
rect 17018 11146 17052 11162
rect 9380 11112 9440 11114
rect 10394 11112 10454 11114
rect 14468 11112 14528 11114
rect 15484 11112 15544 11114
rect 7832 11058 7914 11082
rect 8088 11078 8104 11112
rect 8660 11078 8676 11112
rect 7832 11024 7856 11058
rect 7890 11024 7914 11058
rect 7832 11000 7914 11024
rect 8850 11058 8932 11082
rect 9106 11078 9122 11112
rect 9678 11078 9694 11112
rect 8850 11024 8874 11058
rect 8908 11024 8932 11058
rect 8088 10970 8104 11004
rect 8660 10970 8676 11004
rect 8850 11000 8932 11024
rect 9868 11058 9950 11082
rect 10124 11078 10140 11112
rect 10696 11078 10712 11112
rect 9868 11024 9892 11058
rect 9926 11024 9950 11058
rect 9106 10970 9122 11004
rect 9678 10970 9694 11004
rect 9868 11000 9950 11024
rect 10886 11058 10968 11082
rect 11142 11078 11158 11112
rect 11714 11078 11730 11112
rect 10886 11024 10910 11058
rect 10944 11024 10968 11058
rect 10124 10970 10140 11004
rect 10696 10970 10712 11004
rect 10886 11000 10968 11024
rect 11904 11058 11986 11082
rect 12160 11078 12176 11112
rect 12732 11078 12748 11112
rect 11904 11024 11928 11058
rect 11962 11024 11986 11058
rect 11142 10970 11158 11004
rect 11714 10970 11730 11004
rect 11904 11000 11986 11024
rect 12922 11058 13004 11082
rect 13178 11078 13194 11112
rect 13750 11078 13766 11112
rect 12922 11024 12946 11058
rect 12980 11024 13004 11058
rect 12160 10970 12176 11004
rect 12732 10970 12748 11004
rect 12922 11000 13004 11024
rect 13940 11058 14022 11082
rect 14196 11078 14212 11112
rect 14768 11078 14784 11112
rect 13940 11024 13964 11058
rect 13998 11024 14022 11058
rect 13178 10970 13194 11004
rect 13750 10970 13766 11004
rect 13940 11000 14022 11024
rect 14958 11058 15040 11082
rect 15214 11078 15230 11112
rect 15786 11078 15802 11112
rect 14958 11024 14982 11058
rect 15016 11024 15040 11058
rect 14196 10970 14212 11004
rect 14768 10970 14784 11004
rect 14958 11000 15040 11024
rect 15976 11058 16058 11082
rect 16232 11078 16248 11112
rect 16804 11078 16820 11112
rect 15976 11024 16000 11058
rect 16034 11024 16058 11058
rect 15214 10970 15230 11004
rect 15786 10970 15802 11004
rect 15976 11000 16058 11024
rect 17004 11058 17086 11082
rect 17004 11024 17028 11058
rect 17062 11024 17086 11058
rect 16232 10970 16248 11004
rect 16804 10970 16820 11004
rect 17004 11000 17086 11024
rect 7856 10920 7890 10936
rect 7856 10328 7890 10344
rect 8874 10920 8908 10936
rect 8874 10328 8908 10344
rect 9892 10920 9926 10936
rect 9892 10328 9926 10344
rect 10910 10920 10944 10936
rect 10910 10328 10944 10344
rect 11928 10920 11962 10936
rect 11928 10328 11962 10344
rect 12946 10920 12980 10936
rect 12946 10328 12980 10344
rect 13964 10920 13998 10936
rect 13964 10328 13998 10344
rect 14982 10920 15016 10936
rect 14982 10328 15016 10344
rect 16000 10920 16034 10936
rect 16000 10328 16034 10344
rect 17018 10920 17052 10936
rect 19854 10886 19870 10920
rect 20426 10886 20442 10920
rect 20872 10886 20888 10920
rect 21444 10886 21460 10920
rect 21890 10886 21906 10920
rect 22462 10886 22478 10920
rect 22908 10886 22924 10920
rect 23480 10886 23496 10920
rect 23926 10886 23942 10920
rect 24498 10886 24514 10920
rect 24944 10886 24960 10920
rect 25516 10886 25532 10920
rect 25962 10886 25978 10920
rect 26534 10886 26550 10920
rect 26980 10886 26996 10920
rect 27552 10886 27568 10920
rect 27998 10886 28014 10920
rect 28570 10886 28586 10920
rect 29016 10886 29032 10920
rect 29588 10886 29604 10920
rect 30034 10886 30050 10920
rect 30606 10886 30622 10920
rect 31052 10886 31068 10920
rect 31624 10886 31640 10920
rect 32070 10886 32086 10920
rect 32642 10886 32658 10920
rect 33088 10886 33104 10920
rect 33660 10886 33676 10920
rect 34106 10886 34122 10920
rect 34678 10886 34694 10920
rect 35124 10886 35140 10920
rect 35696 10886 35712 10920
rect 36142 10886 36158 10920
rect 36714 10886 36730 10920
rect 37160 10886 37176 10920
rect 37732 10886 37748 10920
rect 38178 10886 38194 10920
rect 38750 10886 38766 10920
rect 39196 10886 39212 10920
rect 39768 10886 39784 10920
rect 29278 10880 29338 10886
rect 17018 10328 17052 10344
rect 19622 10836 19656 10852
rect 9384 10294 9444 10296
rect 10398 10294 10458 10296
rect 14472 10294 14532 10296
rect 15488 10294 15548 10296
rect 7832 10240 7914 10264
rect 8088 10260 8104 10294
rect 8660 10260 8676 10294
rect 7832 10206 7856 10240
rect 7890 10206 7914 10240
rect 7832 10182 7914 10206
rect 8850 10240 8932 10264
rect 9106 10260 9122 10294
rect 9678 10260 9694 10294
rect 8850 10206 8874 10240
rect 8908 10206 8932 10240
rect 8088 10152 8104 10186
rect 8660 10152 8676 10186
rect 8850 10182 8932 10206
rect 9868 10240 9950 10264
rect 10124 10260 10140 10294
rect 10696 10260 10712 10294
rect 9868 10206 9892 10240
rect 9926 10206 9950 10240
rect 9106 10152 9122 10186
rect 9678 10152 9694 10186
rect 9868 10182 9950 10206
rect 10886 10240 10968 10264
rect 11142 10260 11158 10294
rect 11714 10260 11730 10294
rect 10886 10206 10910 10240
rect 10944 10206 10968 10240
rect 10124 10152 10140 10186
rect 10696 10152 10712 10186
rect 10886 10182 10968 10206
rect 11904 10240 11986 10264
rect 12160 10260 12176 10294
rect 12732 10260 12748 10294
rect 11904 10206 11928 10240
rect 11962 10206 11986 10240
rect 11142 10152 11158 10186
rect 11714 10152 11730 10186
rect 11904 10182 11986 10206
rect 12922 10240 13004 10264
rect 13178 10260 13194 10294
rect 13750 10260 13766 10294
rect 12922 10206 12946 10240
rect 12980 10206 13004 10240
rect 12160 10152 12176 10186
rect 12732 10152 12748 10186
rect 12922 10182 13004 10206
rect 13940 10240 14022 10264
rect 14196 10260 14212 10294
rect 14768 10260 14784 10294
rect 13940 10206 13964 10240
rect 13998 10206 14022 10240
rect 13178 10152 13194 10186
rect 13750 10152 13766 10186
rect 13940 10182 14022 10206
rect 14958 10240 15040 10264
rect 15214 10260 15230 10294
rect 15786 10260 15802 10294
rect 14958 10206 14982 10240
rect 15016 10206 15040 10240
rect 14196 10152 14212 10186
rect 14768 10152 14784 10186
rect 14958 10182 15040 10206
rect 15976 10240 16058 10264
rect 16232 10260 16248 10294
rect 16804 10260 16820 10294
rect 15976 10206 16000 10240
rect 16034 10206 16058 10240
rect 15214 10152 15230 10186
rect 15786 10152 15802 10186
rect 15976 10182 16058 10206
rect 17004 10240 17086 10264
rect 19622 10244 19656 10260
rect 20640 10836 20674 10852
rect 20640 10244 20674 10260
rect 21658 10836 21692 10852
rect 21658 10244 21692 10260
rect 22676 10836 22710 10852
rect 22676 10244 22710 10260
rect 23694 10836 23728 10852
rect 23694 10244 23728 10260
rect 24712 10836 24746 10852
rect 24712 10244 24746 10260
rect 25730 10836 25764 10852
rect 25730 10244 25764 10260
rect 26748 10836 26782 10852
rect 26748 10244 26782 10260
rect 27766 10836 27800 10852
rect 27766 10244 27800 10260
rect 28784 10836 28818 10852
rect 28784 10244 28818 10260
rect 29802 10836 29836 10852
rect 29802 10244 29836 10260
rect 30820 10836 30854 10852
rect 30820 10244 30854 10260
rect 31838 10836 31872 10852
rect 31838 10244 31872 10260
rect 32856 10836 32890 10852
rect 32856 10244 32890 10260
rect 33874 10836 33908 10852
rect 33874 10244 33908 10260
rect 34892 10836 34926 10852
rect 34892 10244 34926 10260
rect 35910 10836 35944 10852
rect 35910 10244 35944 10260
rect 36928 10836 36962 10852
rect 36928 10244 36962 10260
rect 37946 10836 37980 10852
rect 37946 10244 37980 10260
rect 38964 10836 38998 10852
rect 38964 10244 38998 10260
rect 39982 10836 40016 10852
rect 39982 10244 40016 10260
rect 17004 10206 17028 10240
rect 17062 10206 17086 10240
rect 25206 10210 25266 10216
rect 27242 10210 27302 10216
rect 28262 10210 28322 10216
rect 33334 10210 33394 10216
rect 16232 10152 16248 10186
rect 16804 10152 16820 10186
rect 17004 10182 17086 10206
rect 19854 10176 19870 10210
rect 20426 10176 20442 10210
rect 20872 10176 20888 10210
rect 21444 10176 21460 10210
rect 21890 10176 21906 10210
rect 22462 10176 22478 10210
rect 22908 10176 22924 10210
rect 23480 10176 23496 10210
rect 23926 10176 23942 10210
rect 24498 10176 24514 10210
rect 24944 10176 24960 10210
rect 25516 10176 25532 10210
rect 25962 10176 25978 10210
rect 26534 10176 26550 10210
rect 26980 10176 26996 10210
rect 27552 10176 27568 10210
rect 27998 10176 28014 10210
rect 28570 10176 28586 10210
rect 29016 10176 29032 10210
rect 29588 10176 29604 10210
rect 30034 10176 30050 10210
rect 30606 10176 30622 10210
rect 31052 10176 31068 10210
rect 31624 10176 31640 10210
rect 32070 10176 32086 10210
rect 32642 10176 32658 10210
rect 33088 10176 33104 10210
rect 33660 10176 33676 10210
rect 34106 10176 34122 10210
rect 34678 10176 34694 10210
rect 35124 10176 35140 10210
rect 35696 10176 35712 10210
rect 36142 10176 36158 10210
rect 36714 10176 36730 10210
rect 37160 10176 37176 10210
rect 37732 10176 37748 10210
rect 38178 10176 38194 10210
rect 38750 10176 38766 10210
rect 39196 10176 39212 10210
rect 39768 10176 39784 10210
rect 7856 10102 7890 10118
rect 7856 9510 7890 9526
rect 8874 10102 8908 10118
rect 8874 9510 8908 9526
rect 9892 10102 9926 10118
rect 9892 9510 9926 9526
rect 10910 10102 10944 10118
rect 10910 9510 10944 9526
rect 11928 10102 11962 10118
rect 11928 9510 11962 9526
rect 12946 10102 12980 10118
rect 12946 9510 12980 9526
rect 13964 10102 13998 10118
rect 13964 9510 13998 9526
rect 14982 10102 15016 10118
rect 14982 9510 15016 9526
rect 16000 10102 16034 10118
rect 16000 9510 16034 9526
rect 17018 10102 17052 10118
rect 20126 9964 20208 9988
rect 20126 9930 20150 9964
rect 20184 9930 20208 9964
rect 20126 9906 20208 9930
rect 21144 9964 21226 9988
rect 21144 9930 21168 9964
rect 21202 9930 21226 9964
rect 21144 9906 21226 9930
rect 22162 9964 22244 9988
rect 22162 9930 22186 9964
rect 22220 9930 22244 9964
rect 22162 9906 22244 9930
rect 23180 9964 23262 9988
rect 23180 9930 23204 9964
rect 23238 9930 23262 9964
rect 23180 9906 23262 9930
rect 24198 9964 24280 9988
rect 24198 9930 24222 9964
rect 24256 9930 24280 9964
rect 24198 9906 24280 9930
rect 25216 9964 25298 9988
rect 25216 9930 25240 9964
rect 25274 9930 25298 9964
rect 25216 9906 25298 9930
rect 26234 9964 26316 9988
rect 26234 9930 26258 9964
rect 26292 9930 26316 9964
rect 26234 9906 26316 9930
rect 27252 9964 27334 9988
rect 27252 9930 27276 9964
rect 27310 9930 27334 9964
rect 27252 9906 27334 9930
rect 28270 9964 28352 9988
rect 28270 9930 28294 9964
rect 28328 9930 28352 9964
rect 28270 9906 28352 9930
rect 29288 9964 29370 9988
rect 29288 9930 29312 9964
rect 29346 9930 29370 9964
rect 29288 9906 29370 9930
rect 30306 9964 30388 9988
rect 30306 9930 30330 9964
rect 30364 9930 30388 9964
rect 30306 9906 30388 9930
rect 31324 9964 31406 9988
rect 31324 9930 31348 9964
rect 31382 9930 31406 9964
rect 31324 9906 31406 9930
rect 32342 9964 32424 9988
rect 32342 9930 32366 9964
rect 32400 9930 32424 9964
rect 32342 9906 32424 9930
rect 33360 9964 33442 9988
rect 33360 9930 33384 9964
rect 33418 9930 33442 9964
rect 33360 9906 33442 9930
rect 34378 9964 34460 9988
rect 34378 9930 34402 9964
rect 34436 9930 34460 9964
rect 34378 9906 34460 9930
rect 35396 9964 35478 9988
rect 35396 9930 35420 9964
rect 35454 9930 35478 9964
rect 35396 9906 35478 9930
rect 36414 9964 36496 9988
rect 36414 9930 36438 9964
rect 36472 9930 36496 9964
rect 36414 9906 36496 9930
rect 37432 9964 37514 9988
rect 37432 9930 37456 9964
rect 37490 9930 37514 9964
rect 37432 9906 37514 9930
rect 38450 9964 38532 9988
rect 38450 9930 38474 9964
rect 38508 9930 38532 9964
rect 38450 9906 38532 9930
rect 39468 9964 39550 9988
rect 39468 9930 39492 9964
rect 39526 9930 39550 9964
rect 39468 9906 39550 9930
rect 19854 9654 19870 9688
rect 20426 9654 20442 9688
rect 20872 9654 20888 9688
rect 21444 9654 21460 9688
rect 21890 9654 21906 9688
rect 22462 9654 22478 9688
rect 22908 9654 22924 9688
rect 23480 9654 23496 9688
rect 23926 9654 23942 9688
rect 24498 9654 24514 9688
rect 24944 9654 24960 9688
rect 25516 9654 25532 9688
rect 25962 9654 25978 9688
rect 26534 9654 26550 9688
rect 26980 9654 26996 9688
rect 27552 9654 27568 9688
rect 27998 9654 28014 9688
rect 28570 9654 28586 9688
rect 29016 9654 29032 9688
rect 29588 9654 29604 9688
rect 30034 9654 30050 9688
rect 30606 9654 30622 9688
rect 31052 9654 31068 9688
rect 31624 9654 31640 9688
rect 32070 9654 32086 9688
rect 32642 9654 32658 9688
rect 33088 9654 33104 9688
rect 33660 9654 33676 9688
rect 34106 9654 34122 9688
rect 34678 9654 34694 9688
rect 35124 9654 35140 9688
rect 35696 9654 35712 9688
rect 36142 9654 36158 9688
rect 36714 9654 36730 9688
rect 37160 9654 37176 9688
rect 37732 9654 37748 9688
rect 38178 9654 38194 9688
rect 38750 9654 38766 9688
rect 39196 9654 39212 9688
rect 39768 9654 39784 9688
rect 21140 9650 21200 9654
rect 22156 9650 22216 9654
rect 26232 9646 26292 9654
rect 30298 9650 30358 9654
rect 32332 9650 32392 9654
rect 38444 9650 38504 9654
rect 17018 9510 17052 9526
rect 19622 9604 19656 9620
rect 7832 9422 7914 9446
rect 8088 9442 8104 9476
rect 8660 9442 8676 9476
rect 7832 9388 7856 9422
rect 7890 9388 7914 9422
rect 7832 9364 7914 9388
rect 8850 9422 8932 9446
rect 9106 9442 9122 9476
rect 9678 9442 9694 9476
rect 8850 9388 8874 9422
rect 8908 9388 8932 9422
rect 8088 9334 8104 9368
rect 8660 9334 8676 9368
rect 8850 9364 8932 9388
rect 9868 9422 9950 9446
rect 10124 9442 10140 9476
rect 10696 9442 10712 9476
rect 9868 9388 9892 9422
rect 9926 9388 9950 9422
rect 9106 9334 9122 9368
rect 9678 9334 9694 9368
rect 9868 9364 9950 9388
rect 10886 9422 10968 9446
rect 11142 9442 11158 9476
rect 11714 9442 11730 9476
rect 10886 9388 10910 9422
rect 10944 9388 10968 9422
rect 10124 9334 10140 9368
rect 10696 9334 10712 9368
rect 10886 9364 10968 9388
rect 11904 9422 11986 9446
rect 12160 9442 12176 9476
rect 12732 9442 12748 9476
rect 11904 9388 11928 9422
rect 11962 9388 11986 9422
rect 11142 9334 11158 9368
rect 11714 9334 11730 9368
rect 11904 9364 11986 9388
rect 12922 9422 13004 9446
rect 13178 9442 13194 9476
rect 13750 9442 13766 9476
rect 12922 9388 12946 9422
rect 12980 9388 13004 9422
rect 12160 9334 12176 9368
rect 12732 9334 12748 9368
rect 12922 9364 13004 9388
rect 13940 9422 14022 9446
rect 14196 9442 14212 9476
rect 14768 9442 14784 9476
rect 13940 9388 13964 9422
rect 13998 9388 14022 9422
rect 13178 9334 13194 9368
rect 13750 9334 13766 9368
rect 13940 9364 14022 9388
rect 14958 9422 15040 9446
rect 15214 9442 15230 9476
rect 15786 9442 15802 9476
rect 14958 9388 14982 9422
rect 15016 9388 15040 9422
rect 14196 9334 14212 9368
rect 14768 9334 14784 9368
rect 14958 9364 15040 9388
rect 15976 9422 16058 9446
rect 16232 9442 16248 9476
rect 16804 9442 16820 9476
rect 15976 9388 16000 9422
rect 16034 9388 16058 9422
rect 15214 9334 15230 9368
rect 15786 9334 15802 9368
rect 15976 9364 16058 9388
rect 17004 9422 17086 9446
rect 17004 9388 17028 9422
rect 17062 9388 17086 9422
rect 16232 9334 16248 9368
rect 16804 9334 16820 9368
rect 17004 9364 17086 9388
rect 13444 9332 13504 9334
rect 7856 9284 7890 9300
rect 7856 8692 7890 8708
rect 8874 9284 8908 9300
rect 8874 8692 8908 8708
rect 9892 9284 9926 9300
rect 9892 8692 9926 8708
rect 10910 9284 10944 9300
rect 10910 8692 10944 8708
rect 11928 9284 11962 9300
rect 11928 8692 11962 8708
rect 12946 9284 12980 9300
rect 12946 8692 12980 8708
rect 13964 9284 13998 9300
rect 13964 8692 13998 8708
rect 14982 9284 15016 9300
rect 14982 8692 15016 8708
rect 16000 9284 16034 9300
rect 16000 8692 16034 8708
rect 17018 9284 17052 9300
rect 19622 9012 19656 9028
rect 20640 9604 20674 9620
rect 20640 9012 20674 9028
rect 21658 9604 21692 9620
rect 21658 9012 21692 9028
rect 22676 9604 22710 9620
rect 22676 9012 22710 9028
rect 23694 9604 23728 9620
rect 23694 9012 23728 9028
rect 24712 9604 24746 9620
rect 24712 9012 24746 9028
rect 25730 9604 25764 9620
rect 25730 9012 25764 9028
rect 26748 9604 26782 9620
rect 26748 9012 26782 9028
rect 27766 9604 27800 9620
rect 27766 9012 27800 9028
rect 28784 9604 28818 9620
rect 28784 9012 28818 9028
rect 29802 9604 29836 9620
rect 29802 9012 29836 9028
rect 30820 9604 30854 9620
rect 30820 9012 30854 9028
rect 31838 9604 31872 9620
rect 31838 9012 31872 9028
rect 32856 9604 32890 9620
rect 32856 9012 32890 9028
rect 33874 9604 33908 9620
rect 33874 9012 33908 9028
rect 34892 9604 34926 9620
rect 34892 9012 34926 9028
rect 35910 9604 35944 9620
rect 35910 9012 35944 9028
rect 36928 9604 36962 9620
rect 36928 9012 36962 9028
rect 37946 9604 37980 9620
rect 37946 9012 37980 9028
rect 38964 9604 38998 9620
rect 38964 9012 38998 9028
rect 39982 9604 40016 9620
rect 40016 9028 40022 9076
rect 39982 9012 40016 9028
rect 23166 8978 23226 8980
rect 19854 8944 19870 8978
rect 20426 8944 20442 8978
rect 20872 8944 20888 8978
rect 21444 8944 21460 8978
rect 21890 8944 21906 8978
rect 22462 8944 22478 8978
rect 22908 8944 22924 8978
rect 23480 8944 23496 8978
rect 23926 8944 23942 8978
rect 24498 8944 24514 8978
rect 24944 8944 24960 8978
rect 25516 8944 25532 8978
rect 25962 8944 25978 8978
rect 26534 8944 26550 8978
rect 26980 8944 26996 8978
rect 27552 8944 27568 8978
rect 27998 8944 28014 8978
rect 28570 8944 28586 8978
rect 29016 8944 29032 8978
rect 29588 8944 29604 8978
rect 30034 8944 30050 8978
rect 30606 8944 30622 8978
rect 31052 8944 31068 8978
rect 31624 8944 31640 8978
rect 32070 8944 32086 8978
rect 32642 8944 32658 8978
rect 33088 8944 33104 8978
rect 33660 8944 33676 8978
rect 34106 8944 34122 8978
rect 34678 8944 34694 8978
rect 35124 8944 35140 8978
rect 35696 8944 35712 8978
rect 36142 8944 36158 8978
rect 36714 8944 36730 8978
rect 37160 8944 37176 8978
rect 37732 8944 37748 8978
rect 38178 8944 38194 8978
rect 38750 8944 38766 8978
rect 39196 8944 39212 8978
rect 39768 8944 39784 8978
rect 25200 8940 25260 8944
rect 34358 8930 34418 8944
rect 35392 8930 35452 8944
rect 17018 8692 17052 8708
rect 20114 8728 20196 8752
rect 20114 8694 20138 8728
rect 20172 8694 20196 8728
rect 20114 8670 20196 8694
rect 21132 8728 21214 8752
rect 21132 8694 21156 8728
rect 21190 8694 21214 8728
rect 21132 8670 21214 8694
rect 22150 8728 22232 8752
rect 22150 8694 22174 8728
rect 22208 8694 22232 8728
rect 22150 8670 22232 8694
rect 23168 8728 23250 8752
rect 23168 8694 23192 8728
rect 23226 8694 23250 8728
rect 23168 8670 23250 8694
rect 24186 8728 24268 8752
rect 24186 8694 24210 8728
rect 24244 8694 24268 8728
rect 24186 8670 24268 8694
rect 25204 8728 25286 8752
rect 25204 8694 25228 8728
rect 25262 8694 25286 8728
rect 25204 8670 25286 8694
rect 26222 8728 26304 8752
rect 26222 8694 26246 8728
rect 26280 8694 26304 8728
rect 26222 8670 26304 8694
rect 27240 8728 27322 8752
rect 27240 8694 27264 8728
rect 27298 8694 27322 8728
rect 27240 8670 27322 8694
rect 28258 8728 28340 8752
rect 28258 8694 28282 8728
rect 28316 8694 28340 8728
rect 28258 8670 28340 8694
rect 29276 8728 29358 8752
rect 29276 8694 29300 8728
rect 29334 8694 29358 8728
rect 29276 8670 29358 8694
rect 30294 8728 30376 8752
rect 30294 8694 30318 8728
rect 30352 8694 30376 8728
rect 30294 8670 30376 8694
rect 31312 8728 31394 8752
rect 31312 8694 31336 8728
rect 31370 8694 31394 8728
rect 31312 8670 31394 8694
rect 32330 8728 32412 8752
rect 32330 8694 32354 8728
rect 32388 8694 32412 8728
rect 32330 8670 32412 8694
rect 33348 8728 33430 8752
rect 33348 8694 33372 8728
rect 33406 8694 33430 8728
rect 33348 8670 33430 8694
rect 34366 8728 34448 8752
rect 34366 8694 34390 8728
rect 34424 8694 34448 8728
rect 34366 8670 34448 8694
rect 35384 8728 35466 8752
rect 35384 8694 35408 8728
rect 35442 8694 35466 8728
rect 35384 8670 35466 8694
rect 36402 8728 36484 8752
rect 36402 8694 36426 8728
rect 36460 8694 36484 8728
rect 36402 8670 36484 8694
rect 37420 8728 37502 8752
rect 37420 8694 37444 8728
rect 37478 8694 37502 8728
rect 37420 8670 37502 8694
rect 38438 8728 38520 8752
rect 38438 8694 38462 8728
rect 38496 8694 38520 8728
rect 38438 8670 38520 8694
rect 39456 8728 39538 8752
rect 39456 8694 39480 8728
rect 39514 8694 39538 8728
rect 39456 8670 39538 8694
rect 9370 8658 9430 8660
rect 10384 8658 10444 8660
rect 14458 8658 14518 8660
rect 15474 8658 15534 8660
rect 7832 8604 7914 8628
rect 8088 8624 8104 8658
rect 8660 8624 8676 8658
rect 7832 8570 7856 8604
rect 7890 8570 7914 8604
rect 7832 8546 7914 8570
rect 8850 8604 8932 8628
rect 9106 8624 9122 8658
rect 9678 8624 9694 8658
rect 8850 8570 8874 8604
rect 8908 8570 8932 8604
rect 8088 8516 8104 8550
rect 8660 8516 8676 8550
rect 8850 8546 8932 8570
rect 9868 8604 9950 8628
rect 10124 8624 10140 8658
rect 10696 8624 10712 8658
rect 9868 8570 9892 8604
rect 9926 8570 9950 8604
rect 9106 8516 9122 8550
rect 9678 8516 9694 8550
rect 9868 8546 9950 8570
rect 10886 8604 10968 8628
rect 11142 8624 11158 8658
rect 11714 8624 11730 8658
rect 10886 8570 10910 8604
rect 10944 8570 10968 8604
rect 10124 8516 10140 8550
rect 10696 8516 10712 8550
rect 10886 8546 10968 8570
rect 11904 8604 11986 8628
rect 12160 8624 12176 8658
rect 12732 8624 12748 8658
rect 11904 8570 11928 8604
rect 11962 8570 11986 8604
rect 11142 8516 11158 8550
rect 11714 8516 11730 8550
rect 11904 8546 11986 8570
rect 12922 8604 13004 8628
rect 13178 8624 13194 8658
rect 13750 8624 13766 8658
rect 12922 8570 12946 8604
rect 12980 8570 13004 8604
rect 12160 8516 12176 8550
rect 12732 8516 12748 8550
rect 12922 8546 13004 8570
rect 13940 8604 14022 8628
rect 14196 8624 14212 8658
rect 14768 8624 14784 8658
rect 13940 8570 13964 8604
rect 13998 8570 14022 8604
rect 13178 8516 13194 8550
rect 13750 8516 13766 8550
rect 13940 8546 14022 8570
rect 14958 8604 15040 8628
rect 15214 8624 15230 8658
rect 15786 8624 15802 8658
rect 14958 8570 14982 8604
rect 15016 8570 15040 8604
rect 14196 8516 14212 8550
rect 14768 8516 14784 8550
rect 14958 8546 15040 8570
rect 15976 8604 16058 8628
rect 16232 8624 16248 8658
rect 16804 8624 16820 8658
rect 15976 8570 16000 8604
rect 16034 8570 16058 8604
rect 15214 8516 15230 8550
rect 15786 8516 15802 8550
rect 15976 8546 16058 8570
rect 17004 8604 17086 8628
rect 17004 8570 17028 8604
rect 17062 8570 17086 8604
rect 16232 8516 16248 8550
rect 16804 8516 16820 8550
rect 17004 8546 17086 8570
rect 7856 8466 7890 8482
rect 7856 7874 7890 7890
rect 8874 8466 8908 8482
rect 8874 7874 8908 7890
rect 9892 8466 9926 8482
rect 9892 7874 9926 7890
rect 10910 8466 10944 8482
rect 10910 7874 10944 7890
rect 11928 8466 11962 8482
rect 11928 7874 11962 7890
rect 12946 8466 12980 8482
rect 12946 7874 12980 7890
rect 13964 8466 13998 8482
rect 13964 7874 13998 7890
rect 14982 8466 15016 8482
rect 14982 7874 15016 7890
rect 16000 8466 16034 8482
rect 16000 7874 16034 7890
rect 17018 8466 17052 8482
rect 19852 8420 19868 8454
rect 20424 8420 20440 8454
rect 20870 8420 20886 8454
rect 21442 8420 21458 8454
rect 21888 8420 21904 8454
rect 22460 8420 22476 8454
rect 22906 8420 22922 8454
rect 23478 8420 23494 8454
rect 23924 8420 23940 8454
rect 24496 8420 24512 8454
rect 24942 8420 24958 8454
rect 25514 8420 25530 8454
rect 25960 8420 25976 8454
rect 26532 8420 26548 8454
rect 26978 8420 26994 8454
rect 27550 8420 27566 8454
rect 27996 8420 28012 8454
rect 28568 8420 28584 8454
rect 29014 8420 29030 8454
rect 29586 8420 29602 8454
rect 30032 8420 30048 8454
rect 30604 8420 30620 8454
rect 31050 8420 31066 8454
rect 31622 8420 31638 8454
rect 32068 8420 32084 8454
rect 32640 8420 32656 8454
rect 33086 8420 33102 8454
rect 33658 8420 33674 8454
rect 34104 8420 34120 8454
rect 34676 8420 34692 8454
rect 35122 8420 35138 8454
rect 35694 8420 35710 8454
rect 36140 8420 36156 8454
rect 36712 8420 36728 8454
rect 37158 8420 37174 8454
rect 37730 8420 37746 8454
rect 38176 8420 38192 8454
rect 38748 8420 38764 8454
rect 39194 8420 39210 8454
rect 39766 8420 39782 8454
rect 22162 8416 22222 8420
rect 17018 7874 17052 7890
rect 19620 8370 19654 8386
rect 9374 7840 9434 7842
rect 10388 7840 10448 7842
rect 14462 7840 14522 7842
rect 15478 7840 15538 7842
rect 7832 7786 7914 7810
rect 8088 7806 8104 7840
rect 8660 7806 8676 7840
rect 7832 7752 7856 7786
rect 7890 7752 7914 7786
rect 7832 7728 7914 7752
rect 8850 7786 8932 7810
rect 9106 7806 9122 7840
rect 9678 7806 9694 7840
rect 8850 7752 8874 7786
rect 8908 7752 8932 7786
rect 8088 7698 8104 7732
rect 8660 7698 8676 7732
rect 8850 7728 8932 7752
rect 9868 7786 9950 7810
rect 10124 7806 10140 7840
rect 10696 7806 10712 7840
rect 9868 7752 9892 7786
rect 9926 7752 9950 7786
rect 9106 7698 9122 7732
rect 9678 7698 9694 7732
rect 9868 7728 9950 7752
rect 10886 7786 10968 7810
rect 11142 7806 11158 7840
rect 11714 7806 11730 7840
rect 10886 7752 10910 7786
rect 10944 7752 10968 7786
rect 10124 7698 10140 7732
rect 10696 7698 10712 7732
rect 10886 7728 10968 7752
rect 11904 7786 11986 7810
rect 12160 7806 12176 7840
rect 12732 7806 12748 7840
rect 11904 7752 11928 7786
rect 11962 7752 11986 7786
rect 11142 7698 11158 7732
rect 11714 7698 11730 7732
rect 11904 7728 11986 7752
rect 12922 7786 13004 7810
rect 13178 7806 13194 7840
rect 13750 7806 13766 7840
rect 12922 7752 12946 7786
rect 12980 7752 13004 7786
rect 12160 7698 12176 7732
rect 12732 7698 12748 7732
rect 12922 7728 13004 7752
rect 13940 7786 14022 7810
rect 14196 7806 14212 7840
rect 14768 7806 14784 7840
rect 13940 7752 13964 7786
rect 13998 7752 14022 7786
rect 13178 7698 13194 7732
rect 13750 7698 13766 7732
rect 13940 7728 14022 7752
rect 14958 7786 15040 7810
rect 15214 7806 15230 7840
rect 15786 7806 15802 7840
rect 14958 7752 14982 7786
rect 15016 7752 15040 7786
rect 14196 7698 14212 7732
rect 14768 7698 14784 7732
rect 14958 7728 15040 7752
rect 15976 7786 16058 7810
rect 16232 7806 16248 7840
rect 16804 7806 16820 7840
rect 15976 7752 16000 7786
rect 16034 7752 16058 7786
rect 15214 7698 15230 7732
rect 15786 7698 15802 7732
rect 15976 7728 16058 7752
rect 17004 7786 17086 7810
rect 17004 7752 17028 7786
rect 17062 7752 17086 7786
rect 19620 7778 19654 7794
rect 20638 8370 20672 8386
rect 20638 7778 20672 7794
rect 21656 8370 21690 8386
rect 21656 7778 21690 7794
rect 22674 8370 22708 8386
rect 22674 7778 22708 7794
rect 23692 8370 23726 8386
rect 23692 7778 23726 7794
rect 24710 8370 24744 8386
rect 24710 7778 24744 7794
rect 25728 8370 25762 8386
rect 25728 7778 25762 7794
rect 26746 8370 26780 8386
rect 26746 7778 26780 7794
rect 27764 8370 27798 8386
rect 27764 7778 27798 7794
rect 28782 8370 28816 8386
rect 28782 7778 28816 7794
rect 29800 8370 29834 8386
rect 29800 7778 29834 7794
rect 30818 8370 30852 8386
rect 30818 7778 30852 7794
rect 31836 8370 31870 8386
rect 31836 7778 31870 7794
rect 32854 8370 32888 8386
rect 32854 7778 32888 7794
rect 33872 8370 33906 8386
rect 33872 7778 33906 7794
rect 34890 8370 34924 8386
rect 34890 7778 34924 7794
rect 35908 8370 35942 8386
rect 35908 7778 35942 7794
rect 36926 8370 36960 8386
rect 36926 7778 36960 7794
rect 37944 8370 37978 8386
rect 37944 7778 37978 7794
rect 38962 8370 38996 8386
rect 38962 7778 38996 7794
rect 39980 8370 40014 8386
rect 39980 7778 40014 7794
rect 16232 7698 16248 7732
rect 16804 7698 16820 7732
rect 17004 7728 17086 7752
rect 27230 7744 27290 7748
rect 28258 7744 28318 7746
rect 30302 7744 30362 7748
rect 19852 7710 19868 7744
rect 20424 7710 20440 7744
rect 20870 7710 20886 7744
rect 21442 7710 21458 7744
rect 21888 7710 21904 7744
rect 22460 7710 22476 7744
rect 22906 7710 22922 7744
rect 23478 7710 23494 7744
rect 23924 7710 23940 7744
rect 24496 7710 24512 7744
rect 24942 7710 24958 7744
rect 25514 7710 25530 7744
rect 25960 7710 25976 7744
rect 26532 7710 26548 7744
rect 26978 7710 26994 7744
rect 27550 7710 27566 7744
rect 27996 7710 28012 7744
rect 28568 7710 28584 7744
rect 29014 7710 29030 7744
rect 29586 7710 29602 7744
rect 30032 7710 30048 7744
rect 30604 7710 30620 7744
rect 31050 7710 31066 7744
rect 31622 7710 31638 7744
rect 32068 7710 32084 7744
rect 32640 7710 32656 7744
rect 33086 7710 33102 7744
rect 33658 7710 33674 7744
rect 34104 7710 34120 7744
rect 34676 7710 34692 7744
rect 35122 7710 35138 7744
rect 35694 7710 35710 7744
rect 36140 7710 36156 7744
rect 36712 7710 36728 7744
rect 37158 7710 37174 7744
rect 37730 7710 37746 7744
rect 38176 7710 38192 7744
rect 38748 7710 38764 7744
rect 39194 7710 39210 7744
rect 39766 7710 39782 7744
rect 7856 7648 7890 7664
rect 7856 7056 7890 7072
rect 8874 7648 8908 7664
rect 8874 7056 8908 7072
rect 9892 7648 9926 7664
rect 9892 7056 9926 7072
rect 10910 7648 10944 7664
rect 10910 7056 10944 7072
rect 11928 7648 11962 7664
rect 11928 7056 11962 7072
rect 12946 7648 12980 7664
rect 12946 7056 12980 7072
rect 13964 7648 13998 7664
rect 13964 7056 13998 7072
rect 14982 7648 15016 7664
rect 14982 7056 15016 7072
rect 16000 7648 16034 7664
rect 16000 7056 16034 7072
rect 17018 7648 17052 7664
rect 20114 7504 20196 7528
rect 20114 7470 20138 7504
rect 20172 7470 20196 7504
rect 20114 7446 20196 7470
rect 21132 7504 21214 7528
rect 21132 7470 21156 7504
rect 21190 7470 21214 7504
rect 21132 7446 21214 7470
rect 22150 7504 22232 7528
rect 22150 7470 22174 7504
rect 22208 7470 22232 7504
rect 22150 7446 22232 7470
rect 23168 7504 23250 7528
rect 23168 7470 23192 7504
rect 23226 7470 23250 7504
rect 23168 7446 23250 7470
rect 24186 7504 24268 7528
rect 24186 7470 24210 7504
rect 24244 7470 24268 7504
rect 24186 7446 24268 7470
rect 25204 7504 25286 7528
rect 25204 7470 25228 7504
rect 25262 7470 25286 7504
rect 25204 7446 25286 7470
rect 26222 7504 26304 7528
rect 26222 7470 26246 7504
rect 26280 7470 26304 7504
rect 26222 7446 26304 7470
rect 27240 7504 27322 7528
rect 27240 7470 27264 7504
rect 27298 7470 27322 7504
rect 27240 7446 27322 7470
rect 28258 7504 28340 7528
rect 28258 7470 28282 7504
rect 28316 7470 28340 7504
rect 28258 7446 28340 7470
rect 29276 7504 29358 7528
rect 29276 7470 29300 7504
rect 29334 7470 29358 7504
rect 29276 7446 29358 7470
rect 30294 7504 30376 7528
rect 30294 7470 30318 7504
rect 30352 7470 30376 7504
rect 30294 7446 30376 7470
rect 31312 7504 31394 7528
rect 31312 7470 31336 7504
rect 31370 7470 31394 7504
rect 31312 7446 31394 7470
rect 32330 7504 32412 7528
rect 32330 7470 32354 7504
rect 32388 7470 32412 7504
rect 32330 7446 32412 7470
rect 33348 7504 33430 7528
rect 33348 7470 33372 7504
rect 33406 7470 33430 7504
rect 33348 7446 33430 7470
rect 34366 7504 34448 7528
rect 34366 7470 34390 7504
rect 34424 7470 34448 7504
rect 34366 7446 34448 7470
rect 35384 7504 35466 7528
rect 35384 7470 35408 7504
rect 35442 7470 35466 7504
rect 35384 7446 35466 7470
rect 36402 7504 36484 7528
rect 36402 7470 36426 7504
rect 36460 7470 36484 7504
rect 36402 7446 36484 7470
rect 37420 7504 37502 7528
rect 37420 7470 37444 7504
rect 37478 7470 37502 7504
rect 37420 7446 37502 7470
rect 38438 7504 38520 7528
rect 38438 7470 38462 7504
rect 38496 7470 38520 7504
rect 38438 7446 38520 7470
rect 39456 7504 39538 7528
rect 39456 7470 39480 7504
rect 39514 7470 39538 7504
rect 39456 7446 39538 7470
rect 19852 7186 19868 7220
rect 20424 7186 20440 7220
rect 20870 7186 20886 7220
rect 21442 7186 21458 7220
rect 21888 7186 21904 7220
rect 22460 7186 22476 7220
rect 22906 7186 22922 7220
rect 23478 7186 23494 7220
rect 23924 7186 23940 7220
rect 24496 7186 24512 7220
rect 24942 7186 24958 7220
rect 25514 7186 25530 7220
rect 25960 7186 25976 7220
rect 26532 7186 26548 7220
rect 26978 7186 26994 7220
rect 27550 7186 27566 7220
rect 27996 7186 28012 7220
rect 28568 7186 28584 7220
rect 29014 7186 29030 7220
rect 29586 7186 29602 7220
rect 30032 7186 30048 7220
rect 30604 7186 30620 7220
rect 31050 7186 31066 7220
rect 31622 7186 31638 7220
rect 32068 7186 32084 7220
rect 32640 7186 32656 7220
rect 33086 7186 33102 7220
rect 33658 7186 33674 7220
rect 34104 7186 34120 7220
rect 34676 7186 34692 7220
rect 35122 7186 35138 7220
rect 35694 7186 35710 7220
rect 36140 7186 36156 7220
rect 36712 7186 36728 7220
rect 37158 7186 37174 7220
rect 37730 7186 37746 7220
rect 38176 7186 38192 7220
rect 38748 7186 38764 7220
rect 39194 7186 39210 7220
rect 39766 7186 39782 7220
rect 17018 7056 17052 7072
rect 19620 7136 19654 7152
rect 8348 7022 8408 7024
rect 9374 7022 9434 7026
rect 10388 7022 10448 7026
rect 11408 7022 11468 7024
rect 12430 7022 12490 7024
rect 14462 7022 14522 7026
rect 15478 7022 15538 7026
rect 16498 7022 16558 7024
rect 7832 6968 7914 6992
rect 8088 6988 8104 7022
rect 8660 6988 8676 7022
rect 7832 6934 7856 6968
rect 7890 6934 7914 6968
rect 7832 6910 7914 6934
rect 8850 6968 8932 6992
rect 9106 6988 9122 7022
rect 9678 6988 9694 7022
rect 8850 6934 8874 6968
rect 8908 6934 8932 6968
rect 8088 6880 8104 6914
rect 8660 6880 8676 6914
rect 8850 6910 8932 6934
rect 9868 6968 9950 6992
rect 10124 6988 10140 7022
rect 10696 6988 10712 7022
rect 9868 6934 9892 6968
rect 9926 6934 9950 6968
rect 9106 6880 9122 6914
rect 9678 6880 9694 6914
rect 9868 6910 9950 6934
rect 10886 6968 10968 6992
rect 11142 6988 11158 7022
rect 11714 6988 11730 7022
rect 10886 6934 10910 6968
rect 10944 6934 10968 6968
rect 10124 6880 10140 6914
rect 10696 6880 10712 6914
rect 10886 6910 10968 6934
rect 11904 6968 11986 6992
rect 12160 6988 12176 7022
rect 12732 6988 12748 7022
rect 11904 6934 11928 6968
rect 11962 6934 11986 6968
rect 11142 6880 11158 6914
rect 11714 6880 11730 6914
rect 11904 6910 11986 6934
rect 12922 6968 13004 6992
rect 13178 6988 13194 7022
rect 13750 6988 13766 7022
rect 12922 6934 12946 6968
rect 12980 6934 13004 6968
rect 12160 6880 12176 6914
rect 12732 6880 12748 6914
rect 12922 6910 13004 6934
rect 13940 6968 14022 6992
rect 14196 6988 14212 7022
rect 14768 6988 14784 7022
rect 13940 6934 13964 6968
rect 13998 6934 14022 6968
rect 13178 6880 13194 6914
rect 13750 6880 13766 6914
rect 13940 6910 14022 6934
rect 14958 6968 15040 6992
rect 15214 6988 15230 7022
rect 15786 6988 15802 7022
rect 14958 6934 14982 6968
rect 15016 6934 15040 6968
rect 14196 6880 14212 6914
rect 14768 6880 14784 6914
rect 14958 6910 15040 6934
rect 15976 6968 16058 6992
rect 16232 6988 16248 7022
rect 16804 6988 16820 7022
rect 15976 6934 16000 6968
rect 16034 6934 16058 6968
rect 15214 6880 15230 6914
rect 15786 6880 15802 6914
rect 15976 6910 16058 6934
rect 17004 6968 17086 6992
rect 17004 6934 17028 6968
rect 17062 6934 17086 6968
rect 16232 6880 16248 6914
rect 16804 6880 16820 6914
rect 17004 6910 17086 6934
rect 7856 6830 7890 6846
rect 7856 6238 7890 6254
rect 8874 6830 8908 6846
rect 8874 6238 8908 6254
rect 9892 6830 9926 6846
rect 9892 6238 9926 6254
rect 10910 6830 10944 6846
rect 10910 6238 10944 6254
rect 11928 6830 11962 6846
rect 11928 6238 11962 6254
rect 12946 6830 12980 6846
rect 12946 6238 12980 6254
rect 13964 6830 13998 6846
rect 13964 6238 13998 6254
rect 14982 6830 15016 6846
rect 14982 6238 15016 6254
rect 16000 6830 16034 6846
rect 16000 6238 16034 6254
rect 17018 6830 17052 6846
rect 19620 6544 19654 6560
rect 20638 7136 20672 7152
rect 20638 6544 20672 6560
rect 21656 7136 21690 7152
rect 21656 6544 21690 6560
rect 22674 7136 22708 7152
rect 22674 6544 22708 6560
rect 23692 7136 23726 7152
rect 23692 6544 23726 6560
rect 24710 7136 24744 7152
rect 24710 6544 24744 6560
rect 25728 7136 25762 7152
rect 25728 6544 25762 6560
rect 26746 7136 26780 7152
rect 26746 6544 26780 6560
rect 27764 7136 27798 7152
rect 27764 6544 27798 6560
rect 28782 7136 28816 7152
rect 28782 6544 28816 6560
rect 29800 7136 29834 7152
rect 29800 6544 29834 6560
rect 30818 7136 30852 7152
rect 30818 6544 30852 6560
rect 31836 7136 31870 7152
rect 31836 6544 31870 6560
rect 32854 7136 32888 7152
rect 32854 6544 32888 6560
rect 33872 7136 33906 7152
rect 33872 6544 33906 6560
rect 34890 7136 34924 7152
rect 34890 6544 34924 6560
rect 35908 7136 35942 7152
rect 35908 6544 35942 6560
rect 36926 7136 36960 7152
rect 36926 6544 36960 6560
rect 37944 7136 37978 7152
rect 37944 6544 37978 6560
rect 38962 7136 38996 7152
rect 38962 6544 38996 6560
rect 39980 7136 40014 7152
rect 39980 6544 40014 6560
rect 19852 6476 19868 6510
rect 20424 6476 20440 6510
rect 20870 6476 20886 6510
rect 21442 6476 21458 6510
rect 21888 6476 21904 6510
rect 22460 6476 22476 6510
rect 22906 6476 22922 6510
rect 23478 6476 23494 6510
rect 23924 6476 23940 6510
rect 24496 6476 24512 6510
rect 24942 6476 24958 6510
rect 25514 6476 25530 6510
rect 25960 6476 25976 6510
rect 26532 6476 26548 6510
rect 26978 6476 26994 6510
rect 27550 6476 27566 6510
rect 27996 6476 28012 6510
rect 28568 6476 28584 6510
rect 29014 6476 29030 6510
rect 29586 6476 29602 6510
rect 30032 6476 30048 6510
rect 30604 6476 30620 6510
rect 31050 6476 31066 6510
rect 31622 6476 31638 6510
rect 32068 6476 32084 6510
rect 32640 6476 32656 6510
rect 33086 6476 33102 6510
rect 33658 6476 33674 6510
rect 34104 6476 34120 6510
rect 34676 6476 34692 6510
rect 35122 6476 35138 6510
rect 35694 6476 35710 6510
rect 36140 6476 36156 6510
rect 36712 6476 36728 6510
rect 37158 6476 37174 6510
rect 37730 6476 37746 6510
rect 38176 6476 38192 6510
rect 38748 6476 38764 6510
rect 39194 6476 39210 6510
rect 39766 6476 39782 6510
rect 17018 6238 17052 6254
rect 20126 6268 20208 6292
rect 20126 6234 20150 6268
rect 20184 6234 20208 6268
rect 20126 6210 20208 6234
rect 21144 6268 21226 6292
rect 21144 6234 21168 6268
rect 21202 6234 21226 6268
rect 21144 6210 21226 6234
rect 22162 6268 22244 6292
rect 22162 6234 22186 6268
rect 22220 6234 22244 6268
rect 22162 6210 22244 6234
rect 23180 6268 23262 6292
rect 23180 6234 23204 6268
rect 23238 6234 23262 6268
rect 23180 6210 23262 6234
rect 24198 6268 24280 6292
rect 24198 6234 24222 6268
rect 24256 6234 24280 6268
rect 24198 6210 24280 6234
rect 25216 6268 25298 6292
rect 25216 6234 25240 6268
rect 25274 6234 25298 6268
rect 25216 6210 25298 6234
rect 26234 6268 26316 6292
rect 26234 6234 26258 6268
rect 26292 6234 26316 6268
rect 26234 6210 26316 6234
rect 27252 6268 27334 6292
rect 27252 6234 27276 6268
rect 27310 6234 27334 6268
rect 27252 6210 27334 6234
rect 28270 6268 28352 6292
rect 28270 6234 28294 6268
rect 28328 6234 28352 6268
rect 28270 6210 28352 6234
rect 29288 6268 29370 6292
rect 29288 6234 29312 6268
rect 29346 6234 29370 6268
rect 29288 6210 29370 6234
rect 30306 6268 30388 6292
rect 30306 6234 30330 6268
rect 30364 6234 30388 6268
rect 30306 6210 30388 6234
rect 31324 6268 31406 6292
rect 31324 6234 31348 6268
rect 31382 6234 31406 6268
rect 31324 6210 31406 6234
rect 32342 6268 32424 6292
rect 32342 6234 32366 6268
rect 32400 6234 32424 6268
rect 32342 6210 32424 6234
rect 33360 6268 33442 6292
rect 33360 6234 33384 6268
rect 33418 6234 33442 6268
rect 33360 6210 33442 6234
rect 34378 6268 34460 6292
rect 34378 6234 34402 6268
rect 34436 6234 34460 6268
rect 34378 6210 34460 6234
rect 35396 6268 35478 6292
rect 35396 6234 35420 6268
rect 35454 6234 35478 6268
rect 35396 6210 35478 6234
rect 36414 6268 36496 6292
rect 36414 6234 36438 6268
rect 36472 6234 36496 6268
rect 36414 6210 36496 6234
rect 37432 6268 37514 6292
rect 37432 6234 37456 6268
rect 37490 6234 37514 6268
rect 37432 6210 37514 6234
rect 38450 6268 38532 6292
rect 38450 6234 38474 6268
rect 38508 6234 38532 6268
rect 38450 6210 38532 6234
rect 39468 6268 39550 6292
rect 39468 6234 39492 6268
rect 39526 6234 39550 6268
rect 39468 6210 39550 6234
rect 8088 6170 8104 6204
rect 8660 6170 8676 6204
rect 9106 6170 9122 6204
rect 9678 6170 9694 6204
rect 10124 6170 10140 6204
rect 10696 6170 10712 6204
rect 11142 6170 11158 6204
rect 11714 6170 11730 6204
rect 12160 6170 12176 6204
rect 12732 6170 12748 6204
rect 13178 6170 13194 6204
rect 13750 6170 13766 6204
rect 14196 6170 14212 6204
rect 14768 6170 14784 6204
rect 15214 6170 15230 6204
rect 15786 6170 15802 6204
rect 16232 6170 16248 6204
rect 16804 6170 16820 6204
rect 7820 6074 7902 6098
rect 7820 6040 7844 6074
rect 7878 6040 7902 6074
rect 7820 6016 7902 6040
rect 8838 6074 8920 6098
rect 8838 6040 8862 6074
rect 8896 6040 8920 6074
rect 8838 6016 8920 6040
rect 9856 6074 9938 6098
rect 9856 6040 9880 6074
rect 9914 6040 9938 6074
rect 9856 6016 9938 6040
rect 10874 6074 10956 6098
rect 10874 6040 10898 6074
rect 10932 6040 10956 6074
rect 10874 6016 10956 6040
rect 11892 6074 11974 6098
rect 11892 6040 11916 6074
rect 11950 6040 11974 6074
rect 11892 6016 11974 6040
rect 12910 6074 12992 6098
rect 12910 6040 12934 6074
rect 12968 6040 12992 6074
rect 12910 6016 12992 6040
rect 13928 6074 14010 6098
rect 13928 6040 13952 6074
rect 13986 6040 14010 6074
rect 13928 6016 14010 6040
rect 14946 6074 15028 6098
rect 14946 6040 14970 6074
rect 15004 6040 15028 6074
rect 14946 6016 15028 6040
rect 15964 6074 16046 6098
rect 15964 6040 15988 6074
rect 16022 6040 16046 6074
rect 15964 6016 16046 6040
rect 16992 6074 17074 6098
rect 16992 6040 17016 6074
rect 17050 6040 17074 6074
rect 16992 6016 17074 6040
rect 19852 5954 19868 5988
rect 20424 5954 20440 5988
rect 20870 5954 20886 5988
rect 21442 5954 21458 5988
rect 21888 5954 21904 5988
rect 22460 5954 22476 5988
rect 22906 5954 22922 5988
rect 23478 5954 23494 5988
rect 23924 5954 23940 5988
rect 24496 5954 24512 5988
rect 24942 5954 24958 5988
rect 25514 5954 25530 5988
rect 25960 5954 25976 5988
rect 26532 5954 26548 5988
rect 26978 5954 26994 5988
rect 27550 5954 27566 5988
rect 27996 5954 28012 5988
rect 28568 5954 28584 5988
rect 29014 5954 29030 5988
rect 29586 5954 29602 5988
rect 30032 5954 30048 5988
rect 30604 5954 30620 5988
rect 31050 5954 31066 5988
rect 31622 5954 31638 5988
rect 32068 5954 32084 5988
rect 32640 5954 32656 5988
rect 33086 5954 33102 5988
rect 33658 5954 33674 5988
rect 34104 5954 34120 5988
rect 34676 5954 34692 5988
rect 35122 5954 35138 5988
rect 35694 5954 35710 5988
rect 36140 5954 36156 5988
rect 36712 5954 36728 5988
rect 37158 5954 37174 5988
rect 37730 5954 37746 5988
rect 38176 5954 38192 5988
rect 38748 5954 38764 5988
rect 39194 5954 39210 5988
rect 39766 5954 39782 5988
rect 19620 5904 19654 5920
rect 19620 5312 19654 5328
rect 20638 5904 20672 5920
rect 20638 5312 20672 5328
rect 21656 5904 21690 5920
rect 21656 5312 21690 5328
rect 22674 5904 22708 5920
rect 22674 5312 22708 5328
rect 23692 5904 23726 5920
rect 23692 5312 23726 5328
rect 24710 5904 24744 5920
rect 24710 5312 24744 5328
rect 25728 5904 25762 5920
rect 25728 5312 25762 5328
rect 26746 5904 26780 5920
rect 26746 5312 26780 5328
rect 27764 5904 27798 5920
rect 27764 5312 27798 5328
rect 28782 5904 28816 5920
rect 28782 5312 28816 5328
rect 29800 5904 29834 5920
rect 29800 5312 29834 5328
rect 30818 5904 30852 5920
rect 30818 5312 30852 5328
rect 31836 5904 31870 5920
rect 31836 5312 31870 5328
rect 32854 5904 32888 5920
rect 32854 5312 32888 5328
rect 33872 5904 33906 5920
rect 33872 5312 33906 5328
rect 34890 5904 34924 5920
rect 34890 5312 34924 5328
rect 35908 5904 35942 5920
rect 35908 5312 35942 5328
rect 36926 5904 36960 5920
rect 36926 5312 36960 5328
rect 37944 5904 37978 5920
rect 37944 5312 37978 5328
rect 38962 5904 38996 5920
rect 38962 5312 38996 5328
rect 39980 5904 40014 5920
rect 39980 5312 40014 5328
rect 28270 5278 28330 5280
rect 30314 5278 30374 5282
rect 38448 5278 38508 5280
rect 19852 5244 19868 5278
rect 20424 5244 20440 5278
rect 20870 5244 20886 5278
rect 21442 5244 21458 5278
rect 21888 5244 21904 5278
rect 22460 5244 22476 5278
rect 22906 5244 22922 5278
rect 23478 5244 23494 5278
rect 23924 5244 23940 5278
rect 24496 5244 24512 5278
rect 24942 5244 24958 5278
rect 25514 5244 25530 5278
rect 25960 5244 25976 5278
rect 26532 5244 26548 5278
rect 26978 5244 26994 5278
rect 27550 5244 27566 5278
rect 27996 5244 28012 5278
rect 28568 5244 28584 5278
rect 29014 5244 29030 5278
rect 29586 5244 29602 5278
rect 30032 5244 30048 5278
rect 30604 5244 30620 5278
rect 31050 5244 31066 5278
rect 31622 5244 31638 5278
rect 32068 5244 32084 5278
rect 32640 5244 32656 5278
rect 33086 5244 33102 5278
rect 33658 5244 33674 5278
rect 34104 5244 34120 5278
rect 34676 5244 34692 5278
rect 35122 5244 35138 5278
rect 35694 5244 35710 5278
rect 36140 5244 36156 5278
rect 36712 5244 36728 5278
rect 37158 5244 37174 5278
rect 37730 5244 37746 5278
rect 38176 5244 38192 5278
rect 38748 5244 38764 5278
rect 39194 5244 39210 5278
rect 39766 5244 39782 5278
rect 7024 5126 7106 5150
rect 7024 5092 7048 5126
rect 7082 5092 7106 5126
rect 7024 5068 7106 5092
rect 8042 5126 8124 5150
rect 8042 5092 8066 5126
rect 8100 5092 8124 5126
rect 8042 5068 8124 5092
rect 9060 5126 9142 5150
rect 9060 5092 9084 5126
rect 9118 5092 9142 5126
rect 9060 5068 9142 5092
rect 10078 5126 10160 5150
rect 10078 5092 10102 5126
rect 10136 5092 10160 5126
rect 10078 5068 10160 5092
rect 11096 5126 11178 5150
rect 11096 5092 11120 5126
rect 11154 5092 11178 5126
rect 11096 5068 11178 5092
rect 12114 5126 12196 5150
rect 12114 5092 12138 5126
rect 12172 5092 12196 5126
rect 12114 5068 12196 5092
rect 13132 5126 13214 5150
rect 13132 5092 13156 5126
rect 13190 5092 13214 5126
rect 13132 5068 13214 5092
rect 14150 5126 14232 5150
rect 14150 5092 14174 5126
rect 14208 5092 14232 5126
rect 14150 5068 14232 5092
rect 15168 5126 15250 5150
rect 15168 5092 15192 5126
rect 15226 5092 15250 5126
rect 15168 5068 15250 5092
rect 16186 5126 16268 5150
rect 16186 5092 16210 5126
rect 16244 5092 16268 5126
rect 16186 5068 16268 5092
rect 17204 5126 17286 5150
rect 17204 5092 17228 5126
rect 17262 5092 17286 5126
rect 17204 5068 17286 5092
rect 20126 5020 20208 5044
rect 20126 4986 20150 5020
rect 20184 4986 20208 5020
rect 20126 4962 20208 4986
rect 21144 5020 21226 5044
rect 21144 4986 21168 5020
rect 21202 4986 21226 5020
rect 21144 4962 21226 4986
rect 22162 5020 22244 5044
rect 22162 4986 22186 5020
rect 22220 4986 22244 5020
rect 22162 4962 22244 4986
rect 23180 5020 23262 5044
rect 23180 4986 23204 5020
rect 23238 4986 23262 5020
rect 23180 4962 23262 4986
rect 24198 5020 24280 5044
rect 24198 4986 24222 5020
rect 24256 4986 24280 5020
rect 24198 4962 24280 4986
rect 25216 5020 25298 5044
rect 25216 4986 25240 5020
rect 25274 4986 25298 5020
rect 25216 4962 25298 4986
rect 26234 5020 26316 5044
rect 26234 4986 26258 5020
rect 26292 4986 26316 5020
rect 26234 4962 26316 4986
rect 27252 5020 27334 5044
rect 27252 4986 27276 5020
rect 27310 4986 27334 5020
rect 27252 4962 27334 4986
rect 28270 5020 28352 5044
rect 28270 4986 28294 5020
rect 28328 4986 28352 5020
rect 28270 4962 28352 4986
rect 29288 5020 29370 5044
rect 29288 4986 29312 5020
rect 29346 4986 29370 5020
rect 29288 4962 29370 4986
rect 30306 5020 30388 5044
rect 30306 4986 30330 5020
rect 30364 4986 30388 5020
rect 30306 4962 30388 4986
rect 31324 5020 31406 5044
rect 31324 4986 31348 5020
rect 31382 4986 31406 5020
rect 31324 4962 31406 4986
rect 32342 5020 32424 5044
rect 32342 4986 32366 5020
rect 32400 4986 32424 5020
rect 32342 4962 32424 4986
rect 33360 5020 33442 5044
rect 33360 4986 33384 5020
rect 33418 4986 33442 5020
rect 33360 4962 33442 4986
rect 34378 5020 34460 5044
rect 34378 4986 34402 5020
rect 34436 4986 34460 5020
rect 34378 4962 34460 4986
rect 35396 5020 35478 5044
rect 35396 4986 35420 5020
rect 35454 4986 35478 5020
rect 35396 4962 35478 4986
rect 36414 5020 36496 5044
rect 36414 4986 36438 5020
rect 36472 4986 36496 5020
rect 36414 4962 36496 4986
rect 37432 5020 37514 5044
rect 37432 4986 37456 5020
rect 37490 4986 37514 5020
rect 37432 4962 37514 4986
rect 38450 5020 38532 5044
rect 38450 4986 38474 5020
rect 38508 4986 38532 5020
rect 38450 4962 38532 4986
rect 39468 5020 39550 5044
rect 39468 4986 39492 5020
rect 39526 4986 39550 5020
rect 39468 4962 39550 4986
rect 6764 4856 6780 4890
rect 7336 4856 7352 4890
rect 7782 4856 7798 4890
rect 8354 4856 8370 4890
rect 8800 4856 8816 4890
rect 9372 4856 9388 4890
rect 9818 4856 9834 4890
rect 10390 4856 10406 4890
rect 10836 4856 10852 4890
rect 11408 4856 11424 4890
rect 11854 4856 11870 4890
rect 12426 4856 12442 4890
rect 12872 4856 12888 4890
rect 13444 4856 13460 4890
rect 13890 4856 13906 4890
rect 14462 4856 14478 4890
rect 14908 4856 14924 4890
rect 15480 4856 15496 4890
rect 15926 4856 15942 4890
rect 16498 4856 16514 4890
rect 16944 4856 16960 4890
rect 17516 4856 17532 4890
rect 6532 4806 6566 4822
rect 6532 4214 6566 4230
rect 7550 4806 7584 4822
rect 7550 4214 7584 4230
rect 8568 4806 8602 4822
rect 8568 4214 8602 4230
rect 9586 4806 9620 4822
rect 9586 4214 9620 4230
rect 10604 4806 10638 4822
rect 10604 4214 10638 4230
rect 11622 4806 11656 4822
rect 11622 4214 11656 4230
rect 12640 4806 12674 4822
rect 12640 4214 12674 4230
rect 13658 4806 13692 4822
rect 13658 4214 13692 4230
rect 14676 4806 14710 4822
rect 14676 4214 14710 4230
rect 15694 4806 15728 4822
rect 15694 4214 15728 4230
rect 16712 4806 16746 4822
rect 16712 4214 16746 4230
rect 17730 4806 17764 4822
rect 19852 4720 19868 4754
rect 20424 4720 20440 4754
rect 20870 4720 20886 4754
rect 21442 4720 21458 4754
rect 21888 4720 21904 4754
rect 22460 4720 22476 4754
rect 22906 4720 22922 4754
rect 23478 4720 23494 4754
rect 23924 4720 23940 4754
rect 24496 4720 24512 4754
rect 24942 4720 24958 4754
rect 25514 4720 25530 4754
rect 25960 4720 25976 4754
rect 26532 4720 26548 4754
rect 26978 4720 26994 4754
rect 27550 4720 27566 4754
rect 27996 4720 28012 4754
rect 28568 4720 28584 4754
rect 29014 4720 29030 4754
rect 29586 4720 29602 4754
rect 30032 4720 30048 4754
rect 30604 4720 30620 4754
rect 31050 4720 31066 4754
rect 31622 4720 31638 4754
rect 32068 4720 32084 4754
rect 32640 4720 32656 4754
rect 33086 4720 33102 4754
rect 33658 4720 33674 4754
rect 34104 4720 34120 4754
rect 34676 4720 34692 4754
rect 35122 4720 35138 4754
rect 35694 4720 35710 4754
rect 36140 4720 36156 4754
rect 36712 4720 36728 4754
rect 37158 4720 37174 4754
rect 37730 4720 37746 4754
rect 38176 4720 38192 4754
rect 38748 4720 38764 4754
rect 39194 4720 39210 4754
rect 39766 4720 39782 4754
rect 17730 4214 17764 4230
rect 19620 4670 19654 4686
rect 6764 4146 6780 4180
rect 7336 4146 7352 4180
rect 7782 4146 7798 4180
rect 8354 4146 8370 4180
rect 8800 4146 8816 4180
rect 9372 4146 9388 4180
rect 9818 4146 9834 4180
rect 10390 4146 10406 4180
rect 10836 4146 10852 4180
rect 11408 4146 11424 4180
rect 11854 4146 11870 4180
rect 12426 4146 12442 4180
rect 12872 4146 12888 4180
rect 13444 4146 13460 4180
rect 13890 4146 13906 4180
rect 14462 4146 14478 4180
rect 14908 4146 14924 4180
rect 15480 4146 15496 4180
rect 15926 4146 15942 4180
rect 16498 4146 16514 4180
rect 16944 4146 16960 4180
rect 17516 4146 17532 4180
rect 19620 4078 19654 4094
rect 20638 4670 20672 4686
rect 20638 4078 20672 4094
rect 21656 4670 21690 4686
rect 21656 4078 21690 4094
rect 22674 4670 22708 4686
rect 22674 4078 22708 4094
rect 23692 4670 23726 4686
rect 23692 4078 23726 4094
rect 24710 4670 24744 4686
rect 24710 4078 24744 4094
rect 25728 4670 25762 4686
rect 25728 4078 25762 4094
rect 26746 4670 26780 4686
rect 26746 4078 26780 4094
rect 27764 4670 27798 4686
rect 27764 4078 27798 4094
rect 28782 4670 28816 4686
rect 28782 4078 28816 4094
rect 29800 4670 29834 4686
rect 29800 4078 29834 4094
rect 30818 4670 30852 4686
rect 30818 4078 30852 4094
rect 31836 4670 31870 4686
rect 31836 4078 31870 4094
rect 32854 4670 32888 4686
rect 32854 4078 32888 4094
rect 33872 4670 33906 4686
rect 33872 4078 33906 4094
rect 34890 4670 34924 4686
rect 34890 4078 34924 4094
rect 35908 4670 35942 4686
rect 35908 4078 35942 4094
rect 36926 4670 36960 4686
rect 36926 4078 36960 4094
rect 37944 4670 37978 4686
rect 37944 4078 37978 4094
rect 38962 4670 38996 4686
rect 38962 4078 38996 4094
rect 39980 4670 40014 4686
rect 39980 4078 40014 4094
rect 22146 4044 22206 4048
rect 19852 4010 19868 4044
rect 20424 4010 20440 4044
rect 20870 4010 20886 4044
rect 21442 4010 21458 4044
rect 21888 4010 21904 4044
rect 22460 4010 22476 4044
rect 22906 4010 22922 4044
rect 23478 4010 23494 4044
rect 23924 4010 23940 4044
rect 24496 4010 24512 4044
rect 24942 4010 24958 4044
rect 25514 4010 25530 4044
rect 25960 4010 25976 4044
rect 26532 4010 26548 4044
rect 26978 4010 26994 4044
rect 27550 4010 27566 4044
rect 27996 4010 28012 4044
rect 28568 4010 28584 4044
rect 29014 4010 29030 4044
rect 29586 4010 29602 4044
rect 30032 4010 30048 4044
rect 30604 4010 30620 4044
rect 31050 4010 31066 4044
rect 31622 4010 31638 4044
rect 32068 4010 32084 4044
rect 32640 4010 32656 4044
rect 33086 4010 33102 4044
rect 33658 4010 33674 4044
rect 34104 4010 34120 4044
rect 34676 4010 34692 4044
rect 35122 4010 35138 4044
rect 35694 4010 35710 4044
rect 36140 4010 36156 4044
rect 36712 4010 36728 4044
rect 37158 4010 37174 4044
rect 37730 4010 37746 4044
rect 38176 4010 38192 4044
rect 38748 4010 38764 4044
rect 39194 4010 39210 4044
rect 39766 4010 39782 4044
rect 7036 3984 7118 4008
rect 7036 3950 7060 3984
rect 7094 3950 7118 3984
rect 7036 3926 7118 3950
rect 8054 3984 8136 4008
rect 8054 3950 8078 3984
rect 8112 3950 8136 3984
rect 8054 3926 8136 3950
rect 9072 3984 9154 4008
rect 9072 3950 9096 3984
rect 9130 3950 9154 3984
rect 9072 3926 9154 3950
rect 10090 3984 10172 4008
rect 10090 3950 10114 3984
rect 10148 3950 10172 3984
rect 10090 3926 10172 3950
rect 11108 3984 11190 4008
rect 11108 3950 11132 3984
rect 11166 3950 11190 3984
rect 11108 3926 11190 3950
rect 12126 3984 12208 4008
rect 12126 3950 12150 3984
rect 12184 3950 12208 3984
rect 12126 3926 12208 3950
rect 13144 3984 13226 4008
rect 13144 3950 13168 3984
rect 13202 3950 13226 3984
rect 13144 3926 13226 3950
rect 14162 3984 14244 4008
rect 14162 3950 14186 3984
rect 14220 3950 14244 3984
rect 14162 3926 14244 3950
rect 15180 3984 15262 4008
rect 15180 3950 15204 3984
rect 15238 3950 15262 3984
rect 15180 3926 15262 3950
rect 16198 3984 16280 4008
rect 16198 3950 16222 3984
rect 16256 3950 16280 3984
rect 16198 3926 16280 3950
rect 17216 3984 17298 4008
rect 17216 3950 17240 3984
rect 17274 3950 17298 3984
rect 17216 3926 17298 3950
rect 20102 3784 20184 3808
rect 6764 3744 6780 3778
rect 7336 3744 7352 3778
rect 7782 3744 7798 3778
rect 8354 3744 8370 3778
rect 8800 3744 8816 3778
rect 9372 3744 9388 3778
rect 9818 3744 9834 3778
rect 10390 3744 10406 3778
rect 10836 3744 10852 3778
rect 11408 3744 11424 3778
rect 11854 3744 11870 3778
rect 12426 3744 12442 3778
rect 12872 3744 12888 3778
rect 13444 3744 13460 3778
rect 13890 3744 13906 3778
rect 14462 3744 14478 3778
rect 14908 3744 14924 3778
rect 15480 3744 15496 3778
rect 15926 3744 15942 3778
rect 16498 3744 16514 3778
rect 16944 3744 16960 3778
rect 17516 3744 17532 3778
rect 20102 3750 20126 3784
rect 20160 3750 20184 3784
rect 20102 3726 20184 3750
rect 21120 3784 21202 3808
rect 21120 3750 21144 3784
rect 21178 3750 21202 3784
rect 21120 3726 21202 3750
rect 22138 3784 22220 3808
rect 22138 3750 22162 3784
rect 22196 3750 22220 3784
rect 22138 3726 22220 3750
rect 23156 3784 23238 3808
rect 23156 3750 23180 3784
rect 23214 3750 23238 3784
rect 23156 3726 23238 3750
rect 24174 3784 24256 3808
rect 24174 3750 24198 3784
rect 24232 3750 24256 3784
rect 24174 3726 24256 3750
rect 25192 3784 25274 3808
rect 25192 3750 25216 3784
rect 25250 3750 25274 3784
rect 25192 3726 25274 3750
rect 26210 3784 26292 3808
rect 26210 3750 26234 3784
rect 26268 3750 26292 3784
rect 26210 3726 26292 3750
rect 27228 3784 27310 3808
rect 27228 3750 27252 3784
rect 27286 3750 27310 3784
rect 27228 3726 27310 3750
rect 28246 3784 28328 3808
rect 28246 3750 28270 3784
rect 28304 3750 28328 3784
rect 28246 3726 28328 3750
rect 29264 3784 29346 3808
rect 29264 3750 29288 3784
rect 29322 3750 29346 3784
rect 29264 3726 29346 3750
rect 30282 3784 30364 3808
rect 30282 3750 30306 3784
rect 30340 3750 30364 3784
rect 30282 3726 30364 3750
rect 31300 3784 31382 3808
rect 31300 3750 31324 3784
rect 31358 3750 31382 3784
rect 31300 3726 31382 3750
rect 32318 3784 32400 3808
rect 32318 3750 32342 3784
rect 32376 3750 32400 3784
rect 32318 3726 32400 3750
rect 33336 3784 33418 3808
rect 33336 3750 33360 3784
rect 33394 3750 33418 3784
rect 33336 3726 33418 3750
rect 34354 3784 34436 3808
rect 34354 3750 34378 3784
rect 34412 3750 34436 3784
rect 34354 3726 34436 3750
rect 35372 3784 35454 3808
rect 35372 3750 35396 3784
rect 35430 3750 35454 3784
rect 35372 3726 35454 3750
rect 36390 3784 36472 3808
rect 36390 3750 36414 3784
rect 36448 3750 36472 3784
rect 36390 3726 36472 3750
rect 37408 3784 37490 3808
rect 37408 3750 37432 3784
rect 37466 3750 37490 3784
rect 37408 3726 37490 3750
rect 38426 3784 38508 3808
rect 38426 3750 38450 3784
rect 38484 3750 38508 3784
rect 38426 3726 38508 3750
rect 39444 3784 39526 3808
rect 39444 3750 39468 3784
rect 39502 3750 39526 3784
rect 39444 3726 39526 3750
rect 6532 3694 6566 3710
rect 6532 3102 6566 3118
rect 7550 3694 7584 3710
rect 7550 3102 7584 3118
rect 8568 3694 8602 3710
rect 8568 3102 8602 3118
rect 9586 3694 9620 3710
rect 9586 3102 9620 3118
rect 10604 3694 10638 3710
rect 10604 3102 10638 3118
rect 11622 3694 11656 3710
rect 11622 3102 11656 3118
rect 12640 3694 12674 3710
rect 12640 3102 12674 3118
rect 13658 3694 13692 3710
rect 13658 3102 13692 3118
rect 14676 3694 14710 3710
rect 14676 3102 14710 3118
rect 15694 3694 15728 3710
rect 15694 3102 15728 3118
rect 16712 3694 16746 3710
rect 16712 3102 16746 3118
rect 17730 3694 17764 3710
rect 19852 3486 19868 3520
rect 20424 3486 20440 3520
rect 20870 3486 20886 3520
rect 21442 3486 21458 3520
rect 21888 3486 21904 3520
rect 22460 3486 22476 3520
rect 22906 3486 22922 3520
rect 23478 3486 23494 3520
rect 23924 3486 23940 3520
rect 24496 3486 24512 3520
rect 24942 3486 24958 3520
rect 25514 3486 25530 3520
rect 25960 3486 25976 3520
rect 26532 3486 26548 3520
rect 26978 3486 26994 3520
rect 27550 3486 27566 3520
rect 27996 3486 28012 3520
rect 28568 3486 28584 3520
rect 29014 3486 29030 3520
rect 29586 3486 29602 3520
rect 30032 3486 30048 3520
rect 30604 3486 30620 3520
rect 31050 3486 31066 3520
rect 31622 3486 31638 3520
rect 32068 3486 32084 3520
rect 32640 3486 32656 3520
rect 33086 3486 33102 3520
rect 33658 3486 33674 3520
rect 34104 3486 34120 3520
rect 34676 3486 34692 3520
rect 35122 3486 35138 3520
rect 35694 3486 35710 3520
rect 36140 3486 36156 3520
rect 36712 3486 36728 3520
rect 37158 3486 37174 3520
rect 37730 3486 37746 3520
rect 38176 3486 38192 3520
rect 38748 3486 38764 3520
rect 39194 3486 39210 3520
rect 39766 3486 39782 3520
rect 17730 3102 17764 3118
rect 19620 3436 19654 3452
rect 6764 3034 6780 3068
rect 7336 3034 7352 3068
rect 7782 3034 7798 3068
rect 8354 3034 8370 3068
rect 8800 3034 8816 3068
rect 9372 3034 9388 3068
rect 9818 3034 9834 3068
rect 10390 3034 10406 3068
rect 10836 3034 10852 3068
rect 11408 3034 11424 3068
rect 11854 3034 11870 3068
rect 12426 3034 12442 3068
rect 12872 3034 12888 3068
rect 13444 3034 13460 3068
rect 13890 3034 13906 3068
rect 14462 3034 14478 3068
rect 14908 3034 14924 3068
rect 15480 3034 15496 3068
rect 15926 3034 15942 3068
rect 16498 3034 16514 3068
rect 16944 3034 16960 3068
rect 17516 3034 17532 3068
rect 7014 2876 7096 2900
rect 7014 2842 7038 2876
rect 7072 2842 7096 2876
rect 7014 2818 7096 2842
rect 8032 2876 8114 2900
rect 8032 2842 8056 2876
rect 8090 2842 8114 2876
rect 8032 2818 8114 2842
rect 9050 2876 9132 2900
rect 9050 2842 9074 2876
rect 9108 2842 9132 2876
rect 9050 2818 9132 2842
rect 10068 2876 10150 2900
rect 10068 2842 10092 2876
rect 10126 2842 10150 2876
rect 10068 2818 10150 2842
rect 11086 2876 11168 2900
rect 11086 2842 11110 2876
rect 11144 2842 11168 2876
rect 11086 2818 11168 2842
rect 12104 2876 12186 2900
rect 12104 2842 12128 2876
rect 12162 2842 12186 2876
rect 12104 2818 12186 2842
rect 13122 2876 13204 2900
rect 13122 2842 13146 2876
rect 13180 2842 13204 2876
rect 13122 2818 13204 2842
rect 14140 2876 14222 2900
rect 14140 2842 14164 2876
rect 14198 2842 14222 2876
rect 14140 2818 14222 2842
rect 15158 2876 15240 2900
rect 15158 2842 15182 2876
rect 15216 2842 15240 2876
rect 15158 2818 15240 2842
rect 16176 2876 16258 2900
rect 16176 2842 16200 2876
rect 16234 2842 16258 2876
rect 16176 2818 16258 2842
rect 17194 2876 17276 2900
rect 17194 2842 17218 2876
rect 17252 2842 17276 2876
rect 19620 2844 19654 2860
rect 20638 3436 20672 3452
rect 20638 2844 20672 2860
rect 21656 3436 21690 3452
rect 21656 2844 21690 2860
rect 22674 3436 22708 3452
rect 22674 2844 22708 2860
rect 23692 3436 23726 3452
rect 23692 2844 23726 2860
rect 24710 3436 24744 3452
rect 24710 2844 24744 2860
rect 25728 3436 25762 3452
rect 25728 2844 25762 2860
rect 26746 3436 26780 3452
rect 26746 2844 26780 2860
rect 27764 3436 27798 3452
rect 27764 2844 27798 2860
rect 28782 3436 28816 3452
rect 28782 2844 28816 2860
rect 29800 3436 29834 3452
rect 29800 2844 29834 2860
rect 30818 3436 30852 3452
rect 30818 2844 30852 2860
rect 31836 3436 31870 3452
rect 31836 2844 31870 2860
rect 32854 3436 32888 3452
rect 32854 2844 32888 2860
rect 33872 3436 33906 3452
rect 33872 2844 33906 2860
rect 34890 3436 34924 3452
rect 34890 2844 34924 2860
rect 35908 3436 35942 3452
rect 35908 2844 35942 2860
rect 36926 3436 36960 3452
rect 36926 2844 36960 2860
rect 37944 3436 37978 3452
rect 37944 2844 37978 2860
rect 38962 3436 38996 3452
rect 38962 2844 38996 2860
rect 39980 3436 40014 3452
rect 39980 2844 40014 2860
rect 17194 2818 17276 2842
rect 28270 2810 28330 2812
rect 30314 2810 30374 2814
rect 33352 2810 33412 2814
rect 19852 2776 19868 2810
rect 20424 2776 20440 2810
rect 20870 2776 20886 2810
rect 21442 2776 21458 2810
rect 21888 2776 21904 2810
rect 22460 2776 22476 2810
rect 22906 2776 22922 2810
rect 23478 2776 23494 2810
rect 23924 2776 23940 2810
rect 24496 2776 24512 2810
rect 24942 2776 24958 2810
rect 25514 2776 25530 2810
rect 25960 2776 25976 2810
rect 26532 2776 26548 2810
rect 26978 2776 26994 2810
rect 27550 2776 27566 2810
rect 27996 2776 28012 2810
rect 28568 2776 28584 2810
rect 29014 2776 29030 2810
rect 29586 2776 29602 2810
rect 30032 2776 30048 2810
rect 30604 2776 30620 2810
rect 31050 2776 31066 2810
rect 31622 2776 31638 2810
rect 32068 2776 32084 2810
rect 32640 2776 32656 2810
rect 33086 2776 33102 2810
rect 33658 2776 33674 2810
rect 34104 2776 34120 2810
rect 34676 2776 34692 2810
rect 35122 2776 35138 2810
rect 35694 2776 35710 2810
rect 36140 2776 36156 2810
rect 36712 2776 36728 2810
rect 37158 2776 37174 2810
rect 37730 2776 37746 2810
rect 38176 2776 38192 2810
rect 38748 2776 38764 2810
rect 39194 2776 39210 2810
rect 39766 2776 39782 2810
rect 6764 2632 6780 2666
rect 7336 2632 7352 2666
rect 7782 2632 7798 2666
rect 8354 2632 8370 2666
rect 8800 2632 8816 2666
rect 9372 2632 9388 2666
rect 9818 2632 9834 2666
rect 10390 2632 10406 2666
rect 10836 2632 10852 2666
rect 11408 2632 11424 2666
rect 11854 2632 11870 2666
rect 12426 2632 12442 2666
rect 12872 2632 12888 2666
rect 13444 2632 13460 2666
rect 13890 2632 13906 2666
rect 14462 2632 14478 2666
rect 14908 2632 14924 2666
rect 15480 2632 15496 2666
rect 15926 2632 15942 2666
rect 16498 2632 16514 2666
rect 16944 2632 16960 2666
rect 17516 2632 17532 2666
rect 6532 2582 6566 2598
rect 6532 1990 6566 2006
rect 7550 2582 7584 2598
rect 7550 1990 7584 2006
rect 8568 2582 8602 2598
rect 8568 1990 8602 2006
rect 9586 2582 9620 2598
rect 9586 1990 9620 2006
rect 10604 2582 10638 2598
rect 10604 1990 10638 2006
rect 11622 2582 11656 2598
rect 11622 1990 11656 2006
rect 12640 2582 12674 2598
rect 12640 1990 12674 2006
rect 13658 2582 13692 2598
rect 13658 1990 13692 2006
rect 14676 2582 14710 2598
rect 14676 1990 14710 2006
rect 15694 2582 15728 2598
rect 15694 1990 15728 2006
rect 16712 2582 16746 2598
rect 16712 1990 16746 2006
rect 17730 2582 17764 2598
rect 20114 2560 20196 2584
rect 20114 2526 20138 2560
rect 20172 2526 20196 2560
rect 20114 2502 20196 2526
rect 21132 2560 21214 2584
rect 21132 2526 21156 2560
rect 21190 2526 21214 2560
rect 21132 2502 21214 2526
rect 22150 2560 22232 2584
rect 22150 2526 22174 2560
rect 22208 2526 22232 2560
rect 22150 2502 22232 2526
rect 23168 2560 23250 2584
rect 23168 2526 23192 2560
rect 23226 2526 23250 2560
rect 23168 2502 23250 2526
rect 24186 2560 24268 2584
rect 24186 2526 24210 2560
rect 24244 2526 24268 2560
rect 24186 2502 24268 2526
rect 25204 2560 25286 2584
rect 25204 2526 25228 2560
rect 25262 2526 25286 2560
rect 25204 2502 25286 2526
rect 26222 2560 26304 2584
rect 26222 2526 26246 2560
rect 26280 2526 26304 2560
rect 26222 2502 26304 2526
rect 27240 2560 27322 2584
rect 27240 2526 27264 2560
rect 27298 2526 27322 2560
rect 27240 2502 27322 2526
rect 28258 2560 28340 2584
rect 28258 2526 28282 2560
rect 28316 2526 28340 2560
rect 28258 2502 28340 2526
rect 29276 2560 29358 2584
rect 29276 2526 29300 2560
rect 29334 2526 29358 2560
rect 29276 2502 29358 2526
rect 30294 2560 30376 2584
rect 30294 2526 30318 2560
rect 30352 2526 30376 2560
rect 30294 2502 30376 2526
rect 31312 2560 31394 2584
rect 31312 2526 31336 2560
rect 31370 2526 31394 2560
rect 31312 2502 31394 2526
rect 32330 2560 32412 2584
rect 32330 2526 32354 2560
rect 32388 2526 32412 2560
rect 32330 2502 32412 2526
rect 33348 2560 33430 2584
rect 33348 2526 33372 2560
rect 33406 2526 33430 2560
rect 33348 2502 33430 2526
rect 34366 2560 34448 2584
rect 34366 2526 34390 2560
rect 34424 2526 34448 2560
rect 34366 2502 34448 2526
rect 35384 2560 35466 2584
rect 35384 2526 35408 2560
rect 35442 2526 35466 2560
rect 35384 2502 35466 2526
rect 36402 2560 36484 2584
rect 36402 2526 36426 2560
rect 36460 2526 36484 2560
rect 36402 2502 36484 2526
rect 37420 2560 37502 2584
rect 37420 2526 37444 2560
rect 37478 2526 37502 2560
rect 37420 2502 37502 2526
rect 38438 2560 38520 2584
rect 38438 2526 38462 2560
rect 38496 2526 38520 2560
rect 38438 2502 38520 2526
rect 39456 2560 39538 2584
rect 39456 2526 39480 2560
rect 39514 2526 39538 2560
rect 39456 2502 39538 2526
rect 19852 2254 19868 2288
rect 20424 2254 20440 2288
rect 20870 2254 20886 2288
rect 21442 2254 21458 2288
rect 21888 2254 21904 2288
rect 22460 2254 22476 2288
rect 22906 2254 22922 2288
rect 23478 2254 23494 2288
rect 23924 2254 23940 2288
rect 24496 2254 24512 2288
rect 24942 2254 24958 2288
rect 25514 2254 25530 2288
rect 25960 2254 25976 2288
rect 26532 2254 26548 2288
rect 26978 2254 26994 2288
rect 27550 2254 27566 2288
rect 27996 2254 28012 2288
rect 28568 2254 28584 2288
rect 29014 2254 29030 2288
rect 29586 2254 29602 2288
rect 30032 2254 30048 2288
rect 30604 2254 30620 2288
rect 31050 2254 31066 2288
rect 31622 2254 31638 2288
rect 32068 2254 32084 2288
rect 32640 2254 32656 2288
rect 33086 2254 33102 2288
rect 33658 2254 33674 2288
rect 34104 2254 34120 2288
rect 34676 2254 34692 2288
rect 35122 2254 35138 2288
rect 35694 2254 35710 2288
rect 36140 2254 36156 2288
rect 36712 2254 36728 2288
rect 37158 2254 37174 2288
rect 37730 2254 37746 2288
rect 38176 2254 38192 2288
rect 38748 2254 38764 2288
rect 39194 2254 39210 2288
rect 39766 2254 39782 2288
rect 23174 2252 23234 2254
rect 17730 1990 17764 2006
rect 19620 2204 19654 2220
rect 6764 1922 6780 1956
rect 7336 1922 7352 1956
rect 7782 1922 7798 1956
rect 8354 1922 8370 1956
rect 8800 1922 8816 1956
rect 9372 1922 9388 1956
rect 9818 1922 9834 1956
rect 10390 1922 10406 1956
rect 10836 1922 10852 1956
rect 11408 1922 11424 1956
rect 11854 1922 11870 1956
rect 12426 1922 12442 1956
rect 12872 1922 12888 1956
rect 13444 1922 13460 1956
rect 13890 1922 13906 1956
rect 14462 1922 14478 1956
rect 14908 1922 14924 1956
rect 15480 1922 15496 1956
rect 15926 1922 15942 1956
rect 16498 1922 16514 1956
rect 16944 1922 16960 1956
rect 17516 1922 17532 1956
rect 7014 1770 7096 1794
rect 7014 1736 7038 1770
rect 7072 1736 7096 1770
rect 7014 1712 7096 1736
rect 8032 1770 8114 1794
rect 8032 1736 8056 1770
rect 8090 1736 8114 1770
rect 8032 1712 8114 1736
rect 9050 1770 9132 1794
rect 9050 1736 9074 1770
rect 9108 1736 9132 1770
rect 9050 1712 9132 1736
rect 10068 1770 10150 1794
rect 10068 1736 10092 1770
rect 10126 1736 10150 1770
rect 10068 1712 10150 1736
rect 11086 1770 11168 1794
rect 11086 1736 11110 1770
rect 11144 1736 11168 1770
rect 11086 1712 11168 1736
rect 12104 1770 12186 1794
rect 12104 1736 12128 1770
rect 12162 1736 12186 1770
rect 12104 1712 12186 1736
rect 13122 1770 13204 1794
rect 13122 1736 13146 1770
rect 13180 1736 13204 1770
rect 13122 1712 13204 1736
rect 14140 1770 14222 1794
rect 14140 1736 14164 1770
rect 14198 1736 14222 1770
rect 14140 1712 14222 1736
rect 15158 1770 15240 1794
rect 15158 1736 15182 1770
rect 15216 1736 15240 1770
rect 15158 1712 15240 1736
rect 16176 1770 16258 1794
rect 16176 1736 16200 1770
rect 16234 1736 16258 1770
rect 16176 1712 16258 1736
rect 17194 1770 17276 1794
rect 17194 1736 17218 1770
rect 17252 1736 17276 1770
rect 17194 1712 17276 1736
rect 19620 1612 19654 1628
rect 20638 2204 20672 2220
rect 20638 1612 20672 1628
rect 21656 2204 21690 2220
rect 21656 1612 21690 1628
rect 22674 2204 22708 2220
rect 22674 1612 22708 1628
rect 23692 2204 23726 2220
rect 23692 1612 23726 1628
rect 24710 2204 24744 2220
rect 24710 1612 24744 1628
rect 25728 2204 25762 2220
rect 25728 1612 25762 1628
rect 26746 2204 26780 2220
rect 26746 1612 26780 1628
rect 27764 2204 27798 2220
rect 27764 1612 27798 1628
rect 28782 2204 28816 2220
rect 28782 1612 28816 1628
rect 29800 2204 29834 2220
rect 29800 1612 29834 1628
rect 30818 2204 30852 2220
rect 30818 1612 30852 1628
rect 31836 2204 31870 2220
rect 31836 1612 31870 1628
rect 32854 2204 32888 2220
rect 32854 1612 32888 1628
rect 33872 2204 33906 2220
rect 33872 1612 33906 1628
rect 34890 2204 34924 2220
rect 34890 1612 34924 1628
rect 35908 2204 35942 2220
rect 35908 1612 35942 1628
rect 36926 2204 36960 2220
rect 36926 1612 36960 1628
rect 37944 2204 37978 2220
rect 37944 1612 37978 1628
rect 38962 2204 38996 2220
rect 38962 1612 38996 1628
rect 39980 2204 40014 2220
rect 39980 1612 40014 1628
rect 27246 1578 27306 1588
rect 6764 1520 6780 1554
rect 7336 1520 7352 1554
rect 7782 1520 7798 1554
rect 8354 1520 8370 1554
rect 8800 1520 8816 1554
rect 9372 1520 9388 1554
rect 9818 1520 9834 1554
rect 10390 1520 10406 1554
rect 10836 1520 10852 1554
rect 11408 1520 11424 1554
rect 11854 1520 11870 1554
rect 12426 1520 12442 1554
rect 12872 1520 12888 1554
rect 13444 1520 13460 1554
rect 13890 1520 13906 1554
rect 14462 1520 14478 1554
rect 14908 1520 14924 1554
rect 15480 1520 15496 1554
rect 15926 1520 15942 1554
rect 16498 1520 16514 1554
rect 16944 1520 16960 1554
rect 17516 1520 17532 1554
rect 19852 1544 19868 1578
rect 20424 1544 20440 1578
rect 20870 1544 20886 1578
rect 21442 1544 21458 1578
rect 21888 1544 21904 1578
rect 22460 1544 22476 1578
rect 22906 1544 22922 1578
rect 23478 1544 23494 1578
rect 23924 1544 23940 1578
rect 24496 1544 24512 1578
rect 24942 1544 24958 1578
rect 25514 1544 25530 1578
rect 25960 1544 25976 1578
rect 26532 1544 26548 1578
rect 26978 1544 26994 1578
rect 27550 1544 27566 1578
rect 27996 1544 28012 1578
rect 28568 1544 28584 1578
rect 29014 1544 29030 1578
rect 29586 1544 29602 1578
rect 30032 1544 30048 1578
rect 30604 1544 30620 1578
rect 31050 1544 31066 1578
rect 31622 1544 31638 1578
rect 32068 1544 32084 1578
rect 32640 1544 32656 1578
rect 33086 1544 33102 1578
rect 33658 1544 33674 1578
rect 34104 1544 34120 1578
rect 34676 1544 34692 1578
rect 35122 1544 35138 1578
rect 35694 1544 35710 1578
rect 36140 1544 36156 1578
rect 36712 1544 36728 1578
rect 37158 1544 37174 1578
rect 37730 1544 37746 1578
rect 38176 1544 38192 1578
rect 38748 1544 38764 1578
rect 39194 1544 39210 1578
rect 39766 1544 39782 1578
rect 6532 1470 6566 1486
rect 6532 878 6566 894
rect 7550 1470 7584 1486
rect 7550 878 7584 894
rect 8568 1470 8602 1486
rect 8568 878 8602 894
rect 9586 1470 9620 1486
rect 9586 878 9620 894
rect 10604 1470 10638 1486
rect 10604 878 10638 894
rect 11622 1470 11656 1486
rect 11622 878 11656 894
rect 12640 1470 12674 1486
rect 12640 878 12674 894
rect 13658 1470 13692 1486
rect 13658 878 13692 894
rect 14676 1470 14710 1486
rect 14676 878 14710 894
rect 15694 1470 15728 1486
rect 15694 878 15728 894
rect 16712 1470 16746 1486
rect 16712 878 16746 894
rect 17730 1470 17764 1486
rect 20114 1324 20196 1348
rect 20114 1290 20138 1324
rect 20172 1290 20196 1324
rect 20114 1266 20196 1290
rect 21132 1324 21214 1348
rect 21132 1290 21156 1324
rect 21190 1290 21214 1324
rect 21132 1266 21214 1290
rect 22150 1324 22232 1348
rect 22150 1290 22174 1324
rect 22208 1290 22232 1324
rect 22150 1266 22232 1290
rect 23168 1324 23250 1348
rect 23168 1290 23192 1324
rect 23226 1290 23250 1324
rect 23168 1266 23250 1290
rect 24186 1324 24268 1348
rect 24186 1290 24210 1324
rect 24244 1290 24268 1324
rect 24186 1266 24268 1290
rect 25204 1324 25286 1348
rect 25204 1290 25228 1324
rect 25262 1290 25286 1324
rect 25204 1266 25286 1290
rect 26222 1324 26304 1348
rect 26222 1290 26246 1324
rect 26280 1290 26304 1324
rect 26222 1266 26304 1290
rect 27240 1324 27322 1348
rect 27240 1290 27264 1324
rect 27298 1290 27322 1324
rect 27240 1266 27322 1290
rect 28258 1324 28340 1348
rect 28258 1290 28282 1324
rect 28316 1290 28340 1324
rect 28258 1266 28340 1290
rect 29276 1324 29358 1348
rect 29276 1290 29300 1324
rect 29334 1290 29358 1324
rect 29276 1266 29358 1290
rect 30294 1324 30376 1348
rect 30294 1290 30318 1324
rect 30352 1290 30376 1324
rect 30294 1266 30376 1290
rect 31312 1324 31394 1348
rect 31312 1290 31336 1324
rect 31370 1290 31394 1324
rect 31312 1266 31394 1290
rect 32330 1324 32412 1348
rect 32330 1290 32354 1324
rect 32388 1290 32412 1324
rect 32330 1266 32412 1290
rect 33348 1324 33430 1348
rect 33348 1290 33372 1324
rect 33406 1290 33430 1324
rect 33348 1266 33430 1290
rect 34366 1324 34448 1348
rect 34366 1290 34390 1324
rect 34424 1290 34448 1324
rect 34366 1266 34448 1290
rect 35384 1324 35466 1348
rect 35384 1290 35408 1324
rect 35442 1290 35466 1324
rect 35384 1266 35466 1290
rect 36402 1324 36484 1348
rect 36402 1290 36426 1324
rect 36460 1290 36484 1324
rect 36402 1266 36484 1290
rect 37420 1324 37502 1348
rect 37420 1290 37444 1324
rect 37478 1290 37502 1324
rect 37420 1266 37502 1290
rect 38438 1324 38520 1348
rect 38438 1290 38462 1324
rect 38496 1290 38520 1324
rect 38438 1266 38520 1290
rect 39456 1324 39538 1348
rect 39456 1290 39480 1324
rect 39514 1290 39538 1324
rect 39456 1266 39538 1290
rect 19852 1020 19868 1054
rect 20424 1020 20440 1054
rect 20870 1020 20886 1054
rect 21442 1020 21458 1054
rect 21888 1020 21904 1054
rect 22460 1020 22476 1054
rect 22906 1020 22922 1054
rect 23478 1020 23494 1054
rect 23924 1020 23940 1054
rect 24496 1020 24512 1054
rect 24942 1020 24958 1054
rect 25514 1020 25530 1054
rect 25960 1020 25976 1054
rect 26532 1020 26548 1054
rect 26978 1020 26994 1054
rect 27550 1020 27566 1054
rect 27996 1020 28012 1054
rect 28568 1020 28584 1054
rect 29014 1020 29030 1054
rect 29586 1020 29602 1054
rect 30032 1020 30048 1054
rect 30604 1020 30620 1054
rect 31050 1020 31066 1054
rect 31622 1020 31638 1054
rect 32068 1020 32084 1054
rect 32640 1020 32656 1054
rect 33086 1020 33102 1054
rect 33658 1020 33674 1054
rect 34104 1020 34120 1054
rect 34676 1020 34692 1054
rect 35122 1020 35138 1054
rect 35694 1020 35710 1054
rect 36140 1020 36156 1054
rect 36712 1020 36728 1054
rect 37158 1020 37174 1054
rect 37730 1020 37746 1054
rect 38176 1020 38192 1054
rect 38748 1020 38764 1054
rect 39194 1020 39210 1054
rect 39766 1020 39782 1054
rect 23160 1018 23220 1020
rect 17730 878 17764 894
rect 19620 970 19654 986
rect 6764 810 6780 844
rect 7336 810 7352 844
rect 7782 810 7798 844
rect 8354 810 8370 844
rect 8800 810 8816 844
rect 9372 810 9388 844
rect 9818 810 9834 844
rect 10390 810 10406 844
rect 10836 810 10852 844
rect 11408 810 11424 844
rect 11854 810 11870 844
rect 12426 810 12442 844
rect 12872 810 12888 844
rect 13444 810 13460 844
rect 13890 810 13906 844
rect 14462 810 14478 844
rect 14908 810 14924 844
rect 15480 810 15496 844
rect 15926 810 15942 844
rect 16498 810 16514 844
rect 16944 810 16960 844
rect 17516 810 17532 844
rect 7014 428 7096 452
rect 7014 394 7038 428
rect 7072 394 7096 428
rect 7014 370 7096 394
rect 8032 428 8114 452
rect 8032 394 8056 428
rect 8090 394 8114 428
rect 8032 370 8114 394
rect 9050 428 9132 452
rect 9050 394 9074 428
rect 9108 394 9132 428
rect 9050 370 9132 394
rect 10068 428 10150 452
rect 10068 394 10092 428
rect 10126 394 10150 428
rect 10068 370 10150 394
rect 11086 428 11168 452
rect 11086 394 11110 428
rect 11144 394 11168 428
rect 11086 370 11168 394
rect 12104 428 12186 452
rect 12104 394 12128 428
rect 12162 394 12186 428
rect 12104 370 12186 394
rect 13122 428 13204 452
rect 13122 394 13146 428
rect 13180 394 13204 428
rect 13122 370 13204 394
rect 14140 428 14222 452
rect 14140 394 14164 428
rect 14198 394 14222 428
rect 14140 370 14222 394
rect 15158 428 15240 452
rect 15158 394 15182 428
rect 15216 394 15240 428
rect 15158 370 15240 394
rect 16176 428 16258 452
rect 16176 394 16200 428
rect 16234 394 16258 428
rect 16176 370 16258 394
rect 17194 428 17276 452
rect 17194 394 17218 428
rect 17252 394 17276 428
rect 17194 370 17276 394
rect 19620 378 19654 394
rect 20638 970 20672 986
rect 20638 378 20672 394
rect 21656 970 21690 986
rect 21656 378 21690 394
rect 22674 970 22708 986
rect 22674 378 22708 394
rect 23692 970 23726 986
rect 23692 378 23726 394
rect 24710 970 24744 986
rect 24710 378 24744 394
rect 25728 970 25762 986
rect 25728 378 25762 394
rect 26746 970 26780 986
rect 26746 378 26780 394
rect 27764 970 27798 986
rect 27764 378 27798 394
rect 28782 970 28816 986
rect 28782 378 28816 394
rect 29800 970 29834 986
rect 29800 378 29834 394
rect 30818 970 30852 986
rect 30818 378 30852 394
rect 31836 970 31870 986
rect 31836 378 31870 394
rect 32854 970 32888 986
rect 32854 378 32888 394
rect 33872 970 33906 986
rect 33872 378 33906 394
rect 34890 970 34924 986
rect 34890 378 34924 394
rect 35908 970 35942 986
rect 35908 378 35942 394
rect 36926 970 36960 986
rect 36926 378 36960 394
rect 37944 970 37978 986
rect 37944 378 37978 394
rect 38962 970 38996 986
rect 38962 378 38996 394
rect 39980 970 40014 986
rect 39980 378 40014 394
rect 21128 344 21188 346
rect 27240 344 27300 346
rect 29274 344 29334 346
rect 33340 344 33400 350
rect 37416 344 37476 346
rect 38432 344 38492 346
rect 19852 310 19868 344
rect 20424 310 20440 344
rect 20870 310 20886 344
rect 21442 310 21458 344
rect 21888 310 21904 344
rect 22460 310 22476 344
rect 22906 310 22922 344
rect 23478 310 23494 344
rect 23924 310 23940 344
rect 24496 310 24512 344
rect 24942 310 24958 344
rect 25514 310 25530 344
rect 25960 310 25976 344
rect 26532 310 26548 344
rect 26978 310 26994 344
rect 27550 310 27566 344
rect 27996 310 28012 344
rect 28568 310 28584 344
rect 29014 310 29030 344
rect 29586 310 29602 344
rect 30032 310 30048 344
rect 30604 310 30620 344
rect 31050 310 31066 344
rect 31622 310 31638 344
rect 32068 310 32084 344
rect 32640 310 32656 344
rect 33086 310 33102 344
rect 33658 310 33674 344
rect 34104 310 34120 344
rect 34676 310 34692 344
rect 35122 310 35138 344
rect 35694 310 35710 344
rect 36140 310 36156 344
rect 36712 310 36728 344
rect 37158 310 37174 344
rect 37730 310 37746 344
rect 38176 310 38192 344
rect 38748 310 38764 344
rect 39194 310 39210 344
rect 39766 310 39782 344
rect 20126 78 20208 102
rect 20126 44 20150 78
rect 20184 44 20208 78
rect 20126 20 20208 44
rect 21144 78 21226 102
rect 21144 44 21168 78
rect 21202 44 21226 78
rect 21144 20 21226 44
rect 22162 78 22244 102
rect 22162 44 22186 78
rect 22220 44 22244 78
rect 22162 20 22244 44
rect 23180 78 23262 102
rect 23180 44 23204 78
rect 23238 44 23262 78
rect 23180 20 23262 44
rect 24198 78 24280 102
rect 24198 44 24222 78
rect 24256 44 24280 78
rect 24198 20 24280 44
rect 25216 78 25298 102
rect 25216 44 25240 78
rect 25274 44 25298 78
rect 25216 20 25298 44
rect 26234 78 26316 102
rect 26234 44 26258 78
rect 26292 44 26316 78
rect 26234 20 26316 44
rect 27252 78 27334 102
rect 27252 44 27276 78
rect 27310 44 27334 78
rect 27252 20 27334 44
rect 28270 78 28352 102
rect 28270 44 28294 78
rect 28328 44 28352 78
rect 28270 20 28352 44
rect 29288 78 29370 102
rect 29288 44 29312 78
rect 29346 44 29370 78
rect 29288 20 29370 44
rect 30306 78 30388 102
rect 30306 44 30330 78
rect 30364 44 30388 78
rect 30306 20 30388 44
rect 31324 78 31406 102
rect 31324 44 31348 78
rect 31382 44 31406 78
rect 31324 20 31406 44
rect 32342 78 32424 102
rect 32342 44 32366 78
rect 32400 44 32424 78
rect 32342 20 32424 44
rect 33360 78 33442 102
rect 33360 44 33384 78
rect 33418 44 33442 78
rect 33360 20 33442 44
rect 34378 78 34460 102
rect 34378 44 34402 78
rect 34436 44 34460 78
rect 34378 20 34460 44
rect 35396 78 35478 102
rect 35396 44 35420 78
rect 35454 44 35478 78
rect 35396 20 35478 44
rect 36414 78 36496 102
rect 36414 44 36438 78
rect 36472 44 36496 78
rect 36414 20 36496 44
rect 37432 78 37514 102
rect 37432 44 37456 78
rect 37490 44 37514 78
rect 37432 20 37514 44
rect 38450 78 38532 102
rect 38450 44 38474 78
rect 38508 44 38532 78
rect 38450 20 38532 44
rect 39468 78 39550 102
rect 39468 44 39492 78
rect 39526 44 39550 78
rect 39468 20 39550 44
rect 7222 -22 7238 12
rect 7794 -22 7810 12
rect 8240 -22 8256 12
rect 8812 -22 8828 12
rect 9258 -22 9274 12
rect 9830 -22 9846 12
rect 10276 -22 10292 12
rect 10848 -22 10864 12
rect 11294 -22 11310 12
rect 11866 -22 11882 12
rect 12312 -22 12328 12
rect 12884 -22 12900 12
rect 13330 -22 13346 12
rect 13902 -22 13918 12
rect 14348 -22 14364 12
rect 14920 -22 14936 12
rect 15366 -22 15382 12
rect 15938 -22 15954 12
rect 16384 -22 16400 12
rect 16956 -22 16972 12
rect 6990 -72 7024 -56
rect 6990 -664 7024 -648
rect 8008 -72 8042 -56
rect 8008 -664 8042 -648
rect 9026 -72 9060 -56
rect 9026 -664 9060 -648
rect 10044 -72 10078 -56
rect 10044 -664 10078 -648
rect 11062 -72 11096 -56
rect 11062 -664 11096 -648
rect 12080 -72 12114 -56
rect 12080 -664 12114 -648
rect 13098 -72 13132 -56
rect 13098 -664 13132 -648
rect 14116 -72 14150 -56
rect 14116 -664 14150 -648
rect 15134 -72 15168 -56
rect 15134 -664 15168 -648
rect 16152 -72 16186 -56
rect 16152 -664 16186 -648
rect 17170 -72 17204 -56
rect 19852 -212 19868 -178
rect 20424 -212 20440 -178
rect 20870 -212 20886 -178
rect 21442 -212 21458 -178
rect 21888 -212 21904 -178
rect 22460 -212 22476 -178
rect 22906 -212 22922 -178
rect 23478 -212 23494 -178
rect 23924 -212 23940 -178
rect 24496 -212 24512 -178
rect 24942 -212 24958 -178
rect 25514 -212 25530 -178
rect 25960 -212 25976 -178
rect 26532 -212 26548 -178
rect 26978 -212 26994 -178
rect 27550 -212 27566 -178
rect 27996 -212 28012 -178
rect 28568 -212 28584 -178
rect 29014 -212 29030 -178
rect 29586 -212 29602 -178
rect 30032 -212 30048 -178
rect 30604 -212 30620 -178
rect 31050 -212 31066 -178
rect 31622 -212 31638 -178
rect 32068 -212 32084 -178
rect 32640 -212 32656 -178
rect 33086 -212 33102 -178
rect 33658 -212 33674 -178
rect 34104 -212 34120 -178
rect 34676 -212 34692 -178
rect 35122 -212 35138 -178
rect 35694 -212 35710 -178
rect 36140 -212 36156 -178
rect 36712 -212 36728 -178
rect 37158 -212 37174 -178
rect 37730 -212 37746 -178
rect 38176 -212 38192 -178
rect 38748 -212 38764 -178
rect 39194 -212 39210 -178
rect 39766 -212 39782 -178
rect 17170 -664 17204 -648
rect 19620 -262 19654 -246
rect 7222 -732 7238 -698
rect 7794 -732 7810 -698
rect 8240 -732 8256 -698
rect 8812 -732 8828 -698
rect 9258 -732 9274 -698
rect 9830 -732 9846 -698
rect 10276 -732 10292 -698
rect 10848 -732 10864 -698
rect 11294 -732 11310 -698
rect 11866 -732 11882 -698
rect 12312 -732 12328 -698
rect 12884 -732 12900 -698
rect 13330 -732 13346 -698
rect 13902 -732 13918 -698
rect 14348 -732 14364 -698
rect 14920 -732 14936 -698
rect 15366 -732 15382 -698
rect 15938 -732 15954 -698
rect 16384 -732 16400 -698
rect 16956 -732 16972 -698
rect 19620 -854 19654 -838
rect 20638 -262 20672 -246
rect 20638 -854 20672 -838
rect 21656 -262 21690 -246
rect 21656 -854 21690 -838
rect 22674 -262 22708 -246
rect 22674 -854 22708 -838
rect 23692 -262 23726 -246
rect 23692 -854 23726 -838
rect 24710 -262 24744 -246
rect 24710 -854 24744 -838
rect 25728 -262 25762 -246
rect 25728 -854 25762 -838
rect 26746 -262 26780 -246
rect 26746 -854 26780 -838
rect 27764 -262 27798 -246
rect 27764 -854 27798 -838
rect 28782 -262 28816 -246
rect 28782 -854 28816 -838
rect 29800 -262 29834 -246
rect 29800 -854 29834 -838
rect 30818 -262 30852 -246
rect 30818 -854 30852 -838
rect 31836 -262 31870 -246
rect 31836 -854 31870 -838
rect 32854 -262 32888 -246
rect 32854 -854 32888 -838
rect 33872 -262 33906 -246
rect 33872 -854 33906 -838
rect 34890 -262 34924 -246
rect 34890 -854 34924 -838
rect 35908 -262 35942 -246
rect 35908 -854 35942 -838
rect 36926 -262 36960 -246
rect 36926 -854 36960 -838
rect 37944 -262 37978 -246
rect 37944 -854 37978 -838
rect 38962 -262 38996 -246
rect 38962 -854 38996 -838
rect 39980 -262 40014 -246
rect 39980 -854 40014 -838
rect 19852 -922 19868 -888
rect 20424 -922 20440 -888
rect 20870 -922 20886 -888
rect 21442 -922 21458 -888
rect 21888 -922 21904 -888
rect 22460 -922 22476 -888
rect 22906 -922 22922 -888
rect 23478 -922 23494 -888
rect 23924 -922 23940 -888
rect 24496 -922 24512 -888
rect 24942 -922 24958 -888
rect 25514 -922 25530 -888
rect 25960 -922 25976 -888
rect 26532 -922 26548 -888
rect 26978 -922 26994 -888
rect 27550 -922 27566 -888
rect 27996 -922 28012 -888
rect 28568 -922 28584 -888
rect 29014 -922 29030 -888
rect 29586 -922 29602 -888
rect 30032 -922 30048 -888
rect 30604 -922 30620 -888
rect 31050 -922 31066 -888
rect 31622 -922 31638 -888
rect 32068 -922 32084 -888
rect 32640 -922 32656 -888
rect 33086 -922 33102 -888
rect 33658 -922 33674 -888
rect 34104 -922 34120 -888
rect 34676 -922 34692 -888
rect 35122 -922 35138 -888
rect 35694 -922 35710 -888
rect 36140 -922 36156 -888
rect 36712 -922 36728 -888
rect 37158 -922 37174 -888
rect 37730 -922 37746 -888
rect 38176 -922 38192 -888
rect 38748 -922 38764 -888
rect 39194 -922 39210 -888
rect 39766 -922 39782 -888
rect 6824 -1018 6906 -994
rect 6824 -1052 6848 -1018
rect 6882 -1052 6906 -1018
rect 6824 -1076 6906 -1052
rect 7842 -1018 7924 -994
rect 7842 -1052 7866 -1018
rect 7900 -1052 7924 -1018
rect 7842 -1076 7924 -1052
rect 8860 -1018 8942 -994
rect 8860 -1052 8884 -1018
rect 8918 -1052 8942 -1018
rect 8860 -1076 8942 -1052
rect 9878 -1018 9960 -994
rect 9878 -1052 9902 -1018
rect 9936 -1052 9960 -1018
rect 9878 -1076 9960 -1052
rect 10896 -1018 10978 -994
rect 10896 -1052 10920 -1018
rect 10954 -1052 10978 -1018
rect 10896 -1076 10978 -1052
rect 11914 -1018 11996 -994
rect 11914 -1052 11938 -1018
rect 11972 -1052 11996 -1018
rect 11914 -1076 11996 -1052
rect 12932 -1018 13014 -994
rect 12932 -1052 12956 -1018
rect 12990 -1052 13014 -1018
rect 12932 -1076 13014 -1052
rect 13950 -1018 14032 -994
rect 13950 -1052 13974 -1018
rect 14008 -1052 14032 -1018
rect 13950 -1076 14032 -1052
rect 14968 -1018 15050 -994
rect 14968 -1052 14992 -1018
rect 15026 -1052 15050 -1018
rect 14968 -1076 15050 -1052
rect 15986 -1018 16068 -994
rect 15986 -1052 16010 -1018
rect 16044 -1052 16068 -1018
rect 15986 -1076 16068 -1052
rect 17004 -1018 17086 -994
rect 17004 -1052 17028 -1018
rect 17062 -1052 17086 -1018
rect 17004 -1076 17086 -1052
rect 20114 -1100 20196 -1076
rect 20114 -1134 20138 -1100
rect 20172 -1134 20196 -1100
rect 20114 -1158 20196 -1134
rect 21132 -1100 21214 -1076
rect 21132 -1134 21156 -1100
rect 21190 -1134 21214 -1100
rect 21132 -1158 21214 -1134
rect 22150 -1100 22232 -1076
rect 22150 -1134 22174 -1100
rect 22208 -1134 22232 -1100
rect 22150 -1158 22232 -1134
rect 23168 -1100 23250 -1076
rect 23168 -1134 23192 -1100
rect 23226 -1134 23250 -1100
rect 23168 -1158 23250 -1134
rect 24186 -1100 24268 -1076
rect 24186 -1134 24210 -1100
rect 24244 -1134 24268 -1100
rect 24186 -1158 24268 -1134
rect 25204 -1100 25286 -1076
rect 25204 -1134 25228 -1100
rect 25262 -1134 25286 -1100
rect 25204 -1158 25286 -1134
rect 26222 -1100 26304 -1076
rect 26222 -1134 26246 -1100
rect 26280 -1134 26304 -1100
rect 26222 -1158 26304 -1134
rect 27240 -1100 27322 -1076
rect 27240 -1134 27264 -1100
rect 27298 -1134 27322 -1100
rect 27240 -1158 27322 -1134
rect 28258 -1100 28340 -1076
rect 28258 -1134 28282 -1100
rect 28316 -1134 28340 -1100
rect 28258 -1158 28340 -1134
rect 29276 -1100 29358 -1076
rect 29276 -1134 29300 -1100
rect 29334 -1134 29358 -1100
rect 29276 -1158 29358 -1134
rect 30294 -1100 30376 -1076
rect 30294 -1134 30318 -1100
rect 30352 -1134 30376 -1100
rect 30294 -1158 30376 -1134
rect 31312 -1100 31394 -1076
rect 31312 -1134 31336 -1100
rect 31370 -1134 31394 -1100
rect 31312 -1158 31394 -1134
rect 32330 -1100 32412 -1076
rect 32330 -1134 32354 -1100
rect 32388 -1134 32412 -1100
rect 32330 -1158 32412 -1134
rect 33348 -1100 33430 -1076
rect 33348 -1134 33372 -1100
rect 33406 -1134 33430 -1100
rect 33348 -1158 33430 -1134
rect 34366 -1100 34448 -1076
rect 34366 -1134 34390 -1100
rect 34424 -1134 34448 -1100
rect 34366 -1158 34448 -1134
rect 35384 -1100 35466 -1076
rect 35384 -1134 35408 -1100
rect 35442 -1134 35466 -1100
rect 35384 -1158 35466 -1134
rect 36402 -1100 36484 -1076
rect 36402 -1134 36426 -1100
rect 36460 -1134 36484 -1100
rect 36402 -1158 36484 -1134
rect 37420 -1100 37502 -1076
rect 37420 -1134 37444 -1100
rect 37478 -1134 37502 -1100
rect 37420 -1158 37502 -1134
rect 38438 -1100 38520 -1076
rect 38438 -1134 38462 -1100
rect 38496 -1134 38520 -1100
rect 38438 -1158 38520 -1134
rect 39456 -1100 39538 -1076
rect 39456 -1134 39480 -1100
rect 39514 -1134 39538 -1100
rect 39456 -1158 39538 -1134
rect 4718 -2142 4818 -1980
rect 41862 -2142 41962 -1980
<< viali >>
rect 17518 29302 17580 29402
rect 17580 29302 41700 29402
rect 41700 29302 41762 29402
rect 17418 15352 17518 28782
rect 23822 26601 24286 26635
rect 24840 26601 25304 26635
rect 25858 26601 26322 26635
rect 26876 26601 27340 26635
rect 27894 26601 28358 26635
rect 28912 26601 29376 26635
rect 29930 26601 30394 26635
rect 30948 26601 31412 26635
rect 31966 26601 32430 26635
rect 32984 26601 33448 26635
rect 34002 26601 34466 26635
rect 35020 26601 35484 26635
rect 36038 26601 36502 26635
rect 37056 26601 37520 26635
rect 38074 26601 38538 26635
rect 39092 26601 39556 26635
rect 23528 25966 23562 26542
rect 24546 25966 24580 26542
rect 25564 25966 25598 26542
rect 26582 25966 26616 26542
rect 27600 25966 27634 26542
rect 28618 25966 28652 26542
rect 29636 25966 29670 26542
rect 30654 25966 30688 26542
rect 31672 25966 31706 26542
rect 32690 25966 32724 26542
rect 33708 25966 33742 26542
rect 34726 25966 34760 26542
rect 35744 25966 35778 26542
rect 36762 25966 36796 26542
rect 37780 25966 37814 26542
rect 38798 25966 38832 26542
rect 39816 25966 39850 26542
rect 23822 25873 24286 25907
rect 24840 25873 25304 25907
rect 25858 25873 26322 25907
rect 26876 25873 27340 25907
rect 27894 25873 28358 25907
rect 28912 25873 29376 25907
rect 29930 25873 30394 25907
rect 30948 25873 31412 25907
rect 31966 25873 32430 25907
rect 32984 25873 33448 25907
rect 34002 25873 34466 25907
rect 35020 25873 35484 25907
rect 36038 25873 36502 25907
rect 37056 25873 37520 25907
rect 38074 25873 38538 25907
rect 39092 25873 39556 25907
rect 23822 25465 24286 25499
rect 24840 25465 25304 25499
rect 25858 25465 26322 25499
rect 26876 25465 27340 25499
rect 27894 25465 28358 25499
rect 28912 25465 29376 25499
rect 29930 25465 30394 25499
rect 30948 25465 31412 25499
rect 31966 25465 32430 25499
rect 32984 25465 33448 25499
rect 34002 25465 34466 25499
rect 35020 25465 35484 25499
rect 36038 25465 36502 25499
rect 37056 25465 37520 25499
rect 38074 25465 38538 25499
rect 39092 25465 39556 25499
rect 23528 24830 23562 25406
rect 24546 24830 24580 25406
rect 25564 24830 25598 25406
rect 26582 24830 26616 25406
rect 27600 24830 27634 25406
rect 28618 24830 28652 25406
rect 29636 24830 29670 25406
rect 30654 24830 30688 25406
rect 31672 24830 31706 25406
rect 32690 24830 32724 25406
rect 33708 24830 33742 25406
rect 34726 24830 34760 25406
rect 35744 24830 35778 25406
rect 36762 24830 36796 25406
rect 37780 24830 37814 25406
rect 38798 24830 38832 25406
rect 39816 24830 39850 25406
rect 23822 24737 24286 24771
rect 24840 24737 25304 24771
rect 25858 24737 26322 24771
rect 26876 24737 27340 24771
rect 27894 24737 28358 24771
rect 28912 24737 29376 24771
rect 29930 24737 30394 24771
rect 30948 24737 31412 24771
rect 31966 24737 32430 24771
rect 32984 24737 33448 24771
rect 34002 24737 34466 24771
rect 35020 24737 35484 24771
rect 36038 24737 36502 24771
rect 37056 24737 37520 24771
rect 38074 24737 38538 24771
rect 39092 24737 39556 24771
rect 23822 24329 24286 24363
rect 24840 24329 25304 24363
rect 25858 24329 26322 24363
rect 26876 24329 27340 24363
rect 27894 24329 28358 24363
rect 28912 24329 29376 24363
rect 29930 24329 30394 24363
rect 30948 24329 31412 24363
rect 31966 24329 32430 24363
rect 32984 24329 33448 24363
rect 34002 24329 34466 24363
rect 35020 24329 35484 24363
rect 36038 24329 36502 24363
rect 37056 24329 37520 24363
rect 38074 24329 38538 24363
rect 39092 24329 39556 24363
rect 23528 23694 23562 24270
rect 24546 23694 24580 24270
rect 25564 23694 25598 24270
rect 26582 23694 26616 24270
rect 27600 23694 27634 24270
rect 28618 23694 28652 24270
rect 29636 23694 29670 24270
rect 30654 23694 30688 24270
rect 31672 23694 31706 24270
rect 32690 23694 32724 24270
rect 33708 23694 33742 24270
rect 34726 23694 34760 24270
rect 35744 23694 35778 24270
rect 36762 23694 36796 24270
rect 37780 23694 37814 24270
rect 38798 23694 38832 24270
rect 39816 23694 39850 24270
rect 23822 23601 24286 23635
rect 24840 23601 25304 23635
rect 25858 23601 26322 23635
rect 26876 23601 27340 23635
rect 27894 23601 28358 23635
rect 28912 23601 29376 23635
rect 29930 23601 30394 23635
rect 30948 23601 31412 23635
rect 31966 23601 32430 23635
rect 32984 23601 33448 23635
rect 34002 23601 34466 23635
rect 35020 23601 35484 23635
rect 36038 23601 36502 23635
rect 37056 23601 37520 23635
rect 38074 23601 38538 23635
rect 39092 23601 39556 23635
rect 25016 22691 25480 22725
rect 26034 22691 26498 22725
rect 27052 22691 27516 22725
rect 28070 22691 28534 22725
rect 29088 22691 29552 22725
rect 30106 22691 30570 22725
rect 31124 22691 31588 22725
rect 32142 22691 32606 22725
rect 33160 22691 33624 22725
rect 34178 22691 34642 22725
rect 35196 22691 35660 22725
rect 36214 22691 36678 22725
rect 37232 22691 37696 22725
rect 38250 22691 38714 22725
rect 24722 22056 24756 22632
rect 25740 22056 25774 22632
rect 26758 22056 26792 22632
rect 27776 22056 27810 22632
rect 28794 22056 28828 22632
rect 29812 22056 29846 22632
rect 30830 22056 30864 22632
rect 31848 22056 31882 22632
rect 32866 22056 32900 22632
rect 33884 22056 33918 22632
rect 34902 22056 34936 22632
rect 35920 22056 35954 22632
rect 36938 22056 36972 22632
rect 37956 22056 37990 22632
rect 38974 22056 39008 22632
rect 25016 21963 25480 21997
rect 26034 21963 26498 21997
rect 27052 21963 27516 21997
rect 28070 21963 28534 21997
rect 29088 21963 29552 21997
rect 30106 21963 30570 21997
rect 31124 21963 31588 21997
rect 32142 21963 32606 21997
rect 33160 21963 33624 21997
rect 34178 21963 34642 21997
rect 35196 21963 35660 21997
rect 36214 21963 36678 21997
rect 37232 21963 37696 21997
rect 38250 21963 38714 21997
rect 25016 21659 25480 21693
rect 26034 21659 26498 21693
rect 27052 21659 27516 21693
rect 28070 21659 28534 21693
rect 29088 21659 29552 21693
rect 30106 21659 30570 21693
rect 31124 21659 31588 21693
rect 32142 21659 32606 21693
rect 33160 21659 33624 21693
rect 34178 21659 34642 21693
rect 35196 21659 35660 21693
rect 36214 21659 36678 21693
rect 37232 21659 37696 21693
rect 38250 21659 38714 21693
rect 24722 21024 24756 21600
rect 25740 21024 25774 21600
rect 26758 21024 26792 21600
rect 27776 21024 27810 21600
rect 28794 21024 28828 21600
rect 29812 21024 29846 21600
rect 30830 21024 30864 21600
rect 31848 21024 31882 21600
rect 32866 21024 32900 21600
rect 33884 21024 33918 21600
rect 34902 21024 34936 21600
rect 35920 21024 35954 21600
rect 36938 21024 36972 21600
rect 37956 21024 37990 21600
rect 38974 21024 39008 21600
rect 25016 20931 25480 20965
rect 26034 20931 26498 20965
rect 27052 20931 27516 20965
rect 28070 20931 28534 20965
rect 29088 20931 29552 20965
rect 30106 20931 30570 20965
rect 31124 20931 31588 20965
rect 32142 20931 32606 20965
rect 33160 20931 33624 20965
rect 34178 20931 34642 20965
rect 35196 20931 35660 20965
rect 36214 20931 36678 20965
rect 37232 20931 37696 20965
rect 38250 20931 38714 20965
rect 24808 20055 25272 20089
rect 25826 20055 26290 20089
rect 26844 20055 27308 20089
rect 27862 20055 28326 20089
rect 28880 20055 29344 20089
rect 29898 20055 30362 20089
rect 30916 20055 31380 20089
rect 31934 20055 32398 20089
rect 32952 20055 33416 20089
rect 33970 20055 34434 20089
rect 34988 20055 35452 20089
rect 36006 20055 36470 20089
rect 37024 20055 37488 20089
rect 38042 20055 38506 20089
rect 39060 20055 39524 20089
rect 19504 19951 19968 19985
rect 20522 19951 20986 19985
rect 21540 19951 22004 19985
rect 22558 19951 23022 19985
rect 19210 19316 19244 19892
rect 20228 19316 20262 19892
rect 21246 19316 21280 19892
rect 22264 19316 22298 19892
rect 23282 19316 23316 19892
rect 24514 19420 24548 19996
rect 25532 19420 25566 19996
rect 26550 19420 26584 19996
rect 27568 19420 27602 19996
rect 28586 19420 28620 19996
rect 29604 19420 29638 19996
rect 30622 19420 30656 19996
rect 31640 19420 31674 19996
rect 32658 19420 32692 19996
rect 33676 19420 33710 19996
rect 34694 19420 34728 19996
rect 35712 19420 35746 19996
rect 36730 19420 36764 19996
rect 37748 19420 37782 19996
rect 38766 19420 38800 19996
rect 39784 19420 39818 19996
rect 24808 19327 25272 19361
rect 25826 19327 26290 19361
rect 26844 19327 27308 19361
rect 27862 19327 28326 19361
rect 28880 19327 29344 19361
rect 29898 19327 30362 19361
rect 30916 19327 31380 19361
rect 31934 19327 32398 19361
rect 32952 19327 33416 19361
rect 33970 19327 34434 19361
rect 34988 19327 35452 19361
rect 36006 19327 36470 19361
rect 37024 19327 37488 19361
rect 38042 19327 38506 19361
rect 39060 19327 39524 19361
rect 19504 19223 19968 19257
rect 20522 19223 20986 19257
rect 21540 19223 22004 19257
rect 22558 19223 23022 19257
rect 19504 18919 19968 18953
rect 20522 18919 20986 18953
rect 21540 18919 22004 18953
rect 22558 18919 23022 18953
rect 19210 18284 19244 18860
rect 20228 18284 20262 18860
rect 21246 18284 21280 18860
rect 22264 18284 22298 18860
rect 23282 18284 23316 18860
rect 24808 18799 25272 18833
rect 25826 18799 26290 18833
rect 26844 18799 27308 18833
rect 27862 18799 28326 18833
rect 28880 18799 29344 18833
rect 29898 18799 30362 18833
rect 30916 18799 31380 18833
rect 31934 18799 32398 18833
rect 32952 18799 33416 18833
rect 33970 18799 34434 18833
rect 34988 18799 35452 18833
rect 36006 18799 36470 18833
rect 37024 18799 37488 18833
rect 38042 18799 38506 18833
rect 39060 18799 39524 18833
rect 19504 18191 19968 18225
rect 20522 18191 20986 18225
rect 21540 18191 22004 18225
rect 22558 18191 23022 18225
rect 24514 18164 24548 18740
rect 25532 18164 25566 18740
rect 26550 18164 26584 18740
rect 27568 18164 27602 18740
rect 28586 18164 28620 18740
rect 29604 18164 29638 18740
rect 30622 18164 30656 18740
rect 31640 18164 31674 18740
rect 32658 18164 32692 18740
rect 33676 18164 33710 18740
rect 34694 18164 34728 18740
rect 35712 18164 35746 18740
rect 36730 18164 36764 18740
rect 37748 18164 37782 18740
rect 38766 18164 38800 18740
rect 39784 18164 39818 18740
rect 24808 18071 25272 18105
rect 25826 18071 26290 18105
rect 26844 18071 27308 18105
rect 27862 18071 28326 18105
rect 28880 18071 29344 18105
rect 29898 18071 30362 18105
rect 30916 18071 31380 18105
rect 31934 18071 32398 18105
rect 32952 18071 33416 18105
rect 33970 18071 34434 18105
rect 34988 18071 35452 18105
rect 36006 18071 36470 18105
rect 37024 18071 37488 18105
rect 38042 18071 38506 18105
rect 39060 18071 39524 18105
rect 19504 17887 19968 17921
rect 20522 17887 20986 17921
rect 21540 17887 22004 17921
rect 22558 17887 23022 17921
rect 19210 17252 19244 17828
rect 20228 17252 20262 17828
rect 21246 17252 21280 17828
rect 22264 17252 22298 17828
rect 23282 17252 23316 17828
rect 24808 17543 25272 17577
rect 25826 17543 26290 17577
rect 26844 17543 27308 17577
rect 27862 17543 28326 17577
rect 28880 17543 29344 17577
rect 29898 17543 30362 17577
rect 30916 17543 31380 17577
rect 31934 17543 32398 17577
rect 32952 17543 33416 17577
rect 33970 17543 34434 17577
rect 34988 17543 35452 17577
rect 36006 17543 36470 17577
rect 37024 17543 37488 17577
rect 38042 17543 38506 17577
rect 39060 17543 39524 17577
rect 19504 17159 19968 17193
rect 20522 17159 20986 17193
rect 21540 17159 22004 17193
rect 22558 17159 23022 17193
rect 24514 16908 24548 17484
rect 25532 16908 25566 17484
rect 26550 16908 26584 17484
rect 27568 16908 27602 17484
rect 28586 16908 28620 17484
rect 29604 16908 29638 17484
rect 30622 16908 30656 17484
rect 31640 16908 31674 17484
rect 32658 16908 32692 17484
rect 33676 16908 33710 17484
rect 34694 16908 34728 17484
rect 35712 16908 35746 17484
rect 36730 16908 36764 17484
rect 37748 16908 37782 17484
rect 38766 16908 38800 17484
rect 39784 16908 39818 17484
rect 19504 16855 19968 16889
rect 20522 16855 20986 16889
rect 21540 16855 22004 16889
rect 22558 16855 23022 16889
rect 24808 16815 25272 16849
rect 25826 16815 26290 16849
rect 26844 16815 27308 16849
rect 27862 16815 28326 16849
rect 28880 16815 29344 16849
rect 29898 16815 30362 16849
rect 30916 16815 31380 16849
rect 31934 16815 32398 16849
rect 32952 16815 33416 16849
rect 33970 16815 34434 16849
rect 34988 16815 35452 16849
rect 36006 16815 36470 16849
rect 37024 16815 37488 16849
rect 38042 16815 38506 16849
rect 39060 16815 39524 16849
rect 19210 16220 19244 16796
rect 20228 16220 20262 16796
rect 21246 16220 21280 16796
rect 22264 16220 22298 16796
rect 23282 16220 23316 16796
rect 24808 16287 25272 16321
rect 25826 16287 26290 16321
rect 26844 16287 27308 16321
rect 27862 16287 28326 16321
rect 28880 16287 29344 16321
rect 29898 16287 30362 16321
rect 30916 16287 31380 16321
rect 31934 16287 32398 16321
rect 32952 16287 33416 16321
rect 33970 16287 34434 16321
rect 34988 16287 35452 16321
rect 36006 16287 36470 16321
rect 37024 16287 37488 16321
rect 38042 16287 38506 16321
rect 39060 16287 39524 16321
rect 19504 16127 19968 16161
rect 20522 16127 20986 16161
rect 21540 16127 22004 16161
rect 22558 16127 23022 16161
rect 24514 15652 24548 16228
rect 25532 15652 25566 16228
rect 26550 15652 26584 16228
rect 27568 15652 27602 16228
rect 28586 15652 28620 16228
rect 29604 15652 29638 16228
rect 30622 15652 30656 16228
rect 31640 15652 31674 16228
rect 32658 15652 32692 16228
rect 33676 15652 33710 16228
rect 34694 15652 34728 16228
rect 35712 15652 35746 16228
rect 36730 15652 36764 16228
rect 37748 15652 37782 16228
rect 38766 15652 38800 16228
rect 39784 15652 39818 16228
rect 24808 15559 25272 15593
rect 25826 15559 26290 15593
rect 26844 15559 27308 15593
rect 27862 15559 28326 15593
rect 28880 15559 29344 15593
rect 29898 15559 30362 15593
rect 30916 15559 31380 15593
rect 31934 15559 32398 15593
rect 32952 15559 33416 15593
rect 33970 15559 34434 15593
rect 34988 15559 35452 15593
rect 36006 15559 36470 15593
rect 37024 15559 37488 15593
rect 38042 15559 38506 15593
rect 39060 15559 39524 15593
rect 41762 15352 41862 28782
rect 17518 14732 17580 14832
rect 17580 14732 41700 14832
rect 41700 14732 41762 14832
rect 4818 13802 4880 13902
rect 4880 13802 41800 13902
rect 41800 13802 41862 13902
rect 19916 13082 20380 13116
rect 20934 13082 21398 13116
rect 21952 13082 22416 13116
rect 22970 13082 23434 13116
rect 23988 13082 24452 13116
rect 25006 13082 25470 13116
rect 26024 13082 26488 13116
rect 27042 13082 27506 13116
rect 28060 13082 28524 13116
rect 29078 13082 29542 13116
rect 30096 13082 30560 13116
rect 31114 13082 31578 13116
rect 32132 13082 32596 13116
rect 33150 13082 33614 13116
rect 34168 13082 34632 13116
rect 35186 13082 35650 13116
rect 36204 13082 36668 13116
rect 37222 13082 37686 13116
rect 38240 13082 38704 13116
rect 39258 13082 39722 13116
rect -102 842 -40 942
rect -40 842 4240 942
rect 4240 842 4302 942
rect -202 -1773 -102 673
rect 390 480 474 514
rect 648 480 732 514
rect 906 480 990 514
rect 1164 480 1248 514
rect 1422 480 1506 514
rect 1680 480 1764 514
rect 1938 480 2022 514
rect 2196 480 2280 514
rect 2454 480 2538 514
rect 2712 480 2796 514
rect 2970 480 3054 514
rect 3228 480 3312 514
rect 3486 480 3570 514
rect 3744 480 3828 514
rect 286 54 320 430
rect 544 54 578 430
rect 802 54 836 430
rect 1060 54 1094 430
rect 1318 54 1352 430
rect 1576 54 1610 430
rect 1834 54 1868 430
rect 2092 54 2126 430
rect 2350 54 2384 430
rect 2608 54 2642 430
rect 2866 54 2900 430
rect 3124 54 3158 430
rect 3382 54 3416 430
rect 3640 54 3674 430
rect 3898 54 3932 430
rect 390 -30 474 4
rect 648 -30 732 4
rect 906 -30 990 4
rect 1164 -30 1248 4
rect 1422 -30 1506 4
rect 1680 -30 1764 4
rect 1938 -30 2022 4
rect 2196 -30 2280 4
rect 2454 -30 2538 4
rect 2712 -30 2796 4
rect 2970 -30 3054 4
rect 3228 -30 3312 4
rect 3486 -30 3570 4
rect 3744 -30 3828 4
rect 390 -520 474 -486
rect 648 -520 732 -486
rect 906 -520 990 -486
rect 1164 -520 1248 -486
rect 1422 -520 1506 -486
rect 1680 -520 1764 -486
rect 1938 -520 2022 -486
rect 2196 -520 2280 -486
rect 2454 -520 2538 -486
rect 2712 -520 2796 -486
rect 2970 -520 3054 -486
rect 3228 -520 3312 -486
rect 3486 -520 3570 -486
rect 3744 -520 3828 -486
rect 286 -946 320 -570
rect 544 -946 578 -570
rect 802 -946 836 -570
rect 1060 -946 1094 -570
rect 1318 -946 1352 -570
rect 1576 -946 1610 -570
rect 1834 -946 1868 -570
rect 2092 -946 2126 -570
rect 2350 -946 2384 -570
rect 2608 -946 2642 -570
rect 2866 -946 2900 -570
rect 3124 -946 3158 -570
rect 3382 -946 3416 -570
rect 3640 -946 3674 -570
rect 3898 -946 3932 -570
rect 390 -1030 474 -996
rect 648 -1030 732 -996
rect 906 -1030 990 -996
rect 1164 -1030 1248 -996
rect 1422 -1030 1506 -996
rect 1680 -1030 1764 -996
rect 1938 -1030 2022 -996
rect 2196 -1030 2280 -996
rect 2454 -1030 2538 -996
rect 2712 -1030 2796 -996
rect 2970 -1030 3054 -996
rect 3228 -1030 3312 -996
rect 3486 -1030 3570 -996
rect 3744 -1030 3828 -996
rect 4302 -1773 4402 673
rect -102 -2042 -40 -1942
rect -40 -2042 4240 -1942
rect 4240 -2042 4302 -1942
rect 4718 -1250 4818 13010
rect 8150 12606 8614 12640
rect 9168 12606 9632 12640
rect 10186 12606 10650 12640
rect 11204 12606 11668 12640
rect 12222 12606 12686 12640
rect 13240 12606 13704 12640
rect 14258 12606 14722 12640
rect 15276 12606 15740 12640
rect 16294 12606 16758 12640
rect 7856 11980 7890 12556
rect 8874 11980 8908 12556
rect 9892 11980 9926 12556
rect 10910 11980 10944 12556
rect 11928 11980 11962 12556
rect 12946 11980 12980 12556
rect 13964 11980 13998 12556
rect 14982 11980 15016 12556
rect 16000 11980 16034 12556
rect 17018 11980 17052 12556
rect 19622 12456 19656 13032
rect 20640 12456 20674 13032
rect 21658 12456 21692 13032
rect 22676 12456 22710 13032
rect 23694 12456 23728 13032
rect 24712 12456 24746 13032
rect 25730 12456 25764 13032
rect 26748 12456 26782 13032
rect 27766 12456 27800 13032
rect 28784 12456 28818 13032
rect 29802 12456 29836 13032
rect 30820 12456 30854 13032
rect 31838 12456 31872 13032
rect 32856 12456 32890 13032
rect 33874 12456 33908 13032
rect 34892 12456 34926 13032
rect 35910 12456 35944 13032
rect 36928 12456 36962 13032
rect 37946 12456 37980 13032
rect 38964 12456 38998 13032
rect 39982 12456 40016 13032
rect 19916 12372 20380 12406
rect 20934 12372 21398 12406
rect 21952 12372 22416 12406
rect 22970 12372 23434 12406
rect 23988 12372 24452 12406
rect 25006 12372 25470 12406
rect 26024 12372 26488 12406
rect 27042 12372 27506 12406
rect 28060 12372 28524 12406
rect 29078 12372 29542 12406
rect 30096 12372 30560 12406
rect 31114 12372 31578 12406
rect 32132 12372 32596 12406
rect 33150 12372 33614 12406
rect 34168 12372 34632 12406
rect 35186 12372 35650 12406
rect 36204 12372 36668 12406
rect 37222 12372 37686 12406
rect 38240 12372 38704 12406
rect 39258 12372 39722 12406
rect 19916 12264 20380 12298
rect 20934 12264 21398 12298
rect 21952 12264 22416 12298
rect 22970 12264 23434 12298
rect 23988 12264 24452 12298
rect 25006 12264 25470 12298
rect 26024 12264 26488 12298
rect 27042 12264 27506 12298
rect 28060 12264 28524 12298
rect 29078 12264 29542 12298
rect 30096 12264 30560 12298
rect 31114 12264 31578 12298
rect 32132 12264 32596 12298
rect 33150 12264 33614 12298
rect 34168 12264 34632 12298
rect 35186 12264 35650 12298
rect 36204 12264 36668 12298
rect 37222 12264 37686 12298
rect 38240 12264 38704 12298
rect 39258 12264 39722 12298
rect 8150 11896 8614 11930
rect 9168 11896 9632 11930
rect 8150 11788 8614 11822
rect 10186 11896 10650 11930
rect 9168 11788 9632 11822
rect 11204 11896 11668 11930
rect 10186 11788 10650 11822
rect 12222 11896 12686 11930
rect 11204 11788 11668 11822
rect 13240 11896 13704 11930
rect 12222 11788 12686 11822
rect 14258 11896 14722 11930
rect 13240 11788 13704 11822
rect 15276 11896 15740 11930
rect 14258 11788 14722 11822
rect 16294 11896 16758 11930
rect 15276 11788 15740 11822
rect 16294 11788 16758 11822
rect 7856 11162 7890 11738
rect 8874 11162 8908 11738
rect 9892 11162 9926 11738
rect 10910 11162 10944 11738
rect 11928 11162 11962 11738
rect 12946 11162 12980 11738
rect 13964 11162 13998 11738
rect 14982 11162 15016 11738
rect 16000 11162 16034 11738
rect 17018 11162 17052 11738
rect 19622 11638 19656 12214
rect 20640 11638 20674 12214
rect 21658 11638 21692 12214
rect 22676 11638 22710 12214
rect 23694 11638 23728 12214
rect 24712 11638 24746 12214
rect 25730 11638 25764 12214
rect 26748 11638 26782 12214
rect 27766 11638 27800 12214
rect 28784 11638 28818 12214
rect 29802 11638 29836 12214
rect 30820 11638 30854 12214
rect 31838 11638 31872 12214
rect 32856 11638 32890 12214
rect 33874 11638 33908 12214
rect 34892 11638 34926 12214
rect 35910 11638 35944 12214
rect 36928 11638 36962 12214
rect 37946 11638 37980 12214
rect 38964 11638 38998 12214
rect 39982 11638 40016 12214
rect 19916 11554 20380 11588
rect 20934 11554 21398 11588
rect 21952 11554 22416 11588
rect 22970 11554 23434 11588
rect 23988 11554 24452 11588
rect 25006 11554 25470 11588
rect 26024 11554 26488 11588
rect 27042 11554 27506 11588
rect 28060 11554 28524 11588
rect 29078 11554 29542 11588
rect 30096 11554 30560 11588
rect 31114 11554 31578 11588
rect 32132 11554 32596 11588
rect 33150 11554 33614 11588
rect 34168 11554 34632 11588
rect 35186 11554 35650 11588
rect 36204 11554 36668 11588
rect 37222 11554 37686 11588
rect 38240 11554 38704 11588
rect 39258 11554 39722 11588
rect 8150 11078 8614 11112
rect 9168 11078 9632 11112
rect 8150 10970 8614 11004
rect 10186 11078 10650 11112
rect 9168 10970 9632 11004
rect 11204 11078 11668 11112
rect 10186 10970 10650 11004
rect 12222 11078 12686 11112
rect 11204 10970 11668 11004
rect 13240 11078 13704 11112
rect 12222 10970 12686 11004
rect 14258 11078 14722 11112
rect 13240 10970 13704 11004
rect 15276 11078 15740 11112
rect 14258 10970 14722 11004
rect 16294 11078 16758 11112
rect 15276 10970 15740 11004
rect 16294 10970 16758 11004
rect 7856 10344 7890 10920
rect 8874 10344 8908 10920
rect 9892 10344 9926 10920
rect 10910 10344 10944 10920
rect 11928 10344 11962 10920
rect 12946 10344 12980 10920
rect 13964 10344 13998 10920
rect 14982 10344 15016 10920
rect 16000 10344 16034 10920
rect 17018 10344 17052 10920
rect 19916 10886 20380 10920
rect 20934 10886 21398 10920
rect 21952 10886 22416 10920
rect 22970 10886 23434 10920
rect 23988 10886 24452 10920
rect 25006 10886 25470 10920
rect 26024 10886 26488 10920
rect 27042 10886 27506 10920
rect 28060 10886 28524 10920
rect 29078 10886 29542 10920
rect 30096 10886 30560 10920
rect 31114 10886 31578 10920
rect 32132 10886 32596 10920
rect 33150 10886 33614 10920
rect 34168 10886 34632 10920
rect 35186 10886 35650 10920
rect 36204 10886 36668 10920
rect 37222 10886 37686 10920
rect 38240 10886 38704 10920
rect 39258 10886 39722 10920
rect 8150 10260 8614 10294
rect 9168 10260 9632 10294
rect 8150 10152 8614 10186
rect 10186 10260 10650 10294
rect 9168 10152 9632 10186
rect 11204 10260 11668 10294
rect 10186 10152 10650 10186
rect 12222 10260 12686 10294
rect 11204 10152 11668 10186
rect 13240 10260 13704 10294
rect 12222 10152 12686 10186
rect 14258 10260 14722 10294
rect 13240 10152 13704 10186
rect 15276 10260 15740 10294
rect 14258 10152 14722 10186
rect 16294 10260 16758 10294
rect 15276 10152 15740 10186
rect 19622 10260 19656 10836
rect 20640 10260 20674 10836
rect 21658 10260 21692 10836
rect 22676 10260 22710 10836
rect 23694 10260 23728 10836
rect 24712 10260 24746 10836
rect 25730 10260 25764 10836
rect 26748 10260 26782 10836
rect 27766 10260 27800 10836
rect 28784 10260 28818 10836
rect 29802 10260 29836 10836
rect 30820 10260 30854 10836
rect 31838 10260 31872 10836
rect 32856 10260 32890 10836
rect 33874 10260 33908 10836
rect 34892 10260 34926 10836
rect 35910 10260 35944 10836
rect 36928 10260 36962 10836
rect 37946 10260 37980 10836
rect 38964 10260 38998 10836
rect 39982 10260 40016 10836
rect 16294 10152 16758 10186
rect 19916 10176 20380 10210
rect 20934 10176 21398 10210
rect 21952 10176 22416 10210
rect 22970 10176 23434 10210
rect 23988 10176 24452 10210
rect 25006 10176 25470 10210
rect 26024 10176 26488 10210
rect 27042 10176 27506 10210
rect 28060 10176 28524 10210
rect 29078 10176 29542 10210
rect 30096 10176 30560 10210
rect 31114 10176 31578 10210
rect 32132 10176 32596 10210
rect 33150 10176 33614 10210
rect 34168 10176 34632 10210
rect 35186 10176 35650 10210
rect 36204 10176 36668 10210
rect 37222 10176 37686 10210
rect 38240 10176 38704 10210
rect 39258 10176 39722 10210
rect 7856 9526 7890 10102
rect 8874 9526 8908 10102
rect 9892 9526 9926 10102
rect 10910 9526 10944 10102
rect 11928 9526 11962 10102
rect 12946 9526 12980 10102
rect 13964 9526 13998 10102
rect 14982 9526 15016 10102
rect 16000 9526 16034 10102
rect 17018 9526 17052 10102
rect 19916 9654 20380 9688
rect 20934 9654 21398 9688
rect 21952 9654 22416 9688
rect 22970 9654 23434 9688
rect 23988 9654 24452 9688
rect 25006 9654 25470 9688
rect 26024 9654 26488 9688
rect 27042 9654 27506 9688
rect 28060 9654 28524 9688
rect 29078 9654 29542 9688
rect 30096 9654 30560 9688
rect 31114 9654 31578 9688
rect 32132 9654 32596 9688
rect 33150 9654 33614 9688
rect 34168 9654 34632 9688
rect 35186 9654 35650 9688
rect 36204 9654 36668 9688
rect 37222 9654 37686 9688
rect 38240 9654 38704 9688
rect 39258 9654 39722 9688
rect 8150 9442 8614 9476
rect 9168 9442 9632 9476
rect 8150 9334 8614 9368
rect 10186 9442 10650 9476
rect 9168 9334 9632 9368
rect 11204 9442 11668 9476
rect 10186 9334 10650 9368
rect 12222 9442 12686 9476
rect 11204 9334 11668 9368
rect 13240 9442 13704 9476
rect 12222 9334 12686 9368
rect 14258 9442 14722 9476
rect 13240 9334 13704 9368
rect 15276 9442 15740 9476
rect 14258 9334 14722 9368
rect 16294 9442 16758 9476
rect 15276 9334 15740 9368
rect 16294 9334 16758 9368
rect 7856 8708 7890 9284
rect 8874 8708 8908 9284
rect 9892 8708 9926 9284
rect 10910 8708 10944 9284
rect 11928 8708 11962 9284
rect 12946 8708 12980 9284
rect 13964 8708 13998 9284
rect 14982 8708 15016 9284
rect 16000 8708 16034 9284
rect 17018 8708 17052 9284
rect 19622 9028 19656 9604
rect 20640 9028 20674 9604
rect 21658 9028 21692 9604
rect 22676 9028 22710 9604
rect 23694 9028 23728 9604
rect 24712 9028 24746 9604
rect 25730 9028 25764 9604
rect 26748 9028 26782 9604
rect 27766 9028 27800 9604
rect 28784 9028 28818 9604
rect 29802 9028 29836 9604
rect 30820 9028 30854 9604
rect 31838 9028 31872 9604
rect 32856 9028 32890 9604
rect 33874 9028 33908 9604
rect 34892 9028 34926 9604
rect 35910 9028 35944 9604
rect 36928 9028 36962 9604
rect 37946 9028 37980 9604
rect 38964 9028 38998 9604
rect 39982 9028 40016 9604
rect 19916 8944 20380 8978
rect 20934 8944 21398 8978
rect 21952 8944 22416 8978
rect 22970 8944 23434 8978
rect 23988 8944 24452 8978
rect 25006 8944 25470 8978
rect 26024 8944 26488 8978
rect 27042 8944 27506 8978
rect 28060 8944 28524 8978
rect 29078 8944 29542 8978
rect 30096 8944 30560 8978
rect 31114 8944 31578 8978
rect 32132 8944 32596 8978
rect 33150 8944 33614 8978
rect 34168 8944 34632 8978
rect 35186 8944 35650 8978
rect 36204 8944 36668 8978
rect 37222 8944 37686 8978
rect 38240 8944 38704 8978
rect 39258 8944 39722 8978
rect 8150 8624 8614 8658
rect 9168 8624 9632 8658
rect 8150 8516 8614 8550
rect 10186 8624 10650 8658
rect 9168 8516 9632 8550
rect 11204 8624 11668 8658
rect 10186 8516 10650 8550
rect 12222 8624 12686 8658
rect 11204 8516 11668 8550
rect 13240 8624 13704 8658
rect 12222 8516 12686 8550
rect 14258 8624 14722 8658
rect 13240 8516 13704 8550
rect 15276 8624 15740 8658
rect 14258 8516 14722 8550
rect 16294 8624 16758 8658
rect 15276 8516 15740 8550
rect 16294 8516 16758 8550
rect 7856 7890 7890 8466
rect 8874 7890 8908 8466
rect 9892 7890 9926 8466
rect 10910 7890 10944 8466
rect 11928 7890 11962 8466
rect 12946 7890 12980 8466
rect 13964 7890 13998 8466
rect 14982 7890 15016 8466
rect 16000 7890 16034 8466
rect 17018 7890 17052 8466
rect 19914 8420 20378 8454
rect 20932 8420 21396 8454
rect 21950 8420 22414 8454
rect 22968 8420 23432 8454
rect 23986 8420 24450 8454
rect 25004 8420 25468 8454
rect 26022 8420 26486 8454
rect 27040 8420 27504 8454
rect 28058 8420 28522 8454
rect 29076 8420 29540 8454
rect 30094 8420 30558 8454
rect 31112 8420 31576 8454
rect 32130 8420 32594 8454
rect 33148 8420 33612 8454
rect 34166 8420 34630 8454
rect 35184 8420 35648 8454
rect 36202 8420 36666 8454
rect 37220 8420 37684 8454
rect 38238 8420 38702 8454
rect 39256 8420 39720 8454
rect 8150 7806 8614 7840
rect 9168 7806 9632 7840
rect 8150 7698 8614 7732
rect 10186 7806 10650 7840
rect 9168 7698 9632 7732
rect 11204 7806 11668 7840
rect 10186 7698 10650 7732
rect 12222 7806 12686 7840
rect 11204 7698 11668 7732
rect 13240 7806 13704 7840
rect 12222 7698 12686 7732
rect 14258 7806 14722 7840
rect 13240 7698 13704 7732
rect 15276 7806 15740 7840
rect 14258 7698 14722 7732
rect 16294 7806 16758 7840
rect 15276 7698 15740 7732
rect 19620 7794 19654 8370
rect 20638 7794 20672 8370
rect 21656 7794 21690 8370
rect 22674 7794 22708 8370
rect 23692 7794 23726 8370
rect 24710 7794 24744 8370
rect 25728 7794 25762 8370
rect 26746 7794 26780 8370
rect 27764 7794 27798 8370
rect 28782 7794 28816 8370
rect 29800 7794 29834 8370
rect 30818 7794 30852 8370
rect 31836 7794 31870 8370
rect 32854 7794 32888 8370
rect 33872 7794 33906 8370
rect 34890 7794 34924 8370
rect 35908 7794 35942 8370
rect 36926 7794 36960 8370
rect 37944 7794 37978 8370
rect 38962 7794 38996 8370
rect 39980 7794 40014 8370
rect 16294 7698 16758 7732
rect 19914 7710 20378 7744
rect 20932 7710 21396 7744
rect 21950 7710 22414 7744
rect 22968 7710 23432 7744
rect 23986 7710 24450 7744
rect 25004 7710 25468 7744
rect 26022 7710 26486 7744
rect 27040 7710 27504 7744
rect 28058 7710 28522 7744
rect 29076 7710 29540 7744
rect 30094 7710 30558 7744
rect 31112 7710 31576 7744
rect 32130 7710 32594 7744
rect 33148 7710 33612 7744
rect 34166 7710 34630 7744
rect 35184 7710 35648 7744
rect 36202 7710 36666 7744
rect 37220 7710 37684 7744
rect 38238 7710 38702 7744
rect 39256 7710 39720 7744
rect 7856 7072 7890 7648
rect 8874 7072 8908 7648
rect 9892 7072 9926 7648
rect 10910 7072 10944 7648
rect 11928 7072 11962 7648
rect 12946 7072 12980 7648
rect 13964 7072 13998 7648
rect 14982 7072 15016 7648
rect 16000 7072 16034 7648
rect 17018 7072 17052 7648
rect 19914 7186 20378 7220
rect 20932 7186 21396 7220
rect 21950 7186 22414 7220
rect 22968 7186 23432 7220
rect 23986 7186 24450 7220
rect 25004 7186 25468 7220
rect 26022 7186 26486 7220
rect 27040 7186 27504 7220
rect 28058 7186 28522 7220
rect 29076 7186 29540 7220
rect 30094 7186 30558 7220
rect 31112 7186 31576 7220
rect 32130 7186 32594 7220
rect 33148 7186 33612 7220
rect 34166 7186 34630 7220
rect 35184 7186 35648 7220
rect 36202 7186 36666 7220
rect 37220 7186 37684 7220
rect 38238 7186 38702 7220
rect 39256 7186 39720 7220
rect 8150 6988 8614 7022
rect 9168 6988 9632 7022
rect 8150 6880 8614 6914
rect 10186 6988 10650 7022
rect 9168 6880 9632 6914
rect 11204 6988 11668 7022
rect 10186 6880 10650 6914
rect 12222 6988 12686 7022
rect 11204 6880 11668 6914
rect 13240 6988 13704 7022
rect 12222 6880 12686 6914
rect 14258 6988 14722 7022
rect 13240 6880 13704 6914
rect 15276 6988 15740 7022
rect 14258 6880 14722 6914
rect 16294 6988 16758 7022
rect 15276 6880 15740 6914
rect 16294 6880 16758 6914
rect 7856 6254 7890 6830
rect 8874 6254 8908 6830
rect 9892 6254 9926 6830
rect 10910 6254 10944 6830
rect 11928 6254 11962 6830
rect 12946 6254 12980 6830
rect 13964 6254 13998 6830
rect 14982 6254 15016 6830
rect 16000 6254 16034 6830
rect 17018 6254 17052 6830
rect 19620 6560 19654 7136
rect 20638 6560 20672 7136
rect 21656 6560 21690 7136
rect 22674 6560 22708 7136
rect 23692 6560 23726 7136
rect 24710 6560 24744 7136
rect 25728 6560 25762 7136
rect 26746 6560 26780 7136
rect 27764 6560 27798 7136
rect 28782 6560 28816 7136
rect 29800 6560 29834 7136
rect 30818 6560 30852 7136
rect 31836 6560 31870 7136
rect 32854 6560 32888 7136
rect 33872 6560 33906 7136
rect 34890 6560 34924 7136
rect 35908 6560 35942 7136
rect 36926 6560 36960 7136
rect 37944 6560 37978 7136
rect 38962 6560 38996 7136
rect 39980 6560 40014 7136
rect 19914 6476 20378 6510
rect 20932 6476 21396 6510
rect 21950 6476 22414 6510
rect 22968 6476 23432 6510
rect 23986 6476 24450 6510
rect 25004 6476 25468 6510
rect 26022 6476 26486 6510
rect 27040 6476 27504 6510
rect 28058 6476 28522 6510
rect 29076 6476 29540 6510
rect 30094 6476 30558 6510
rect 31112 6476 31576 6510
rect 32130 6476 32594 6510
rect 33148 6476 33612 6510
rect 34166 6476 34630 6510
rect 35184 6476 35648 6510
rect 36202 6476 36666 6510
rect 37220 6476 37684 6510
rect 38238 6476 38702 6510
rect 39256 6476 39720 6510
rect 8150 6170 8614 6204
rect 9168 6170 9632 6204
rect 10186 6170 10650 6204
rect 11204 6170 11668 6204
rect 12222 6170 12686 6204
rect 13240 6170 13704 6204
rect 14258 6170 14722 6204
rect 15276 6170 15740 6204
rect 16294 6170 16758 6204
rect 19914 5954 20378 5988
rect 20932 5954 21396 5988
rect 21950 5954 22414 5988
rect 22968 5954 23432 5988
rect 23986 5954 24450 5988
rect 25004 5954 25468 5988
rect 26022 5954 26486 5988
rect 27040 5954 27504 5988
rect 28058 5954 28522 5988
rect 29076 5954 29540 5988
rect 30094 5954 30558 5988
rect 31112 5954 31576 5988
rect 32130 5954 32594 5988
rect 33148 5954 33612 5988
rect 34166 5954 34630 5988
rect 35184 5954 35648 5988
rect 36202 5954 36666 5988
rect 37220 5954 37684 5988
rect 38238 5954 38702 5988
rect 39256 5954 39720 5988
rect 19620 5328 19654 5904
rect 20638 5328 20672 5904
rect 21656 5328 21690 5904
rect 22674 5328 22708 5904
rect 23692 5328 23726 5904
rect 24710 5328 24744 5904
rect 25728 5328 25762 5904
rect 26746 5328 26780 5904
rect 27764 5328 27798 5904
rect 28782 5328 28816 5904
rect 29800 5328 29834 5904
rect 30818 5328 30852 5904
rect 31836 5328 31870 5904
rect 32854 5328 32888 5904
rect 33872 5328 33906 5904
rect 34890 5328 34924 5904
rect 35908 5328 35942 5904
rect 36926 5328 36960 5904
rect 37944 5328 37978 5904
rect 38962 5328 38996 5904
rect 39980 5328 40014 5904
rect 19914 5244 20378 5278
rect 20932 5244 21396 5278
rect 21950 5244 22414 5278
rect 22968 5244 23432 5278
rect 23986 5244 24450 5278
rect 25004 5244 25468 5278
rect 26022 5244 26486 5278
rect 27040 5244 27504 5278
rect 28058 5244 28522 5278
rect 29076 5244 29540 5278
rect 30094 5244 30558 5278
rect 31112 5244 31576 5278
rect 32130 5244 32594 5278
rect 33148 5244 33612 5278
rect 34166 5244 34630 5278
rect 35184 5244 35648 5278
rect 36202 5244 36666 5278
rect 37220 5244 37684 5278
rect 38238 5244 38702 5278
rect 39256 5244 39720 5278
rect 6826 4856 7290 4890
rect 7844 4856 8308 4890
rect 8862 4856 9326 4890
rect 9880 4856 10344 4890
rect 10898 4856 11362 4890
rect 11916 4856 12380 4890
rect 12934 4856 13398 4890
rect 13952 4856 14416 4890
rect 14970 4856 15434 4890
rect 15988 4856 16452 4890
rect 17006 4856 17470 4890
rect 6532 4230 6566 4806
rect 7550 4230 7584 4806
rect 8568 4230 8602 4806
rect 9586 4230 9620 4806
rect 10604 4230 10638 4806
rect 11622 4230 11656 4806
rect 12640 4230 12674 4806
rect 13658 4230 13692 4806
rect 14676 4230 14710 4806
rect 15694 4230 15728 4806
rect 16712 4230 16746 4806
rect 17730 4230 17764 4806
rect 19914 4720 20378 4754
rect 20932 4720 21396 4754
rect 21950 4720 22414 4754
rect 22968 4720 23432 4754
rect 23986 4720 24450 4754
rect 25004 4720 25468 4754
rect 26022 4720 26486 4754
rect 27040 4720 27504 4754
rect 28058 4720 28522 4754
rect 29076 4720 29540 4754
rect 30094 4720 30558 4754
rect 31112 4720 31576 4754
rect 32130 4720 32594 4754
rect 33148 4720 33612 4754
rect 34166 4720 34630 4754
rect 35184 4720 35648 4754
rect 36202 4720 36666 4754
rect 37220 4720 37684 4754
rect 38238 4720 38702 4754
rect 39256 4720 39720 4754
rect 6826 4146 7290 4180
rect 7844 4146 8308 4180
rect 8862 4146 9326 4180
rect 9880 4146 10344 4180
rect 10898 4146 11362 4180
rect 11916 4146 12380 4180
rect 12934 4146 13398 4180
rect 13952 4146 14416 4180
rect 14970 4146 15434 4180
rect 15988 4146 16452 4180
rect 17006 4146 17470 4180
rect 19620 4094 19654 4670
rect 20638 4094 20672 4670
rect 21656 4094 21690 4670
rect 22674 4094 22708 4670
rect 23692 4094 23726 4670
rect 24710 4094 24744 4670
rect 25728 4094 25762 4670
rect 26746 4094 26780 4670
rect 27764 4094 27798 4670
rect 28782 4094 28816 4670
rect 29800 4094 29834 4670
rect 30818 4094 30852 4670
rect 31836 4094 31870 4670
rect 32854 4094 32888 4670
rect 33872 4094 33906 4670
rect 34890 4094 34924 4670
rect 35908 4094 35942 4670
rect 36926 4094 36960 4670
rect 37944 4094 37978 4670
rect 38962 4094 38996 4670
rect 39980 4094 40014 4670
rect 19914 4010 20378 4044
rect 20932 4010 21396 4044
rect 21950 4010 22414 4044
rect 22968 4010 23432 4044
rect 23986 4010 24450 4044
rect 25004 4010 25468 4044
rect 26022 4010 26486 4044
rect 27040 4010 27504 4044
rect 28058 4010 28522 4044
rect 29076 4010 29540 4044
rect 30094 4010 30558 4044
rect 31112 4010 31576 4044
rect 32130 4010 32594 4044
rect 33148 4010 33612 4044
rect 34166 4010 34630 4044
rect 35184 4010 35648 4044
rect 36202 4010 36666 4044
rect 37220 4010 37684 4044
rect 38238 4010 38702 4044
rect 39256 4010 39720 4044
rect 6826 3744 7290 3778
rect 7844 3744 8308 3778
rect 8862 3744 9326 3778
rect 9880 3744 10344 3778
rect 10898 3744 11362 3778
rect 11916 3744 12380 3778
rect 12934 3744 13398 3778
rect 13952 3744 14416 3778
rect 14970 3744 15434 3778
rect 15988 3744 16452 3778
rect 17006 3744 17470 3778
rect 6532 3118 6566 3694
rect 7550 3118 7584 3694
rect 8568 3118 8602 3694
rect 9586 3118 9620 3694
rect 10604 3118 10638 3694
rect 11622 3118 11656 3694
rect 12640 3118 12674 3694
rect 13658 3118 13692 3694
rect 14676 3118 14710 3694
rect 15694 3118 15728 3694
rect 16712 3118 16746 3694
rect 17730 3118 17764 3694
rect 19914 3486 20378 3520
rect 20932 3486 21396 3520
rect 21950 3486 22414 3520
rect 22968 3486 23432 3520
rect 23986 3486 24450 3520
rect 25004 3486 25468 3520
rect 26022 3486 26486 3520
rect 27040 3486 27504 3520
rect 28058 3486 28522 3520
rect 29076 3486 29540 3520
rect 30094 3486 30558 3520
rect 31112 3486 31576 3520
rect 32130 3486 32594 3520
rect 33148 3486 33612 3520
rect 34166 3486 34630 3520
rect 35184 3486 35648 3520
rect 36202 3486 36666 3520
rect 37220 3486 37684 3520
rect 38238 3486 38702 3520
rect 39256 3486 39720 3520
rect 6826 3034 7290 3068
rect 7844 3034 8308 3068
rect 8862 3034 9326 3068
rect 9880 3034 10344 3068
rect 10898 3034 11362 3068
rect 11916 3034 12380 3068
rect 12934 3034 13398 3068
rect 13952 3034 14416 3068
rect 14970 3034 15434 3068
rect 15988 3034 16452 3068
rect 17006 3034 17470 3068
rect 19620 2860 19654 3436
rect 20638 2860 20672 3436
rect 21656 2860 21690 3436
rect 22674 2860 22708 3436
rect 23692 2860 23726 3436
rect 24710 2860 24744 3436
rect 25728 2860 25762 3436
rect 26746 2860 26780 3436
rect 27764 2860 27798 3436
rect 28782 2860 28816 3436
rect 29800 2860 29834 3436
rect 30818 2860 30852 3436
rect 31836 2860 31870 3436
rect 32854 2860 32888 3436
rect 33872 2860 33906 3436
rect 34890 2860 34924 3436
rect 35908 2860 35942 3436
rect 36926 2860 36960 3436
rect 37944 2860 37978 3436
rect 38962 2860 38996 3436
rect 39980 2860 40014 3436
rect 19914 2776 20378 2810
rect 20932 2776 21396 2810
rect 21950 2776 22414 2810
rect 22968 2776 23432 2810
rect 23986 2776 24450 2810
rect 25004 2776 25468 2810
rect 26022 2776 26486 2810
rect 27040 2776 27504 2810
rect 28058 2776 28522 2810
rect 29076 2776 29540 2810
rect 30094 2776 30558 2810
rect 31112 2776 31576 2810
rect 32130 2776 32594 2810
rect 33148 2776 33612 2810
rect 34166 2776 34630 2810
rect 35184 2776 35648 2810
rect 36202 2776 36666 2810
rect 37220 2776 37684 2810
rect 38238 2776 38702 2810
rect 39256 2776 39720 2810
rect 6826 2632 7290 2666
rect 7844 2632 8308 2666
rect 8862 2632 9326 2666
rect 9880 2632 10344 2666
rect 10898 2632 11362 2666
rect 11916 2632 12380 2666
rect 12934 2632 13398 2666
rect 13952 2632 14416 2666
rect 14970 2632 15434 2666
rect 15988 2632 16452 2666
rect 17006 2632 17470 2666
rect 6532 2006 6566 2582
rect 7550 2006 7584 2582
rect 8568 2006 8602 2582
rect 9586 2006 9620 2582
rect 10604 2006 10638 2582
rect 11622 2006 11656 2582
rect 12640 2006 12674 2582
rect 13658 2006 13692 2582
rect 14676 2006 14710 2582
rect 15694 2006 15728 2582
rect 16712 2006 16746 2582
rect 17730 2006 17764 2582
rect 19914 2254 20378 2288
rect 20932 2254 21396 2288
rect 21950 2254 22414 2288
rect 22968 2254 23432 2288
rect 23986 2254 24450 2288
rect 25004 2254 25468 2288
rect 26022 2254 26486 2288
rect 27040 2254 27504 2288
rect 28058 2254 28522 2288
rect 29076 2254 29540 2288
rect 30094 2254 30558 2288
rect 31112 2254 31576 2288
rect 32130 2254 32594 2288
rect 33148 2254 33612 2288
rect 34166 2254 34630 2288
rect 35184 2254 35648 2288
rect 36202 2254 36666 2288
rect 37220 2254 37684 2288
rect 38238 2254 38702 2288
rect 39256 2254 39720 2288
rect 6826 1922 7290 1956
rect 7844 1922 8308 1956
rect 8862 1922 9326 1956
rect 9880 1922 10344 1956
rect 10898 1922 11362 1956
rect 11916 1922 12380 1956
rect 12934 1922 13398 1956
rect 13952 1922 14416 1956
rect 14970 1922 15434 1956
rect 15988 1922 16452 1956
rect 17006 1922 17470 1956
rect 19620 1628 19654 2204
rect 20638 1628 20672 2204
rect 21656 1628 21690 2204
rect 22674 1628 22708 2204
rect 23692 1628 23726 2204
rect 24710 1628 24744 2204
rect 25728 1628 25762 2204
rect 26746 1628 26780 2204
rect 27764 1628 27798 2204
rect 28782 1628 28816 2204
rect 29800 1628 29834 2204
rect 30818 1628 30852 2204
rect 31836 1628 31870 2204
rect 32854 1628 32888 2204
rect 33872 1628 33906 2204
rect 34890 1628 34924 2204
rect 35908 1628 35942 2204
rect 36926 1628 36960 2204
rect 37944 1628 37978 2204
rect 38962 1628 38996 2204
rect 39980 1628 40014 2204
rect 6826 1520 7290 1554
rect 7844 1520 8308 1554
rect 8862 1520 9326 1554
rect 9880 1520 10344 1554
rect 10898 1520 11362 1554
rect 11916 1520 12380 1554
rect 12934 1520 13398 1554
rect 13952 1520 14416 1554
rect 14970 1520 15434 1554
rect 15988 1520 16452 1554
rect 17006 1520 17470 1554
rect 19914 1544 20378 1578
rect 20932 1544 21396 1578
rect 21950 1544 22414 1578
rect 22968 1544 23432 1578
rect 23986 1544 24450 1578
rect 25004 1544 25468 1578
rect 26022 1544 26486 1578
rect 27040 1544 27504 1578
rect 28058 1544 28522 1578
rect 29076 1544 29540 1578
rect 30094 1544 30558 1578
rect 31112 1544 31576 1578
rect 32130 1544 32594 1578
rect 33148 1544 33612 1578
rect 34166 1544 34630 1578
rect 35184 1544 35648 1578
rect 36202 1544 36666 1578
rect 37220 1544 37684 1578
rect 38238 1544 38702 1578
rect 39256 1544 39720 1578
rect 6532 894 6566 1470
rect 7550 894 7584 1470
rect 8568 894 8602 1470
rect 9586 894 9620 1470
rect 10604 894 10638 1470
rect 11622 894 11656 1470
rect 12640 894 12674 1470
rect 13658 894 13692 1470
rect 14676 894 14710 1470
rect 15694 894 15728 1470
rect 16712 894 16746 1470
rect 17730 894 17764 1470
rect 19914 1020 20378 1054
rect 20932 1020 21396 1054
rect 21950 1020 22414 1054
rect 22968 1020 23432 1054
rect 23986 1020 24450 1054
rect 25004 1020 25468 1054
rect 26022 1020 26486 1054
rect 27040 1020 27504 1054
rect 28058 1020 28522 1054
rect 29076 1020 29540 1054
rect 30094 1020 30558 1054
rect 31112 1020 31576 1054
rect 32130 1020 32594 1054
rect 33148 1020 33612 1054
rect 34166 1020 34630 1054
rect 35184 1020 35648 1054
rect 36202 1020 36666 1054
rect 37220 1020 37684 1054
rect 38238 1020 38702 1054
rect 39256 1020 39720 1054
rect 6826 810 7290 844
rect 7844 810 8308 844
rect 8862 810 9326 844
rect 9880 810 10344 844
rect 10898 810 11362 844
rect 11916 810 12380 844
rect 12934 810 13398 844
rect 13952 810 14416 844
rect 14970 810 15434 844
rect 15988 810 16452 844
rect 17006 810 17470 844
rect 19620 394 19654 970
rect 20638 394 20672 970
rect 21656 394 21690 970
rect 22674 394 22708 970
rect 23692 394 23726 970
rect 24710 394 24744 970
rect 25728 394 25762 970
rect 26746 394 26780 970
rect 27764 394 27798 970
rect 28782 394 28816 970
rect 29800 394 29834 970
rect 30818 394 30852 970
rect 31836 394 31870 970
rect 32854 394 32888 970
rect 33872 394 33906 970
rect 34890 394 34924 970
rect 35908 394 35942 970
rect 36926 394 36960 970
rect 37944 394 37978 970
rect 38962 394 38996 970
rect 39980 394 40014 970
rect 19914 310 20378 344
rect 20932 310 21396 344
rect 21950 310 22414 344
rect 22968 310 23432 344
rect 23986 310 24450 344
rect 25004 310 25468 344
rect 26022 310 26486 344
rect 27040 310 27504 344
rect 28058 310 28522 344
rect 29076 310 29540 344
rect 30094 310 30558 344
rect 31112 310 31576 344
rect 32130 310 32594 344
rect 33148 310 33612 344
rect 34166 310 34630 344
rect 35184 310 35648 344
rect 36202 310 36666 344
rect 37220 310 37684 344
rect 38238 310 38702 344
rect 39256 310 39720 344
rect 7284 -22 7748 12
rect 8302 -22 8766 12
rect 9320 -22 9784 12
rect 10338 -22 10802 12
rect 11356 -22 11820 12
rect 12374 -22 12838 12
rect 13392 -22 13856 12
rect 14410 -22 14874 12
rect 15428 -22 15892 12
rect 16446 -22 16910 12
rect 6990 -648 7024 -72
rect 8008 -648 8042 -72
rect 9026 -648 9060 -72
rect 10044 -648 10078 -72
rect 11062 -648 11096 -72
rect 12080 -648 12114 -72
rect 13098 -648 13132 -72
rect 14116 -648 14150 -72
rect 15134 -648 15168 -72
rect 16152 -648 16186 -72
rect 17170 -648 17204 -72
rect 19914 -212 20378 -178
rect 20932 -212 21396 -178
rect 21950 -212 22414 -178
rect 22968 -212 23432 -178
rect 23986 -212 24450 -178
rect 25004 -212 25468 -178
rect 26022 -212 26486 -178
rect 27040 -212 27504 -178
rect 28058 -212 28522 -178
rect 29076 -212 29540 -178
rect 30094 -212 30558 -178
rect 31112 -212 31576 -178
rect 32130 -212 32594 -178
rect 33148 -212 33612 -178
rect 34166 -212 34630 -178
rect 35184 -212 35648 -178
rect 36202 -212 36666 -178
rect 37220 -212 37684 -178
rect 38238 -212 38702 -178
rect 39256 -212 39720 -178
rect 7284 -732 7748 -698
rect 8302 -732 8766 -698
rect 9320 -732 9784 -698
rect 10338 -732 10802 -698
rect 11356 -732 11820 -698
rect 12374 -732 12838 -698
rect 13392 -732 13856 -698
rect 14410 -732 14874 -698
rect 15428 -732 15892 -698
rect 16446 -732 16910 -698
rect 19620 -838 19654 -262
rect 20638 -838 20672 -262
rect 21656 -838 21690 -262
rect 22674 -838 22708 -262
rect 23692 -838 23726 -262
rect 24710 -838 24744 -262
rect 25728 -838 25762 -262
rect 26746 -838 26780 -262
rect 27764 -838 27798 -262
rect 28782 -838 28816 -262
rect 29800 -838 29834 -262
rect 30818 -838 30852 -262
rect 31836 -838 31870 -262
rect 32854 -838 32888 -262
rect 33872 -838 33906 -262
rect 34890 -838 34924 -262
rect 35908 -838 35942 -262
rect 36926 -838 36960 -262
rect 37944 -838 37978 -262
rect 38962 -838 38996 -262
rect 39980 -838 40014 -262
rect 19914 -922 20378 -888
rect 20932 -922 21396 -888
rect 21950 -922 22414 -888
rect 22968 -922 23432 -888
rect 23986 -922 24450 -888
rect 25004 -922 25468 -888
rect 26022 -922 26486 -888
rect 27040 -922 27504 -888
rect 28058 -922 28522 -888
rect 29076 -922 29540 -888
rect 30094 -922 30558 -888
rect 31112 -922 31576 -888
rect 32130 -922 32594 -888
rect 33148 -922 33612 -888
rect 34166 -922 34630 -888
rect 35184 -922 35648 -888
rect 36202 -922 36666 -888
rect 37220 -922 37684 -888
rect 38238 -922 38702 -888
rect 39256 -922 39720 -888
rect 41862 -1250 41962 13010
rect 4818 -2142 4880 -2042
rect 4880 -2142 41800 -2042
rect 41800 -2142 41862 -2042
<< metal1 >>
rect 17412 29402 41868 29408
rect 17412 29302 17518 29402
rect 41762 29302 41868 29402
rect 17412 29296 41868 29302
rect 17412 28782 17524 29296
rect 18124 28996 18134 29296
rect 41146 28996 41156 29296
rect 17412 15352 17418 28782
rect 17518 15352 17524 28782
rect 21038 28914 37918 28946
rect 21038 28700 21101 28914
rect 37886 28700 37918 28914
rect 21038 28678 21088 28700
rect 21148 28678 21524 28700
rect 21584 28678 21962 28700
rect 22022 28678 22396 28700
rect 22456 28680 37918 28700
rect 41756 28782 41868 29296
rect 22456 28678 25392 28680
rect 25552 27204 25612 28680
rect 27588 27204 27648 28680
rect 28092 27204 28152 28680
rect 28600 27204 28660 28680
rect 29112 27204 29172 28680
rect 29626 27204 29686 28680
rect 31658 27204 31718 28680
rect 33698 27204 33758 28680
rect 34188 27204 34248 28680
rect 34708 27204 34768 28680
rect 35216 27204 35276 28680
rect 35730 27204 35790 28680
rect 37766 27204 37826 28680
rect 25552 27144 37826 27204
rect 25020 26938 25026 26998
rect 25086 26938 25092 26998
rect 23514 26722 24592 26782
rect 23514 26542 23574 26722
rect 24018 26641 24078 26722
rect 23810 26635 24298 26641
rect 23810 26601 23822 26635
rect 24286 26601 24298 26635
rect 23810 26595 24298 26601
rect 23514 26502 23528 26542
rect 23522 25966 23528 26502
rect 23562 26502 23574 26542
rect 24532 26542 24592 26722
rect 25026 26641 25086 26938
rect 25552 26752 25612 27144
rect 26102 26938 26108 26998
rect 26168 26938 26174 26998
rect 27060 26938 27066 26998
rect 27126 26938 27132 26998
rect 25546 26692 25552 26752
rect 25612 26692 25618 26752
rect 24828 26635 25316 26641
rect 24828 26601 24840 26635
rect 25304 26601 25316 26635
rect 24828 26595 25316 26601
rect 24532 26516 24546 26542
rect 23562 25966 23568 26502
rect 24540 26002 24546 26516
rect 23522 25954 23568 25966
rect 24534 25966 24546 26002
rect 24580 26516 24592 26542
rect 25552 26542 25612 26692
rect 26108 26641 26168 26938
rect 27066 26641 27126 26938
rect 27588 26752 27648 27144
rect 27582 26692 27588 26752
rect 27648 26692 27654 26752
rect 25846 26635 26334 26641
rect 25846 26601 25858 26635
rect 26322 26601 26334 26635
rect 25846 26595 26334 26601
rect 26864 26635 27352 26641
rect 26864 26601 26876 26635
rect 27340 26601 27352 26635
rect 26864 26595 27352 26601
rect 27066 26592 27126 26595
rect 25552 26518 25564 26542
rect 24580 26002 24586 26516
rect 25558 26006 25564 26518
rect 24580 25966 24594 26002
rect 23810 25907 24298 25913
rect 23810 25873 23822 25907
rect 24286 25873 24298 25907
rect 23810 25867 24298 25873
rect 24534 25820 24594 25966
rect 25554 25966 25564 26006
rect 25598 26518 25612 26542
rect 26576 26542 26622 26554
rect 25598 26006 25604 26518
rect 25598 25966 25614 26006
rect 26576 25994 26582 26542
rect 25038 25913 25098 25914
rect 24828 25907 25316 25913
rect 24828 25873 24840 25907
rect 25304 25873 25316 25907
rect 24828 25867 25316 25873
rect 23364 25760 23370 25820
rect 23430 25760 23436 25820
rect 24528 25760 24534 25820
rect 24594 25760 24600 25820
rect 23234 25556 23240 25616
rect 23300 25556 23306 25616
rect 21226 23372 21232 23432
rect 21292 23372 21298 23432
rect 19054 20056 20276 20116
rect 19054 18140 19114 20056
rect 19196 19892 19256 20056
rect 19708 19991 19768 20056
rect 19492 19985 19980 19991
rect 19492 19951 19504 19985
rect 19968 19951 19980 19985
rect 19492 19945 19980 19951
rect 19196 19842 19210 19892
rect 19204 19316 19210 19842
rect 19244 19842 19256 19892
rect 20216 19892 20276 20056
rect 20510 19985 20998 19991
rect 20510 19951 20522 19985
rect 20986 19951 20998 19985
rect 20510 19945 20998 19951
rect 19244 19316 19250 19842
rect 20216 19840 20228 19892
rect 19204 19304 19250 19316
rect 20222 19316 20228 19840
rect 20262 19840 20276 19892
rect 21232 19892 21292 23372
rect 23240 23000 23300 25556
rect 23370 23146 23430 25760
rect 24528 25556 24534 25616
rect 24594 25556 24600 25616
rect 23810 25499 24298 25505
rect 23810 25465 23822 25499
rect 24286 25465 24298 25499
rect 23810 25459 24298 25465
rect 23522 25406 23568 25418
rect 23522 24866 23528 25406
rect 23516 24830 23528 24866
rect 23562 24866 23568 25406
rect 24534 25406 24594 25556
rect 25038 25505 25098 25867
rect 24828 25499 25316 25505
rect 24828 25465 24840 25499
rect 25304 25465 25316 25499
rect 24828 25459 25316 25465
rect 25038 25456 25098 25459
rect 24534 25368 24546 25406
rect 23562 24830 23576 24866
rect 24540 24860 24546 25368
rect 23516 24680 23576 24830
rect 24534 24830 24546 24860
rect 24580 25368 24594 25406
rect 25554 25406 25614 25966
rect 26570 25966 26582 25994
rect 26616 25994 26622 26542
rect 27588 26542 27648 26692
rect 28092 26641 28152 27144
rect 27882 26635 28370 26641
rect 27882 26601 27894 26635
rect 28358 26601 28370 26635
rect 27882 26595 28370 26601
rect 27588 26518 27600 26542
rect 27594 26024 27600 26518
rect 26616 25966 26630 25994
rect 25846 25907 26334 25913
rect 25846 25873 25858 25907
rect 26322 25873 26334 25907
rect 25846 25867 26334 25873
rect 26570 25716 26630 25966
rect 27578 25966 27600 26024
rect 27634 26518 27648 26542
rect 28600 26542 28660 27144
rect 29112 26641 29172 27144
rect 29626 26754 29686 27144
rect 30124 26938 30130 26998
rect 30190 26938 30196 26998
rect 31142 26938 31148 26998
rect 31208 26938 31214 26998
rect 29620 26694 29626 26754
rect 29686 26694 29692 26754
rect 28900 26635 29388 26641
rect 28900 26601 28912 26635
rect 29376 26601 29388 26635
rect 28900 26595 29388 26601
rect 27634 26024 27640 26518
rect 28600 26472 28618 26542
rect 27634 25966 27642 26024
rect 26864 25907 27352 25913
rect 26864 25873 26876 25907
rect 27340 25873 27352 25907
rect 26864 25867 27352 25873
rect 26564 25656 26570 25716
rect 26630 25656 26636 25716
rect 25846 25499 26334 25505
rect 25846 25465 25858 25499
rect 26322 25465 26334 25499
rect 25846 25459 26334 25465
rect 26864 25499 27352 25505
rect 26864 25465 26876 25499
rect 27340 25465 27352 25499
rect 26864 25459 27352 25465
rect 24580 24860 24586 25368
rect 25554 25366 25564 25406
rect 24580 24830 24594 24860
rect 25558 24856 25564 25366
rect 23810 24771 24298 24777
rect 23810 24737 23822 24771
rect 24286 24737 24298 24771
rect 23810 24731 24298 24737
rect 24028 24680 24088 24731
rect 24534 24680 24594 24830
rect 25550 24830 25564 24856
rect 25598 25366 25614 25406
rect 26576 25406 26622 25418
rect 25598 24856 25604 25366
rect 25598 24830 25610 24856
rect 26576 24850 26582 25406
rect 25020 24777 25080 24784
rect 24828 24771 25316 24777
rect 24828 24737 24840 24771
rect 25304 24737 25316 24771
rect 24828 24731 25316 24737
rect 23516 24620 24594 24680
rect 24528 24476 24588 24478
rect 23518 24416 24588 24476
rect 23518 24270 23578 24416
rect 24028 24369 24088 24416
rect 23810 24363 24298 24369
rect 23810 24329 23822 24363
rect 24286 24329 24298 24363
rect 23810 24323 24298 24329
rect 23518 24238 23528 24270
rect 23522 23694 23528 24238
rect 23562 24238 23578 24270
rect 24528 24270 24588 24416
rect 25020 24466 25080 24731
rect 25020 24369 25080 24406
rect 25550 24684 25610 24830
rect 26568 24830 26582 24850
rect 26616 24850 26622 25406
rect 27578 25406 27642 25966
rect 28612 25966 28618 26472
rect 28652 26472 28660 26542
rect 29626 26542 29686 26694
rect 30130 26641 30190 26938
rect 31148 26641 31208 26938
rect 31658 26754 31718 27144
rect 32166 26938 32172 26998
rect 32232 26938 32238 26998
rect 33178 26938 33184 26998
rect 33244 26938 33250 26998
rect 31650 26694 31656 26754
rect 31716 26694 31722 26754
rect 29918 26635 30406 26641
rect 29918 26601 29930 26635
rect 30394 26601 30406 26635
rect 29918 26595 30406 26601
rect 30936 26635 31424 26641
rect 30936 26601 30948 26635
rect 31412 26601 31424 26635
rect 30936 26595 31424 26601
rect 29626 26502 29636 26542
rect 28652 25966 28658 26472
rect 29630 26020 29636 26502
rect 28612 25954 28658 25966
rect 29614 25966 29636 26020
rect 29670 26502 29686 26542
rect 30648 26542 30694 26554
rect 29670 26020 29676 26502
rect 29670 25966 29678 26020
rect 30648 26006 30654 26542
rect 27882 25907 28370 25913
rect 27882 25873 27894 25907
rect 28358 25873 28370 25907
rect 27882 25867 28370 25873
rect 28900 25907 29388 25913
rect 28900 25873 28912 25907
rect 29376 25873 29388 25907
rect 28900 25867 29388 25873
rect 28600 25656 28606 25716
rect 28666 25656 28672 25716
rect 27882 25499 28370 25505
rect 27882 25465 27894 25499
rect 28358 25465 28370 25499
rect 27882 25459 28370 25465
rect 27578 25376 27600 25406
rect 27594 24858 27600 25376
rect 26616 24830 26628 24850
rect 26048 24777 26108 24778
rect 25846 24771 26334 24777
rect 25846 24737 25858 24771
rect 26322 24737 26334 24771
rect 25846 24731 26334 24737
rect 26048 24684 26108 24731
rect 26568 24684 26628 24830
rect 27586 24830 27600 24858
rect 27634 25376 27642 25406
rect 28606 25406 28666 25656
rect 28900 25499 29388 25505
rect 28900 25465 28912 25499
rect 29376 25465 29388 25499
rect 28900 25459 29388 25465
rect 27634 24858 27640 25376
rect 28606 25368 28618 25406
rect 28612 24866 28618 25368
rect 27634 24856 27646 24858
rect 27634 24830 27650 24856
rect 27076 24777 27136 24782
rect 26864 24771 27352 24777
rect 26864 24737 26876 24771
rect 27340 24737 27352 24771
rect 26864 24731 27352 24737
rect 27076 24684 27136 24731
rect 25550 24682 27136 24684
rect 27586 24682 27650 24830
rect 28604 24830 28618 24866
rect 28652 25368 28666 25406
rect 29614 25406 29678 25966
rect 30644 25966 30654 26006
rect 30688 26006 30694 26542
rect 31658 26542 31718 26694
rect 32172 26641 32232 26938
rect 33184 26641 33244 26938
rect 33698 26756 33758 27144
rect 33692 26696 33698 26756
rect 33758 26696 33764 26756
rect 31954 26635 32442 26641
rect 31954 26601 31966 26635
rect 32430 26601 32442 26635
rect 31954 26595 32442 26601
rect 32972 26635 33460 26641
rect 32972 26601 32984 26635
rect 33448 26601 33460 26635
rect 32972 26595 33460 26601
rect 31658 26502 31672 26542
rect 31666 26022 31672 26502
rect 30688 25966 30704 26006
rect 30132 25913 30192 25916
rect 29918 25907 30406 25913
rect 29918 25873 29930 25907
rect 30394 25873 30406 25907
rect 29918 25867 30406 25873
rect 30132 25505 30192 25867
rect 30644 25820 30704 25966
rect 31656 25966 31672 26022
rect 31706 26502 31718 26542
rect 32684 26542 32730 26554
rect 31706 26022 31712 26502
rect 31706 25966 31720 26022
rect 32684 26004 32690 26542
rect 31150 25913 31210 25922
rect 30936 25907 31424 25913
rect 30936 25873 30948 25907
rect 31412 25873 31424 25907
rect 30936 25867 31424 25873
rect 30638 25760 30644 25820
rect 30704 25760 30710 25820
rect 30634 25556 30640 25616
rect 30700 25556 30706 25616
rect 29918 25499 30406 25505
rect 29918 25465 29930 25499
rect 30394 25465 30406 25499
rect 29918 25459 30406 25465
rect 30132 25458 30192 25459
rect 29614 25372 29636 25406
rect 28652 24866 28658 25368
rect 29630 24866 29636 25372
rect 28652 24830 28668 24866
rect 27882 24771 28370 24777
rect 27882 24737 27894 24771
rect 28358 24737 28370 24771
rect 27882 24731 28370 24737
rect 25550 24624 27076 24682
rect 24828 24363 25316 24369
rect 24828 24329 24840 24363
rect 25304 24329 25316 24363
rect 24828 24323 25316 24329
rect 24528 24238 24546 24270
rect 23562 23694 23568 24238
rect 24540 23736 24546 24238
rect 23522 23682 23568 23694
rect 24528 23694 24546 23736
rect 24580 24238 24588 24270
rect 25550 24270 25610 24624
rect 27580 24622 27586 24682
rect 27646 24622 27652 24682
rect 27076 24616 27136 24622
rect 26562 24520 26568 24584
rect 26632 24520 26638 24584
rect 26052 24406 26058 24466
rect 26118 24406 26124 24466
rect 26568 24426 26632 24520
rect 26058 24369 26118 24406
rect 25846 24363 26334 24369
rect 25846 24329 25858 24363
rect 26322 24329 26334 24363
rect 25846 24323 26334 24329
rect 24580 23736 24586 24238
rect 25550 24218 25564 24270
rect 24580 23694 24592 23736
rect 25558 23730 25564 24218
rect 23810 23635 24298 23641
rect 23810 23601 23822 23635
rect 24286 23601 24298 23635
rect 23810 23595 24298 23601
rect 24528 23486 24592 23694
rect 25550 23694 25564 23730
rect 25598 24218 25610 24270
rect 26568 24270 26634 24426
rect 27064 24406 27070 24466
rect 27130 24406 27136 24466
rect 27070 24369 27130 24406
rect 26864 24363 27352 24369
rect 26864 24329 26876 24363
rect 27340 24329 27352 24363
rect 26864 24323 27352 24329
rect 27070 24322 27130 24323
rect 26568 24220 26582 24270
rect 25598 23730 25604 24218
rect 25598 23694 25610 23730
rect 26576 23718 26582 24220
rect 24828 23635 25316 23641
rect 24828 23601 24840 23635
rect 25304 23601 25316 23635
rect 24828 23595 25316 23601
rect 24084 23426 24592 23486
rect 23364 23086 23370 23146
rect 23430 23086 23436 23146
rect 23240 22940 23660 23000
rect 23600 20128 23660 22940
rect 23720 20678 23726 20738
rect 23786 20678 23792 20738
rect 22250 20060 23460 20120
rect 23594 20068 23600 20128
rect 23660 20068 23666 20128
rect 21528 19985 22016 19991
rect 21528 19951 21540 19985
rect 22004 19951 22016 19985
rect 21528 19945 22016 19951
rect 20262 19316 20268 19840
rect 20222 19304 20268 19316
rect 21232 19316 21246 19892
rect 21280 19316 21292 19892
rect 22250 19892 22310 20060
rect 22762 19991 22822 20060
rect 22546 19985 23034 19991
rect 22546 19951 22558 19985
rect 23022 19951 23034 19985
rect 22546 19945 23034 19951
rect 22250 19844 22264 19892
rect 19492 19257 19980 19263
rect 19492 19223 19504 19257
rect 19968 19223 19980 19257
rect 19492 19217 19980 19223
rect 20510 19257 20998 19263
rect 20510 19223 20522 19257
rect 20986 19223 20998 19257
rect 20510 19217 20998 19223
rect 20716 19174 20776 19217
rect 20710 19114 20716 19174
rect 20776 19114 20782 19174
rect 20818 19002 20824 19062
rect 20884 19002 20890 19062
rect 20824 18959 20884 19002
rect 19492 18953 19980 18959
rect 19492 18919 19504 18953
rect 19968 18919 19980 18953
rect 19492 18913 19980 18919
rect 20510 18953 20998 18959
rect 20510 18919 20522 18953
rect 20986 18919 20998 18953
rect 20510 18913 20998 18919
rect 19204 18860 19250 18872
rect 19204 18342 19210 18860
rect 19194 18284 19210 18342
rect 19244 18342 19250 18860
rect 20222 18860 20268 18872
rect 19244 18284 19254 18342
rect 20222 18334 20228 18860
rect 19048 18080 19054 18140
rect 19114 18080 19120 18140
rect 18928 17052 18988 17058
rect 19054 17052 19114 18080
rect 19194 18030 19254 18284
rect 20214 18284 20228 18334
rect 20262 18334 20268 18860
rect 21232 18860 21292 19316
rect 22258 19316 22264 19844
rect 22298 19844 22310 19892
rect 23268 19892 23328 20060
rect 23268 19846 23282 19892
rect 22298 19316 22304 19844
rect 22258 19304 22304 19316
rect 23276 19316 23282 19846
rect 23316 19846 23328 19892
rect 23316 19316 23322 19846
rect 23276 19304 23322 19316
rect 21528 19257 22016 19263
rect 21528 19223 21540 19257
rect 22004 19223 22016 19257
rect 21528 19217 22016 19223
rect 22546 19257 23034 19263
rect 22546 19223 22558 19257
rect 23022 19223 23034 19257
rect 22546 19217 23034 19223
rect 21608 19062 21668 19217
rect 21732 19114 21738 19174
rect 21798 19114 21804 19174
rect 21602 19002 21608 19062
rect 21668 19002 21674 19062
rect 21738 18959 21798 19114
rect 21528 18953 22016 18959
rect 21528 18919 21540 18953
rect 22004 18919 22016 18953
rect 21528 18913 22016 18919
rect 22546 18953 23034 18959
rect 22546 18919 22558 18953
rect 23022 18919 23034 18953
rect 22546 18913 23034 18919
rect 20262 18284 20274 18334
rect 19492 18225 19980 18231
rect 19492 18191 19504 18225
rect 19968 18191 19980 18225
rect 19492 18185 19980 18191
rect 19696 18030 19756 18185
rect 20214 18030 20274 18284
rect 21232 18284 21246 18860
rect 21280 18284 21292 18860
rect 22258 18860 22304 18872
rect 22258 18370 22264 18860
rect 20510 18225 20998 18231
rect 20510 18191 20522 18225
rect 20986 18191 20998 18225
rect 20510 18185 20998 18191
rect 19194 17970 20214 18030
rect 20274 17970 20280 18030
rect 19194 17828 19254 17970
rect 19696 17927 19756 17970
rect 19492 17921 19980 17927
rect 19492 17887 19504 17921
rect 19968 17887 19980 17921
rect 19492 17881 19980 17887
rect 19194 17768 19210 17828
rect 19204 17252 19210 17768
rect 19244 17768 19254 17828
rect 20214 17828 20274 17970
rect 20724 17927 20784 18185
rect 20510 17921 20998 17927
rect 20510 17887 20522 17921
rect 20986 17887 20998 17921
rect 20510 17881 20998 17887
rect 19244 17252 19250 17768
rect 20214 17764 20228 17828
rect 19204 17240 19250 17252
rect 20222 17252 20228 17764
rect 20262 17764 20274 17828
rect 21232 17828 21292 18284
rect 22248 18284 22264 18370
rect 22298 18370 22304 18860
rect 23276 18860 23322 18872
rect 22298 18284 22308 18370
rect 23276 18330 23282 18860
rect 21528 18225 22016 18231
rect 21528 18191 21540 18225
rect 22004 18191 22016 18225
rect 21528 18185 22016 18191
rect 21742 17927 21802 18185
rect 22248 18140 22308 18284
rect 23268 18284 23282 18330
rect 23316 18330 23322 18860
rect 23316 18284 23328 18330
rect 22546 18225 23034 18231
rect 22546 18191 22558 18225
rect 23022 18191 23034 18225
rect 22546 18185 23034 18191
rect 22762 18140 22822 18185
rect 23268 18140 23328 18284
rect 22242 18080 22248 18140
rect 22308 18080 23328 18140
rect 21528 17921 22016 17927
rect 21528 17887 21540 17921
rect 22004 17887 22016 17921
rect 21528 17881 22016 17887
rect 20262 17252 20268 17764
rect 20222 17240 20268 17252
rect 21232 17252 21246 17828
rect 21280 17252 21292 17828
rect 22248 17828 22308 18080
rect 22762 17927 22822 18080
rect 22546 17921 23034 17927
rect 22546 17887 22558 17921
rect 23022 17887 23034 17921
rect 22546 17881 23034 17887
rect 22248 17772 22264 17828
rect 19492 17193 19980 17199
rect 19492 17159 19504 17193
rect 19968 17159 19980 17193
rect 19492 17153 19980 17159
rect 20510 17193 20998 17199
rect 20510 17159 20522 17193
rect 20986 17159 20998 17193
rect 20510 17153 20998 17159
rect 20730 17106 20790 17153
rect 18988 16992 20278 17052
rect 20724 17046 20730 17106
rect 20790 17046 20796 17106
rect 18928 16986 18988 16992
rect 19192 16796 19252 16992
rect 19700 16895 19760 16992
rect 19492 16889 19980 16895
rect 19492 16855 19504 16889
rect 19968 16855 19980 16889
rect 19492 16849 19980 16855
rect 19192 16744 19210 16796
rect 19204 16220 19210 16744
rect 19244 16744 19252 16796
rect 20218 16796 20278 16992
rect 20830 16946 20836 17006
rect 20896 16946 20902 17006
rect 20836 16895 20896 16946
rect 20510 16889 20998 16895
rect 20510 16855 20522 16889
rect 20986 16855 20998 16889
rect 20510 16849 20998 16855
rect 20218 16748 20228 16796
rect 19244 16220 19250 16744
rect 19204 16208 19250 16220
rect 20222 16220 20228 16748
rect 20262 16748 20278 16796
rect 21232 16796 21292 17252
rect 22258 17252 22264 17772
rect 22298 17772 22308 17828
rect 23268 17828 23328 18080
rect 23400 18030 23460 20060
rect 23394 17970 23400 18030
rect 23460 17970 23466 18030
rect 23268 17792 23282 17828
rect 22298 17252 22304 17772
rect 22258 17240 22304 17252
rect 23276 17252 23282 17792
rect 23316 17792 23328 17828
rect 23316 17252 23322 17792
rect 23276 17240 23322 17252
rect 21528 17193 22016 17199
rect 21528 17159 21540 17193
rect 22004 17159 22016 17193
rect 21528 17153 22016 17159
rect 22546 17193 23034 17199
rect 22546 17159 22558 17193
rect 23022 17159 23034 17193
rect 22546 17153 23034 17159
rect 21622 17006 21682 17153
rect 21734 17046 21740 17106
rect 21800 17046 21806 17106
rect 23400 17052 23460 17970
rect 23586 17842 23592 17902
rect 23652 17842 23658 17902
rect 21616 16946 21622 17006
rect 21682 16946 21688 17006
rect 21740 16895 21800 17046
rect 22248 16992 23460 17052
rect 21528 16889 22016 16895
rect 21528 16855 21540 16889
rect 22004 16855 22016 16889
rect 21528 16849 22016 16855
rect 20262 16220 20268 16748
rect 21232 16722 21246 16796
rect 20222 16208 20268 16220
rect 21240 16220 21246 16722
rect 21280 16722 21292 16796
rect 22248 16796 22308 16992
rect 22750 16895 22810 16992
rect 22546 16889 23034 16895
rect 22546 16855 22558 16889
rect 23022 16855 23034 16889
rect 22546 16849 23034 16855
rect 22248 16766 22264 16796
rect 21280 16220 21286 16722
rect 22258 16302 22264 16766
rect 21240 16208 21286 16220
rect 22250 16220 22264 16302
rect 22298 16766 22308 16796
rect 23268 16796 23328 16992
rect 22298 16302 22304 16766
rect 23268 16728 23282 16796
rect 22298 16220 22310 16302
rect 21728 16167 21788 16171
rect 19492 16161 19980 16167
rect 19492 16127 19504 16161
rect 19968 16127 19980 16161
rect 19492 16121 19980 16127
rect 20510 16161 20998 16167
rect 20510 16127 20522 16161
rect 20986 16127 20998 16161
rect 20510 16121 20998 16127
rect 21528 16161 22016 16167
rect 21528 16127 21540 16161
rect 22004 16127 22016 16161
rect 21528 16121 22016 16127
rect 18442 15996 18502 16002
rect 20722 15996 20782 16121
rect 18502 15936 20782 15996
rect 18442 15930 18502 15936
rect 18582 15820 18642 15826
rect 21728 15820 21788 16121
rect 18642 15760 21788 15820
rect 18582 15754 18642 15760
rect 19482 15646 19542 15652
rect 22250 15646 22310 16220
rect 23276 16220 23282 16728
rect 23316 16728 23328 16796
rect 23316 16220 23322 16728
rect 23276 16208 23322 16220
rect 22546 16161 23034 16167
rect 22546 16127 22558 16161
rect 23022 16127 23034 16161
rect 22546 16121 23034 16127
rect 19542 15586 22310 15646
rect 19482 15580 19542 15586
rect 18322 15496 18382 15502
rect 23592 15496 23652 17842
rect 23726 16750 23786 20678
rect 23836 20068 23842 20128
rect 23902 20068 23908 20128
rect 23842 18006 23902 20068
rect 24084 19164 24144 23426
rect 24528 23296 24592 23426
rect 24522 23232 24528 23296
rect 24592 23232 24598 23296
rect 24352 23146 24412 23152
rect 24352 20210 24412 23086
rect 25030 23040 25090 23595
rect 25550 23544 25610 23694
rect 26566 23694 26582 23718
rect 26616 24224 26634 24270
rect 27586 24270 27650 24622
rect 28080 24474 28140 24731
rect 28604 24584 28668 24830
rect 29620 24830 29636 24866
rect 29670 25372 29678 25406
rect 30640 25406 30700 25556
rect 31150 25505 31210 25867
rect 30936 25499 31424 25505
rect 30936 25465 30948 25499
rect 31412 25465 31424 25499
rect 30936 25459 31424 25465
rect 30640 25380 30654 25406
rect 29670 24866 29676 25372
rect 29670 24864 29680 24866
rect 29670 24830 29684 24864
rect 28900 24771 29388 24777
rect 28900 24737 28912 24771
rect 29376 24737 29388 24771
rect 28900 24731 29388 24737
rect 28438 24520 28444 24584
rect 28508 24520 28668 24584
rect 29104 24474 29164 24731
rect 29620 24682 29684 24830
rect 30648 24830 30654 25380
rect 30688 25380 30700 25406
rect 31656 25406 31720 25966
rect 32678 25966 32690 26004
rect 32724 26004 32730 26542
rect 33698 26542 33758 26696
rect 34188 26641 34248 27144
rect 34708 26756 34768 27144
rect 34702 26696 34708 26756
rect 34768 26696 34774 26756
rect 33990 26635 34478 26641
rect 33990 26601 34002 26635
rect 34466 26601 34478 26635
rect 33990 26595 34478 26601
rect 33698 26504 33708 26542
rect 33702 26006 33708 26504
rect 32724 25966 32738 26004
rect 32166 25913 32226 25919
rect 31954 25907 32442 25913
rect 31954 25873 31966 25907
rect 32430 25873 32442 25907
rect 31954 25867 32442 25873
rect 32166 25505 32226 25867
rect 32678 25820 32738 25966
rect 33694 25966 33708 26006
rect 33742 26504 33758 26542
rect 34708 26542 34768 26696
rect 35216 26641 35276 27144
rect 35730 26756 35790 27144
rect 36236 26938 36242 26998
rect 36302 26938 36308 26998
rect 37248 26938 37254 26998
rect 37314 26938 37320 26998
rect 35724 26696 35730 26756
rect 35790 26696 35796 26756
rect 35008 26635 35496 26641
rect 35008 26601 35020 26635
rect 35484 26601 35496 26635
rect 35008 26595 35496 26601
rect 35216 26592 35276 26595
rect 33742 26006 33748 26504
rect 34708 26472 34726 26542
rect 33742 25966 33758 26006
rect 33178 25913 33238 25919
rect 32972 25907 33460 25913
rect 32972 25873 32984 25907
rect 33448 25873 33460 25907
rect 32972 25867 33460 25873
rect 32672 25760 32678 25820
rect 32738 25760 32744 25820
rect 33178 25616 33238 25867
rect 32670 25556 32676 25616
rect 32736 25556 32742 25616
rect 33172 25556 33178 25616
rect 33238 25556 33244 25616
rect 31954 25499 32442 25505
rect 31954 25465 31966 25499
rect 32430 25465 32442 25499
rect 31954 25459 32442 25465
rect 32166 25456 32226 25459
rect 30688 24830 30694 25380
rect 31656 25374 31672 25406
rect 31666 24878 31672 25374
rect 30648 24818 30694 24830
rect 31658 24830 31672 24878
rect 31706 25374 31720 25406
rect 32676 25406 32736 25556
rect 33178 25505 33238 25556
rect 32972 25499 33460 25505
rect 32972 25465 32984 25499
rect 33448 25465 33460 25499
rect 32972 25459 33460 25465
rect 33178 25456 33238 25459
rect 32676 25374 32690 25406
rect 31706 24878 31712 25374
rect 31706 24876 31718 24878
rect 31706 24830 31722 24876
rect 32684 24860 32690 25374
rect 30132 24777 30192 24784
rect 29918 24771 30406 24777
rect 29918 24737 29930 24771
rect 30394 24737 30406 24771
rect 29918 24731 30406 24737
rect 30936 24771 31424 24777
rect 30936 24737 30948 24771
rect 31412 24737 31424 24771
rect 30936 24731 31424 24737
rect 29614 24622 29620 24682
rect 29680 24622 29686 24682
rect 28074 24414 28080 24474
rect 28140 24414 28146 24474
rect 29098 24414 29104 24474
rect 29164 24414 29170 24474
rect 27882 24363 28370 24369
rect 27882 24329 27894 24363
rect 28358 24329 28370 24363
rect 27882 24323 28370 24329
rect 28900 24363 29388 24369
rect 28900 24329 28912 24363
rect 29376 24329 29388 24363
rect 28900 24323 29388 24329
rect 26616 24220 26632 24224
rect 27586 24222 27600 24270
rect 26616 23718 26622 24220
rect 27594 23720 27600 24222
rect 26616 23694 26630 23718
rect 25846 23635 26334 23641
rect 25846 23601 25858 23635
rect 26322 23601 26334 23635
rect 25846 23595 26334 23601
rect 25544 23484 25550 23544
rect 25610 23484 25616 23544
rect 26072 23040 26132 23595
rect 26566 23434 26630 23694
rect 27586 23694 27600 23720
rect 27634 24222 27650 24270
rect 28612 24270 28658 24282
rect 27634 23720 27640 24222
rect 28612 23750 28618 24270
rect 27634 23718 27646 23720
rect 27634 23694 27650 23718
rect 26864 23635 27352 23641
rect 26864 23601 26876 23635
rect 27340 23601 27352 23635
rect 26864 23595 27352 23601
rect 26560 23370 26566 23434
rect 26630 23370 26636 23434
rect 27072 23040 27132 23595
rect 27586 23544 27650 23694
rect 28606 23694 28618 23750
rect 28652 23750 28658 24270
rect 29620 24270 29684 24622
rect 30132 24474 30192 24731
rect 30126 24414 30132 24474
rect 30192 24414 30198 24474
rect 30132 24369 30192 24414
rect 31160 24369 31220 24731
rect 31658 24680 31722 24830
rect 32678 24830 32690 24860
rect 32724 25374 32736 25406
rect 33694 25406 33758 25966
rect 34720 25966 34726 26472
rect 34760 26472 34768 26542
rect 35730 26542 35790 26696
rect 36242 26641 36302 26938
rect 37254 26641 37314 26938
rect 37766 26756 37826 27144
rect 38266 26938 38272 26998
rect 38332 26938 38338 26998
rect 37760 26696 37766 26756
rect 37826 26696 37832 26756
rect 36026 26635 36514 26641
rect 36026 26601 36038 26635
rect 36502 26601 36514 26635
rect 36026 26595 36514 26601
rect 37044 26635 37532 26641
rect 37044 26601 37056 26635
rect 37520 26601 37532 26635
rect 37044 26595 37532 26601
rect 35730 26514 35744 26542
rect 34760 25966 34766 26472
rect 35738 26014 35744 26514
rect 34720 25954 34766 25966
rect 35730 25966 35744 26014
rect 35778 26514 35790 26542
rect 36756 26542 36802 26554
rect 35778 26014 35784 26514
rect 35778 25966 35790 26014
rect 36756 25998 36762 26542
rect 33990 25907 34478 25913
rect 33990 25873 34002 25907
rect 34466 25873 34478 25907
rect 33990 25867 34478 25873
rect 35008 25907 35496 25913
rect 35008 25873 35020 25907
rect 35484 25873 35496 25907
rect 35008 25867 35496 25873
rect 34706 25656 34712 25716
rect 34772 25656 34778 25716
rect 34192 25556 34198 25616
rect 34258 25556 34264 25616
rect 34198 25505 34258 25556
rect 33990 25499 34478 25505
rect 33990 25465 34002 25499
rect 34466 25465 34478 25499
rect 33990 25459 34478 25465
rect 32724 24860 32730 25374
rect 33694 25358 33708 25406
rect 33702 24874 33708 25358
rect 32724 24830 32738 24860
rect 32178 24777 32238 24789
rect 31954 24771 32442 24777
rect 31954 24737 31966 24771
rect 32430 24737 32442 24771
rect 31954 24731 32442 24737
rect 31652 24620 31658 24680
rect 31718 24620 31724 24680
rect 29918 24363 30406 24369
rect 29918 24329 29930 24363
rect 30394 24329 30406 24363
rect 29918 24323 30406 24329
rect 30936 24363 31424 24369
rect 30936 24329 30948 24363
rect 31412 24329 31424 24363
rect 30936 24323 31424 24329
rect 31160 24316 31220 24323
rect 29620 24210 29636 24270
rect 28652 23694 28666 23750
rect 29630 23728 29636 24210
rect 28108 23641 28168 23644
rect 27882 23635 28370 23641
rect 27882 23601 27894 23635
rect 28358 23601 28370 23635
rect 27882 23595 28370 23601
rect 28108 23544 28168 23595
rect 28606 23544 28666 23694
rect 29620 23694 29636 23728
rect 29670 24210 29684 24270
rect 30648 24270 30694 24282
rect 29670 23728 29676 24210
rect 29670 23726 29680 23728
rect 30648 23726 30654 24270
rect 29670 23694 29684 23726
rect 28900 23635 29388 23641
rect 28900 23601 28912 23635
rect 29376 23601 29388 23635
rect 28900 23595 29388 23601
rect 27580 23484 27586 23544
rect 27646 23484 27652 23544
rect 28102 23484 28108 23544
rect 28168 23484 28174 23544
rect 28600 23484 28606 23544
rect 28666 23484 28672 23544
rect 29080 23540 29140 23595
rect 29620 23548 29684 23694
rect 30638 23694 30654 23726
rect 30688 23726 30694 24270
rect 31658 24270 31722 24620
rect 32178 24369 32238 24731
rect 32678 24582 32738 24830
rect 33694 24830 33708 24874
rect 33742 25358 33758 25406
rect 34712 25406 34772 25656
rect 35218 25556 35224 25616
rect 35284 25556 35290 25616
rect 35730 25612 35790 25966
rect 36746 25966 36762 25998
rect 36796 25998 36802 26542
rect 37766 26542 37826 26696
rect 38272 26641 38332 26938
rect 38786 26704 39866 26764
rect 38062 26635 38550 26641
rect 38062 26601 38074 26635
rect 38538 26601 38550 26635
rect 38062 26595 38550 26601
rect 37766 26510 37780 26542
rect 37774 26004 37780 26510
rect 36796 25966 36806 25998
rect 36026 25907 36514 25913
rect 36026 25873 36038 25907
rect 36502 25873 36514 25907
rect 36026 25867 36514 25873
rect 36746 25716 36806 25966
rect 37770 25966 37780 26004
rect 37814 26510 37826 26542
rect 38786 26542 38846 26704
rect 39288 26641 39348 26704
rect 39080 26635 39568 26641
rect 39080 26601 39092 26635
rect 39556 26601 39568 26635
rect 39080 26595 39568 26601
rect 38786 26512 38798 26542
rect 37814 26004 37820 26510
rect 38792 26006 38798 26512
rect 37814 25966 37830 26004
rect 37044 25907 37532 25913
rect 37044 25873 37056 25907
rect 37520 25873 37532 25907
rect 37044 25867 37532 25873
rect 36740 25656 36746 25716
rect 36806 25656 36812 25716
rect 37770 25618 37830 25966
rect 38786 25966 38798 26006
rect 38832 26512 38846 26542
rect 39806 26542 39866 26704
rect 38832 26006 38838 26512
rect 39806 26496 39816 26542
rect 38832 25966 38846 26006
rect 38250 25913 38310 25925
rect 38062 25907 38550 25913
rect 38062 25873 38074 25907
rect 38538 25873 38550 25907
rect 38062 25867 38550 25873
rect 37770 25612 37834 25618
rect 35224 25505 35284 25556
rect 35724 25552 35730 25612
rect 35790 25552 35796 25612
rect 36238 25552 36244 25612
rect 36304 25552 36310 25612
rect 36742 25552 36748 25612
rect 36808 25552 36814 25612
rect 37248 25552 37254 25612
rect 37314 25552 37320 25612
rect 37770 25552 37774 25612
rect 35008 25499 35496 25505
rect 35008 25465 35020 25499
rect 35484 25465 35496 25499
rect 35008 25459 35496 25465
rect 34712 25382 34726 25406
rect 33742 24874 33748 25358
rect 33742 24872 33754 24874
rect 33742 24830 33758 24872
rect 33178 24777 33238 24785
rect 32972 24771 33460 24777
rect 32972 24737 32984 24771
rect 33448 24737 33460 24771
rect 32972 24731 33460 24737
rect 32672 24522 32678 24582
rect 32738 24522 32744 24582
rect 33178 24369 33238 24731
rect 33694 24680 33758 24830
rect 34720 24830 34726 25382
rect 34760 25382 34772 25406
rect 35730 25406 35790 25552
rect 36244 25505 36304 25552
rect 36026 25499 36514 25505
rect 36026 25465 36038 25499
rect 36502 25465 36514 25499
rect 36026 25459 36514 25465
rect 34760 24830 34766 25382
rect 35730 25362 35744 25406
rect 35738 24866 35744 25362
rect 34720 24818 34766 24830
rect 35730 24830 35744 24866
rect 35778 25362 35790 25406
rect 36748 25406 36808 25552
rect 37254 25505 37314 25552
rect 37770 25546 37834 25552
rect 37044 25499 37532 25505
rect 37044 25465 37056 25499
rect 37520 25465 37532 25499
rect 37044 25459 37532 25465
rect 36748 25378 36762 25406
rect 35778 24866 35784 25362
rect 36756 24900 36762 25378
rect 35778 24830 35790 24866
rect 33990 24771 34478 24777
rect 33990 24737 34002 24771
rect 34466 24737 34478 24771
rect 33990 24731 34478 24737
rect 35008 24771 35496 24777
rect 35008 24737 35020 24771
rect 35484 24737 35496 24771
rect 35008 24731 35496 24737
rect 35730 24680 35790 24830
rect 36746 24830 36762 24900
rect 36796 25378 36808 25406
rect 37770 25406 37830 25546
rect 38250 25505 38310 25867
rect 38786 25820 38846 25966
rect 39810 25966 39816 26496
rect 39850 26496 39866 26542
rect 39850 25966 39856 26496
rect 39810 25954 39856 25966
rect 39080 25907 39568 25913
rect 39080 25873 39092 25907
rect 39556 25873 39568 25907
rect 39080 25867 39568 25873
rect 38780 25760 38786 25820
rect 38846 25760 38852 25820
rect 40030 25760 40036 25820
rect 40096 25760 40102 25820
rect 38790 25544 39860 25604
rect 38062 25499 38550 25505
rect 38062 25465 38074 25499
rect 38538 25465 38550 25499
rect 38062 25459 38550 25465
rect 36796 24900 36802 25378
rect 37770 25370 37780 25406
rect 36796 24830 36806 24900
rect 37774 24862 37780 25370
rect 36026 24771 36514 24777
rect 36026 24737 36038 24771
rect 36502 24737 36514 24771
rect 36026 24731 36514 24737
rect 36232 24680 36292 24731
rect 33688 24620 33694 24680
rect 33754 24620 33760 24680
rect 34188 24620 34194 24680
rect 34254 24620 34260 24680
rect 34702 24620 34708 24680
rect 34768 24620 34774 24680
rect 35226 24620 35232 24680
rect 35292 24620 35298 24680
rect 35724 24620 35730 24680
rect 35790 24620 35796 24680
rect 36226 24620 36232 24680
rect 36292 24620 36298 24680
rect 36746 24678 36806 24830
rect 37764 24830 37780 24862
rect 37814 25370 37830 25406
rect 38790 25406 38850 25544
rect 39296 25505 39356 25544
rect 39080 25499 39568 25505
rect 39080 25465 39092 25499
rect 39556 25465 39568 25499
rect 39080 25459 39568 25465
rect 38790 25378 38798 25406
rect 37814 24862 37820 25370
rect 37814 24860 37824 24862
rect 38792 24860 38798 25378
rect 37814 24830 37828 24860
rect 37254 24777 37314 24784
rect 37044 24771 37532 24777
rect 37044 24737 37056 24771
rect 37520 24737 37532 24771
rect 37044 24731 37532 24737
rect 37254 24678 37314 24731
rect 37764 24678 37828 24830
rect 38786 24830 38798 24860
rect 38832 25378 38850 25406
rect 39800 25406 39860 25544
rect 38832 24860 38838 25378
rect 39800 25372 39816 25406
rect 38832 24830 38846 24860
rect 38250 24777 38310 24783
rect 38062 24771 38550 24777
rect 38062 24737 38074 24771
rect 38538 24737 38550 24771
rect 38062 24731 38550 24737
rect 31954 24363 32442 24369
rect 31954 24329 31966 24363
rect 32430 24329 32442 24363
rect 31954 24323 32442 24329
rect 32972 24363 33460 24369
rect 32972 24329 32984 24363
rect 33448 24329 33460 24363
rect 32972 24323 33460 24329
rect 33178 24322 33238 24323
rect 31658 24230 31672 24270
rect 31666 23754 31672 24230
rect 30688 23694 30702 23726
rect 29918 23635 30406 23641
rect 29918 23601 29930 23635
rect 30394 23601 30406 23635
rect 29918 23595 30406 23601
rect 24462 22980 24468 23040
rect 24528 22980 24534 23040
rect 25024 22980 25030 23040
rect 25090 22980 25096 23040
rect 26066 22980 26072 23040
rect 26132 22980 26138 23040
rect 27066 22980 27072 23040
rect 27132 22980 27138 23040
rect 24468 20398 24528 22980
rect 29080 22942 29140 23480
rect 29588 23544 29684 23548
rect 29588 23542 29620 23544
rect 29680 23484 29686 23544
rect 30074 23484 30080 23544
rect 30140 23484 30146 23544
rect 29588 22942 29648 23482
rect 30080 22942 30140 23484
rect 30234 23040 30294 23595
rect 30638 23292 30702 23694
rect 31656 23694 31672 23754
rect 31706 24230 31722 24270
rect 32684 24270 32730 24282
rect 31706 23754 31712 24230
rect 31706 23694 31716 23754
rect 32684 23730 32690 24270
rect 30936 23635 31424 23641
rect 30936 23601 30948 23635
rect 31412 23601 31424 23635
rect 30936 23595 31424 23601
rect 30638 23222 30702 23228
rect 31124 23546 31184 23552
rect 30228 22980 30234 23040
rect 30294 22980 30300 23040
rect 31124 22942 31184 23486
rect 31244 23040 31304 23595
rect 31656 23544 31716 23694
rect 32674 23694 32690 23730
rect 32724 23730 32730 24270
rect 33694 24270 33758 24620
rect 34194 24369 34254 24620
rect 33990 24363 34478 24369
rect 33990 24329 34002 24363
rect 34466 24329 34478 24363
rect 33990 24323 34478 24329
rect 33694 24218 33708 24270
rect 33702 23736 33708 24218
rect 32724 23694 32738 23730
rect 31954 23635 32442 23641
rect 31954 23601 31966 23635
rect 32430 23601 32442 23635
rect 31954 23595 32442 23601
rect 31650 23484 31656 23544
rect 31716 23484 31722 23544
rect 32186 23040 32246 23595
rect 32674 23150 32738 23694
rect 33694 23694 33708 23736
rect 33742 24218 33758 24270
rect 34708 24270 34768 24620
rect 35232 24369 35292 24620
rect 35008 24363 35496 24369
rect 35008 24329 35020 24363
rect 35484 24329 35496 24363
rect 35008 24323 35496 24329
rect 33742 23736 33748 24218
rect 34708 24216 34726 24270
rect 34720 24140 34726 24216
rect 33742 23734 33754 23736
rect 33742 23694 33758 23734
rect 32972 23635 33460 23641
rect 32972 23601 32984 23635
rect 33448 23601 33460 23635
rect 32972 23595 33460 23601
rect 33168 23546 33228 23552
rect 33694 23546 33758 23694
rect 34712 23694 34726 24140
rect 34760 24216 34768 24270
rect 35730 24270 35790 24620
rect 36740 24618 36746 24678
rect 36806 24618 36812 24678
rect 37248 24618 37254 24678
rect 37314 24618 37320 24678
rect 37758 24618 37764 24678
rect 37824 24618 37830 24678
rect 36230 24406 36236 24466
rect 36296 24406 36302 24466
rect 37242 24406 37248 24466
rect 37308 24406 37314 24466
rect 36236 24369 36296 24406
rect 37248 24369 37308 24406
rect 36026 24363 36514 24369
rect 36026 24329 36038 24363
rect 36502 24329 36514 24363
rect 36026 24323 36514 24329
rect 37044 24363 37532 24369
rect 37044 24329 37056 24363
rect 37520 24329 37532 24363
rect 37044 24323 37532 24329
rect 35730 24216 35744 24270
rect 34760 24140 34766 24216
rect 34760 23694 34772 24140
rect 35738 23724 35744 24216
rect 34190 23641 34250 23650
rect 33990 23635 34478 23641
rect 33990 23601 34002 23635
rect 34466 23601 34478 23635
rect 33990 23595 34478 23601
rect 32668 23086 32674 23150
rect 32738 23086 32744 23150
rect 31238 22980 31244 23040
rect 31304 22980 31310 23040
rect 32180 22980 32186 23040
rect 32246 22980 32252 23040
rect 33168 22942 33228 23486
rect 33662 23542 33758 23546
rect 33662 23540 33694 23542
rect 33754 23482 33760 23542
rect 34190 23536 34250 23595
rect 34712 23546 34772 23694
rect 35730 23694 35744 23724
rect 35778 24216 35790 24270
rect 36756 24270 36802 24282
rect 35778 23724 35784 24216
rect 36756 23728 36762 24270
rect 35778 23722 35790 23724
rect 35778 23694 35794 23722
rect 35190 23641 35250 23644
rect 35008 23635 35496 23641
rect 35008 23601 35020 23635
rect 35484 23601 35496 23635
rect 35008 23595 35496 23601
rect 33662 22942 33722 23480
rect 34190 22942 34250 23476
rect 34678 23540 34772 23546
rect 34738 23538 34772 23540
rect 34678 23478 34712 23480
rect 34678 23472 34772 23478
rect 35190 23536 35250 23595
rect 35730 23540 35794 23694
rect 36746 23694 36762 23728
rect 36796 23728 36802 24270
rect 37764 24270 37828 24618
rect 38250 24466 38310 24731
rect 38786 24582 38846 24830
rect 39810 24830 39816 25372
rect 39850 25372 39860 25406
rect 39850 24830 39856 25372
rect 39810 24818 39856 24830
rect 39080 24771 39568 24777
rect 39080 24737 39092 24771
rect 39556 24737 39568 24771
rect 39080 24731 39568 24737
rect 38780 24522 38786 24582
rect 38846 24522 38852 24582
rect 38788 24468 38848 24470
rect 38244 24406 38250 24466
rect 38310 24406 38316 24466
rect 38788 24408 39860 24468
rect 38250 24369 38310 24406
rect 38062 24363 38550 24369
rect 38062 24329 38074 24363
rect 38538 24329 38550 24363
rect 38062 24323 38550 24329
rect 38250 24320 38310 24323
rect 37764 24224 37780 24270
rect 36796 23694 36810 23728
rect 37774 23724 37780 24224
rect 36026 23635 36514 23641
rect 36026 23601 36038 23635
rect 36502 23601 36514 23635
rect 36026 23595 36514 23601
rect 35724 23480 35730 23540
rect 35790 23480 35796 23540
rect 34678 22942 34738 23472
rect 35190 22942 35250 23476
rect 36746 23434 36810 23694
rect 37764 23694 37780 23724
rect 37814 24224 37828 24270
rect 38788 24270 38848 24408
rect 39292 24369 39352 24408
rect 39080 24363 39568 24369
rect 39080 24329 39092 24363
rect 39556 24329 39568 24363
rect 39080 24323 39568 24329
rect 38788 24244 38798 24270
rect 37814 23724 37820 24224
rect 38792 23782 38798 24244
rect 37814 23722 37824 23724
rect 37814 23694 37828 23722
rect 37044 23635 37532 23641
rect 37044 23601 37056 23635
rect 37520 23601 37532 23635
rect 37044 23595 37532 23601
rect 37764 23540 37828 23694
rect 38780 23694 38798 23782
rect 38832 24244 38848 24270
rect 39800 24270 39860 24408
rect 38832 23782 38838 24244
rect 39800 24220 39816 24270
rect 38832 23694 38840 23782
rect 38062 23635 38550 23641
rect 38062 23601 38074 23635
rect 38538 23601 38550 23635
rect 38062 23595 38550 23601
rect 37758 23480 37764 23540
rect 37824 23480 37830 23540
rect 36740 23370 36746 23434
rect 36810 23370 36816 23434
rect 38780 23146 38840 23694
rect 39810 23694 39816 24220
rect 39850 24220 39860 24270
rect 39850 23694 39856 24220
rect 39810 23682 39856 23694
rect 39080 23635 39568 23641
rect 39080 23601 39092 23635
rect 39556 23601 39568 23635
rect 39080 23595 39568 23601
rect 40036 23302 40096 25760
rect 40032 23296 40096 23302
rect 40032 23226 40096 23232
rect 38774 23086 38780 23146
rect 38840 23086 38846 23146
rect 26744 22882 36984 22942
rect 24576 22778 24582 22838
rect 24642 22778 24648 22838
rect 24582 20864 24642 22778
rect 25004 22725 25492 22731
rect 25004 22691 25016 22725
rect 25480 22691 25492 22725
rect 25004 22685 25492 22691
rect 26022 22725 26510 22731
rect 26022 22691 26034 22725
rect 26498 22691 26510 22725
rect 26022 22685 26510 22691
rect 24716 22632 24762 22644
rect 24716 22086 24722 22632
rect 24708 22056 24722 22086
rect 24756 22086 24762 22632
rect 25734 22632 25780 22644
rect 24756 22056 24768 22086
rect 25734 22080 25740 22632
rect 24708 21904 24768 22056
rect 25726 22056 25740 22080
rect 25774 22080 25780 22632
rect 26744 22632 26804 22882
rect 27754 22778 27760 22838
rect 27820 22778 27826 22838
rect 27040 22725 27528 22731
rect 27040 22691 27052 22725
rect 27516 22691 27528 22725
rect 27040 22685 27528 22691
rect 25774 22056 25786 22080
rect 25004 21997 25492 22003
rect 25004 21963 25016 21997
rect 25480 21963 25492 21997
rect 25004 21957 25492 21963
rect 25220 21904 25280 21957
rect 25726 21904 25786 22056
rect 26744 22056 26758 22632
rect 26792 22056 26804 22632
rect 27760 22632 27820 22778
rect 28058 22725 28546 22731
rect 28058 22691 28070 22725
rect 28534 22691 28546 22725
rect 28058 22685 28546 22691
rect 27760 22568 27776 22632
rect 26022 21997 26510 22003
rect 26022 21963 26034 21997
rect 26498 21963 26510 21997
rect 26022 21957 26510 21963
rect 24708 21902 25786 21904
rect 24708 21844 25726 21902
rect 25720 21842 25726 21844
rect 25786 21842 25792 21902
rect 26230 21794 26290 21957
rect 26224 21734 26230 21794
rect 26290 21734 26296 21794
rect 26230 21699 26290 21734
rect 25004 21693 25492 21699
rect 25004 21659 25016 21693
rect 25480 21659 25492 21693
rect 25004 21653 25492 21659
rect 26022 21693 26510 21699
rect 26022 21659 26034 21693
rect 26498 21659 26510 21693
rect 26022 21653 26510 21659
rect 24716 21600 24762 21612
rect 24716 21080 24722 21600
rect 24708 21024 24722 21080
rect 24756 21080 24762 21600
rect 25734 21600 25780 21612
rect 24756 21024 24768 21080
rect 25734 21054 25740 21600
rect 24708 20864 24768 21024
rect 25722 21024 25740 21054
rect 25774 21054 25780 21600
rect 26744 21600 26804 22056
rect 27770 22056 27776 22568
rect 27810 22568 27820 22632
rect 28782 22632 28842 22882
rect 29076 22725 29564 22731
rect 29076 22691 29088 22725
rect 29552 22691 29564 22725
rect 29076 22685 29564 22691
rect 30094 22725 30582 22731
rect 30094 22691 30106 22725
rect 30570 22691 30582 22725
rect 30094 22685 30582 22691
rect 27810 22056 27816 22568
rect 27770 22044 27816 22056
rect 28782 22056 28794 22632
rect 28828 22056 28842 22632
rect 29806 22632 29852 22644
rect 29806 22120 29812 22632
rect 27250 22003 27310 22009
rect 27040 21997 27528 22003
rect 27040 21963 27052 21997
rect 27516 21963 27528 21997
rect 27040 21957 27528 21963
rect 28058 21997 28546 22003
rect 28058 21963 28070 21997
rect 28534 21963 28546 21997
rect 28058 21957 28546 21963
rect 27250 21800 27310 21957
rect 27754 21842 27760 21902
rect 27820 21842 27826 21902
rect 27250 21794 27312 21800
rect 27250 21734 27252 21794
rect 27250 21728 27312 21734
rect 27250 21699 27310 21728
rect 27040 21693 27528 21699
rect 27040 21659 27052 21693
rect 27516 21659 27528 21693
rect 27040 21653 27528 21659
rect 25774 21024 25782 21054
rect 25004 20965 25492 20971
rect 25004 20931 25016 20965
rect 25480 20931 25492 20965
rect 25004 20925 25492 20931
rect 25210 20864 25270 20925
rect 25722 20870 25782 21024
rect 26744 21024 26758 21600
rect 26792 21024 26804 21600
rect 27760 21600 27820 21842
rect 28272 21800 28332 21957
rect 28270 21794 28332 21800
rect 28330 21734 28332 21794
rect 28270 21728 28332 21734
rect 28272 21699 28332 21728
rect 28058 21693 28546 21699
rect 28058 21659 28070 21693
rect 28534 21659 28546 21693
rect 28058 21653 28546 21659
rect 28272 21646 28332 21653
rect 27760 21554 27776 21600
rect 26022 20965 26510 20971
rect 26022 20931 26034 20965
rect 26498 20931 26510 20965
rect 26022 20925 26510 20931
rect 25716 20864 25722 20870
rect 24582 20810 25722 20864
rect 25782 20810 25788 20870
rect 24582 20804 25788 20810
rect 26228 20736 26288 20925
rect 26228 20670 26288 20676
rect 26744 20528 26804 21024
rect 27770 21024 27776 21554
rect 27810 21554 27820 21600
rect 28782 21600 28842 22056
rect 29802 22056 29812 22120
rect 29846 22120 29852 22632
rect 30820 22632 30880 22882
rect 31822 22778 31828 22838
rect 31888 22778 31894 22838
rect 31112 22725 31600 22731
rect 31112 22691 31124 22725
rect 31588 22691 31600 22725
rect 31112 22685 31600 22691
rect 29846 22056 29862 22120
rect 29076 21997 29564 22003
rect 29076 21963 29088 21997
rect 29552 21963 29564 21997
rect 29076 21957 29564 21963
rect 29292 21800 29352 21957
rect 29802 21902 29862 22056
rect 30820 22056 30830 22632
rect 30864 22056 30880 22632
rect 31828 22632 31888 22778
rect 32130 22725 32618 22731
rect 32130 22691 32142 22725
rect 32606 22691 32618 22725
rect 32130 22685 32618 22691
rect 31828 22558 31848 22632
rect 30308 22003 30368 22005
rect 30094 21997 30582 22003
rect 30094 21963 30106 21997
rect 30570 21963 30582 21997
rect 30094 21957 30582 21963
rect 29796 21842 29802 21902
rect 29862 21842 29868 21902
rect 29292 21794 29354 21800
rect 29292 21734 29294 21794
rect 29292 21728 29354 21734
rect 30308 21794 30368 21957
rect 29292 21699 29352 21728
rect 30308 21699 30368 21734
rect 29076 21693 29564 21699
rect 29076 21659 29088 21693
rect 29552 21659 29564 21693
rect 29076 21653 29564 21659
rect 30094 21693 30582 21699
rect 30094 21659 30106 21693
rect 30570 21659 30582 21693
rect 30094 21653 30582 21659
rect 27810 21024 27816 21554
rect 27770 21012 27816 21024
rect 28782 21024 28794 21600
rect 28828 21024 28842 21600
rect 29806 21600 29852 21612
rect 29806 21090 29812 21600
rect 27242 20971 27302 20974
rect 27040 20965 27528 20971
rect 27040 20931 27052 20965
rect 27516 20931 27528 20965
rect 27040 20925 27528 20931
rect 28058 20965 28546 20971
rect 28058 20931 28070 20965
rect 28534 20931 28546 20965
rect 28058 20925 28546 20931
rect 27242 20732 27302 20925
rect 28274 20740 28334 20925
rect 28274 20674 28334 20680
rect 27242 20666 27302 20672
rect 28782 20528 28842 21024
rect 29802 21024 29812 21090
rect 29846 21090 29852 21600
rect 30820 21600 30880 22056
rect 31842 22056 31848 22558
rect 31882 22056 31888 22632
rect 31842 22044 31888 22056
rect 32856 22632 32916 22882
rect 33148 22725 33636 22731
rect 33148 22691 33160 22725
rect 33624 22691 33636 22725
rect 33148 22685 33636 22691
rect 34166 22725 34654 22731
rect 34166 22691 34178 22725
rect 34642 22691 34654 22725
rect 34166 22685 34654 22691
rect 32856 22056 32866 22632
rect 32900 22056 32916 22632
rect 33878 22632 33924 22644
rect 33878 22120 33884 22632
rect 31112 21997 31600 22003
rect 31112 21963 31124 21997
rect 31588 21963 31600 21997
rect 31112 21957 31600 21963
rect 32130 21997 32618 22003
rect 32130 21963 32142 21997
rect 32606 21963 32618 21997
rect 32130 21957 32618 21963
rect 31324 21800 31384 21957
rect 31822 21842 31828 21902
rect 31888 21842 31894 21902
rect 31324 21794 31386 21800
rect 31324 21734 31326 21794
rect 31324 21728 31386 21734
rect 31324 21699 31384 21728
rect 31112 21693 31600 21699
rect 31112 21659 31124 21693
rect 31588 21659 31600 21693
rect 31112 21653 31600 21659
rect 29846 21024 29862 21090
rect 29076 20965 29564 20971
rect 29076 20931 29088 20965
rect 29552 20931 29564 20965
rect 29076 20925 29564 20931
rect 29272 20740 29332 20925
rect 29802 20870 29862 21024
rect 30820 21024 30830 21600
rect 30864 21024 30880 21600
rect 31828 21600 31888 21842
rect 32334 21800 32394 21957
rect 32334 21794 32396 21800
rect 32334 21734 32336 21794
rect 32334 21728 32396 21734
rect 32334 21699 32394 21728
rect 32130 21693 32618 21699
rect 32130 21659 32142 21693
rect 32606 21659 32618 21693
rect 32130 21653 32618 21659
rect 31828 21538 31848 21600
rect 31842 21116 31848 21538
rect 30316 20971 30376 20984
rect 30094 20965 30582 20971
rect 30094 20931 30106 20965
rect 30570 20931 30582 20965
rect 30094 20925 30582 20931
rect 29796 20810 29802 20870
rect 29862 20810 29868 20870
rect 29272 20674 29332 20680
rect 30316 20740 30376 20925
rect 30316 20674 30376 20680
rect 30820 20528 30880 21024
rect 31838 21024 31848 21116
rect 31882 21116 31888 21600
rect 32856 21600 32916 22056
rect 33870 22056 33884 22120
rect 33918 22120 33924 22632
rect 34886 22632 34946 22882
rect 35898 22778 35904 22838
rect 35964 22778 35970 22838
rect 35184 22725 35672 22731
rect 35184 22691 35196 22725
rect 35660 22691 35672 22725
rect 35184 22685 35672 22691
rect 34886 22222 34902 22632
rect 34896 22128 34902 22222
rect 33918 22056 33930 22120
rect 33356 22003 33416 22005
rect 33148 21997 33636 22003
rect 33148 21963 33160 21997
rect 33624 21963 33636 21997
rect 33148 21957 33636 21963
rect 33356 21800 33416 21957
rect 33870 21902 33930 22056
rect 34886 22056 34902 22128
rect 34936 22222 34946 22632
rect 35904 22632 35964 22778
rect 36202 22725 36690 22731
rect 36202 22691 36214 22725
rect 36678 22691 36690 22725
rect 36202 22685 36690 22691
rect 35904 22568 35920 22632
rect 34936 22128 34942 22222
rect 34936 22056 34946 22128
rect 34370 22003 34430 22005
rect 34166 21997 34654 22003
rect 34166 21963 34178 21997
rect 34642 21963 34654 21997
rect 34166 21957 34654 21963
rect 33864 21842 33870 21902
rect 33930 21842 33936 21902
rect 34370 21800 34430 21957
rect 33356 21794 33418 21800
rect 33356 21734 33358 21794
rect 33356 21728 33418 21734
rect 34370 21794 34432 21800
rect 34370 21734 34372 21794
rect 34370 21728 34432 21734
rect 33356 21699 33416 21728
rect 34370 21699 34430 21728
rect 33148 21693 33636 21699
rect 33148 21659 33160 21693
rect 33624 21659 33636 21693
rect 33148 21653 33636 21659
rect 34166 21693 34654 21699
rect 34166 21659 34178 21693
rect 34642 21659 34654 21693
rect 34166 21653 34654 21659
rect 31882 21024 31898 21116
rect 31320 20971 31380 20974
rect 31112 20965 31600 20971
rect 31112 20931 31124 20965
rect 31588 20931 31600 20965
rect 31112 20925 31600 20931
rect 31320 20736 31380 20925
rect 31320 20670 31380 20676
rect 31838 20620 31898 21024
rect 32856 21024 32866 21600
rect 32900 21024 32916 21600
rect 33878 21600 33924 21612
rect 33878 21106 33884 21600
rect 32336 20971 32396 20978
rect 32130 20965 32618 20971
rect 32130 20931 32142 20965
rect 32606 20931 32618 20965
rect 32130 20925 32618 20931
rect 32336 20736 32396 20925
rect 32336 20670 32396 20676
rect 31628 20560 31898 20620
rect 26744 20468 31120 20528
rect 31180 20468 31186 20528
rect 24468 20338 28636 20398
rect 24346 20150 24352 20210
rect 24412 20150 24418 20210
rect 25512 20150 25518 20210
rect 25578 20150 25584 20210
rect 24078 19104 24084 19164
rect 24144 19104 24150 19164
rect 23836 17946 23842 18006
rect 23902 17946 23908 18006
rect 23832 17732 23838 17792
rect 23898 17732 23904 17792
rect 23720 16690 23726 16750
rect 23786 16690 23792 16750
rect 18382 15436 23652 15496
rect 18322 15430 18382 15436
rect 3048 14898 14318 14958
rect 3048 14410 3114 14898
rect 3342 14702 14318 14898
rect 17412 14838 17524 15352
rect 19376 15234 19436 15240
rect 23838 15234 23898 17732
rect 24084 15492 24144 19104
rect 24214 19006 24220 19066
rect 24280 19006 24286 19066
rect 24078 15432 24084 15492
rect 24144 15432 24150 15492
rect 24220 15362 24280 19006
rect 24352 16542 24412 20150
rect 24796 20089 25284 20095
rect 24796 20055 24808 20089
rect 25272 20055 25284 20089
rect 24796 20049 25284 20055
rect 24508 19996 24554 20008
rect 24508 19456 24514 19996
rect 24500 19420 24514 19456
rect 24548 19456 24554 19996
rect 25518 19996 25578 20150
rect 25814 20089 26302 20095
rect 25814 20055 25826 20089
rect 26290 20055 26302 20089
rect 25814 20049 26302 20055
rect 25518 19970 25532 19996
rect 24548 19420 24560 19456
rect 25526 19444 25532 19970
rect 24500 19262 24560 19420
rect 25516 19420 25532 19444
rect 25566 19970 25578 19996
rect 26534 19996 26594 20338
rect 27548 20150 27554 20210
rect 27614 20150 27620 20210
rect 26832 20089 27320 20095
rect 26832 20055 26844 20089
rect 27308 20055 27320 20089
rect 26832 20049 27320 20055
rect 25566 19444 25572 19970
rect 26534 19950 26550 19996
rect 26544 19444 26550 19950
rect 25566 19420 25576 19444
rect 24796 19361 25284 19367
rect 24796 19327 24808 19361
rect 25272 19327 25284 19361
rect 24796 19321 25284 19327
rect 25014 19262 25074 19321
rect 25516 19262 25576 19420
rect 26536 19420 26550 19444
rect 26584 19950 26594 19996
rect 27554 19996 27614 20150
rect 28056 20146 28062 20210
rect 28126 20146 28132 20210
rect 28062 20095 28126 20146
rect 27850 20089 28338 20095
rect 27850 20055 27862 20089
rect 28326 20055 28338 20089
rect 27850 20049 28338 20055
rect 27554 19972 27568 19996
rect 26584 19444 26590 19950
rect 26584 19420 26596 19444
rect 25814 19361 26302 19367
rect 25814 19327 25826 19361
rect 26290 19327 26302 19361
rect 25814 19321 26302 19327
rect 24500 19202 25576 19262
rect 26006 18960 26066 19321
rect 26536 19262 26596 19420
rect 27562 19420 27568 19972
rect 27602 19972 27614 19996
rect 28576 19996 28636 20338
rect 29080 20095 29140 20468
rect 28868 20089 29356 20095
rect 28868 20055 28880 20089
rect 29344 20055 29356 20089
rect 28868 20049 29356 20055
rect 27602 19420 27608 19972
rect 28576 19942 28586 19996
rect 28580 19448 28586 19942
rect 27562 19408 27608 19420
rect 28572 19420 28586 19448
rect 28620 19942 28636 19996
rect 29588 19996 29648 20468
rect 30080 20095 30140 20468
rect 31118 20095 31178 20468
rect 29886 20089 30374 20095
rect 29886 20055 29898 20089
rect 30362 20055 30374 20089
rect 29886 20049 30374 20055
rect 30904 20089 31392 20095
rect 30904 20055 30916 20089
rect 31380 20055 31392 20089
rect 30904 20049 31392 20055
rect 28620 19448 28626 19942
rect 28620 19420 28632 19448
rect 26832 19361 27320 19367
rect 26832 19327 26844 19361
rect 27308 19327 27320 19361
rect 26832 19321 27320 19327
rect 27850 19361 28338 19367
rect 27850 19327 27862 19361
rect 28326 19327 28338 19361
rect 27850 19321 28338 19327
rect 26530 19202 26536 19262
rect 26596 19202 26602 19262
rect 27044 19208 27104 19321
rect 28050 19208 28110 19321
rect 28572 19262 28632 19420
rect 29588 19420 29604 19996
rect 29638 19420 29648 19996
rect 30616 19996 30662 20008
rect 30616 19444 30622 19996
rect 28868 19361 29356 19367
rect 28868 19327 28880 19361
rect 29344 19327 29356 19361
rect 28868 19321 29356 19327
rect 29082 19266 29142 19321
rect 29588 19266 29648 19420
rect 30608 19420 30622 19444
rect 30656 19444 30662 19996
rect 31628 19996 31688 20560
rect 32856 20528 32916 21024
rect 33870 21024 33884 21106
rect 33918 21106 33924 21600
rect 34886 21600 34946 22056
rect 35914 22056 35920 22568
rect 35954 22568 35964 22632
rect 36924 22632 36984 22882
rect 39094 22778 39100 22838
rect 39160 22778 39166 22838
rect 37220 22725 37708 22731
rect 37220 22691 37232 22725
rect 37696 22691 37708 22725
rect 37220 22685 37708 22691
rect 38238 22725 38726 22731
rect 38238 22691 38250 22725
rect 38714 22691 38726 22725
rect 38238 22685 38726 22691
rect 35954 22056 35960 22568
rect 35914 22044 35960 22056
rect 36924 22056 36938 22632
rect 36972 22056 36984 22632
rect 37950 22632 37996 22644
rect 37950 22132 37956 22632
rect 35402 22003 35462 22005
rect 36412 22003 36472 22005
rect 35184 21997 35672 22003
rect 35184 21963 35196 21997
rect 35660 21963 35672 21997
rect 35184 21957 35672 21963
rect 36202 21997 36690 22003
rect 36202 21963 36214 21997
rect 36678 21963 36690 21997
rect 36202 21957 36690 21963
rect 35402 21800 35462 21957
rect 35900 21842 35906 21902
rect 35966 21842 35972 21902
rect 35402 21794 35464 21800
rect 35402 21734 35404 21794
rect 35402 21728 35464 21734
rect 35402 21699 35462 21728
rect 35184 21693 35672 21699
rect 35184 21659 35196 21693
rect 35660 21659 35672 21693
rect 35184 21653 35672 21659
rect 33918 21024 33930 21106
rect 33148 20965 33636 20971
rect 33148 20931 33160 20965
rect 33624 20931 33636 20965
rect 33148 20925 33636 20931
rect 33340 20736 33400 20925
rect 33870 20870 33930 21024
rect 34886 21024 34902 21600
rect 34936 21024 34946 21600
rect 35906 21600 35966 21842
rect 36412 21800 36472 21957
rect 36412 21794 36474 21800
rect 36412 21734 36414 21794
rect 36412 21728 36474 21734
rect 36412 21699 36472 21728
rect 36202 21693 36690 21699
rect 36202 21659 36214 21693
rect 36678 21659 36690 21693
rect 36202 21653 36690 21659
rect 35906 21532 35920 21600
rect 34166 20965 34654 20971
rect 34166 20931 34178 20965
rect 34642 20931 34654 20965
rect 34166 20925 34654 20931
rect 33864 20810 33870 20870
rect 33930 20810 33936 20870
rect 33340 20670 33400 20676
rect 34372 20740 34432 20925
rect 34372 20674 34432 20680
rect 32130 20268 32136 20332
rect 32200 20268 32206 20332
rect 32136 20210 32200 20268
rect 32856 20238 32916 20468
rect 34886 20628 34946 21024
rect 35914 21024 35920 21532
rect 35954 21532 35966 21600
rect 36924 21600 36984 22056
rect 37942 22056 37956 22132
rect 37990 22132 37996 22632
rect 38968 22632 39014 22644
rect 37990 22056 38002 22132
rect 38968 22082 38974 22632
rect 37220 21997 37708 22003
rect 37220 21963 37232 21997
rect 37696 21963 37708 21997
rect 37220 21957 37708 21963
rect 37434 21800 37494 21957
rect 37942 21904 38002 22056
rect 38958 22056 38974 22082
rect 39008 22082 39014 22632
rect 39008 22056 39018 22082
rect 38238 21997 38726 22003
rect 38238 21963 38250 21997
rect 38714 21963 38726 21997
rect 38238 21957 38726 21963
rect 38464 21904 38524 21957
rect 38958 21904 39018 22056
rect 37942 21902 39018 21904
rect 37936 21842 37942 21902
rect 38002 21844 39018 21902
rect 38002 21842 38008 21844
rect 37434 21794 37496 21800
rect 37434 21734 37436 21794
rect 37434 21728 37496 21734
rect 37434 21699 37494 21728
rect 37220 21693 37708 21699
rect 37220 21659 37232 21693
rect 37696 21659 37708 21693
rect 37220 21653 37708 21659
rect 38238 21693 38726 21699
rect 38238 21659 38250 21693
rect 38714 21659 38726 21693
rect 38238 21653 38726 21659
rect 35954 21024 35960 21532
rect 35914 21012 35960 21024
rect 36924 21024 36938 21600
rect 36972 21024 36984 21600
rect 37950 21600 37996 21612
rect 37950 21100 37956 21600
rect 35388 20971 35448 20974
rect 35184 20965 35672 20971
rect 35184 20931 35196 20965
rect 35660 20931 35672 20965
rect 35184 20925 35672 20931
rect 36202 20965 36690 20971
rect 36202 20931 36214 20965
rect 36678 20931 36690 20965
rect 36202 20925 36690 20931
rect 35388 20736 35448 20925
rect 35388 20670 35448 20676
rect 36416 20736 36476 20925
rect 36416 20670 36476 20676
rect 36924 20628 36984 21024
rect 37938 21024 37956 21100
rect 37990 21100 37996 21600
rect 38968 21600 39014 21612
rect 37990 21024 37998 21100
rect 38968 21096 38974 21600
rect 37436 20971 37496 20974
rect 37220 20965 37708 20971
rect 37220 20931 37232 20965
rect 37696 20931 37708 20965
rect 37220 20925 37708 20931
rect 37436 20736 37496 20925
rect 37938 20874 37998 21024
rect 38958 21024 38974 21096
rect 39008 21096 39014 21600
rect 39008 21024 39018 21096
rect 38238 20965 38726 20971
rect 38238 20931 38250 20965
rect 38714 20931 38726 20965
rect 38238 20925 38726 20931
rect 38426 20874 38486 20925
rect 38958 20874 39018 21024
rect 39100 20874 39160 22778
rect 37936 20870 39160 20874
rect 37932 20810 37938 20870
rect 37998 20814 39160 20870
rect 37998 20810 38004 20814
rect 39888 20678 39894 20738
rect 39954 20678 39960 20738
rect 37436 20670 37496 20676
rect 34886 20568 36984 20628
rect 34886 20238 34946 20568
rect 38748 20452 38754 20512
rect 38814 20452 38820 20512
rect 36194 20268 36200 20332
rect 36264 20268 36270 20332
rect 37218 20268 37224 20332
rect 37288 20268 37294 20332
rect 38230 20268 38236 20332
rect 38300 20268 38306 20332
rect 32132 20146 32138 20210
rect 32202 20146 32208 20210
rect 32856 20178 35250 20238
rect 36200 20214 36264 20268
rect 32136 20095 32200 20146
rect 33168 20095 33228 20178
rect 31922 20089 32410 20095
rect 31922 20055 31934 20089
rect 32398 20055 32410 20089
rect 31922 20049 32410 20055
rect 32940 20089 33428 20095
rect 32940 20055 32952 20089
rect 33416 20055 33428 20089
rect 32940 20049 33428 20055
rect 30656 19420 30668 19444
rect 29886 19361 30374 19367
rect 29886 19327 29898 19361
rect 30362 19327 30374 19361
rect 29886 19321 30374 19327
rect 30102 19266 30162 19321
rect 30608 19266 30668 19420
rect 31628 19420 31640 19996
rect 31674 19420 31688 19996
rect 32652 19996 32698 20008
rect 32652 19498 32658 19996
rect 30904 19361 31392 19367
rect 30904 19327 30916 19361
rect 31380 19327 31392 19361
rect 30904 19321 31392 19327
rect 31112 19266 31172 19321
rect 26536 19066 26596 19202
rect 27044 19148 28110 19208
rect 28566 19202 28572 19262
rect 28632 19202 28638 19262
rect 28908 19204 28914 19264
rect 28974 19204 28980 19264
rect 29082 19206 31172 19266
rect 31628 19264 31688 19420
rect 32646 19420 32658 19498
rect 32692 19498 32698 19996
rect 33662 19996 33722 20178
rect 34190 20095 34250 20178
rect 33958 20089 34446 20095
rect 33958 20055 33970 20089
rect 34434 20055 34446 20089
rect 33958 20049 34446 20055
rect 34190 20048 34250 20049
rect 32692 19420 32706 19498
rect 31922 19361 32410 19367
rect 31922 19327 31934 19361
rect 32398 19327 32410 19361
rect 31922 19321 32410 19327
rect 26530 19006 26536 19066
rect 26596 19006 26602 19066
rect 27044 18960 27104 19148
rect 27550 19008 27556 19068
rect 27616 19008 27622 19068
rect 25516 18896 25522 18956
rect 25582 18896 25588 18956
rect 26006 18900 27104 18960
rect 27556 18956 27616 19008
rect 24796 18833 25284 18839
rect 24796 18799 24808 18833
rect 25272 18799 25284 18833
rect 24796 18793 25284 18799
rect 24508 18740 24554 18752
rect 24508 18200 24514 18740
rect 24504 18164 24514 18200
rect 24548 18200 24554 18740
rect 25522 18740 25582 18896
rect 26006 18839 26066 18900
rect 27044 18839 27104 18900
rect 27550 18896 27556 18956
rect 27616 18896 27622 18956
rect 25814 18833 26302 18839
rect 25814 18799 25826 18833
rect 26290 18799 26302 18833
rect 25814 18793 26302 18799
rect 26832 18833 27320 18839
rect 26832 18799 26844 18833
rect 27308 18799 27320 18833
rect 26832 18793 27320 18799
rect 25522 18714 25532 18740
rect 24548 18164 24564 18200
rect 25526 18188 25532 18714
rect 24504 18006 24564 18164
rect 25520 18164 25532 18188
rect 25566 18714 25582 18740
rect 26544 18740 26590 18752
rect 25566 18188 25572 18714
rect 26544 18190 26550 18740
rect 25566 18164 25580 18188
rect 24796 18105 25284 18111
rect 24796 18071 24808 18105
rect 25272 18071 25284 18105
rect 24796 18065 25284 18071
rect 25018 18006 25078 18065
rect 25520 18006 25580 18164
rect 26538 18164 26550 18190
rect 26584 18190 26590 18740
rect 27556 18740 27616 18896
rect 28050 18839 28110 19148
rect 28914 18950 28974 19204
rect 28572 18890 28974 18950
rect 27850 18833 28338 18839
rect 27850 18799 27862 18833
rect 28326 18799 28338 18833
rect 27850 18793 28338 18799
rect 27556 18718 27568 18740
rect 26584 18164 26598 18190
rect 26000 18111 26060 18112
rect 25814 18105 26302 18111
rect 25814 18071 25826 18105
rect 26290 18071 26302 18105
rect 25814 18065 26302 18071
rect 24504 17946 25580 18006
rect 24504 17792 24564 17946
rect 24498 17732 24504 17792
rect 24564 17732 24570 17792
rect 24502 17622 25578 17682
rect 24502 17484 24562 17622
rect 25016 17583 25076 17622
rect 24796 17577 25284 17583
rect 24796 17543 24808 17577
rect 25272 17543 25284 17577
rect 24796 17537 25284 17543
rect 24502 17450 24514 17484
rect 24508 16908 24514 17450
rect 24548 17450 24562 17484
rect 25518 17484 25578 17622
rect 26000 17583 26060 18065
rect 26538 17902 26598 18164
rect 27562 18164 27568 18718
rect 27602 18718 27616 18740
rect 28572 18740 28632 18890
rect 28868 18833 29356 18839
rect 28868 18799 28880 18833
rect 29344 18799 29356 18833
rect 28868 18793 29356 18799
rect 27602 18164 27608 18718
rect 28572 18682 28586 18740
rect 28580 18194 28586 18682
rect 27562 18152 27608 18164
rect 28574 18164 28586 18194
rect 28620 18682 28632 18740
rect 29588 18740 29648 19206
rect 31622 19204 31628 19264
rect 31688 19204 31694 19264
rect 32646 19068 32706 19420
rect 33662 19420 33676 19996
rect 33710 19420 33722 19996
rect 32940 19361 33428 19367
rect 32940 19327 32952 19361
rect 33416 19327 33428 19361
rect 32940 19321 33428 19327
rect 33156 19266 33216 19321
rect 33662 19266 33722 19420
rect 34678 19996 34738 20178
rect 35190 20095 35250 20178
rect 35694 20150 35700 20210
rect 35760 20150 35766 20210
rect 34976 20089 35464 20095
rect 34976 20055 34988 20089
rect 35452 20055 35464 20089
rect 34976 20049 35464 20055
rect 35190 20042 35250 20049
rect 34678 19420 34694 19996
rect 34728 19420 34738 19996
rect 35700 19996 35760 20150
rect 36200 20095 36264 20150
rect 37224 20095 37288 20268
rect 37728 20150 37734 20210
rect 37794 20150 37800 20210
rect 35994 20089 36482 20095
rect 35994 20055 36006 20089
rect 36470 20055 36482 20089
rect 35994 20049 36482 20055
rect 37012 20089 37500 20095
rect 37012 20055 37024 20089
rect 37488 20055 37500 20089
rect 37012 20049 37500 20055
rect 35700 19968 35712 19996
rect 33958 19361 34446 19367
rect 33958 19327 33970 19361
rect 34434 19327 34446 19361
rect 33958 19321 34446 19327
rect 34182 19266 34242 19321
rect 34678 19266 34738 19420
rect 35706 19420 35712 19968
rect 35746 19968 35760 19996
rect 36724 19996 36770 20008
rect 35746 19420 35752 19968
rect 36724 19444 36730 19996
rect 35706 19408 35752 19420
rect 36716 19420 36730 19444
rect 36764 19444 36770 19996
rect 37734 19996 37794 20150
rect 38236 20095 38300 20268
rect 38754 20214 38814 20452
rect 38754 20154 39830 20214
rect 38030 20089 38518 20095
rect 38030 20055 38042 20089
rect 38506 20055 38518 20089
rect 38030 20049 38518 20055
rect 37734 19972 37748 19996
rect 36764 19420 36776 19444
rect 34976 19361 35464 19367
rect 34976 19327 34988 19361
rect 35452 19327 35464 19361
rect 34976 19321 35464 19327
rect 35994 19361 36482 19367
rect 35994 19327 36006 19361
rect 36470 19327 36482 19361
rect 35994 19321 36482 19327
rect 35194 19266 35254 19321
rect 33156 19206 35254 19266
rect 32640 19008 32646 19068
rect 32706 19008 32712 19068
rect 30606 18894 30612 18954
rect 30672 18894 30678 18954
rect 32640 18894 32646 18954
rect 32706 18894 32712 18954
rect 29886 18833 30374 18839
rect 29886 18799 29898 18833
rect 30362 18799 30374 18833
rect 29886 18793 30374 18799
rect 29588 18696 29604 18740
rect 28620 18194 28626 18682
rect 29598 18194 29604 18696
rect 28620 18164 28634 18194
rect 27038 18111 27098 18112
rect 28044 18111 28104 18112
rect 26832 18105 27320 18111
rect 26832 18071 26844 18105
rect 27308 18071 27320 18105
rect 26832 18065 27320 18071
rect 27850 18105 28338 18111
rect 27850 18071 27862 18105
rect 28326 18071 28338 18105
rect 27850 18065 28338 18071
rect 26538 17836 26598 17842
rect 26532 17638 26538 17698
rect 26598 17638 26604 17698
rect 25814 17577 26302 17583
rect 25814 17543 25826 17577
rect 26290 17543 26302 17577
rect 25814 17537 26302 17543
rect 25518 17462 25532 17484
rect 24548 16908 24554 17450
rect 25526 16936 25532 17462
rect 24508 16896 24554 16908
rect 25520 16908 25532 16936
rect 25566 17462 25578 17484
rect 26538 17484 26598 17638
rect 27038 17583 27098 18065
rect 28044 17583 28104 18065
rect 28574 17902 28634 18164
rect 29590 18164 29604 18194
rect 29638 18696 29648 18740
rect 30612 18740 30672 18894
rect 30904 18833 31392 18839
rect 30904 18799 30916 18833
rect 31380 18799 31392 18833
rect 30904 18793 31392 18799
rect 31922 18833 32410 18839
rect 31922 18799 31934 18833
rect 32398 18799 32410 18833
rect 31922 18793 32410 18799
rect 30612 18712 30622 18740
rect 29638 18194 29644 18696
rect 29638 18164 29650 18194
rect 28868 18105 29356 18111
rect 28868 18071 28880 18105
rect 29344 18071 29356 18105
rect 28868 18065 29356 18071
rect 29094 18010 29154 18065
rect 29590 18010 29650 18164
rect 30616 18164 30622 18712
rect 30656 18712 30672 18740
rect 31634 18740 31680 18752
rect 30656 18164 30662 18712
rect 31634 18188 31640 18740
rect 30616 18152 30662 18164
rect 31628 18164 31640 18188
rect 31674 18188 31680 18740
rect 32646 18740 32706 18894
rect 32940 18833 33428 18839
rect 32940 18799 32952 18833
rect 33416 18799 33428 18833
rect 32940 18793 33428 18799
rect 33958 18833 34446 18839
rect 33958 18799 33970 18833
rect 34434 18799 34446 18833
rect 33958 18793 34446 18799
rect 32646 18710 32658 18740
rect 32652 18192 32658 18710
rect 31674 18164 31688 18188
rect 29886 18105 30374 18111
rect 29886 18071 29898 18105
rect 30362 18071 30374 18105
rect 29886 18065 30374 18071
rect 30904 18105 31392 18111
rect 30904 18071 30916 18105
rect 31380 18071 31392 18105
rect 30904 18065 31392 18071
rect 30106 18010 30166 18065
rect 29094 17950 30166 18010
rect 28568 17842 28574 17902
rect 28634 17842 28640 17902
rect 28566 17740 28572 17800
rect 28632 17740 28638 17800
rect 28572 17698 28632 17740
rect 28566 17638 28572 17698
rect 28632 17638 28638 17698
rect 26832 17577 27320 17583
rect 26832 17543 26844 17577
rect 27308 17543 27320 17577
rect 26832 17537 27320 17543
rect 27850 17577 28338 17583
rect 27850 17543 27862 17577
rect 28326 17543 28338 17577
rect 27850 17537 28338 17543
rect 25566 16936 25572 17462
rect 26538 17460 26550 17484
rect 25566 16908 25580 16936
rect 24796 16849 25284 16855
rect 24796 16815 24808 16849
rect 25272 16815 25284 16849
rect 24796 16809 25284 16815
rect 25520 16750 25580 16908
rect 26544 16908 26550 17460
rect 26584 17460 26598 17484
rect 27562 17484 27608 17496
rect 26584 16908 26590 17460
rect 27562 16932 27568 17484
rect 26544 16896 26590 16908
rect 27556 16908 27568 16932
rect 27602 16932 27608 17484
rect 28572 17484 28632 17638
rect 28868 17577 29356 17583
rect 28868 17543 28880 17577
rect 29344 17543 29356 17577
rect 28868 17537 29356 17543
rect 28572 17456 28586 17484
rect 27602 16908 27616 16932
rect 28580 16927 28586 17456
rect 26012 16855 26072 16862
rect 27050 16855 27110 16862
rect 25814 16849 26302 16855
rect 25814 16815 25826 16849
rect 26290 16815 26302 16849
rect 25814 16809 26302 16815
rect 26832 16849 27320 16855
rect 26832 16815 26844 16849
rect 27308 16815 27320 16849
rect 26832 16809 27320 16815
rect 25514 16690 25520 16750
rect 25580 16690 25586 16750
rect 24346 16482 24352 16542
rect 24412 16482 24418 16542
rect 24502 16384 25578 16444
rect 24502 16228 24562 16384
rect 25016 16327 25076 16384
rect 24796 16321 25284 16327
rect 24796 16287 24808 16321
rect 25272 16287 25284 16321
rect 24796 16281 25284 16287
rect 24502 16190 24514 16228
rect 24508 15652 24514 16190
rect 24548 16190 24562 16228
rect 25518 16228 25578 16384
rect 26012 16327 26072 16809
rect 26528 16380 26534 16440
rect 26594 16380 26600 16440
rect 25814 16321 26302 16327
rect 25814 16287 25826 16321
rect 26290 16287 26302 16321
rect 25814 16281 26302 16287
rect 25518 16202 25532 16228
rect 24548 15652 24554 16190
rect 25526 15678 25532 16202
rect 24508 15640 24554 15652
rect 25516 15652 25532 15678
rect 25566 16202 25578 16228
rect 26534 16228 26594 16380
rect 27050 16327 27110 16809
rect 27556 16750 27616 16908
rect 28574 16908 28586 16927
rect 28620 17456 28632 17484
rect 29590 17484 29650 17950
rect 30602 17946 30608 18006
rect 30668 17946 30674 18006
rect 29886 17577 30374 17583
rect 29886 17543 29898 17577
rect 30362 17543 30374 17577
rect 29886 17537 30374 17543
rect 28620 16927 28626 17456
rect 29590 17446 29604 17484
rect 29598 16942 29604 17446
rect 28620 16908 28634 16927
rect 28056 16855 28116 16862
rect 27850 16849 28338 16855
rect 27850 16815 27862 16849
rect 28326 16815 28338 16849
rect 27850 16809 28338 16815
rect 27550 16690 27556 16750
rect 27616 16690 27622 16750
rect 27556 16642 27616 16690
rect 27550 16582 27556 16642
rect 27616 16582 27622 16642
rect 28056 16592 28116 16809
rect 28574 16758 28634 16908
rect 29588 16908 29604 16942
rect 29638 17446 29650 17484
rect 30608 17484 30668 17946
rect 31110 17844 31170 18065
rect 31628 18006 31688 18164
rect 32646 18164 32658 18192
rect 32692 18710 32706 18740
rect 33670 18740 33716 18752
rect 32692 18192 32698 18710
rect 33670 18192 33676 18740
rect 32692 18164 32706 18192
rect 32140 18111 32200 18118
rect 31922 18105 32410 18111
rect 31922 18071 31934 18105
rect 32398 18071 32410 18105
rect 31922 18065 32410 18071
rect 31622 17946 31628 18006
rect 31688 17946 31694 18006
rect 32140 17844 32200 18065
rect 31110 17784 32200 17844
rect 31110 17583 31170 17784
rect 31622 17640 31628 17700
rect 31688 17640 31694 17700
rect 30904 17577 31392 17583
rect 30904 17543 30916 17577
rect 31380 17543 31392 17577
rect 30904 17537 31392 17543
rect 31110 17532 31170 17537
rect 30608 17460 30622 17484
rect 29638 16942 29644 17446
rect 29638 16908 29648 16942
rect 30616 16938 30622 17460
rect 28868 16849 29356 16855
rect 28868 16815 28880 16849
rect 29344 16815 29356 16849
rect 28868 16809 29356 16815
rect 29092 16758 29152 16809
rect 29588 16758 29648 16908
rect 30610 16908 30622 16938
rect 30656 17460 30668 17484
rect 31628 17484 31688 17640
rect 32140 17583 32200 17784
rect 32646 17700 32706 18164
rect 33664 18164 33676 18192
rect 33710 18192 33716 18740
rect 34678 18740 34738 19206
rect 35696 18894 35702 18954
rect 35762 18894 35768 18954
rect 34976 18833 35464 18839
rect 34976 18799 34988 18833
rect 35452 18799 35464 18833
rect 34976 18793 35464 18799
rect 34678 18720 34694 18740
rect 34688 18192 34694 18720
rect 33710 18164 33724 18192
rect 33152 18111 33212 18118
rect 32940 18105 33428 18111
rect 32940 18071 32952 18105
rect 33416 18071 33428 18105
rect 32940 18065 33428 18071
rect 32640 17640 32646 17700
rect 32706 17640 32712 17700
rect 33152 17583 33212 18065
rect 33664 18006 33724 18164
rect 34678 18164 34694 18192
rect 34728 18720 34738 18740
rect 35702 18740 35762 18894
rect 36202 18839 36262 19321
rect 36716 19262 36776 19420
rect 37742 19420 37748 19972
rect 37782 19972 37794 19996
rect 38754 19996 38814 20154
rect 39268 20095 39328 20154
rect 39048 20089 39536 20095
rect 39048 20055 39060 20089
rect 39524 20055 39536 20089
rect 39048 20049 39536 20055
rect 37782 19420 37788 19972
rect 38754 19960 38766 19996
rect 38760 19448 38766 19960
rect 37742 19408 37788 19420
rect 38752 19420 38766 19448
rect 38800 19960 38814 19996
rect 39770 19996 39830 20154
rect 39770 19972 39784 19996
rect 38800 19448 38806 19960
rect 38800 19420 38812 19448
rect 38232 19367 38292 19373
rect 37012 19361 37500 19367
rect 37012 19327 37024 19361
rect 37488 19327 37500 19361
rect 37012 19321 37500 19327
rect 38030 19361 38518 19367
rect 38030 19327 38042 19361
rect 38506 19327 38518 19361
rect 38030 19321 38518 19327
rect 36710 19202 36716 19262
rect 36776 19202 36782 19262
rect 37226 18839 37286 19321
rect 37730 18894 37736 18954
rect 37796 18894 37802 18954
rect 35994 18833 36482 18839
rect 35994 18799 36006 18833
rect 36470 18799 36482 18833
rect 35994 18793 36482 18799
rect 37012 18833 37500 18839
rect 37012 18799 37024 18833
rect 37488 18799 37500 18833
rect 37012 18793 37500 18799
rect 34728 18192 34734 18720
rect 35702 18712 35712 18740
rect 34728 18164 34738 18192
rect 33958 18105 34446 18111
rect 33958 18071 33970 18105
rect 34434 18071 34446 18105
rect 33958 18065 34446 18071
rect 34182 18008 34242 18065
rect 34678 18008 34738 18164
rect 35706 18164 35712 18712
rect 35746 18712 35762 18740
rect 36724 18740 36770 18752
rect 35746 18164 35752 18712
rect 36724 18200 36730 18740
rect 35706 18152 35752 18164
rect 36714 18164 36730 18200
rect 36764 18200 36770 18740
rect 37736 18740 37796 18894
rect 38232 18839 38292 19321
rect 38752 19262 38812 19420
rect 39778 19420 39784 19972
rect 39818 19972 39830 19996
rect 39818 19420 39824 19972
rect 39778 19408 39824 19420
rect 39048 19361 39536 19367
rect 39048 19327 39060 19361
rect 39524 19327 39536 19361
rect 39048 19321 39536 19327
rect 38746 19202 38752 19262
rect 38812 19202 38818 19262
rect 38754 18900 39830 18960
rect 38030 18833 38518 18839
rect 38030 18799 38042 18833
rect 38506 18799 38518 18833
rect 38030 18793 38518 18799
rect 37736 18716 37748 18740
rect 36764 18164 36774 18200
rect 37742 18192 37748 18716
rect 36196 18111 36256 18112
rect 34976 18105 35464 18111
rect 34976 18071 34988 18105
rect 35452 18071 35464 18105
rect 34976 18065 35464 18071
rect 35994 18105 36482 18111
rect 35994 18071 36006 18105
rect 36470 18071 36482 18105
rect 35994 18065 36482 18071
rect 35194 18008 35254 18065
rect 33658 17946 33664 18006
rect 33724 17946 33730 18006
rect 34182 17948 35254 18008
rect 33656 17640 33662 17700
rect 33722 17640 33728 17700
rect 31922 17577 32410 17583
rect 31922 17543 31934 17577
rect 32398 17543 32410 17577
rect 31922 17537 32410 17543
rect 32940 17577 33428 17583
rect 32940 17543 32952 17577
rect 33416 17543 33428 17577
rect 32940 17537 33428 17543
rect 31628 17462 31640 17484
rect 30656 16938 30662 17460
rect 30656 16908 30670 16938
rect 29886 16849 30374 16855
rect 29886 16815 29898 16849
rect 30362 16815 30374 16849
rect 29886 16809 30374 16815
rect 30104 16758 30164 16809
rect 28568 16698 28574 16758
rect 28634 16698 28640 16758
rect 29092 16698 30164 16758
rect 30370 16698 30376 16758
rect 30436 16698 30442 16758
rect 30610 16752 30670 16908
rect 31634 16908 31640 17462
rect 31674 17462 31688 17484
rect 32652 17484 32698 17496
rect 31674 16908 31680 17462
rect 32652 16934 32658 17484
rect 31634 16896 31680 16908
rect 32646 16908 32658 16934
rect 32692 16934 32698 17484
rect 33662 17484 33722 17640
rect 33958 17577 34446 17583
rect 33958 17543 33970 17577
rect 34434 17543 34446 17577
rect 33958 17537 34446 17543
rect 33662 17458 33676 17484
rect 32692 16908 32706 16934
rect 30904 16849 31392 16855
rect 30904 16815 30916 16849
rect 31380 16815 31392 16849
rect 30904 16809 31392 16815
rect 31922 16849 32410 16855
rect 31922 16815 31934 16849
rect 32398 16815 32410 16849
rect 31922 16809 32410 16815
rect 28056 16532 28832 16592
rect 28056 16327 28116 16532
rect 28562 16380 28568 16440
rect 28628 16380 28634 16440
rect 28772 16428 28832 16532
rect 26832 16321 27320 16327
rect 26832 16287 26844 16321
rect 27308 16287 27320 16321
rect 26832 16281 27320 16287
rect 27850 16321 28338 16327
rect 27850 16287 27862 16321
rect 28326 16287 28338 16321
rect 27850 16281 28338 16287
rect 26534 16202 26550 16228
rect 25566 15678 25572 16202
rect 25566 15652 25576 15678
rect 24796 15593 25284 15599
rect 24796 15559 24808 15593
rect 25272 15559 25284 15593
rect 24796 15553 25284 15559
rect 25516 15492 25576 15652
rect 26544 15652 26550 16202
rect 26584 16202 26594 16228
rect 27562 16228 27608 16240
rect 26584 15652 26590 16202
rect 27562 15674 27568 16228
rect 26544 15640 26590 15652
rect 27552 15652 27568 15674
rect 27602 15674 27608 16228
rect 28568 16228 28628 16380
rect 28766 16368 28772 16428
rect 28832 16368 28838 16428
rect 28868 16321 29356 16327
rect 28868 16287 28880 16321
rect 29344 16287 29356 16321
rect 28868 16281 29356 16287
rect 28568 16198 28586 16228
rect 28580 15688 28586 16198
rect 27602 15652 27612 15674
rect 25814 15593 26302 15599
rect 25814 15559 25826 15593
rect 26290 15559 26302 15593
rect 25814 15553 26302 15559
rect 26832 15593 27320 15599
rect 26832 15559 26844 15593
rect 27308 15559 27320 15593
rect 26832 15553 27320 15559
rect 25510 15432 25516 15492
rect 25576 15432 25582 15492
rect 26024 15378 26084 15553
rect 27048 15378 27108 15553
rect 27552 15492 27612 15652
rect 28574 15652 28586 15688
rect 28620 16198 28628 16228
rect 29588 16228 29648 16698
rect 30376 16488 30436 16698
rect 30604 16692 30610 16752
rect 30670 16692 30676 16752
rect 31106 16630 31166 16809
rect 32134 16630 32194 16809
rect 32646 16752 32706 16908
rect 33670 16908 33676 17458
rect 33710 17458 33722 17484
rect 34678 17484 34738 17948
rect 35692 17842 35698 17902
rect 35758 17842 35764 17902
rect 34976 17577 35464 17583
rect 34976 17543 34988 17577
rect 35452 17543 35464 17577
rect 34976 17537 35464 17543
rect 33710 16908 33716 17458
rect 34678 17454 34694 17484
rect 34688 16940 34694 17454
rect 33670 16896 33716 16908
rect 34676 16908 34694 16940
rect 34728 17454 34738 17484
rect 35698 17484 35758 17842
rect 36196 17583 36256 18065
rect 36560 17960 36566 18020
rect 36626 17960 36632 18020
rect 36566 17700 36626 17960
rect 36714 17910 36774 18164
rect 37734 18164 37748 18192
rect 37782 18716 37796 18740
rect 38754 18740 38814 18900
rect 39268 18839 39328 18900
rect 39048 18833 39536 18839
rect 39048 18799 39060 18833
rect 39524 18799 39536 18833
rect 39048 18793 39536 18799
rect 37782 18192 37788 18716
rect 38754 18706 38766 18740
rect 38760 18204 38766 18706
rect 37782 18164 37794 18192
rect 37220 18111 37280 18112
rect 37012 18105 37500 18111
rect 37012 18071 37024 18105
rect 37488 18071 37500 18105
rect 37012 18065 37500 18071
rect 36708 17850 36714 17910
rect 36774 17850 36780 17910
rect 36560 17640 36566 17700
rect 36626 17640 36632 17700
rect 36712 17642 36718 17702
rect 36778 17642 36784 17702
rect 35994 17577 36482 17583
rect 35994 17543 36006 17577
rect 36470 17543 36482 17577
rect 35994 17537 36482 17543
rect 34728 16940 34734 17454
rect 35698 17452 35712 17484
rect 35706 16940 35712 17452
rect 34728 16908 34736 16940
rect 32940 16849 33428 16855
rect 32940 16815 32952 16849
rect 33416 16815 33428 16849
rect 32940 16809 33428 16815
rect 33958 16849 34446 16855
rect 33958 16815 33970 16849
rect 34434 16815 34446 16849
rect 33958 16809 34446 16815
rect 32640 16692 32646 16752
rect 32706 16692 32712 16752
rect 31106 16570 32194 16630
rect 32638 16582 32644 16642
rect 32704 16582 32710 16642
rect 30376 16428 31684 16488
rect 29886 16321 30374 16327
rect 29886 16287 29898 16321
rect 30362 16287 30374 16321
rect 29886 16281 30374 16287
rect 30904 16321 31392 16327
rect 30904 16287 30916 16321
rect 31380 16287 31392 16321
rect 30904 16281 31392 16287
rect 28620 15688 28626 16198
rect 29588 16170 29604 16228
rect 28620 15652 28634 15688
rect 29598 15684 29604 16170
rect 27850 15593 28338 15599
rect 27850 15559 27862 15593
rect 28326 15559 28338 15593
rect 27850 15553 28338 15559
rect 27546 15432 27552 15492
rect 27612 15432 27618 15492
rect 28054 15378 28114 15553
rect 24214 15302 24220 15362
rect 24280 15302 24286 15362
rect 26024 15318 28114 15378
rect 19372 15174 19376 15234
rect 19436 15174 23898 15234
rect 19376 15168 19436 15174
rect 19256 15116 19316 15122
rect 24220 15116 24280 15302
rect 19316 15056 24280 15116
rect 19256 15050 19316 15056
rect 18810 14998 18870 15004
rect 26024 14998 26084 15318
rect 28054 15108 28114 15318
rect 28574 15222 28634 15652
rect 29588 15652 29604 15684
rect 29638 16170 29648 16228
rect 30616 16228 30662 16240
rect 29638 15684 29644 16170
rect 30616 15696 30622 16228
rect 29638 15652 29648 15684
rect 28868 15593 29356 15599
rect 28868 15559 28880 15593
rect 29344 15559 29356 15593
rect 28868 15553 29356 15559
rect 29092 15498 29152 15553
rect 29588 15498 29648 15652
rect 30610 15652 30622 15696
rect 30656 15696 30662 16228
rect 31624 16228 31684 16428
rect 32134 16428 32194 16570
rect 32134 16327 32194 16368
rect 31922 16321 32410 16327
rect 31922 16287 31934 16321
rect 32398 16287 32410 16321
rect 31922 16281 32410 16287
rect 31624 16176 31640 16228
rect 30656 15652 30670 15696
rect 29886 15593 30374 15599
rect 29886 15559 29898 15593
rect 30362 15559 30374 15593
rect 29886 15553 30374 15559
rect 30104 15498 30164 15553
rect 30610 15498 30670 15652
rect 31634 15652 31640 16176
rect 31674 16176 31684 16228
rect 32644 16228 32704 16582
rect 33150 16428 33210 16809
rect 34180 16756 34240 16809
rect 34676 16756 34736 16908
rect 35700 16908 35712 16940
rect 35746 17452 35758 17484
rect 36718 17484 36778 17642
rect 37220 17583 37280 18065
rect 37734 17800 37794 18164
rect 38754 18164 38766 18204
rect 38800 18706 38814 18740
rect 39770 18740 39830 18900
rect 39770 18718 39784 18740
rect 38800 18204 38806 18706
rect 38800 18164 38814 18204
rect 38226 18111 38286 18118
rect 38030 18105 38518 18111
rect 38030 18071 38042 18105
rect 38506 18071 38518 18105
rect 38030 18065 38518 18071
rect 37728 17740 37734 17800
rect 37794 17740 37800 17800
rect 38226 17583 38286 18065
rect 38754 17910 38814 18164
rect 39778 18164 39784 18718
rect 39818 18718 39830 18740
rect 39818 18164 39824 18718
rect 39778 18152 39824 18164
rect 39048 18105 39536 18111
rect 39048 18071 39060 18105
rect 39524 18071 39536 18105
rect 39048 18065 39536 18071
rect 39894 17910 39954 20678
rect 40036 20510 40096 23226
rect 40324 20810 40330 20870
rect 40390 20810 40396 20870
rect 40036 20444 40096 20450
rect 40172 20150 40178 20210
rect 40238 20150 40244 20210
rect 40012 19008 40018 19068
rect 40078 19008 40084 19068
rect 38748 17850 38754 17910
rect 38814 17850 38820 17910
rect 39888 17850 39894 17910
rect 39954 17850 39960 17910
rect 38746 17642 38752 17702
rect 38812 17642 38818 17702
rect 37012 17577 37500 17583
rect 37012 17543 37024 17577
rect 37488 17543 37500 17577
rect 37012 17537 37500 17543
rect 38030 17577 38518 17583
rect 38030 17543 38042 17577
rect 38506 17543 38518 17577
rect 38030 17537 38518 17543
rect 36718 17464 36730 17484
rect 35746 16940 35752 17452
rect 35746 16908 35760 16940
rect 34976 16849 35464 16855
rect 34976 16815 34988 16849
rect 35452 16815 35464 16849
rect 34976 16809 35464 16815
rect 35192 16756 35252 16809
rect 34180 16696 35252 16756
rect 35700 16754 35760 16908
rect 36724 16908 36730 17464
rect 36764 17464 36778 17484
rect 37742 17484 37788 17496
rect 36764 16908 36770 17464
rect 37742 16936 37748 17484
rect 36724 16896 36770 16908
rect 37736 16908 37748 16936
rect 37782 16936 37788 17484
rect 38752 17484 38812 17642
rect 39048 17577 39536 17583
rect 39048 17543 39060 17577
rect 39524 17543 39536 17577
rect 39048 17537 39536 17543
rect 38752 17460 38766 17484
rect 38760 16944 38766 17460
rect 37782 16908 37796 16936
rect 36208 16855 36268 16862
rect 37232 16855 37292 16862
rect 35994 16849 36482 16855
rect 35994 16815 36006 16849
rect 36470 16815 36482 16849
rect 35994 16809 36482 16815
rect 37012 16849 37500 16855
rect 37012 16815 37024 16849
rect 37488 16815 37500 16849
rect 37012 16809 37500 16815
rect 33150 16362 33210 16368
rect 32940 16321 33428 16327
rect 32940 16287 32952 16321
rect 33416 16287 33428 16321
rect 32940 16281 33428 16287
rect 33958 16321 34446 16327
rect 33958 16287 33970 16321
rect 34434 16287 34446 16321
rect 33958 16281 34446 16287
rect 31674 15652 31680 16176
rect 32644 16164 32658 16228
rect 31634 15640 31680 15652
rect 32652 15652 32658 16164
rect 32692 16164 32704 16228
rect 33670 16228 33716 16240
rect 32692 15652 32698 16164
rect 33670 15680 33676 16228
rect 32652 15640 32698 15652
rect 33662 15652 33676 15680
rect 33710 15680 33716 16228
rect 34676 16228 34736 16696
rect 35694 16694 35700 16754
rect 35760 16694 35766 16754
rect 36208 16434 36268 16809
rect 36208 16428 36270 16434
rect 36208 16368 36210 16428
rect 36716 16380 36722 16440
rect 36782 16380 36788 16440
rect 36208 16362 36270 16368
rect 36208 16327 36268 16362
rect 34976 16321 35464 16327
rect 34976 16287 34988 16321
rect 35452 16287 35464 16321
rect 34976 16281 35464 16287
rect 35994 16321 36482 16327
rect 35994 16287 36006 16321
rect 36470 16287 36482 16321
rect 35994 16281 36482 16287
rect 34676 16190 34694 16228
rect 34688 15682 34694 16190
rect 33710 15652 33722 15680
rect 30904 15593 31392 15599
rect 30904 15559 30916 15593
rect 31380 15559 31392 15593
rect 30904 15553 31392 15559
rect 31922 15593 32410 15599
rect 31922 15559 31934 15593
rect 32398 15559 32410 15593
rect 31922 15553 32410 15559
rect 32940 15593 33428 15599
rect 32940 15559 32952 15593
rect 33416 15559 33428 15593
rect 32940 15553 33428 15559
rect 31120 15498 31180 15553
rect 33146 15498 33206 15553
rect 33662 15498 33722 15652
rect 34676 15652 34694 15682
rect 34728 16190 34736 16228
rect 35706 16228 35752 16240
rect 34728 15682 34734 16190
rect 34728 15652 34736 15682
rect 35706 15678 35712 16228
rect 33958 15593 34446 15599
rect 33958 15559 33970 15593
rect 34434 15559 34446 15593
rect 33958 15553 34446 15559
rect 34180 15498 34240 15553
rect 34676 15498 34736 15652
rect 35704 15652 35712 15678
rect 35746 15678 35752 16228
rect 36722 16228 36782 16380
rect 37232 16327 37292 16809
rect 37736 16754 37796 16908
rect 38752 16908 38766 16944
rect 38800 17460 38812 17484
rect 39778 17484 39824 17496
rect 38800 16944 38806 17460
rect 38800 16908 38812 16944
rect 39778 16932 39784 17484
rect 38238 16855 38298 16868
rect 38030 16849 38518 16855
rect 38030 16815 38042 16849
rect 38506 16815 38518 16849
rect 38030 16809 38518 16815
rect 37730 16694 37736 16754
rect 37796 16694 37802 16754
rect 38238 16327 38298 16809
rect 38752 16750 38812 16908
rect 39768 16908 39784 16932
rect 39818 16932 39824 17484
rect 39818 16908 39828 16932
rect 39048 16849 39536 16855
rect 39048 16815 39060 16849
rect 39524 16815 39536 16849
rect 39048 16809 39536 16815
rect 39266 16750 39326 16809
rect 39768 16750 39828 16908
rect 38752 16690 39828 16750
rect 39894 16642 39954 17850
rect 40018 17702 40078 19008
rect 40012 17642 40018 17702
rect 40078 17642 40084 17702
rect 39888 16582 39894 16642
rect 39954 16582 39960 16642
rect 38750 16380 38756 16440
rect 38816 16380 38822 16440
rect 37012 16321 37500 16327
rect 37012 16287 37024 16321
rect 37488 16287 37500 16321
rect 37012 16281 37500 16287
rect 38030 16321 38518 16327
rect 38030 16287 38042 16321
rect 38506 16287 38518 16321
rect 38030 16281 38518 16287
rect 36722 16202 36730 16228
rect 35746 15652 35764 15678
rect 34976 15593 35464 15599
rect 34976 15559 34988 15593
rect 35452 15559 35464 15593
rect 34976 15553 35464 15559
rect 35192 15498 35252 15553
rect 29092 15438 35252 15498
rect 35704 15492 35764 15652
rect 36724 15652 36730 16202
rect 36764 16202 36782 16228
rect 37742 16228 37788 16240
rect 36764 15652 36770 16202
rect 37742 15674 37748 16228
rect 36724 15640 36770 15652
rect 37740 15652 37748 15674
rect 37782 15674 37788 16228
rect 38756 16228 38816 16380
rect 39048 16321 39536 16327
rect 39048 16287 39060 16321
rect 39524 16287 39536 16321
rect 39048 16281 39536 16287
rect 38756 16198 38766 16228
rect 38760 15690 38766 16198
rect 37782 15652 37800 15674
rect 36212 15599 36272 15606
rect 35994 15593 36482 15599
rect 35994 15559 36006 15593
rect 36470 15559 36482 15593
rect 35994 15553 36482 15559
rect 37012 15593 37500 15599
rect 37012 15559 37024 15593
rect 37488 15559 37500 15593
rect 37012 15553 37500 15559
rect 35698 15432 35704 15492
rect 35764 15432 35770 15492
rect 36212 15380 36272 15553
rect 37232 15380 37292 15553
rect 37740 15492 37800 15652
rect 38754 15652 38766 15690
rect 38800 16198 38816 16228
rect 39778 16228 39824 16240
rect 38800 15690 38806 16198
rect 38800 15652 38814 15690
rect 39778 15678 39784 16228
rect 38030 15593 38518 15599
rect 38030 15559 38042 15593
rect 38506 15559 38518 15593
rect 38030 15553 38518 15559
rect 37734 15432 37740 15492
rect 37800 15432 37806 15492
rect 38234 15380 38294 15553
rect 38754 15496 38814 15652
rect 39770 15652 39784 15678
rect 39818 15678 39824 16228
rect 39818 15652 39830 15678
rect 39048 15593 39536 15599
rect 39048 15559 39060 15593
rect 39524 15559 39536 15593
rect 39048 15553 39536 15559
rect 39268 15496 39328 15553
rect 39770 15496 39830 15652
rect 38754 15436 39830 15496
rect 36212 15320 38294 15380
rect 28568 15162 28574 15222
rect 28634 15162 28640 15222
rect 36212 15108 36272 15320
rect 40178 15222 40238 20150
rect 40330 18954 40390 20810
rect 40324 18894 40330 18954
rect 40390 18894 40396 18954
rect 41756 15352 41762 28782
rect 41862 15352 41868 28782
rect 40172 15162 40178 15222
rect 40238 15162 40244 15222
rect 28054 15048 36272 15108
rect 18870 14938 26084 14998
rect 18810 14932 18870 14938
rect 41756 14838 41868 15352
rect 17412 14832 41868 14838
rect 17412 14732 17518 14832
rect 41762 14732 41868 14832
rect 17412 14726 41868 14732
rect 14174 14410 14318 14702
rect 3048 14102 14318 14410
rect 3048 13908 15400 14102
rect 3048 13902 41968 13908
rect 3048 13802 4818 13902
rect 41862 13802 41968 13902
rect 3048 13796 41968 13802
rect 3048 13780 15398 13796
rect 4712 13010 4824 13780
rect 18928 13722 18988 13728
rect 19250 13672 19256 13732
rect 19316 13672 19322 13732
rect 19376 13724 19436 13730
rect 18316 13526 18322 13586
rect 18382 13526 18388 13586
rect 18436 13528 18442 13588
rect 18502 13528 18508 13588
rect 18576 13546 18582 13606
rect 18642 13546 18648 13606
rect 18804 13562 18810 13622
rect 18870 13562 18876 13622
rect 18184 13398 18190 13458
rect 18250 13398 18256 13458
rect 4712 12860 4718 13010
rect 4662 12790 4718 12860
rect 4818 12860 4824 13010
rect 4818 12790 5100 12860
rect 15472 12800 15478 12860
rect 15538 12800 15544 12860
rect 4662 1198 4704 12790
rect 4962 1198 5100 12790
rect 15478 12756 15538 12800
rect 7844 12696 15538 12756
rect 7844 12556 7904 12696
rect 8354 12646 8414 12696
rect 8138 12640 8626 12646
rect 8138 12606 8150 12640
rect 8614 12606 8626 12640
rect 8138 12600 8626 12606
rect 7844 12526 7856 12556
rect 7850 11998 7856 12526
rect 7840 11980 7856 11998
rect 7890 12526 7904 12556
rect 8860 12556 8920 12696
rect 9362 12646 9422 12696
rect 10390 12646 10450 12696
rect 9156 12640 9644 12646
rect 9156 12606 9168 12640
rect 9632 12606 9644 12640
rect 9156 12600 9644 12606
rect 10174 12640 10662 12646
rect 10174 12606 10186 12640
rect 10650 12606 10662 12640
rect 10174 12600 10662 12606
rect 8860 12532 8874 12556
rect 7890 11998 7896 12526
rect 8868 12002 8874 12532
rect 7890 11980 7900 11998
rect 7840 11738 7900 11980
rect 8860 11980 8874 12002
rect 8908 12532 8920 12556
rect 9886 12556 9932 12568
rect 8908 12002 8914 12532
rect 9886 12004 9892 12556
rect 8908 11980 8920 12002
rect 8138 11930 8626 11936
rect 8138 11896 8150 11930
rect 8614 11896 8626 11930
rect 8138 11890 8626 11896
rect 8354 11828 8414 11890
rect 8138 11822 8626 11828
rect 8138 11788 8150 11822
rect 8614 11788 8626 11822
rect 8138 11782 8626 11788
rect 7840 11708 7856 11738
rect 7850 11184 7856 11708
rect 7842 11162 7856 11184
rect 7890 11708 7900 11738
rect 8860 11738 8920 11980
rect 9880 11980 9892 12004
rect 9926 12004 9932 12556
rect 10898 12556 10958 12696
rect 11404 12646 11464 12696
rect 12418 12646 12478 12696
rect 11192 12640 11680 12646
rect 11192 12606 11204 12640
rect 11668 12606 11680 12640
rect 11192 12600 11680 12606
rect 12210 12640 12698 12646
rect 12210 12606 12222 12640
rect 12686 12606 12698 12640
rect 12210 12600 12698 12606
rect 10898 12518 10910 12556
rect 9926 11980 9940 12004
rect 10904 12000 10910 12518
rect 9156 11930 9644 11936
rect 9156 11896 9168 11930
rect 9632 11896 9644 11930
rect 9156 11890 9644 11896
rect 9358 11828 9418 11890
rect 9156 11822 9644 11828
rect 9156 11788 9168 11822
rect 9632 11788 9644 11822
rect 9156 11782 9644 11788
rect 8860 11712 8874 11738
rect 7890 11184 7896 11708
rect 8868 11188 8874 11712
rect 7890 11162 7902 11184
rect 7842 10920 7902 11162
rect 8862 11162 8874 11188
rect 8908 11712 8920 11738
rect 9880 11738 9940 11980
rect 10898 11980 10910 12000
rect 10944 12518 10958 12556
rect 11922 12556 11968 12568
rect 12934 12556 12994 12696
rect 13450 12646 13510 12696
rect 14456 12646 14516 12696
rect 13228 12640 13716 12646
rect 13228 12606 13240 12640
rect 13704 12606 13716 12640
rect 13228 12600 13716 12606
rect 14246 12640 14734 12646
rect 14246 12606 14258 12640
rect 14722 12606 14734 12640
rect 14246 12600 14734 12606
rect 10944 12000 10950 12518
rect 11922 12008 11928 12556
rect 10944 11980 10958 12000
rect 10174 11930 10662 11936
rect 10174 11896 10186 11930
rect 10650 11896 10662 11930
rect 10174 11890 10662 11896
rect 10388 11828 10448 11890
rect 10174 11822 10662 11828
rect 10174 11788 10186 11822
rect 10650 11788 10662 11822
rect 10174 11782 10662 11788
rect 9880 11714 9892 11738
rect 8908 11188 8914 11712
rect 9886 11190 9892 11714
rect 8908 11162 8922 11188
rect 8138 11112 8626 11118
rect 8138 11078 8150 11112
rect 8614 11078 8626 11112
rect 8138 11072 8626 11078
rect 8354 11010 8414 11072
rect 8138 11004 8626 11010
rect 8138 10970 8150 11004
rect 8614 10970 8626 11004
rect 8138 10964 8626 10970
rect 7842 10894 7856 10920
rect 7850 10356 7856 10894
rect 7842 10344 7856 10356
rect 7890 10894 7902 10920
rect 8862 10920 8922 11162
rect 9882 11162 9892 11190
rect 9926 11714 9940 11738
rect 10898 11738 10958 11980
rect 11918 11980 11928 12008
rect 11962 12008 11968 12556
rect 12932 12522 12946 12556
rect 12934 12510 12946 12522
rect 11962 11980 11978 12008
rect 12940 12000 12946 12510
rect 11192 11930 11680 11936
rect 11192 11896 11204 11930
rect 11668 11896 11680 11930
rect 11192 11890 11680 11896
rect 11390 11828 11450 11890
rect 11192 11822 11680 11828
rect 11192 11788 11204 11822
rect 11668 11788 11680 11822
rect 11192 11782 11680 11788
rect 9926 11190 9932 11714
rect 10898 11710 10910 11738
rect 9926 11162 9942 11190
rect 10904 11186 10910 11710
rect 9156 11112 9644 11118
rect 9156 11078 9168 11112
rect 9632 11078 9644 11112
rect 9156 11072 9644 11078
rect 9370 11010 9430 11072
rect 9156 11004 9644 11010
rect 9156 10970 9168 11004
rect 9632 10970 9644 11004
rect 9156 10964 9644 10970
rect 8862 10898 8874 10920
rect 7890 10356 7896 10894
rect 8868 10360 8874 10898
rect 7890 10344 7902 10356
rect 7842 10102 7902 10344
rect 8862 10344 8874 10360
rect 8908 10898 8922 10920
rect 9882 10920 9942 11162
rect 10900 11162 10910 11186
rect 10944 11710 10958 11738
rect 11918 11738 11978 11980
rect 12930 11980 12946 12000
rect 12980 12510 12994 12556
rect 13958 12556 14004 12568
rect 12980 12000 12986 12510
rect 13958 12000 13964 12556
rect 12980 11980 12990 12000
rect 12210 11930 12698 11936
rect 12210 11896 12222 11930
rect 12686 11896 12698 11930
rect 12210 11890 12698 11896
rect 12420 11828 12480 11890
rect 12210 11822 12698 11828
rect 12210 11788 12222 11822
rect 12686 11788 12698 11822
rect 12210 11782 12698 11788
rect 11918 11718 11928 11738
rect 10944 11186 10950 11710
rect 11922 11194 11928 11718
rect 10944 11162 10960 11186
rect 10174 11112 10662 11118
rect 10174 11078 10186 11112
rect 10650 11078 10662 11112
rect 10174 11072 10662 11078
rect 10388 11010 10448 11072
rect 10174 11004 10662 11010
rect 10174 10970 10186 11004
rect 10650 10970 10662 11004
rect 10174 10964 10662 10970
rect 9882 10900 9892 10920
rect 8908 10360 8914 10898
rect 9886 10362 9892 10900
rect 8908 10344 8922 10360
rect 8138 10294 8626 10300
rect 8138 10260 8150 10294
rect 8614 10260 8626 10294
rect 8138 10254 8626 10260
rect 8348 10192 8408 10254
rect 8138 10186 8626 10192
rect 8138 10152 8150 10186
rect 8614 10152 8626 10186
rect 8138 10146 8626 10152
rect 7842 10066 7856 10102
rect 7850 9544 7856 10066
rect 7842 9526 7856 9544
rect 7890 10066 7902 10102
rect 8862 10102 8922 10344
rect 9882 10344 9892 10362
rect 9926 10900 9942 10920
rect 10900 10920 10960 11162
rect 11920 11162 11928 11194
rect 11962 11718 11978 11738
rect 12930 11738 12990 11980
rect 13952 11980 13964 12000
rect 13998 12000 14004 12556
rect 14968 12556 15028 12696
rect 15478 12646 15538 12696
rect 16998 12666 17004 12726
rect 17064 12666 17070 12726
rect 15264 12640 15752 12646
rect 15264 12606 15276 12640
rect 15740 12606 15752 12640
rect 15264 12600 15752 12606
rect 16282 12640 16770 12646
rect 16282 12606 16294 12640
rect 16758 12606 16770 12640
rect 16282 12600 16770 12606
rect 14968 12520 14982 12556
rect 14976 12000 14982 12520
rect 13998 11980 14012 12000
rect 13228 11930 13716 11936
rect 13228 11896 13240 11930
rect 13704 11896 13716 11930
rect 13228 11890 13716 11896
rect 13436 11828 13496 11890
rect 13228 11822 13716 11828
rect 13228 11788 13240 11822
rect 13704 11788 13716 11822
rect 13228 11782 13716 11788
rect 11962 11194 11968 11718
rect 12930 11710 12946 11738
rect 11962 11162 11980 11194
rect 12940 11186 12946 11710
rect 11192 11112 11680 11118
rect 11192 11078 11204 11112
rect 11668 11078 11680 11112
rect 11192 11072 11680 11078
rect 11390 11010 11450 11072
rect 11192 11004 11680 11010
rect 11192 10970 11204 11004
rect 11668 10970 11680 11004
rect 11192 10964 11680 10970
rect 9926 10362 9932 10900
rect 10900 10896 10910 10920
rect 9926 10344 9942 10362
rect 10904 10358 10910 10896
rect 9156 10294 9644 10300
rect 9156 10260 9168 10294
rect 9632 10260 9644 10294
rect 9156 10254 9644 10260
rect 9370 10192 9430 10254
rect 9156 10186 9644 10192
rect 9156 10152 9168 10186
rect 9632 10152 9644 10186
rect 9156 10146 9644 10152
rect 8862 10070 8874 10102
rect 7890 9544 7896 10066
rect 8868 9548 8874 10070
rect 7890 9526 7902 9544
rect 7842 9284 7902 9526
rect 8862 9526 8874 9548
rect 8908 10070 8922 10102
rect 9882 10102 9942 10344
rect 10900 10344 10910 10358
rect 10944 10896 10960 10920
rect 11920 10920 11980 11162
rect 12932 11162 12946 11186
rect 12980 11710 12990 11738
rect 13952 11738 14012 11980
rect 14972 11980 14982 12000
rect 15016 12520 15028 12556
rect 15994 12556 16040 12568
rect 15016 12000 15022 12520
rect 15994 12004 16000 12556
rect 15016 11980 15032 12000
rect 14246 11930 14734 11936
rect 14246 11896 14258 11930
rect 14722 11896 14734 11930
rect 14246 11890 14734 11896
rect 14458 11828 14518 11890
rect 14246 11822 14734 11828
rect 14246 11788 14258 11822
rect 14722 11788 14734 11822
rect 14246 11782 14734 11788
rect 13952 11710 13964 11738
rect 12980 11186 12986 11710
rect 13958 11186 13964 11710
rect 12980 11162 12992 11186
rect 12210 11112 12698 11118
rect 12210 11078 12222 11112
rect 12686 11078 12698 11112
rect 12210 11072 12698 11078
rect 12420 11010 12480 11072
rect 12210 11004 12698 11010
rect 12210 10970 12222 11004
rect 12686 10970 12698 11004
rect 12210 10964 12698 10970
rect 11920 10904 11928 10920
rect 10944 10358 10950 10896
rect 11922 10366 11928 10904
rect 10944 10344 10960 10358
rect 10174 10294 10662 10300
rect 10174 10260 10186 10294
rect 10650 10260 10662 10294
rect 10174 10254 10662 10260
rect 10382 10192 10442 10254
rect 10174 10186 10662 10192
rect 10174 10152 10186 10186
rect 10650 10152 10662 10186
rect 10174 10146 10662 10152
rect 9882 10072 9892 10102
rect 8908 9548 8914 10070
rect 9886 9550 9892 10072
rect 8908 9526 8922 9548
rect 8138 9476 8626 9482
rect 8138 9442 8150 9476
rect 8614 9442 8626 9476
rect 8138 9436 8626 9442
rect 8346 9374 8406 9436
rect 8138 9368 8626 9374
rect 8138 9334 8150 9368
rect 8614 9334 8626 9368
rect 8138 9328 8626 9334
rect 7842 9254 7856 9284
rect 7850 8724 7856 9254
rect 7842 8708 7856 8724
rect 7890 9254 7902 9284
rect 8862 9284 8922 9526
rect 9882 9526 9892 9550
rect 9926 10072 9942 10102
rect 10900 10102 10960 10344
rect 11920 10344 11928 10366
rect 11962 10904 11980 10920
rect 12932 10920 12992 11162
rect 13954 11162 13964 11186
rect 13998 11710 14012 11738
rect 14972 11738 15032 11980
rect 15988 11980 16000 12004
rect 16034 12004 16040 12556
rect 17004 12556 17064 12666
rect 17004 12520 17018 12556
rect 16034 11980 16048 12004
rect 17012 12000 17018 12520
rect 15264 11930 15752 11936
rect 15264 11896 15276 11930
rect 15740 11896 15752 11930
rect 15264 11890 15752 11896
rect 15470 11828 15530 11890
rect 15264 11822 15752 11828
rect 15264 11788 15276 11822
rect 15740 11788 15752 11822
rect 15264 11782 15752 11788
rect 14972 11710 14982 11738
rect 13998 11186 14004 11710
rect 14976 11186 14982 11710
rect 13998 11162 14014 11186
rect 13228 11112 13716 11118
rect 13228 11078 13240 11112
rect 13704 11078 13716 11112
rect 13228 11072 13716 11078
rect 13436 11010 13496 11072
rect 13228 11004 13716 11010
rect 13228 10970 13240 11004
rect 13704 10970 13716 11004
rect 13228 10964 13716 10970
rect 11962 10366 11968 10904
rect 12932 10896 12946 10920
rect 11962 10344 11980 10366
rect 12940 10358 12946 10896
rect 11192 10294 11680 10300
rect 11192 10260 11204 10294
rect 11668 10260 11680 10294
rect 11192 10254 11680 10260
rect 11384 10192 11444 10254
rect 11192 10186 11680 10192
rect 11192 10152 11204 10186
rect 11668 10152 11680 10186
rect 11192 10146 11680 10152
rect 9926 9550 9932 10072
rect 10900 10068 10910 10102
rect 9926 9526 9942 9550
rect 10904 9546 10910 10068
rect 9156 9476 9644 9482
rect 9156 9442 9168 9476
rect 9632 9442 9644 9476
rect 9156 9436 9644 9442
rect 9364 9374 9424 9436
rect 9156 9368 9644 9374
rect 9156 9334 9168 9368
rect 9632 9334 9644 9368
rect 9156 9328 9644 9334
rect 8862 9258 8874 9284
rect 7890 8724 7896 9254
rect 8868 8728 8874 9258
rect 7890 8708 7902 8724
rect 7842 8466 7902 8708
rect 8862 8708 8874 8728
rect 8908 9258 8922 9284
rect 9882 9284 9942 9526
rect 10900 9526 10910 9546
rect 10944 10068 10960 10102
rect 11920 10102 11980 10344
rect 12932 10344 12946 10358
rect 12980 10896 12992 10920
rect 13954 10920 14014 11162
rect 14974 11162 14982 11186
rect 15016 11710 15032 11738
rect 15988 11738 16048 11980
rect 17010 11980 17018 12000
rect 17052 12520 17064 12556
rect 17052 12000 17058 12520
rect 17052 11980 17070 12000
rect 16282 11930 16770 11936
rect 16282 11896 16294 11930
rect 16758 11896 16770 11930
rect 16282 11890 16770 11896
rect 16490 11828 16550 11890
rect 16282 11822 16770 11828
rect 16282 11788 16294 11822
rect 16758 11788 16770 11822
rect 16282 11782 16770 11788
rect 15988 11714 16000 11738
rect 15016 11186 15022 11710
rect 15994 11190 16000 11714
rect 15016 11162 15034 11186
rect 14246 11112 14734 11118
rect 14246 11078 14258 11112
rect 14722 11078 14734 11112
rect 14246 11072 14734 11078
rect 14458 11010 14518 11072
rect 14246 11004 14734 11010
rect 14246 10970 14258 11004
rect 14722 10970 14734 11004
rect 14246 10964 14734 10970
rect 13954 10896 13964 10920
rect 12980 10358 12986 10896
rect 13958 10358 13964 10896
rect 12980 10344 12992 10358
rect 12210 10294 12698 10300
rect 12210 10260 12222 10294
rect 12686 10260 12698 10294
rect 12210 10254 12698 10260
rect 12414 10192 12474 10254
rect 12210 10186 12698 10192
rect 12210 10152 12222 10186
rect 12686 10152 12698 10186
rect 12210 10146 12698 10152
rect 11920 10076 11928 10102
rect 10944 9546 10950 10068
rect 11922 9554 11928 10076
rect 10944 9526 10960 9546
rect 10174 9476 10662 9482
rect 10174 9442 10186 9476
rect 10650 9442 10662 9476
rect 10174 9436 10662 9442
rect 10380 9374 10440 9436
rect 10174 9368 10662 9374
rect 10174 9334 10186 9368
rect 10650 9334 10662 9368
rect 10174 9328 10662 9334
rect 9882 9260 9892 9284
rect 8908 8728 8914 9258
rect 9886 8730 9892 9260
rect 8908 8708 8922 8728
rect 8138 8658 8626 8664
rect 8138 8624 8150 8658
rect 8614 8624 8626 8658
rect 8138 8618 8626 8624
rect 8348 8556 8408 8618
rect 8138 8550 8626 8556
rect 8138 8516 8150 8550
rect 8614 8516 8626 8550
rect 8138 8510 8626 8516
rect 7842 8434 7856 8466
rect 7850 7912 7856 8434
rect 7842 7890 7856 7912
rect 7890 8434 7902 8466
rect 8862 8466 8922 8708
rect 9882 8708 9892 8730
rect 9926 9260 9942 9284
rect 10900 9284 10960 9526
rect 11920 9526 11928 9554
rect 11962 10076 11980 10102
rect 12932 10102 12992 10344
rect 13954 10344 13964 10358
rect 13998 10896 14014 10920
rect 14974 10920 15034 11162
rect 15990 11162 16000 11190
rect 16034 11714 16048 11738
rect 17010 11738 17070 11980
rect 16034 11190 16040 11714
rect 17010 11710 17018 11738
rect 16034 11162 16050 11190
rect 15264 11112 15752 11118
rect 15264 11078 15276 11112
rect 15740 11078 15752 11112
rect 15264 11072 15752 11078
rect 15470 11010 15530 11072
rect 15264 11004 15752 11010
rect 15264 10970 15276 11004
rect 15740 10970 15752 11004
rect 15264 10964 15752 10970
rect 14974 10896 14982 10920
rect 13998 10358 14004 10896
rect 14976 10358 14982 10896
rect 13998 10344 14014 10358
rect 13228 10294 13716 10300
rect 13228 10260 13240 10294
rect 13704 10260 13716 10294
rect 13228 10254 13716 10260
rect 13430 10192 13490 10254
rect 13228 10186 13716 10192
rect 13228 10152 13240 10186
rect 13704 10152 13716 10186
rect 13228 10146 13716 10152
rect 11962 9554 11968 10076
rect 12932 10068 12946 10102
rect 11962 9526 11980 9554
rect 12940 9546 12946 10068
rect 11192 9476 11680 9482
rect 11192 9442 11204 9476
rect 11668 9442 11680 9476
rect 11192 9436 11680 9442
rect 11382 9374 11442 9436
rect 11192 9368 11680 9374
rect 11192 9334 11204 9368
rect 11668 9334 11680 9368
rect 11192 9328 11680 9334
rect 9926 8730 9932 9260
rect 10900 9256 10910 9284
rect 9926 8708 9942 8730
rect 10904 8726 10910 9256
rect 9156 8658 9644 8664
rect 9156 8624 9168 8658
rect 9632 8624 9644 8658
rect 9156 8618 9644 8624
rect 9362 8556 9422 8618
rect 9156 8550 9644 8556
rect 9156 8516 9168 8550
rect 9632 8516 9644 8550
rect 9156 8510 9644 8516
rect 8862 8438 8874 8466
rect 7890 7912 7896 8434
rect 8868 7916 8874 8438
rect 7890 7890 7902 7912
rect 7842 7648 7902 7890
rect 8862 7890 8874 7916
rect 8908 8438 8922 8466
rect 9882 8466 9942 8708
rect 10900 8708 10910 8726
rect 10944 9256 10960 9284
rect 11920 9284 11980 9526
rect 12932 9526 12946 9546
rect 12980 10068 12992 10102
rect 13954 10102 14014 10344
rect 14974 10344 14982 10358
rect 15016 10896 15034 10920
rect 15990 10920 16050 11162
rect 17012 11162 17018 11710
rect 17052 11710 17070 11738
rect 17052 11186 17058 11710
rect 17052 11162 17072 11186
rect 16282 11112 16770 11118
rect 16282 11078 16294 11112
rect 16758 11078 16770 11112
rect 16282 11072 16770 11078
rect 16490 11010 16550 11072
rect 16282 11004 16770 11010
rect 16282 10970 16294 11004
rect 16758 10970 16770 11004
rect 16282 10964 16770 10970
rect 15990 10900 16000 10920
rect 15016 10358 15022 10896
rect 15994 10362 16000 10900
rect 15016 10344 15034 10358
rect 14246 10294 14734 10300
rect 14246 10260 14258 10294
rect 14722 10260 14734 10294
rect 14246 10254 14734 10260
rect 14452 10192 14512 10254
rect 14246 10186 14734 10192
rect 14246 10152 14258 10186
rect 14722 10152 14734 10186
rect 14246 10146 14734 10152
rect 13954 10068 13964 10102
rect 12980 9546 12986 10068
rect 13958 9546 13964 10068
rect 12980 9526 12992 9546
rect 12210 9476 12698 9482
rect 12210 9442 12222 9476
rect 12686 9442 12698 9476
rect 12210 9436 12698 9442
rect 12412 9374 12472 9436
rect 12210 9368 12698 9374
rect 12210 9334 12222 9368
rect 12686 9334 12698 9368
rect 12210 9328 12698 9334
rect 11920 9264 11928 9284
rect 10944 8726 10950 9256
rect 11922 8734 11928 9264
rect 10944 8708 10960 8726
rect 10174 8658 10662 8664
rect 10174 8624 10186 8658
rect 10650 8624 10662 8658
rect 10174 8618 10662 8624
rect 10382 8556 10442 8618
rect 10174 8550 10662 8556
rect 10174 8516 10186 8550
rect 10650 8516 10662 8550
rect 10174 8510 10662 8516
rect 9882 8440 9892 8466
rect 8908 7916 8914 8438
rect 9886 7918 9892 8440
rect 8908 7890 8922 7916
rect 8138 7840 8626 7846
rect 8138 7806 8150 7840
rect 8614 7806 8626 7840
rect 8138 7800 8626 7806
rect 8350 7738 8410 7800
rect 8138 7732 8626 7738
rect 8138 7698 8150 7732
rect 8614 7698 8626 7732
rect 8138 7692 8626 7698
rect 7842 7622 7856 7648
rect 7850 7094 7856 7622
rect 7842 7072 7856 7094
rect 7890 7622 7902 7648
rect 8862 7648 8922 7890
rect 9882 7890 9892 7918
rect 9926 8440 9942 8466
rect 10900 8466 10960 8708
rect 11920 8708 11928 8734
rect 11962 9264 11980 9284
rect 12932 9284 12992 9526
rect 13954 9526 13964 9546
rect 13998 10068 14014 10102
rect 14974 10102 15034 10344
rect 15990 10344 16000 10362
rect 16034 10900 16050 10920
rect 17012 10920 17072 11162
rect 16034 10362 16040 10900
rect 16034 10344 16050 10362
rect 15264 10294 15752 10300
rect 15264 10260 15276 10294
rect 15740 10260 15752 10294
rect 15264 10254 15752 10260
rect 15464 10192 15524 10254
rect 15264 10186 15752 10192
rect 15264 10152 15276 10186
rect 15740 10152 15752 10186
rect 15264 10146 15752 10152
rect 14974 10068 14982 10102
rect 13998 9546 14004 10068
rect 14976 9546 14982 10068
rect 13998 9526 14014 9546
rect 13228 9476 13716 9482
rect 13228 9442 13240 9476
rect 13704 9442 13716 9476
rect 13228 9436 13716 9442
rect 13428 9374 13488 9436
rect 13228 9368 13716 9374
rect 13228 9334 13240 9368
rect 13704 9334 13716 9368
rect 13228 9328 13716 9334
rect 11962 8734 11968 9264
rect 12932 9256 12946 9284
rect 11962 8708 11980 8734
rect 12940 8726 12946 9256
rect 11192 8658 11680 8664
rect 11192 8624 11204 8658
rect 11668 8624 11680 8658
rect 11192 8618 11680 8624
rect 11384 8556 11444 8618
rect 11192 8550 11680 8556
rect 11192 8516 11204 8550
rect 11668 8516 11680 8550
rect 11192 8510 11680 8516
rect 9926 7918 9932 8440
rect 10900 8436 10910 8466
rect 9926 7890 9942 7918
rect 10904 7914 10910 8436
rect 9156 7840 9644 7846
rect 9156 7806 9168 7840
rect 9632 7806 9644 7840
rect 9156 7800 9644 7806
rect 9364 7738 9424 7800
rect 9156 7732 9644 7738
rect 9156 7698 9168 7732
rect 9632 7698 9644 7732
rect 9156 7692 9644 7698
rect 8862 7626 8874 7648
rect 7890 7094 7896 7622
rect 8868 7098 8874 7626
rect 7890 7072 7902 7094
rect 7842 6830 7902 7072
rect 8862 7072 8874 7098
rect 8908 7626 8922 7648
rect 9882 7648 9942 7890
rect 10900 7890 10910 7914
rect 10944 8436 10960 8466
rect 11920 8466 11980 8708
rect 12932 8708 12946 8726
rect 12980 9256 12992 9284
rect 13954 9284 14014 9526
rect 14974 9526 14982 9546
rect 15016 10068 15034 10102
rect 15990 10102 16050 10344
rect 17012 10344 17018 10920
rect 17052 10896 17072 10920
rect 17052 10358 17058 10896
rect 17052 10344 17072 10358
rect 16282 10294 16770 10300
rect 16282 10260 16294 10294
rect 16758 10260 16770 10294
rect 16282 10254 16770 10260
rect 16484 10192 16544 10254
rect 16282 10186 16770 10192
rect 16282 10152 16294 10186
rect 16758 10152 16770 10186
rect 16282 10146 16770 10152
rect 15990 10072 16000 10102
rect 15016 9546 15022 10068
rect 15994 9550 16000 10072
rect 15016 9526 15034 9546
rect 14246 9476 14734 9482
rect 14246 9442 14258 9476
rect 14722 9442 14734 9476
rect 14246 9436 14734 9442
rect 14450 9374 14510 9436
rect 14246 9368 14734 9374
rect 14246 9334 14258 9368
rect 14722 9334 14734 9368
rect 14246 9328 14734 9334
rect 13954 9256 13964 9284
rect 12980 8726 12986 9256
rect 13958 8726 13964 9256
rect 12980 8708 12992 8726
rect 12210 8658 12698 8664
rect 12210 8624 12222 8658
rect 12686 8624 12698 8658
rect 12210 8618 12698 8624
rect 12414 8556 12474 8618
rect 12210 8550 12698 8556
rect 12210 8516 12222 8550
rect 12686 8516 12698 8550
rect 12210 8510 12698 8516
rect 11920 8444 11928 8466
rect 10944 7914 10950 8436
rect 11922 7922 11928 8444
rect 10944 7890 10960 7914
rect 10174 7840 10662 7846
rect 10174 7806 10186 7840
rect 10650 7806 10662 7840
rect 10174 7800 10662 7806
rect 10384 7738 10444 7800
rect 10174 7732 10662 7738
rect 10174 7698 10186 7732
rect 10650 7698 10662 7732
rect 10174 7692 10662 7698
rect 9882 7628 9892 7648
rect 8908 7098 8914 7626
rect 9886 7100 9892 7628
rect 8908 7072 8922 7098
rect 8138 7022 8626 7028
rect 8138 6988 8150 7022
rect 8614 6988 8626 7022
rect 8138 6982 8626 6988
rect 8352 6920 8412 6982
rect 8138 6914 8626 6920
rect 8138 6880 8150 6914
rect 8614 6880 8626 6914
rect 8138 6874 8626 6880
rect 7842 6804 7856 6830
rect 7850 6254 7856 6804
rect 7890 6804 7902 6830
rect 8862 6830 8922 7072
rect 9882 7072 9892 7100
rect 9926 7628 9942 7648
rect 10900 7648 10960 7890
rect 11920 7890 11928 7922
rect 11962 8444 11980 8466
rect 12932 8466 12992 8708
rect 13954 8708 13964 8726
rect 13998 9256 14014 9284
rect 14974 9284 15034 9526
rect 15990 9526 16000 9550
rect 16034 10072 16050 10102
rect 17012 10102 17072 10344
rect 16034 9550 16040 10072
rect 16034 9526 16050 9550
rect 15264 9476 15752 9482
rect 15264 9442 15276 9476
rect 15740 9442 15752 9476
rect 15264 9436 15752 9442
rect 15462 9374 15522 9436
rect 15264 9368 15752 9374
rect 15264 9334 15276 9368
rect 15740 9334 15752 9368
rect 15264 9328 15752 9334
rect 14974 9256 14982 9284
rect 13998 8726 14004 9256
rect 14976 8726 14982 9256
rect 13998 8708 14014 8726
rect 13228 8658 13716 8664
rect 13228 8624 13240 8658
rect 13704 8624 13716 8658
rect 13228 8618 13716 8624
rect 13430 8556 13490 8618
rect 13228 8550 13716 8556
rect 13228 8516 13240 8550
rect 13704 8516 13716 8550
rect 13228 8510 13716 8516
rect 11962 7922 11968 8444
rect 12932 8436 12946 8466
rect 11962 7890 11980 7922
rect 12940 7914 12946 8436
rect 11192 7840 11680 7846
rect 11192 7806 11204 7840
rect 11668 7806 11680 7840
rect 11192 7800 11680 7806
rect 11386 7738 11446 7800
rect 11192 7732 11680 7738
rect 11192 7698 11204 7732
rect 11668 7698 11680 7732
rect 11192 7692 11680 7698
rect 9926 7100 9932 7628
rect 10900 7624 10910 7648
rect 9926 7072 9942 7100
rect 10904 7096 10910 7624
rect 9156 7022 9644 7028
rect 9156 6988 9168 7022
rect 9632 6988 9644 7022
rect 9156 6982 9644 6988
rect 9366 6920 9426 6982
rect 9156 6914 9644 6920
rect 9156 6880 9168 6914
rect 9632 6880 9644 6914
rect 9156 6874 9644 6880
rect 8862 6808 8874 6830
rect 7890 6254 7896 6804
rect 7850 6242 7896 6254
rect 8868 6254 8874 6808
rect 8908 6808 8922 6830
rect 9882 6830 9942 7072
rect 10900 7072 10910 7096
rect 10944 7624 10960 7648
rect 11920 7648 11980 7890
rect 12932 7890 12946 7914
rect 12980 8436 12992 8466
rect 13954 8466 14014 8708
rect 14974 8708 14982 8726
rect 15016 9256 15034 9284
rect 15990 9284 16050 9526
rect 17012 9526 17018 10102
rect 17052 10068 17072 10102
rect 17052 9546 17058 10068
rect 17052 9526 17072 9546
rect 16282 9476 16770 9482
rect 16282 9442 16294 9476
rect 16758 9442 16770 9476
rect 16282 9436 16770 9442
rect 16482 9374 16542 9436
rect 16282 9368 16770 9374
rect 16282 9334 16294 9368
rect 16758 9334 16770 9368
rect 16282 9328 16770 9334
rect 15990 9260 16000 9284
rect 15016 8726 15022 9256
rect 15994 8730 16000 9260
rect 15016 8708 15034 8726
rect 14246 8658 14734 8664
rect 14246 8624 14258 8658
rect 14722 8624 14734 8658
rect 14246 8618 14734 8624
rect 14452 8556 14512 8618
rect 14246 8550 14734 8556
rect 14246 8516 14258 8550
rect 14722 8516 14734 8550
rect 14246 8510 14734 8516
rect 13954 8436 13964 8466
rect 12980 7914 12986 8436
rect 13958 7914 13964 8436
rect 12980 7890 12992 7914
rect 12210 7840 12698 7846
rect 12210 7806 12222 7840
rect 12686 7806 12698 7840
rect 12210 7800 12698 7806
rect 12416 7738 12476 7800
rect 12210 7732 12698 7738
rect 12210 7698 12222 7732
rect 12686 7698 12698 7732
rect 12210 7692 12698 7698
rect 11920 7632 11928 7648
rect 10944 7096 10950 7624
rect 11922 7104 11928 7632
rect 10944 7072 10960 7096
rect 10174 7022 10662 7028
rect 10174 6988 10186 7022
rect 10650 6988 10662 7022
rect 10174 6982 10662 6988
rect 10386 6920 10446 6982
rect 10174 6914 10662 6920
rect 10174 6880 10186 6914
rect 10650 6880 10662 6914
rect 10174 6874 10662 6880
rect 9882 6810 9892 6830
rect 8908 6254 8914 6808
rect 9886 6300 9892 6810
rect 8868 6242 8914 6254
rect 9876 6254 9892 6300
rect 9926 6810 9942 6830
rect 10900 6830 10960 7072
rect 11920 7072 11928 7104
rect 11962 7632 11980 7648
rect 12932 7648 12992 7890
rect 13954 7890 13964 7914
rect 13998 8436 14014 8466
rect 14974 8466 15034 8708
rect 15990 8708 16000 8730
rect 16034 9260 16050 9284
rect 17012 9284 17072 9526
rect 16034 8730 16040 9260
rect 16034 8708 16050 8730
rect 15264 8658 15752 8664
rect 15264 8624 15276 8658
rect 15740 8624 15752 8658
rect 15264 8618 15752 8624
rect 15464 8556 15524 8618
rect 15264 8550 15752 8556
rect 15264 8516 15276 8550
rect 15740 8516 15752 8550
rect 15264 8510 15752 8516
rect 14974 8436 14982 8466
rect 13998 7914 14004 8436
rect 14976 7914 14982 8436
rect 13998 7890 14014 7914
rect 13228 7840 13716 7846
rect 13228 7806 13240 7840
rect 13704 7806 13716 7840
rect 13228 7800 13716 7806
rect 13432 7738 13492 7800
rect 13228 7732 13716 7738
rect 13228 7698 13240 7732
rect 13704 7698 13716 7732
rect 13228 7692 13716 7698
rect 11962 7104 11968 7632
rect 12932 7624 12946 7648
rect 11962 7072 11980 7104
rect 12940 7096 12946 7624
rect 11192 7022 11680 7028
rect 11192 6988 11204 7022
rect 11668 6988 11680 7022
rect 11192 6982 11680 6988
rect 11388 6920 11448 6982
rect 11192 6914 11680 6920
rect 11192 6880 11204 6914
rect 11668 6880 11680 6914
rect 11192 6874 11680 6880
rect 9926 6300 9932 6810
rect 10900 6806 10910 6830
rect 9926 6254 9936 6300
rect 8138 6204 8626 6210
rect 8138 6170 8150 6204
rect 8614 6170 8626 6204
rect 8138 6164 8626 6170
rect 9156 6204 9644 6210
rect 9156 6170 9168 6204
rect 9632 6170 9644 6204
rect 9156 6164 9644 6170
rect 9876 6080 9936 6254
rect 10904 6254 10910 6806
rect 10944 6806 10960 6830
rect 11920 6830 11980 7072
rect 12932 7072 12946 7096
rect 12980 7624 12992 7648
rect 13954 7648 14014 7890
rect 14974 7890 14982 7914
rect 15016 8436 15034 8466
rect 15990 8466 16050 8708
rect 17012 8708 17018 9284
rect 17052 9256 17072 9284
rect 17052 8726 17058 9256
rect 17052 8708 17072 8726
rect 16282 8658 16770 8664
rect 16282 8624 16294 8658
rect 16758 8624 16770 8658
rect 16282 8618 16770 8624
rect 16484 8556 16544 8618
rect 16282 8550 16770 8556
rect 16282 8516 16294 8550
rect 16758 8516 16770 8550
rect 16282 8510 16770 8516
rect 15990 8440 16000 8466
rect 15016 7914 15022 8436
rect 15994 7918 16000 8440
rect 15016 7890 15034 7914
rect 14246 7840 14734 7846
rect 14246 7806 14258 7840
rect 14722 7806 14734 7840
rect 14246 7800 14734 7806
rect 14454 7738 14514 7800
rect 14246 7732 14734 7738
rect 14246 7698 14258 7732
rect 14722 7698 14734 7732
rect 14246 7692 14734 7698
rect 13954 7624 13964 7648
rect 12980 7096 12986 7624
rect 13958 7096 13964 7624
rect 12980 7072 12992 7096
rect 12210 7022 12698 7028
rect 12210 6988 12222 7022
rect 12686 6988 12698 7022
rect 12210 6982 12698 6988
rect 12418 6920 12478 6982
rect 12210 6914 12698 6920
rect 12210 6880 12222 6914
rect 12686 6880 12698 6914
rect 12210 6874 12698 6880
rect 11920 6814 11928 6830
rect 10944 6254 10950 6806
rect 11922 6302 11928 6814
rect 10904 6242 10950 6254
rect 11914 6254 11928 6302
rect 11962 6814 11980 6830
rect 12932 6830 12992 7072
rect 13954 7072 13964 7096
rect 13998 7624 14014 7648
rect 14974 7648 15034 7890
rect 15990 7890 16000 7918
rect 16034 8440 16050 8466
rect 17012 8466 17072 8708
rect 16034 7918 16040 8440
rect 16034 7890 16050 7918
rect 15264 7840 15752 7846
rect 15264 7806 15276 7840
rect 15740 7806 15752 7840
rect 15264 7800 15752 7806
rect 15466 7738 15526 7800
rect 15264 7732 15752 7738
rect 15264 7698 15276 7732
rect 15740 7698 15752 7732
rect 15264 7692 15752 7698
rect 14974 7624 14982 7648
rect 13998 7096 14004 7624
rect 14976 7096 14982 7624
rect 13998 7072 14014 7096
rect 13228 7022 13716 7028
rect 13228 6988 13240 7022
rect 13704 6988 13716 7022
rect 13228 6982 13716 6988
rect 13434 6920 13494 6982
rect 13228 6914 13716 6920
rect 13228 6880 13240 6914
rect 13704 6880 13716 6914
rect 13228 6874 13716 6880
rect 11962 6302 11968 6814
rect 12932 6806 12946 6830
rect 11962 6254 11974 6302
rect 10174 6204 10662 6210
rect 10174 6170 10186 6204
rect 10650 6170 10662 6204
rect 10174 6164 10662 6170
rect 11192 6204 11680 6210
rect 11192 6170 11204 6204
rect 11668 6170 11680 6204
rect 11192 6164 11680 6170
rect 11914 6080 11974 6254
rect 12940 6254 12946 6806
rect 12980 6806 12992 6830
rect 13954 6830 14014 7072
rect 14974 7072 14982 7096
rect 15016 7624 15034 7648
rect 15990 7648 16050 7890
rect 17012 7890 17018 8466
rect 17052 8436 17072 8466
rect 17052 7914 17058 8436
rect 17052 7890 17072 7914
rect 16282 7840 16770 7846
rect 16282 7806 16294 7840
rect 16758 7806 16770 7840
rect 16282 7800 16770 7806
rect 16486 7738 16546 7800
rect 16282 7732 16770 7738
rect 16282 7698 16294 7732
rect 16758 7698 16770 7732
rect 16282 7692 16770 7698
rect 15990 7628 16000 7648
rect 15016 7096 15022 7624
rect 15994 7100 16000 7628
rect 15016 7072 15034 7096
rect 14246 7022 14734 7028
rect 14246 6988 14258 7022
rect 14722 6988 14734 7022
rect 14246 6982 14734 6988
rect 14456 6920 14516 6982
rect 14246 6914 14734 6920
rect 14246 6880 14258 6914
rect 14722 6880 14734 6914
rect 14246 6874 14734 6880
rect 13954 6806 13964 6830
rect 12980 6254 12986 6806
rect 13958 6298 13964 6806
rect 12940 6242 12986 6254
rect 13950 6254 13964 6298
rect 13998 6806 14014 6830
rect 14974 6830 15034 7072
rect 15990 7072 16000 7100
rect 16034 7628 16050 7648
rect 17012 7648 17072 7890
rect 16034 7100 16040 7628
rect 16034 7072 16050 7100
rect 15264 7022 15752 7028
rect 15264 6988 15276 7022
rect 15740 6988 15752 7022
rect 15264 6982 15752 6988
rect 15468 6920 15528 6982
rect 15264 6914 15752 6920
rect 15264 6880 15276 6914
rect 15740 6880 15752 6914
rect 15264 6874 15752 6880
rect 14974 6806 14982 6830
rect 13998 6298 14004 6806
rect 13998 6254 14010 6298
rect 12210 6204 12698 6210
rect 12210 6170 12222 6204
rect 12686 6170 12698 6204
rect 12210 6164 12698 6170
rect 13228 6204 13716 6210
rect 13228 6170 13240 6204
rect 13704 6170 13716 6204
rect 13228 6164 13716 6170
rect 13950 6080 14010 6254
rect 14976 6254 14982 6806
rect 15016 6806 15034 6830
rect 15990 6830 16050 7072
rect 17012 7072 17018 7648
rect 17052 7624 17072 7648
rect 17052 7096 17058 7624
rect 17052 7072 17072 7096
rect 16282 7022 16770 7028
rect 16282 6988 16294 7022
rect 16758 6988 16770 7022
rect 16282 6982 16770 6988
rect 16488 6920 16548 6982
rect 16282 6914 16770 6920
rect 16282 6880 16294 6914
rect 16758 6880 16770 6914
rect 16282 6874 16770 6880
rect 15990 6810 16000 6830
rect 15016 6254 15022 6806
rect 15994 6296 16000 6810
rect 14976 6242 15022 6254
rect 15986 6254 16000 6296
rect 16034 6810 16050 6830
rect 17012 6830 17072 7072
rect 16034 6296 16040 6810
rect 17012 6308 17018 6830
rect 16034 6254 16046 6296
rect 14246 6204 14734 6210
rect 14246 6170 14258 6204
rect 14722 6170 14734 6204
rect 14246 6164 14734 6170
rect 15264 6204 15752 6210
rect 15264 6170 15276 6204
rect 15740 6170 15752 6204
rect 15264 6164 15752 6170
rect 15986 6080 16046 6254
rect 17006 6254 17018 6308
rect 17052 6806 17072 6830
rect 17052 6308 17058 6806
rect 17052 6254 17066 6308
rect 18190 6258 18250 13398
rect 16282 6204 16770 6210
rect 16282 6170 16294 6204
rect 16758 6170 16770 6204
rect 16282 6164 16770 6170
rect 16500 6080 16560 6164
rect 17006 6080 17066 6254
rect 18184 6198 18190 6258
rect 18250 6198 18256 6258
rect 9876 6020 18170 6080
rect 13636 5272 13642 5332
rect 13702 5272 13708 5332
rect 7532 5186 7592 5192
rect 11606 5126 11612 5186
rect 11672 5126 11678 5186
rect 6372 4998 6378 5058
rect 6438 4998 6444 5058
rect 6378 2826 6438 4998
rect 7532 4994 7592 5126
rect 9050 4998 9056 5058
rect 9116 4998 9122 5058
rect 10082 4998 10088 5058
rect 10148 4998 10154 5058
rect 6516 4934 7592 4994
rect 6516 4806 6576 4934
rect 7024 4896 7084 4934
rect 6814 4890 7302 4896
rect 6814 4856 6826 4890
rect 7290 4856 7302 4890
rect 6814 4850 7302 4856
rect 6516 4760 6532 4806
rect 6526 4230 6532 4760
rect 6566 4760 6576 4806
rect 7532 4806 7592 4934
rect 9056 4896 9116 4998
rect 10088 4896 10148 4998
rect 7832 4890 8320 4896
rect 7832 4856 7844 4890
rect 8308 4856 8320 4890
rect 7832 4850 8320 4856
rect 8850 4890 9338 4896
rect 8850 4856 8862 4890
rect 9326 4856 9338 4890
rect 8850 4850 9338 4856
rect 9868 4890 10356 4896
rect 9868 4856 9880 4890
rect 10344 4856 10356 4890
rect 9868 4850 10356 4856
rect 10886 4890 11374 4896
rect 10886 4856 10898 4890
rect 11362 4856 11374 4890
rect 10886 4850 11374 4856
rect 7532 4766 7550 4806
rect 6566 4230 6572 4760
rect 6526 4218 6572 4230
rect 7544 4230 7550 4766
rect 7584 4766 7592 4806
rect 8562 4806 8608 4818
rect 7584 4230 7590 4766
rect 8562 4294 8568 4806
rect 7544 4218 7590 4230
rect 8554 4230 8568 4294
rect 8602 4294 8608 4806
rect 9580 4806 9626 4818
rect 8602 4230 8614 4294
rect 9580 4276 9586 4806
rect 6814 4180 7302 4186
rect 6814 4146 6826 4180
rect 7290 4146 7302 4180
rect 6814 4140 7302 4146
rect 7832 4180 8320 4186
rect 7832 4146 7844 4180
rect 8308 4146 8320 4180
rect 7832 4140 8320 4146
rect 8036 4096 8096 4140
rect 8030 4036 8036 4096
rect 8096 4036 8102 4096
rect 7530 3932 7536 3992
rect 7596 3932 7602 3992
rect 7536 3890 7596 3932
rect 6516 3830 7596 3890
rect 6516 3694 6576 3830
rect 7020 3784 7080 3830
rect 6814 3778 7302 3784
rect 6814 3744 6826 3778
rect 7290 3744 7302 3778
rect 6814 3738 7302 3744
rect 6516 3648 6532 3694
rect 6526 3118 6532 3648
rect 6566 3648 6576 3694
rect 7536 3694 7596 3830
rect 8554 3888 8614 4230
rect 9572 4230 9586 4276
rect 9620 4276 9626 4806
rect 10598 4806 10644 4818
rect 10598 4292 10604 4806
rect 9620 4230 9632 4276
rect 8850 4180 9338 4186
rect 8850 4146 8862 4180
rect 9326 4146 9338 4180
rect 8850 4140 9338 4146
rect 9054 4036 9060 4096
rect 9120 4036 9126 4096
rect 7832 3778 8320 3784
rect 7832 3744 7844 3778
rect 8308 3744 8320 3778
rect 7832 3738 8320 3744
rect 6566 3118 6572 3648
rect 6526 3106 6572 3118
rect 7536 3118 7550 3694
rect 7584 3118 7596 3694
rect 6814 3068 7302 3074
rect 6814 3034 6826 3068
rect 7290 3034 7302 3068
rect 6814 3028 7302 3034
rect 6372 2766 6378 2826
rect 6438 2766 6444 2826
rect 4662 1148 4718 1198
rect 4712 1022 4718 1148
rect -210 986 4718 1022
rect 4818 1148 5100 1198
rect 4818 1022 4824 1148
rect 4818 986 4968 1022
rect -210 896 -156 986
rect 4924 896 4968 986
rect -210 842 -102 896
rect 4302 842 4718 896
rect -210 838 4718 842
rect -208 836 4408 838
rect -208 673 -96 836
rect -8 688 -2 748
rect 58 688 64 748
rect -208 -1773 -202 673
rect -102 -1773 -96 673
rect -2 -1218 58 688
rect 136 564 142 624
rect 202 564 208 624
rect 272 620 332 836
rect 404 620 464 836
rect 784 688 790 748
rect 850 688 856 748
rect 142 -1092 202 564
rect 272 560 464 620
rect 272 430 332 560
rect 404 520 464 560
rect 378 514 486 520
rect 378 480 390 514
rect 474 480 486 514
rect 378 474 486 480
rect 636 514 744 520
rect 636 480 648 514
rect 732 480 744 514
rect 636 474 744 480
rect 272 54 286 430
rect 320 54 332 430
rect 538 430 584 442
rect 538 80 544 430
rect 272 -244 332 54
rect 532 54 544 80
rect 578 80 584 430
rect 790 430 850 688
rect 1172 624 1232 836
rect 1304 624 1364 836
rect 1432 624 1492 836
rect 1172 564 1492 624
rect 1812 564 1818 624
rect 1878 564 1884 624
rect 2332 564 2338 624
rect 2398 564 2404 624
rect 2724 622 2784 836
rect 2856 622 2916 836
rect 2984 622 3044 836
rect 3360 688 3366 748
rect 3426 688 3432 748
rect 1172 520 1232 564
rect 1304 562 1492 564
rect 894 514 1002 520
rect 894 480 906 514
rect 990 480 1002 514
rect 894 474 1002 480
rect 1152 514 1260 520
rect 1152 480 1164 514
rect 1248 480 1260 514
rect 1152 474 1260 480
rect 790 382 802 430
rect 578 54 592 80
rect 378 4 486 10
rect 378 -30 390 4
rect 474 -30 486 4
rect 378 -36 486 -30
rect 404 -244 464 -36
rect 272 -304 464 -244
rect 272 -570 332 -304
rect 404 -480 464 -304
rect 532 -358 592 54
rect 796 54 802 382
rect 836 382 850 430
rect 1054 430 1100 442
rect 836 54 842 382
rect 1054 102 1060 430
rect 796 42 842 54
rect 1050 54 1060 102
rect 1094 102 1100 430
rect 1304 430 1364 562
rect 1432 520 1492 562
rect 1410 514 1518 520
rect 1410 480 1422 514
rect 1506 480 1518 514
rect 1410 474 1518 480
rect 1668 514 1776 520
rect 1668 480 1680 514
rect 1764 480 1776 514
rect 1668 474 1776 480
rect 1094 54 1110 102
rect 636 4 744 10
rect 636 -30 648 4
rect 732 -30 744 4
rect 636 -36 744 -30
rect 894 4 1002 10
rect 894 -30 906 4
rect 990 -30 1002 4
rect 894 -36 1002 -30
rect 662 -110 722 -36
rect 920 -108 980 -36
rect 656 -170 662 -110
rect 722 -170 728 -110
rect 914 -168 920 -108
rect 980 -168 986 -108
rect 526 -418 532 -358
rect 592 -418 598 -358
rect 662 -480 722 -170
rect 784 -300 790 -240
rect 850 -300 856 -240
rect 378 -486 486 -480
rect 378 -520 390 -486
rect 474 -520 486 -486
rect 378 -526 486 -520
rect 636 -486 744 -480
rect 636 -520 648 -486
rect 732 -520 744 -486
rect 636 -526 744 -520
rect 272 -946 286 -570
rect 320 -946 332 -570
rect 538 -570 584 -558
rect 538 -902 544 -570
rect 272 -1090 332 -946
rect 532 -946 544 -902
rect 578 -902 584 -570
rect 790 -570 850 -300
rect 920 -480 980 -168
rect 1050 -358 1110 54
rect 1304 54 1318 430
rect 1352 54 1364 430
rect 1570 430 1616 442
rect 1570 104 1576 430
rect 1152 4 1260 10
rect 1152 -30 1164 4
rect 1248 -30 1260 4
rect 1152 -36 1260 -30
rect 1172 -242 1232 -36
rect 1304 -242 1364 54
rect 1564 54 1576 104
rect 1610 104 1616 430
rect 1818 430 1878 564
rect 1926 514 2034 520
rect 1926 480 1938 514
rect 2022 480 2034 514
rect 1926 474 2034 480
rect 2184 514 2292 520
rect 2184 480 2196 514
rect 2280 480 2292 514
rect 2184 474 2292 480
rect 1818 386 1834 430
rect 1610 54 1624 104
rect 1410 4 1518 10
rect 1410 -30 1422 4
rect 1506 -30 1518 4
rect 1410 -36 1518 -30
rect 1172 -244 1364 -242
rect 1434 -244 1494 -36
rect 1564 -240 1624 54
rect 1828 54 1834 386
rect 1868 386 1878 430
rect 2086 430 2132 442
rect 1868 54 1874 386
rect 2086 110 2092 430
rect 1828 42 1874 54
rect 2080 54 2092 110
rect 2126 110 2132 430
rect 2338 430 2398 564
rect 2724 562 3044 622
rect 2724 520 2784 562
rect 2856 560 3044 562
rect 2442 514 2550 520
rect 2442 480 2454 514
rect 2538 480 2550 514
rect 2442 474 2550 480
rect 2700 514 2808 520
rect 2700 480 2712 514
rect 2796 480 2808 514
rect 2700 474 2808 480
rect 2338 390 2350 430
rect 2126 54 2140 110
rect 1668 4 1776 10
rect 1668 -30 1680 4
rect 1764 -30 1776 4
rect 1668 -36 1776 -30
rect 1926 4 2034 10
rect 1926 -30 1938 4
rect 2022 -30 2034 4
rect 1926 -36 2034 -30
rect 1692 -110 1752 -36
rect 1952 -110 2012 -36
rect 1686 -170 1692 -110
rect 1752 -170 1758 -110
rect 1946 -170 1952 -110
rect 2012 -170 2018 -110
rect 1172 -302 1494 -244
rect 1558 -300 1564 -240
rect 1624 -300 1630 -240
rect 1044 -418 1050 -358
rect 1110 -418 1116 -358
rect 1172 -480 1232 -302
rect 1304 -304 1494 -302
rect 894 -486 1002 -480
rect 894 -520 906 -486
rect 990 -520 1002 -486
rect 894 -526 1002 -520
rect 1152 -486 1260 -480
rect 1152 -520 1164 -486
rect 1248 -520 1260 -486
rect 1152 -526 1260 -520
rect 790 -620 802 -570
rect 578 -946 592 -902
rect 378 -996 486 -990
rect 378 -1030 390 -996
rect 474 -1030 486 -996
rect 378 -1036 486 -1030
rect 398 -1090 458 -1036
rect 136 -1152 142 -1092
rect 202 -1152 208 -1092
rect 272 -1150 458 -1090
rect 532 -1092 592 -946
rect 796 -946 802 -620
rect 836 -620 850 -570
rect 1054 -570 1100 -558
rect 836 -946 842 -620
rect 1054 -910 1060 -570
rect 796 -958 842 -946
rect 1048 -946 1060 -910
rect 1094 -910 1100 -570
rect 1304 -570 1364 -304
rect 1434 -480 1494 -304
rect 1692 -480 1752 -170
rect 1816 -418 1822 -358
rect 1882 -418 1888 -358
rect 1410 -486 1518 -480
rect 1410 -520 1422 -486
rect 1506 -520 1518 -486
rect 1410 -526 1518 -520
rect 1668 -486 1776 -480
rect 1668 -520 1680 -486
rect 1764 -520 1776 -486
rect 1668 -526 1776 -520
rect 1094 -946 1108 -910
rect 636 -996 744 -990
rect 636 -1030 648 -996
rect 732 -1030 744 -996
rect 636 -1036 744 -1030
rect 894 -996 1002 -990
rect 894 -1030 906 -996
rect 990 -1030 1002 -996
rect 894 -1036 1002 -1030
rect 1048 -1092 1108 -946
rect 1304 -946 1318 -570
rect 1352 -946 1364 -570
rect 1570 -570 1616 -558
rect 1570 -888 1576 -570
rect 1152 -996 1260 -990
rect 1152 -1030 1164 -996
rect 1248 -1030 1260 -996
rect 1152 -1036 1260 -1030
rect 1170 -1092 1230 -1036
rect 1304 -1092 1364 -946
rect 1560 -946 1576 -888
rect 1610 -888 1616 -570
rect 1822 -570 1882 -418
rect 1952 -480 2012 -170
rect 2080 -240 2140 54
rect 2344 54 2350 390
rect 2384 390 2398 430
rect 2602 430 2648 442
rect 2384 54 2390 390
rect 2602 120 2608 430
rect 2344 42 2390 54
rect 2598 54 2608 120
rect 2642 120 2648 430
rect 2856 430 2916 560
rect 2984 520 3044 560
rect 2958 514 3066 520
rect 2958 480 2970 514
rect 3054 480 3066 514
rect 2958 474 3066 480
rect 3216 514 3324 520
rect 3216 480 3228 514
rect 3312 480 3324 514
rect 3216 474 3324 480
rect 2642 54 2658 120
rect 2184 4 2292 10
rect 2184 -30 2196 4
rect 2280 -30 2292 4
rect 2184 -36 2292 -30
rect 2442 4 2550 10
rect 2442 -30 2454 4
rect 2538 -30 2550 4
rect 2442 -36 2550 -30
rect 2208 -110 2268 -36
rect 2466 -110 2526 -36
rect 2202 -170 2208 -110
rect 2268 -170 2274 -110
rect 2460 -170 2466 -110
rect 2526 -170 2532 -110
rect 2074 -300 2080 -240
rect 2140 -300 2146 -240
rect 2208 -480 2268 -170
rect 2330 -418 2336 -358
rect 2396 -418 2402 -358
rect 1926 -486 2034 -480
rect 1926 -520 1938 -486
rect 2022 -520 2034 -486
rect 1926 -526 2034 -520
rect 2184 -486 2292 -480
rect 2184 -520 2196 -486
rect 2280 -520 2292 -486
rect 2184 -526 2292 -520
rect 1822 -616 1834 -570
rect 1610 -946 1620 -888
rect 1410 -996 1518 -990
rect 1410 -1030 1422 -996
rect 1506 -1030 1518 -996
rect 1410 -1036 1518 -1030
rect 1432 -1092 1492 -1036
rect -8 -1278 -2 -1218
rect 58 -1278 64 -1218
rect 272 -1352 332 -1150
rect 398 -1352 458 -1150
rect 526 -1152 532 -1092
rect 592 -1152 598 -1092
rect 1042 -1152 1048 -1092
rect 1108 -1152 1114 -1092
rect 1170 -1152 1492 -1092
rect 1170 -1352 1230 -1152
rect 1304 -1352 1364 -1152
rect 1432 -1352 1492 -1152
rect 1560 -1218 1620 -946
rect 1828 -946 1834 -616
rect 1868 -616 1882 -570
rect 2086 -570 2132 -558
rect 1868 -946 1874 -616
rect 2086 -894 2092 -570
rect 1828 -958 1874 -946
rect 2082 -946 2092 -894
rect 2126 -894 2132 -570
rect 2336 -570 2396 -418
rect 2466 -480 2526 -170
rect 2598 -240 2658 54
rect 2856 54 2866 430
rect 2900 54 2916 430
rect 3118 430 3164 442
rect 3118 126 3124 430
rect 2700 4 2808 10
rect 2700 -30 2712 4
rect 2796 -30 2808 4
rect 2700 -36 2808 -30
rect 2592 -300 2598 -240
rect 2658 -300 2664 -240
rect 2724 -244 2784 -36
rect 2856 -244 2916 54
rect 3112 54 3124 126
rect 3158 126 3164 430
rect 3366 430 3426 688
rect 3758 624 3818 836
rect 3882 624 3942 836
rect 4128 688 4134 748
rect 4194 688 4200 748
rect 3758 564 3942 624
rect 3992 564 3998 624
rect 4058 564 4064 624
rect 3758 520 3818 564
rect 3474 514 3582 520
rect 3474 480 3486 514
rect 3570 480 3582 514
rect 3474 474 3582 480
rect 3732 514 3840 520
rect 3732 480 3744 514
rect 3828 480 3840 514
rect 3732 474 3840 480
rect 3366 370 3382 430
rect 3158 54 3172 126
rect 2958 4 3066 10
rect 2958 -30 2970 4
rect 3054 -30 3066 4
rect 2958 -36 3066 -30
rect 2724 -246 2916 -244
rect 2986 -246 3046 -36
rect 2724 -304 3046 -246
rect 2724 -480 2784 -304
rect 2856 -306 3046 -304
rect 2442 -486 2550 -480
rect 2442 -520 2454 -486
rect 2538 -520 2550 -486
rect 2442 -526 2550 -520
rect 2700 -486 2808 -480
rect 2700 -520 2712 -486
rect 2796 -520 2808 -486
rect 2700 -526 2808 -520
rect 2336 -616 2350 -570
rect 2126 -946 2142 -894
rect 1668 -996 1776 -990
rect 1668 -1030 1680 -996
rect 1764 -1030 1776 -996
rect 1668 -1036 1776 -1030
rect 1926 -996 2034 -990
rect 1926 -1030 1938 -996
rect 2022 -1030 2034 -996
rect 1926 -1036 2034 -1030
rect 2082 -1218 2142 -946
rect 2344 -946 2350 -616
rect 2384 -616 2396 -570
rect 2602 -570 2648 -558
rect 2384 -946 2390 -616
rect 2602 -890 2608 -570
rect 2344 -958 2390 -946
rect 2596 -946 2608 -890
rect 2642 -890 2648 -570
rect 2856 -570 2916 -306
rect 2986 -480 3046 -306
rect 3112 -358 3172 54
rect 3376 54 3382 370
rect 3416 370 3426 430
rect 3634 430 3680 442
rect 3416 54 3422 370
rect 3634 102 3640 430
rect 3376 42 3422 54
rect 3626 54 3640 102
rect 3674 102 3680 430
rect 3882 430 3942 564
rect 3674 54 3686 102
rect 3216 4 3324 10
rect 3216 -30 3228 4
rect 3312 -30 3324 4
rect 3216 -36 3324 -30
rect 3474 4 3582 10
rect 3474 -30 3486 4
rect 3570 -30 3582 4
rect 3474 -36 3582 -30
rect 3242 -110 3302 -36
rect 3502 -110 3562 -36
rect 3236 -170 3242 -110
rect 3302 -170 3308 -110
rect 3496 -170 3502 -110
rect 3562 -170 3568 -110
rect 3106 -418 3112 -358
rect 3172 -418 3178 -358
rect 3242 -480 3302 -170
rect 3362 -300 3368 -240
rect 3428 -300 3434 -240
rect 2958 -486 3066 -480
rect 2958 -520 2970 -486
rect 3054 -520 3066 -486
rect 2958 -526 3066 -520
rect 3216 -486 3324 -480
rect 3216 -520 3228 -486
rect 3312 -520 3324 -486
rect 3216 -526 3324 -520
rect 2642 -946 2656 -890
rect 2184 -996 2292 -990
rect 2184 -1030 2196 -996
rect 2280 -1030 2292 -996
rect 2184 -1036 2292 -1030
rect 2442 -996 2550 -990
rect 2442 -1030 2454 -996
rect 2538 -1030 2550 -996
rect 2442 -1036 2550 -1030
rect 2596 -1218 2656 -946
rect 2856 -946 2866 -570
rect 2900 -946 2916 -570
rect 3118 -570 3164 -558
rect 3118 -902 3124 -570
rect 2700 -996 2808 -990
rect 2700 -1030 2712 -996
rect 2796 -1030 2808 -996
rect 2700 -1036 2808 -1030
rect 2722 -1094 2782 -1036
rect 2856 -1094 2916 -946
rect 3112 -946 3124 -902
rect 3158 -902 3164 -570
rect 3368 -570 3428 -300
rect 3502 -480 3562 -170
rect 3626 -358 3686 54
rect 3882 54 3898 430
rect 3932 54 3942 430
rect 3732 4 3840 10
rect 3732 -30 3744 4
rect 3828 -30 3840 4
rect 3732 -36 3840 -30
rect 3754 -240 3814 -36
rect 3882 -240 3942 54
rect 3754 -300 3942 -240
rect 3620 -418 3626 -358
rect 3686 -418 3692 -358
rect 3754 -480 3814 -300
rect 3474 -486 3582 -480
rect 3474 -520 3486 -486
rect 3570 -520 3582 -486
rect 3474 -526 3582 -520
rect 3732 -486 3840 -480
rect 3732 -520 3744 -486
rect 3828 -520 3840 -486
rect 3732 -526 3840 -520
rect 3368 -632 3382 -570
rect 3158 -946 3172 -902
rect 2958 -996 3066 -990
rect 2958 -1030 2970 -996
rect 3054 -1030 3066 -996
rect 2958 -1036 3066 -1030
rect 2984 -1094 3044 -1036
rect 3112 -1092 3172 -946
rect 3376 -946 3382 -632
rect 3416 -632 3428 -570
rect 3634 -570 3680 -558
rect 3416 -946 3422 -632
rect 3634 -906 3640 -570
rect 3376 -958 3422 -946
rect 3626 -946 3640 -906
rect 3674 -906 3680 -570
rect 3882 -570 3942 -300
rect 3674 -946 3686 -906
rect 3216 -996 3324 -990
rect 3216 -1030 3228 -996
rect 3312 -1030 3324 -996
rect 3216 -1036 3324 -1030
rect 3474 -996 3582 -990
rect 3474 -1030 3486 -996
rect 3570 -1030 3582 -996
rect 3474 -1036 3582 -1030
rect 3626 -1092 3686 -946
rect 3882 -946 3898 -570
rect 3932 -946 3942 -570
rect 3732 -996 3840 -990
rect 3732 -1030 3744 -996
rect 3828 -1030 3840 -996
rect 3732 -1036 3840 -1030
rect 3752 -1092 3812 -1036
rect 3882 -1092 3942 -946
rect 3998 -1092 4058 564
rect 2722 -1154 3044 -1094
rect 3106 -1152 3112 -1092
rect 3172 -1152 3178 -1092
rect 3620 -1152 3626 -1092
rect 3686 -1152 3692 -1092
rect 3752 -1152 3942 -1092
rect 3992 -1152 3998 -1092
rect 4058 -1152 4064 -1092
rect 1554 -1278 1560 -1218
rect 1620 -1278 1626 -1218
rect 2076 -1278 2082 -1218
rect 2142 -1278 2148 -1218
rect 2590 -1278 2596 -1218
rect 2656 -1278 2662 -1218
rect 2722 -1352 2782 -1154
rect 2856 -1352 2916 -1154
rect 2984 -1352 3044 -1154
rect 3752 -1352 3812 -1152
rect 3882 -1352 3942 -1152
rect 4134 -1218 4194 688
rect 4296 673 4408 836
rect 4128 -1278 4134 -1218
rect 4194 -1278 4200 -1218
rect 204 -1402 3996 -1352
rect 204 -1506 258 -1402
rect 3950 -1506 3996 -1402
rect 204 -1550 3996 -1506
rect -208 -1936 -96 -1773
rect 504 -1936 514 -1636
rect 3686 -1936 3696 -1636
rect 4296 -1773 4302 673
rect 4402 -1773 4408 673
rect 4296 -1936 4408 -1773
rect -208 -1942 4408 -1936
rect -208 -2042 -102 -1942
rect 4302 -2042 4408 -1942
rect -208 -2048 4408 -2042
rect 4712 -1250 4718 838
rect 4818 838 4968 896
rect 4818 -1250 4824 838
rect 6378 700 6438 2766
rect 6814 2666 7302 2672
rect 6814 2632 6826 2666
rect 7290 2632 7302 2666
rect 6814 2626 7302 2632
rect 6526 2582 6572 2594
rect 6526 2040 6532 2582
rect 6520 2006 6532 2040
rect 6566 2040 6572 2582
rect 7536 2582 7596 3118
rect 8554 3694 8614 3828
rect 9060 3784 9120 4036
rect 9572 3992 9632 4230
rect 10590 4230 10604 4292
rect 10638 4292 10644 4806
rect 11612 4806 11672 5126
rect 13142 4998 13148 5058
rect 13208 4998 13214 5058
rect 13148 4896 13208 4998
rect 11904 4890 12392 4896
rect 11904 4856 11916 4890
rect 12380 4856 12392 4890
rect 11904 4850 12392 4856
rect 12922 4890 13410 4896
rect 12922 4856 12934 4890
rect 13398 4856 13410 4890
rect 12922 4850 13410 4856
rect 11612 4742 11622 4806
rect 10638 4230 10650 4292
rect 9868 4180 10356 4186
rect 9868 4146 9880 4180
rect 10344 4146 10356 4180
rect 9868 4140 10356 4146
rect 10086 4036 10092 4096
rect 10152 4036 10158 4096
rect 9566 3932 9572 3992
rect 9632 3932 9638 3992
rect 10092 3784 10152 4036
rect 10590 3888 10650 4230
rect 11616 4230 11622 4742
rect 11656 4742 11672 4806
rect 12634 4806 12680 4818
rect 11656 4230 11662 4742
rect 12634 4302 12640 4806
rect 11616 4218 11662 4230
rect 12622 4230 12640 4302
rect 12674 4302 12680 4806
rect 13642 4806 13702 5272
rect 15666 5126 15672 5186
rect 15732 5126 15738 5186
rect 17850 5126 17856 5186
rect 17916 5126 17922 5186
rect 14138 4998 14144 5058
rect 14204 4998 14210 5058
rect 14144 4896 14204 4998
rect 13940 4890 14428 4896
rect 13940 4856 13952 4890
rect 14416 4856 14428 4890
rect 13940 4850 14428 4856
rect 14958 4890 15446 4896
rect 14958 4856 14970 4890
rect 15434 4856 15446 4890
rect 14958 4850 15446 4856
rect 14144 4848 14204 4850
rect 15672 4818 15732 5126
rect 15976 4890 16464 4896
rect 15976 4856 15988 4890
rect 16452 4856 16464 4890
rect 15976 4850 16464 4856
rect 16994 4890 17482 4896
rect 16994 4856 17006 4890
rect 17470 4856 17482 4890
rect 16994 4850 17482 4856
rect 12674 4230 12682 4302
rect 10886 4180 11374 4186
rect 10886 4146 10898 4180
rect 11362 4146 11374 4180
rect 10886 4140 11374 4146
rect 11904 4180 12392 4186
rect 11904 4146 11916 4180
rect 12380 4146 12392 4180
rect 11904 4140 12392 4146
rect 11092 4096 11152 4140
rect 12112 4096 12172 4140
rect 11086 4036 11092 4096
rect 11152 4036 11158 4096
rect 12106 4036 12112 4096
rect 12172 4036 12178 4096
rect 11602 3932 11608 3992
rect 11668 3932 11674 3992
rect 8850 3778 9338 3784
rect 8850 3744 8862 3778
rect 9326 3744 9338 3778
rect 8850 3738 9338 3744
rect 9868 3778 10356 3784
rect 9868 3744 9880 3778
rect 10344 3744 10356 3778
rect 9868 3738 10356 3744
rect 8554 3118 8568 3694
rect 8602 3118 8614 3694
rect 9580 3694 9626 3706
rect 9580 3156 9586 3694
rect 7832 3068 8320 3074
rect 7832 3034 7844 3068
rect 8308 3034 8320 3068
rect 7832 3028 8320 3034
rect 8028 2826 8088 3028
rect 8022 2766 8028 2826
rect 8088 2766 8094 2826
rect 8028 2672 8088 2766
rect 7832 2666 8320 2672
rect 7832 2632 7844 2666
rect 8308 2632 8320 2666
rect 7832 2626 8320 2632
rect 7536 2510 7550 2582
rect 6566 2006 6580 2040
rect 7544 2036 7550 2510
rect 6520 1874 6580 2006
rect 7540 2006 7550 2036
rect 7584 2510 7596 2582
rect 8554 2582 8614 3118
rect 9566 3118 9586 3156
rect 9620 3118 9626 3694
rect 8850 3068 9338 3074
rect 8850 3034 8862 3068
rect 9326 3034 9338 3068
rect 8850 3028 9338 3034
rect 9566 2946 9626 3118
rect 10590 3694 10650 3828
rect 10886 3778 11374 3784
rect 10886 3744 10898 3778
rect 11362 3744 11374 3778
rect 10886 3738 11374 3744
rect 10590 3118 10604 3694
rect 10638 3118 10650 3694
rect 9868 3068 10356 3074
rect 9868 3034 9880 3068
rect 10344 3034 10356 3068
rect 9868 3028 10356 3034
rect 9560 2886 9566 2946
rect 9626 2886 9632 2946
rect 8850 2666 9338 2672
rect 8850 2632 8862 2666
rect 9326 2632 9338 2666
rect 8850 2626 9338 2632
rect 7584 2036 7590 2510
rect 7584 2006 7600 2036
rect 6814 1956 7302 1962
rect 6814 1922 6826 1956
rect 7290 1922 7302 1956
rect 6814 1916 7302 1922
rect 7012 1874 7072 1916
rect 7540 1874 7600 2006
rect 8554 2006 8568 2582
rect 8602 2006 8614 2582
rect 9566 2582 9626 2886
rect 9868 2666 10356 2672
rect 9868 2632 9880 2666
rect 10344 2632 10356 2666
rect 9868 2626 10356 2632
rect 9566 2512 9586 2582
rect 7832 1956 8320 1962
rect 7832 1922 7844 1956
rect 8308 1922 8320 1956
rect 7832 1916 8320 1922
rect 6520 1814 7600 1874
rect 7540 1774 7600 1814
rect 8554 1882 8614 2006
rect 9580 2006 9586 2512
rect 9620 2006 9626 2582
rect 9580 1994 9626 2006
rect 10590 2582 10650 3118
rect 11608 3694 11668 3932
rect 12622 3888 12682 4230
rect 13642 4230 13658 4806
rect 13692 4230 13702 4806
rect 14670 4806 14716 4818
rect 14670 4292 14676 4806
rect 12922 4180 13410 4186
rect 12922 4146 12934 4180
rect 13398 4146 13410 4180
rect 12922 4140 13410 4146
rect 13126 4036 13132 4096
rect 13192 4036 13198 4096
rect 12616 3828 12622 3888
rect 12682 3828 12688 3888
rect 11904 3778 12392 3784
rect 11904 3744 11916 3778
rect 12380 3744 12392 3778
rect 11904 3738 12392 3744
rect 11608 3118 11622 3694
rect 11656 3118 11668 3694
rect 10886 3068 11374 3074
rect 10886 3034 10898 3068
rect 11362 3034 11374 3068
rect 10886 3028 11374 3034
rect 11098 2826 11158 3028
rect 11092 2766 11098 2826
rect 11158 2766 11164 2826
rect 11098 2672 11158 2766
rect 10886 2666 11374 2672
rect 10886 2632 10898 2666
rect 11362 2632 11374 2666
rect 10886 2626 11374 2632
rect 10590 2006 10604 2582
rect 10638 2006 10650 2582
rect 11608 2582 11668 3118
rect 12622 3694 12682 3828
rect 13132 3784 13192 4036
rect 13642 3992 13702 4230
rect 14656 4230 14676 4292
rect 14710 4230 14716 4806
rect 15672 4806 15734 4818
rect 15672 4774 15694 4806
rect 13940 4180 14428 4186
rect 13940 4146 13952 4180
rect 14416 4146 14428 4180
rect 13940 4140 14428 4146
rect 14142 4096 14202 4102
rect 13636 3932 13642 3992
rect 13702 3932 13708 3992
rect 14142 3784 14202 4036
rect 14656 3888 14716 4230
rect 15688 4230 15694 4774
rect 15728 4230 15734 4806
rect 16706 4806 16752 4818
rect 16706 4264 16712 4806
rect 15688 4218 15734 4230
rect 16700 4230 16712 4264
rect 16746 4264 16752 4806
rect 17724 4806 17770 4818
rect 17724 4284 17730 4806
rect 16746 4230 16760 4264
rect 14958 4180 15446 4186
rect 14958 4146 14970 4180
rect 15434 4146 15446 4180
rect 14958 4140 15446 4146
rect 15976 4180 16464 4186
rect 15976 4146 15988 4180
rect 16452 4146 16464 4180
rect 15976 4140 16464 4146
rect 15156 4096 15216 4140
rect 16174 4096 16234 4140
rect 15150 4036 15156 4096
rect 15216 4036 15222 4096
rect 16174 4030 16234 4036
rect 16700 4002 16760 4230
rect 17716 4230 17730 4284
rect 17764 4284 17770 4806
rect 17764 4230 17776 4284
rect 16994 4180 17482 4186
rect 16994 4146 17006 4180
rect 17470 4146 17482 4180
rect 16994 4140 17482 4146
rect 17204 4002 17264 4140
rect 17716 4002 17776 4230
rect 15672 3932 15678 3992
rect 15738 3932 15744 3992
rect 16700 3942 17776 4002
rect 12922 3778 13410 3784
rect 12922 3744 12934 3778
rect 13398 3744 13410 3778
rect 12922 3738 13410 3744
rect 13940 3778 14428 3784
rect 13940 3744 13952 3778
rect 14416 3744 14428 3778
rect 13940 3738 14428 3744
rect 12622 3118 12640 3694
rect 12674 3118 12682 3694
rect 13652 3694 13698 3706
rect 13652 3174 13658 3694
rect 11904 3068 12392 3074
rect 11904 3034 11916 3068
rect 12380 3034 12392 3068
rect 11904 3028 12392 3034
rect 12106 2826 12166 3028
rect 12100 2766 12106 2826
rect 12166 2766 12172 2826
rect 12106 2672 12166 2766
rect 11904 2666 12392 2672
rect 11904 2632 11916 2666
rect 12380 2632 12392 2666
rect 11904 2626 12392 2632
rect 11608 2476 11622 2582
rect 11616 2068 11622 2476
rect 8850 1956 9338 1962
rect 8850 1922 8862 1956
rect 9326 1922 9338 1956
rect 8850 1916 9338 1922
rect 9868 1956 10356 1962
rect 9868 1922 9880 1956
rect 10344 1922 10356 1956
rect 9868 1916 10356 1922
rect 7534 1714 7540 1774
rect 7600 1714 7606 1774
rect 8028 1602 8034 1662
rect 8094 1602 8100 1662
rect 8034 1560 8094 1602
rect 6814 1554 7302 1560
rect 6814 1520 6826 1554
rect 7290 1520 7302 1554
rect 6814 1514 7302 1520
rect 7832 1554 8320 1560
rect 7832 1520 7844 1554
rect 8308 1520 8320 1554
rect 7832 1514 8320 1520
rect 6526 1470 6572 1482
rect 6526 936 6532 1470
rect 6516 894 6532 936
rect 6566 936 6572 1470
rect 7544 1470 7590 1482
rect 6566 894 6576 936
rect 7544 930 7550 1470
rect 6516 750 6576 894
rect 7534 894 7550 930
rect 7584 930 7590 1470
rect 8554 1470 8614 1822
rect 9058 1662 9118 1916
rect 9570 1714 9576 1774
rect 9636 1714 9642 1774
rect 9052 1602 9058 1662
rect 9118 1602 9124 1662
rect 8850 1554 9338 1560
rect 8850 1520 8862 1554
rect 9326 1520 9338 1554
rect 8850 1514 9338 1520
rect 8554 1368 8568 1470
rect 7584 894 7594 930
rect 6814 844 7302 850
rect 6814 810 6826 844
rect 7290 810 7302 844
rect 6814 804 7302 810
rect 7020 750 7080 804
rect 7534 750 7594 894
rect 8562 894 8568 1368
rect 8602 1368 8614 1470
rect 9576 1470 9636 1714
rect 10090 1662 10150 1916
rect 10590 1882 10650 2006
rect 11612 2006 11622 2068
rect 11656 2476 11668 2582
rect 12622 2582 12682 3118
rect 13642 3118 13658 3174
rect 13692 3174 13698 3694
rect 14656 3694 14716 3828
rect 14958 3778 15446 3784
rect 14958 3744 14970 3778
rect 15434 3744 15446 3778
rect 14958 3738 15446 3744
rect 13692 3118 13702 3174
rect 12922 3068 13410 3074
rect 12922 3034 12934 3068
rect 13398 3034 13410 3068
rect 12922 3028 13410 3034
rect 13642 2946 13702 3118
rect 14656 3118 14676 3694
rect 14710 3118 14716 3694
rect 13940 3068 14428 3074
rect 13940 3034 13952 3068
rect 14416 3034 14428 3068
rect 13940 3028 14428 3034
rect 13636 2886 13642 2946
rect 13702 2886 13708 2946
rect 12922 2666 13410 2672
rect 12922 2632 12934 2666
rect 13398 2632 13410 2666
rect 12922 2626 13410 2632
rect 11656 2068 11662 2476
rect 11656 2006 11672 2068
rect 10886 1956 11374 1962
rect 10886 1922 10898 1956
rect 11362 1922 11374 1956
rect 10886 1916 11374 1922
rect 10084 1602 10090 1662
rect 10150 1602 10156 1662
rect 9868 1554 10356 1560
rect 9868 1520 9880 1554
rect 10344 1520 10356 1554
rect 9868 1514 10356 1520
rect 9576 1430 9586 1470
rect 8602 894 8608 1368
rect 8562 882 8608 894
rect 9580 894 9586 1430
rect 9620 1430 9636 1470
rect 10590 1470 10650 1822
rect 11612 1774 11672 2006
rect 12622 2006 12640 2582
rect 12674 2006 12682 2582
rect 13642 2582 13702 2886
rect 13940 2666 14428 2672
rect 13940 2632 13952 2666
rect 14416 2632 14428 2666
rect 13940 2626 14428 2632
rect 13642 2540 13658 2582
rect 11904 1956 12392 1962
rect 11904 1922 11916 1956
rect 12380 1922 12392 1956
rect 11904 1916 12392 1922
rect 12622 1882 12682 2006
rect 13652 2006 13658 2540
rect 13692 2540 13702 2582
rect 14656 2582 14716 3118
rect 15678 3694 15738 3932
rect 16700 3888 16760 3942
rect 15976 3778 16464 3784
rect 15976 3744 15988 3778
rect 16452 3744 16464 3778
rect 15976 3738 16464 3744
rect 15678 3118 15694 3694
rect 15728 3118 15738 3694
rect 14958 3068 15446 3074
rect 14958 3034 14970 3068
rect 15434 3034 15446 3068
rect 14958 3028 15446 3034
rect 15168 2826 15228 3028
rect 15162 2766 15168 2826
rect 15228 2766 15234 2826
rect 15168 2672 15228 2766
rect 14958 2666 15446 2672
rect 14958 2632 14970 2666
rect 15434 2632 15446 2666
rect 14958 2626 15446 2632
rect 13692 2006 13698 2540
rect 13652 1994 13698 2006
rect 14656 2006 14676 2582
rect 14710 2006 14716 2582
rect 15678 2582 15738 3118
rect 16700 3694 16760 3828
rect 17204 3784 17264 3942
rect 16994 3778 17482 3784
rect 16994 3744 17006 3778
rect 17470 3744 17482 3778
rect 16994 3738 17482 3744
rect 16700 3118 16712 3694
rect 16746 3118 16760 3694
rect 15976 3068 16464 3074
rect 15976 3034 15988 3068
rect 16452 3034 16464 3068
rect 15976 3028 16464 3034
rect 16194 2826 16254 3028
rect 16700 2882 16760 3118
rect 17716 3694 17776 3942
rect 17716 3118 17730 3694
rect 17764 3118 17776 3694
rect 16994 3068 17482 3074
rect 16994 3034 17006 3068
rect 17470 3034 17482 3068
rect 16994 3028 17482 3034
rect 17200 2882 17260 3028
rect 17716 2882 17776 3118
rect 17856 2946 17916 5126
rect 17970 4036 17976 4096
rect 18036 4036 18042 4096
rect 17850 2886 17856 2946
rect 17916 2886 17922 2946
rect 16188 2766 16194 2826
rect 16254 2766 16260 2826
rect 16700 2822 17776 2882
rect 16194 2672 16254 2766
rect 15976 2666 16464 2672
rect 15976 2632 15988 2666
rect 16452 2632 16464 2666
rect 15976 2626 16464 2632
rect 15678 2526 15694 2582
rect 15688 2052 15694 2526
rect 12922 1956 13410 1962
rect 12922 1922 12934 1956
rect 13398 1922 13410 1956
rect 12922 1916 13410 1922
rect 13940 1956 14428 1962
rect 13940 1922 13952 1956
rect 14416 1922 14428 1956
rect 13940 1916 14428 1922
rect 11606 1714 11612 1774
rect 11672 1714 11678 1774
rect 11084 1602 11090 1662
rect 11150 1602 11156 1662
rect 12104 1602 12110 1662
rect 12170 1602 12176 1662
rect 11090 1560 11150 1602
rect 12110 1560 12170 1602
rect 10886 1554 11374 1560
rect 10886 1520 10898 1554
rect 11362 1520 11374 1554
rect 10886 1514 11374 1520
rect 11904 1554 12392 1560
rect 11904 1520 11916 1554
rect 12380 1520 12392 1554
rect 11904 1514 12392 1520
rect 10590 1432 10604 1470
rect 9620 894 9626 1430
rect 9580 882 9626 894
rect 10598 894 10604 1432
rect 10638 1432 10650 1470
rect 11616 1470 11662 1482
rect 10638 894 10644 1432
rect 11616 954 11622 1470
rect 10598 882 10644 894
rect 11614 894 11622 954
rect 11656 954 11662 1470
rect 12622 1470 12682 1822
rect 13130 1662 13190 1916
rect 13640 1714 13646 1774
rect 13706 1714 13712 1774
rect 13124 1602 13130 1662
rect 13190 1602 13196 1662
rect 12922 1554 13410 1560
rect 12922 1520 12934 1554
rect 13398 1520 13410 1554
rect 12922 1514 13410 1520
rect 12622 1410 12640 1470
rect 11656 894 11674 954
rect 7832 844 8320 850
rect 7832 810 7844 844
rect 8308 810 8320 844
rect 7832 804 8320 810
rect 8850 844 9338 850
rect 8850 810 8862 844
rect 9326 810 9338 844
rect 8850 804 9338 810
rect 9868 844 10356 850
rect 9868 810 9880 844
rect 10344 810 10356 844
rect 9868 804 10356 810
rect 10886 844 11374 850
rect 10886 810 10898 844
rect 11362 810 11374 844
rect 10886 804 11374 810
rect 6372 640 6378 700
rect 6438 640 6444 700
rect 6516 690 7594 750
rect 9048 700 9108 804
rect 10080 700 10140 804
rect 7534 570 7594 690
rect 9042 640 9048 700
rect 9108 640 9114 700
rect 10074 640 10080 700
rect 10140 640 10146 700
rect 11614 570 11674 894
rect 12634 894 12640 1410
rect 12674 1410 12682 1470
rect 13646 1470 13706 1714
rect 14140 1662 14200 1916
rect 14140 1596 14200 1602
rect 14656 1882 14716 2006
rect 15682 2006 15694 2052
rect 15728 2526 15738 2582
rect 16700 2582 16760 2822
rect 17200 2672 17260 2822
rect 16994 2666 17482 2672
rect 16994 2632 17006 2666
rect 17470 2632 17482 2666
rect 16994 2626 17482 2632
rect 15728 2052 15734 2526
rect 15728 2006 15742 2052
rect 14958 1956 15446 1962
rect 14958 1922 14970 1956
rect 15434 1922 15446 1956
rect 14958 1916 15446 1922
rect 13940 1554 14428 1560
rect 13940 1520 13952 1554
rect 14416 1520 14428 1554
rect 13940 1514 14428 1520
rect 13646 1424 13658 1470
rect 12674 894 12680 1410
rect 12634 882 12680 894
rect 13652 894 13658 1424
rect 13692 1424 13706 1470
rect 14656 1470 14716 1822
rect 15682 1774 15742 2006
rect 16700 2006 16712 2582
rect 16746 2006 16760 2582
rect 15976 1956 16464 1962
rect 15976 1922 15988 1956
rect 16452 1922 16464 1956
rect 15976 1916 16464 1922
rect 16700 1882 16760 2006
rect 17716 2582 17776 2822
rect 17716 2006 17730 2582
rect 17764 2006 17776 2582
rect 16994 1956 17482 1962
rect 16994 1922 17006 1956
rect 17470 1922 17482 1956
rect 16994 1916 17482 1922
rect 16694 1822 16700 1882
rect 16760 1822 16766 1882
rect 15676 1714 15682 1774
rect 15742 1714 15748 1774
rect 16700 1770 16760 1822
rect 17208 1770 17268 1916
rect 17716 1770 17776 2006
rect 16700 1710 17776 1770
rect 16172 1662 16232 1668
rect 15148 1602 15154 1662
rect 15214 1602 15220 1662
rect 15154 1560 15214 1602
rect 16172 1560 16232 1602
rect 14958 1554 15446 1560
rect 14958 1520 14970 1554
rect 15434 1520 15446 1554
rect 14958 1514 15446 1520
rect 15976 1554 16464 1560
rect 15976 1520 15988 1554
rect 16452 1520 16464 1554
rect 15976 1514 16464 1520
rect 14656 1428 14676 1470
rect 13692 894 13698 1424
rect 13652 882 13698 894
rect 14670 894 14676 1428
rect 14710 894 14716 1470
rect 15688 1470 15734 1482
rect 15688 922 15694 1470
rect 14670 882 14716 894
rect 15674 894 15694 922
rect 15728 894 15734 1470
rect 16700 1470 16760 1710
rect 17208 1560 17268 1710
rect 16994 1554 17482 1560
rect 16994 1520 17006 1554
rect 17470 1520 17482 1554
rect 16994 1514 17482 1520
rect 16700 1406 16712 1470
rect 11904 844 12392 850
rect 11904 810 11916 844
rect 12380 810 12392 844
rect 11904 804 12392 810
rect 12922 844 13410 850
rect 12922 810 12934 844
rect 13398 810 13410 844
rect 12922 804 13410 810
rect 13940 844 14428 850
rect 13940 810 13952 844
rect 14416 810 14428 844
rect 13940 804 14428 810
rect 14958 844 15446 850
rect 14958 810 14970 844
rect 15434 810 15446 844
rect 14958 804 15446 810
rect 13140 700 13200 804
rect 14136 700 14196 804
rect 13134 640 13140 700
rect 13200 640 13206 700
rect 14130 640 14136 700
rect 14196 640 14202 700
rect 15674 570 15734 894
rect 16706 894 16712 1406
rect 16746 1406 16760 1470
rect 17716 1470 17776 1710
rect 17716 1428 17730 1470
rect 16746 894 16752 1406
rect 16706 882 16752 894
rect 17724 894 17730 1428
rect 17764 1428 17776 1470
rect 17764 894 17770 1428
rect 17724 882 17770 894
rect 15976 844 16464 850
rect 15976 810 15988 844
rect 16452 810 16464 844
rect 15976 804 16464 810
rect 16994 844 17482 850
rect 16994 810 17006 844
rect 17470 810 17482 844
rect 16994 804 17482 810
rect 17856 570 17916 2886
rect 17976 1662 18036 4036
rect 17970 1602 17976 1662
rect 18036 1602 18042 1662
rect 11608 510 11614 570
rect 11674 510 11680 570
rect 15668 510 15674 570
rect 15734 510 15740 570
rect 17850 510 17856 570
rect 17916 510 17922 570
rect 7534 504 7594 510
rect 6942 104 17212 164
rect 6976 -72 7036 104
rect 7476 18 7536 104
rect 7272 12 7760 18
rect 7272 -22 7284 12
rect 7748 -22 7760 12
rect 7272 -28 7760 -22
rect 6976 -106 6990 -72
rect 6984 -648 6990 -106
rect 7024 -106 7036 -72
rect 7998 -72 8058 104
rect 8496 18 8556 104
rect 9530 18 9590 104
rect 10552 18 10612 104
rect 11542 18 11602 104
rect 8290 12 8778 18
rect 8290 -22 8302 12
rect 8766 -22 8778 12
rect 8290 -28 8778 -22
rect 9308 12 9796 18
rect 9308 -22 9320 12
rect 9784 -22 9796 12
rect 9308 -28 9796 -22
rect 10326 12 10814 18
rect 10326 -22 10338 12
rect 10802 -22 10814 12
rect 10326 -28 10814 -22
rect 11344 12 11832 18
rect 11344 -22 11356 12
rect 11820 -22 11832 12
rect 11344 -28 11832 -22
rect 7024 -648 7030 -106
rect 7998 -116 8008 -72
rect 6984 -660 7030 -648
rect 8002 -648 8008 -116
rect 8042 -116 8058 -72
rect 9020 -72 9066 -60
rect 8042 -648 8048 -116
rect 9020 -590 9026 -72
rect 8002 -660 8048 -648
rect 9012 -648 9026 -590
rect 9060 -590 9066 -72
rect 10038 -72 10084 -60
rect 9060 -648 9072 -590
rect 10038 -614 10044 -72
rect 7272 -698 7760 -692
rect 7272 -732 7284 -698
rect 7748 -732 7760 -698
rect 7272 -738 7760 -732
rect 8290 -698 8778 -692
rect 8290 -732 8302 -698
rect 8766 -732 8778 -698
rect 8290 -738 8778 -732
rect 9012 -796 9072 -648
rect 10030 -648 10044 -614
rect 10078 -614 10084 -72
rect 11056 -72 11102 -60
rect 11056 -602 11062 -72
rect 10078 -648 10090 -614
rect 9308 -698 9796 -692
rect 9308 -732 9320 -698
rect 9784 -732 9796 -698
rect 9308 -738 9796 -732
rect 9006 -856 9012 -796
rect 9072 -856 9078 -796
rect 4712 -2036 4824 -1250
rect 9012 -1350 9072 -856
rect 10030 -908 10090 -648
rect 11050 -648 11062 -602
rect 11096 -602 11102 -72
rect 12066 -72 12126 104
rect 12576 18 12636 104
rect 13566 18 13626 104
rect 14598 18 14658 104
rect 15602 18 15662 104
rect 12362 12 12850 18
rect 12362 -22 12374 12
rect 12838 -22 12850 12
rect 12362 -28 12850 -22
rect 13380 12 13868 18
rect 13380 -22 13392 12
rect 13856 -22 13868 12
rect 13380 -28 13868 -22
rect 14398 12 14886 18
rect 14398 -22 14410 12
rect 14874 -22 14886 12
rect 14398 -28 14886 -22
rect 15416 12 15904 18
rect 15416 -22 15428 12
rect 15892 -22 15904 12
rect 15416 -28 15904 -22
rect 12576 -30 12636 -28
rect 14598 -30 14658 -28
rect 12066 -114 12080 -72
rect 11096 -648 11110 -602
rect 10326 -698 10814 -692
rect 10326 -732 10338 -698
rect 10802 -732 10814 -698
rect 10326 -738 10814 -732
rect 11050 -796 11110 -648
rect 12074 -648 12080 -114
rect 12114 -114 12126 -72
rect 13092 -72 13138 -60
rect 12114 -648 12120 -114
rect 13092 -602 13098 -72
rect 12074 -660 12120 -648
rect 13086 -648 13098 -602
rect 13132 -602 13138 -72
rect 14110 -72 14156 -60
rect 13132 -648 13146 -602
rect 14110 -610 14116 -72
rect 11344 -698 11832 -692
rect 11344 -732 11356 -698
rect 11820 -732 11832 -698
rect 11344 -738 11832 -732
rect 12362 -698 12850 -692
rect 12362 -732 12374 -698
rect 12838 -732 12850 -698
rect 12362 -738 12850 -732
rect 13086 -796 13146 -648
rect 14104 -648 14116 -610
rect 14150 -610 14156 -72
rect 15128 -72 15174 -60
rect 14150 -648 14164 -610
rect 15128 -616 15134 -72
rect 13380 -698 13868 -692
rect 13380 -732 13392 -698
rect 13856 -732 13868 -698
rect 13380 -738 13868 -732
rect 11044 -856 11050 -796
rect 11110 -856 11116 -796
rect 13080 -856 13086 -796
rect 13146 -856 13152 -796
rect 10024 -968 10030 -908
rect 10090 -968 10096 -908
rect 11050 -1350 11110 -856
rect 13086 -1350 13146 -856
rect 14104 -908 14164 -648
rect 15122 -648 15134 -616
rect 15168 -616 15174 -72
rect 16142 -72 16202 104
rect 16622 18 16682 104
rect 16434 12 16922 18
rect 16434 -22 16446 12
rect 16910 -22 16922 12
rect 16434 -28 16922 -22
rect 16142 -140 16152 -72
rect 15168 -648 15182 -616
rect 14398 -698 14886 -692
rect 14398 -732 14410 -698
rect 14874 -732 14886 -698
rect 14398 -738 14886 -732
rect 15122 -796 15182 -648
rect 16146 -648 16152 -140
rect 16186 -140 16202 -72
rect 17152 -72 17212 104
rect 17152 -112 17170 -72
rect 16186 -648 16192 -140
rect 16146 -660 16192 -648
rect 17164 -648 17170 -112
rect 17204 -112 17212 -72
rect 17204 -648 17210 -112
rect 17164 -660 17210 -648
rect 15416 -698 15904 -692
rect 15416 -732 15428 -698
rect 15892 -732 15904 -698
rect 15416 -738 15904 -732
rect 16434 -698 16922 -692
rect 16434 -732 16446 -698
rect 16910 -732 16922 -698
rect 16434 -738 16922 -732
rect 15116 -856 15122 -796
rect 15182 -856 15188 -796
rect 14098 -968 14104 -908
rect 14164 -968 14170 -908
rect 15122 -1350 15182 -856
rect 18110 -908 18170 6020
rect 18322 5186 18382 13526
rect 18316 5126 18322 5186
rect 18382 5126 18388 5186
rect 18442 5058 18502 13528
rect 18436 4998 18442 5058
rect 18502 4998 18508 5058
rect 18582 4096 18642 13546
rect 18694 13408 18700 13468
rect 18760 13408 18766 13468
rect 18700 7340 18760 13408
rect 18810 12726 18870 13562
rect 18804 12666 18810 12726
rect 18870 12666 18876 12726
rect 18928 9806 18988 13662
rect 19256 12860 19316 13672
rect 19250 12800 19256 12860
rect 19316 12800 19322 12860
rect 19046 11442 19052 11502
rect 19112 11442 19118 11502
rect 18926 9800 18988 9806
rect 18986 9740 18988 9800
rect 18926 9734 18988 9740
rect 18694 7280 18700 7340
rect 18760 7280 18766 7340
rect 18576 4036 18582 4096
rect 18642 4036 18648 4096
rect 18928 3738 18988 9734
rect 19052 8806 19112 11442
rect 19258 11106 19264 11166
rect 19324 11106 19330 11166
rect 19154 9846 19160 9906
rect 19220 9846 19226 9906
rect 19046 8746 19052 8806
rect 19112 8746 19118 8806
rect 19160 3888 19220 9846
rect 19264 8570 19324 11106
rect 19376 8684 19436 13664
rect 19482 13588 19542 13594
rect 19482 11044 19542 13528
rect 30288 13232 30294 13238
rect 19608 13178 30294 13232
rect 30354 13232 30360 13238
rect 35392 13232 35398 13238
rect 30354 13178 35398 13232
rect 35458 13232 35464 13238
rect 39458 13232 39518 13238
rect 35458 13178 39458 13232
rect 19608 13172 39458 13178
rect 39518 13172 40030 13232
rect 19608 13032 19668 13172
rect 20130 13122 20190 13172
rect 21140 13122 21200 13172
rect 19904 13116 20392 13122
rect 19904 13082 19916 13116
rect 20380 13082 20392 13116
rect 19904 13076 20392 13082
rect 20922 13116 21410 13122
rect 20922 13082 20934 13116
rect 21398 13082 21410 13116
rect 20922 13076 21410 13082
rect 21140 13070 21200 13076
rect 19608 12456 19622 13032
rect 19656 12456 19668 13032
rect 20634 13032 20680 13044
rect 20634 12490 20640 13032
rect 19608 12214 19668 12456
rect 20626 12456 20640 12490
rect 20674 12490 20680 13032
rect 21646 13032 21706 13172
rect 22170 13122 22230 13172
rect 23182 13122 23242 13172
rect 21940 13116 22428 13122
rect 21940 13082 21952 13116
rect 22416 13082 22428 13116
rect 21940 13076 22428 13082
rect 22958 13116 23446 13122
rect 22958 13082 22970 13116
rect 23434 13082 23446 13116
rect 22958 13076 23446 13082
rect 23182 13070 23242 13076
rect 20674 12456 20686 12490
rect 19904 12406 20392 12412
rect 19904 12372 19916 12406
rect 20380 12372 20392 12406
rect 19904 12366 20392 12372
rect 20120 12304 20180 12366
rect 19904 12298 20392 12304
rect 19904 12264 19916 12298
rect 20380 12264 20392 12298
rect 19904 12258 20392 12264
rect 20120 12252 20180 12258
rect 19608 11638 19622 12214
rect 19656 11638 19668 12214
rect 19608 11166 19668 11638
rect 20626 12214 20686 12456
rect 21646 12456 21658 13032
rect 21692 12456 21706 13032
rect 22670 13032 22716 13044
rect 22670 12502 22676 13032
rect 21126 12412 21186 12414
rect 20922 12406 21410 12412
rect 20922 12372 20934 12406
rect 21398 12372 21410 12406
rect 20922 12366 21410 12372
rect 21126 12304 21186 12366
rect 20922 12298 21410 12304
rect 20922 12264 20934 12298
rect 21398 12264 21410 12298
rect 20922 12258 21410 12264
rect 20626 11638 20640 12214
rect 20674 11638 20686 12214
rect 21646 12214 21706 12456
rect 22660 12456 22676 12502
rect 22710 12502 22716 13032
rect 23678 13032 23738 13172
rect 24194 13122 24254 13172
rect 25194 13122 25254 13172
rect 23976 13116 24464 13122
rect 23976 13082 23988 13116
rect 24452 13082 24464 13116
rect 23976 13076 24464 13082
rect 24994 13116 25482 13122
rect 24994 13082 25006 13116
rect 25470 13082 25482 13116
rect 24994 13076 25482 13082
rect 22710 12456 22720 12502
rect 22138 12412 22198 12420
rect 21940 12406 22428 12412
rect 21940 12372 21952 12406
rect 22416 12372 22428 12406
rect 21940 12366 22428 12372
rect 22138 12304 22198 12366
rect 21940 12298 22428 12304
rect 21940 12264 21952 12298
rect 22416 12264 22428 12298
rect 21940 12258 22428 12264
rect 21646 12156 21658 12214
rect 19904 11588 20392 11594
rect 19904 11554 19916 11588
rect 20380 11554 20392 11588
rect 19904 11548 20392 11554
rect 20626 11502 20686 11638
rect 21652 11638 21658 12156
rect 21692 12156 21706 12214
rect 22660 12214 22720 12456
rect 23678 12456 23694 13032
rect 23728 12456 23738 13032
rect 24706 13032 24752 13044
rect 24706 12496 24712 13032
rect 22958 12406 23446 12412
rect 22958 12372 22970 12406
rect 23434 12372 23446 12406
rect 22958 12366 23446 12372
rect 23160 12304 23220 12366
rect 22958 12298 23446 12304
rect 22958 12264 22970 12298
rect 23434 12264 23446 12298
rect 22958 12258 23446 12264
rect 23160 12252 23220 12258
rect 21692 11638 21698 12156
rect 21652 11626 21698 11638
rect 22660 11638 22676 12214
rect 22710 11638 22720 12214
rect 23678 12214 23738 12456
rect 24696 12456 24712 12496
rect 24746 12496 24752 13032
rect 25716 13032 25776 13172
rect 26228 13122 26288 13172
rect 27240 13122 27300 13172
rect 26012 13116 26500 13122
rect 26012 13082 26024 13116
rect 26488 13082 26500 13116
rect 26012 13076 26500 13082
rect 27030 13116 27518 13122
rect 27030 13082 27042 13116
rect 27506 13082 27518 13116
rect 27030 13076 27518 13082
rect 24746 12456 24756 12496
rect 23976 12406 24464 12412
rect 23976 12372 23988 12406
rect 24452 12372 24464 12406
rect 23976 12366 24464 12372
rect 24172 12304 24232 12366
rect 23976 12298 24464 12304
rect 23976 12264 23988 12298
rect 24452 12264 24464 12298
rect 23976 12258 24464 12264
rect 24172 12252 24232 12258
rect 23678 12152 23694 12214
rect 20922 11588 21410 11594
rect 20922 11554 20934 11588
rect 21398 11554 21410 11588
rect 20922 11548 21410 11554
rect 21940 11588 22428 11594
rect 21940 11554 21952 11588
rect 22416 11554 22428 11588
rect 21940 11548 22428 11554
rect 22660 11500 22720 11638
rect 23688 11638 23694 12152
rect 23728 12152 23738 12214
rect 24696 12214 24756 12456
rect 25716 12456 25730 13032
rect 25764 12456 25776 13032
rect 26742 13032 26788 13044
rect 26742 12496 26748 13032
rect 24994 12406 25482 12412
rect 24994 12372 25006 12406
rect 25470 12372 25482 12406
rect 24994 12366 25482 12372
rect 25202 12304 25262 12366
rect 24994 12298 25482 12304
rect 24994 12264 25006 12298
rect 25470 12264 25482 12298
rect 24994 12258 25482 12264
rect 25202 12252 25262 12258
rect 23728 11638 23734 12152
rect 23688 11626 23734 11638
rect 24696 11638 24712 12214
rect 24746 11638 24756 12214
rect 25716 12214 25776 12456
rect 26734 12456 26748 12496
rect 26782 12496 26788 13032
rect 27752 13032 27812 13172
rect 28264 13122 28324 13172
rect 29276 13122 29336 13172
rect 28048 13116 28536 13122
rect 28048 13082 28060 13116
rect 28524 13082 28536 13116
rect 28048 13076 28536 13082
rect 29066 13116 29554 13122
rect 29066 13082 29078 13116
rect 29542 13082 29554 13116
rect 29066 13076 29554 13082
rect 26782 12456 26794 12496
rect 26208 12412 26268 12414
rect 26012 12406 26500 12412
rect 26012 12372 26024 12406
rect 26488 12372 26500 12406
rect 26012 12366 26500 12372
rect 26208 12304 26268 12366
rect 26012 12298 26500 12304
rect 26012 12264 26024 12298
rect 26488 12264 26500 12298
rect 26012 12258 26500 12264
rect 25716 12172 25730 12214
rect 22958 11588 23446 11594
rect 22958 11554 22970 11588
rect 23434 11554 23446 11588
rect 22958 11548 23446 11554
rect 23976 11588 24464 11594
rect 23976 11554 23988 11588
rect 24452 11554 24464 11588
rect 23976 11548 24464 11554
rect 24696 11500 24756 11638
rect 25724 11638 25730 12172
rect 25764 12172 25776 12214
rect 26734 12214 26794 12456
rect 27752 12456 27766 13032
rect 27800 12456 27812 13032
rect 28778 13032 28824 13044
rect 28778 12502 28784 13032
rect 27230 12412 27290 12414
rect 27030 12406 27518 12412
rect 27030 12372 27042 12406
rect 27506 12372 27518 12406
rect 27030 12366 27518 12372
rect 27230 12304 27290 12366
rect 27030 12298 27518 12304
rect 27030 12264 27042 12298
rect 27506 12264 27518 12298
rect 27030 12258 27518 12264
rect 25764 11638 25770 12172
rect 25724 11626 25770 11638
rect 26734 11638 26748 12214
rect 26782 11638 26794 12214
rect 27752 12214 27812 12456
rect 28772 12456 28784 12502
rect 28818 12502 28824 13032
rect 29784 13032 29844 13172
rect 30298 13122 30358 13172
rect 31310 13122 31370 13172
rect 30084 13116 30572 13122
rect 30084 13082 30096 13116
rect 30560 13082 30572 13116
rect 30084 13076 30572 13082
rect 31102 13116 31590 13122
rect 31102 13082 31114 13116
rect 31578 13082 31590 13116
rect 31102 13076 31590 13082
rect 31310 13070 31370 13076
rect 28818 12456 28832 12502
rect 28048 12406 28536 12412
rect 28048 12372 28060 12406
rect 28524 12372 28536 12406
rect 28048 12366 28536 12372
rect 28254 12304 28314 12366
rect 28048 12298 28536 12304
rect 28048 12264 28060 12298
rect 28524 12264 28536 12298
rect 28048 12258 28536 12264
rect 28254 12252 28314 12258
rect 27752 12164 27766 12214
rect 24994 11588 25482 11594
rect 24994 11554 25006 11588
rect 25470 11554 25482 11588
rect 24994 11548 25482 11554
rect 26012 11588 26500 11594
rect 26012 11554 26024 11588
rect 26488 11554 26500 11588
rect 26012 11548 26500 11554
rect 26734 11500 26794 11638
rect 27760 11638 27766 12164
rect 27800 12164 27812 12214
rect 28772 12214 28832 12456
rect 29784 12456 29802 13032
rect 29836 12456 29844 13032
rect 30814 13032 30860 13044
rect 30814 12502 30820 13032
rect 29260 12412 29320 12414
rect 29066 12406 29554 12412
rect 29066 12372 29078 12406
rect 29542 12372 29554 12406
rect 29066 12366 29554 12372
rect 29260 12304 29320 12366
rect 29066 12298 29554 12304
rect 29066 12264 29078 12298
rect 29542 12264 29554 12298
rect 29066 12258 29554 12264
rect 27800 11638 27806 12164
rect 27760 11626 27806 11638
rect 28772 11638 28784 12214
rect 28818 11638 28832 12214
rect 29784 12214 29844 12456
rect 30806 12456 30820 12502
rect 30854 12502 30860 13032
rect 31822 13032 31882 13172
rect 32334 13122 32394 13172
rect 33352 13122 33412 13172
rect 32120 13116 32608 13122
rect 32120 13082 32132 13116
rect 32596 13082 32608 13116
rect 32120 13076 32608 13082
rect 33138 13116 33626 13122
rect 33138 13082 33150 13116
rect 33614 13082 33626 13116
rect 33138 13076 33626 13082
rect 32334 13070 32394 13076
rect 30854 12456 30866 12502
rect 30284 12412 30344 12420
rect 30084 12406 30572 12412
rect 30084 12372 30096 12406
rect 30560 12372 30572 12406
rect 30084 12366 30572 12372
rect 30284 12304 30344 12366
rect 30084 12298 30572 12304
rect 30084 12264 30096 12298
rect 30560 12264 30572 12298
rect 30084 12258 30572 12264
rect 29784 12166 29802 12214
rect 27030 11588 27518 11594
rect 27030 11554 27042 11588
rect 27506 11554 27518 11588
rect 27030 11548 27518 11554
rect 28048 11588 28536 11594
rect 28048 11554 28060 11588
rect 28524 11554 28536 11588
rect 28048 11548 28536 11554
rect 28772 11500 28832 11638
rect 29796 11638 29802 12166
rect 29836 12166 29844 12214
rect 30806 12214 30866 12456
rect 31822 12456 31838 13032
rect 31872 12456 31882 13032
rect 32850 13032 32896 13044
rect 32850 12502 32856 13032
rect 31306 12412 31366 12414
rect 31102 12406 31590 12412
rect 31102 12372 31114 12406
rect 31578 12372 31590 12406
rect 31102 12366 31590 12372
rect 31306 12304 31366 12366
rect 31102 12298 31590 12304
rect 31102 12264 31114 12298
rect 31578 12264 31590 12298
rect 31102 12258 31590 12264
rect 29836 11638 29842 12166
rect 29796 11626 29842 11638
rect 30806 11638 30820 12214
rect 30854 11638 30866 12214
rect 31822 12214 31882 12456
rect 32842 12456 32856 12502
rect 32890 12502 32896 13032
rect 33858 13032 33918 13172
rect 34374 13122 34434 13172
rect 35398 13122 35458 13172
rect 34156 13116 34644 13122
rect 34156 13082 34168 13116
rect 34632 13082 34644 13116
rect 34156 13076 34644 13082
rect 35174 13116 35662 13122
rect 35174 13082 35186 13116
rect 35650 13082 35662 13116
rect 35174 13076 35662 13082
rect 32890 12456 32902 12502
rect 32318 12412 32378 12414
rect 32120 12406 32608 12412
rect 32120 12372 32132 12406
rect 32596 12372 32608 12406
rect 32120 12366 32608 12372
rect 32318 12304 32378 12366
rect 32120 12298 32608 12304
rect 32120 12264 32132 12298
rect 32596 12264 32608 12298
rect 32120 12258 32608 12264
rect 31822 12164 31838 12214
rect 29066 11588 29554 11594
rect 29066 11554 29078 11588
rect 29542 11554 29554 11588
rect 29066 11548 29554 11554
rect 30084 11588 30572 11594
rect 30084 11554 30096 11588
rect 30560 11554 30572 11588
rect 30084 11548 30572 11554
rect 30806 11500 30866 11638
rect 31832 11638 31838 12164
rect 31872 12164 31882 12214
rect 32842 12214 32902 12456
rect 33858 12456 33874 13032
rect 33908 12456 33918 13032
rect 34886 13032 34932 13044
rect 34886 12526 34892 13032
rect 33138 12406 33626 12412
rect 33138 12372 33150 12406
rect 33614 12372 33626 12406
rect 33138 12366 33626 12372
rect 33330 12304 33390 12366
rect 33138 12298 33626 12304
rect 33138 12264 33150 12298
rect 33614 12264 33626 12298
rect 33138 12258 33626 12264
rect 33330 12252 33390 12258
rect 31872 11638 31878 12164
rect 31832 11626 31878 11638
rect 32842 11638 32856 12214
rect 32890 11638 32902 12214
rect 33858 12214 33918 12456
rect 34880 12456 34892 12526
rect 34926 12526 34932 13032
rect 35894 13032 35954 13172
rect 36416 13122 36476 13172
rect 37428 13122 37488 13172
rect 36192 13116 36680 13122
rect 36192 13082 36204 13116
rect 36668 13082 36680 13116
rect 36192 13076 36680 13082
rect 37210 13116 37698 13122
rect 37210 13082 37222 13116
rect 37686 13082 37698 13116
rect 37210 13076 37698 13082
rect 34926 12456 34940 12526
rect 34354 12412 34414 12420
rect 34156 12406 34644 12412
rect 34156 12372 34168 12406
rect 34632 12372 34644 12406
rect 34156 12366 34644 12372
rect 34354 12304 34414 12366
rect 34156 12298 34644 12304
rect 34156 12264 34168 12298
rect 34632 12264 34644 12298
rect 34156 12258 34644 12264
rect 33858 12190 33874 12214
rect 31102 11588 31590 11594
rect 31102 11554 31114 11588
rect 31578 11554 31590 11588
rect 31102 11548 31590 11554
rect 32120 11588 32608 11594
rect 32120 11554 32132 11588
rect 32596 11554 32608 11588
rect 32120 11548 32608 11554
rect 32842 11500 32902 11638
rect 33868 11638 33874 12190
rect 33908 12190 33918 12214
rect 34880 12214 34940 12456
rect 35894 12456 35910 13032
rect 35944 12456 35954 13032
rect 36922 13032 36968 13044
rect 36922 12566 36928 13032
rect 35174 12406 35662 12412
rect 35174 12372 35186 12406
rect 35650 12372 35662 12406
rect 35174 12366 35662 12372
rect 35376 12304 35436 12366
rect 35174 12298 35662 12304
rect 35174 12264 35186 12298
rect 35650 12264 35662 12298
rect 35174 12258 35662 12264
rect 35376 12246 35436 12258
rect 33908 11638 33914 12190
rect 33868 11626 33914 11638
rect 34880 11638 34892 12214
rect 34926 11638 34940 12214
rect 35894 12214 35954 12456
rect 36914 12456 36928 12566
rect 36962 12566 36968 13032
rect 37932 13032 37992 13172
rect 38438 13122 38498 13172
rect 39456 13166 39518 13172
rect 39456 13122 39516 13166
rect 38228 13116 38716 13122
rect 38228 13082 38240 13116
rect 38704 13082 38716 13116
rect 38228 13076 38716 13082
rect 39246 13116 39734 13122
rect 39246 13082 39258 13116
rect 39722 13082 39734 13116
rect 39246 13076 39734 13082
rect 36962 12456 36974 12566
rect 36394 12412 36454 12414
rect 36192 12406 36680 12412
rect 36192 12372 36204 12406
rect 36668 12372 36680 12406
rect 36192 12366 36680 12372
rect 36394 12304 36454 12366
rect 36192 12298 36680 12304
rect 36192 12264 36204 12298
rect 36668 12264 36680 12298
rect 36192 12258 36680 12264
rect 35894 12172 35910 12214
rect 33138 11588 33626 11594
rect 33138 11554 33150 11588
rect 33614 11554 33626 11588
rect 33138 11548 33626 11554
rect 34156 11588 34644 11594
rect 34156 11554 34168 11588
rect 34632 11554 34644 11588
rect 34156 11548 34644 11554
rect 34880 11500 34940 11638
rect 35904 11638 35910 12172
rect 35944 12172 35954 12214
rect 36914 12214 36974 12456
rect 37932 12456 37946 13032
rect 37980 12456 37992 13032
rect 38958 13032 39004 13044
rect 38958 12516 38964 13032
rect 37424 12412 37484 12426
rect 37210 12406 37698 12412
rect 37210 12372 37222 12406
rect 37686 12372 37698 12406
rect 37210 12366 37698 12372
rect 37424 12304 37484 12366
rect 37210 12298 37698 12304
rect 37210 12264 37222 12298
rect 37686 12264 37698 12298
rect 37210 12258 37698 12264
rect 35944 11638 35950 12172
rect 35904 11626 35950 11638
rect 36914 11638 36928 12214
rect 36962 11638 36974 12214
rect 37932 12214 37992 12456
rect 38950 12456 38964 12516
rect 38998 12516 39004 13032
rect 39970 13032 40030 13172
rect 38998 12456 39010 12516
rect 38436 12412 38496 12426
rect 38228 12406 38716 12412
rect 38228 12372 38240 12406
rect 38704 12372 38716 12406
rect 38228 12366 38716 12372
rect 38436 12304 38496 12366
rect 38228 12298 38716 12304
rect 38228 12264 38240 12298
rect 38704 12264 38716 12298
rect 38228 12258 38716 12264
rect 37932 12172 37946 12214
rect 35174 11588 35662 11594
rect 35174 11554 35186 11588
rect 35650 11554 35662 11588
rect 35174 11548 35662 11554
rect 36192 11588 36680 11594
rect 36192 11554 36204 11588
rect 36668 11554 36680 11588
rect 36192 11548 36680 11554
rect 36914 11500 36974 11638
rect 37940 11638 37946 12172
rect 37980 12172 37992 12214
rect 38950 12214 39010 12456
rect 39970 12456 39982 13032
rect 40016 12456 40030 13032
rect 39246 12406 39734 12412
rect 39246 12372 39258 12406
rect 39722 12372 39734 12406
rect 39246 12366 39734 12372
rect 39436 12304 39496 12366
rect 39970 12364 40030 12456
rect 41856 13010 41968 13796
rect 39970 12304 40750 12364
rect 39246 12298 39734 12304
rect 39246 12264 39258 12298
rect 39722 12264 39734 12298
rect 39246 12258 39734 12264
rect 39436 12252 39496 12258
rect 37980 11638 37986 12172
rect 37940 11626 37986 11638
rect 38950 11638 38964 12214
rect 38998 11638 39010 12214
rect 39970 12214 40030 12304
rect 39970 12164 39982 12214
rect 37210 11588 37698 11594
rect 37210 11554 37222 11588
rect 37686 11554 37698 11588
rect 37210 11548 37698 11554
rect 38228 11588 38716 11594
rect 38228 11554 38240 11588
rect 38704 11554 38716 11588
rect 38228 11548 38716 11554
rect 38950 11500 39010 11638
rect 39976 11638 39982 12164
rect 40016 12164 40030 12214
rect 40016 11638 40022 12164
rect 39976 11626 40022 11638
rect 39246 11588 39734 11594
rect 39246 11554 39258 11588
rect 39722 11554 39734 11588
rect 39246 11548 39734 11554
rect 20686 11442 40628 11500
rect 20626 11440 40628 11442
rect 20626 11436 20686 11440
rect 21634 11226 21640 11286
rect 21700 11226 21706 11286
rect 23674 11226 23680 11286
rect 23740 11226 23746 11286
rect 25714 11226 25720 11286
rect 25780 11226 25786 11286
rect 27744 11226 27750 11286
rect 27810 11226 27816 11286
rect 29784 11226 29790 11286
rect 29850 11226 29856 11286
rect 31816 11226 31822 11286
rect 31882 11226 31888 11286
rect 33856 11226 33862 11286
rect 33922 11226 33928 11286
rect 35892 11226 35898 11286
rect 35958 11226 35964 11286
rect 37926 11226 37932 11286
rect 37992 11226 37998 11286
rect 19602 11106 19608 11166
rect 19668 11106 19674 11166
rect 21126 11100 21132 11160
rect 21192 11100 21198 11160
rect 19476 10984 19482 11044
rect 19542 10984 19548 11044
rect 19482 8910 19542 10984
rect 21132 10926 21192 11100
rect 19904 10920 20392 10926
rect 19904 10886 19916 10920
rect 20380 10886 20392 10920
rect 19904 10880 20392 10886
rect 20922 10920 21410 10926
rect 20922 10886 20934 10920
rect 21398 10886 21410 10920
rect 20922 10880 21410 10886
rect 19616 10836 19662 10848
rect 20634 10836 20680 10848
rect 21640 10836 21700 11226
rect 22146 11160 22206 11166
rect 22146 10926 22206 11100
rect 23168 11160 23228 11166
rect 23168 10926 23228 11100
rect 21940 10920 22428 10926
rect 21940 10886 21952 10920
rect 22416 10886 22428 10920
rect 21940 10880 22428 10886
rect 22958 10920 23446 10926
rect 22958 10886 22970 10920
rect 23434 10886 23446 10920
rect 22958 10880 23446 10886
rect 22670 10836 22716 10848
rect 19608 10802 19622 10836
rect 19616 10310 19622 10802
rect 19608 10260 19622 10310
rect 19656 10802 19668 10836
rect 19656 10310 19662 10802
rect 20626 10788 20640 10836
rect 19656 10260 19668 10310
rect 20634 10296 20640 10788
rect 19608 10122 19668 10260
rect 20626 10260 20640 10296
rect 20674 10788 20686 10836
rect 20674 10296 20680 10788
rect 21640 10768 21658 10836
rect 21652 10324 21658 10768
rect 20674 10260 20686 10296
rect 19904 10210 20392 10216
rect 19904 10176 19916 10210
rect 20380 10176 20392 10210
rect 19904 10170 20392 10176
rect 20110 10122 20170 10170
rect 20626 10122 20686 10260
rect 21644 10260 21658 10324
rect 21692 10804 21704 10836
rect 21692 10768 21700 10804
rect 21692 10324 21698 10768
rect 21692 10260 21704 10324
rect 22670 10306 22676 10836
rect 22666 10288 22676 10306
rect 22664 10260 22676 10288
rect 22710 10306 22716 10836
rect 23680 10836 23740 11226
rect 24182 11160 24242 11166
rect 24180 11100 24182 11106
rect 25208 11160 25268 11166
rect 24180 11094 24242 11100
rect 25206 11100 25208 11106
rect 25206 11094 25268 11100
rect 24180 10926 24240 11094
rect 24690 10984 24696 11044
rect 24756 10984 24762 11044
rect 23976 10920 24464 10926
rect 23976 10886 23988 10920
rect 24452 10886 24464 10920
rect 23976 10880 24464 10886
rect 23680 10782 23694 10836
rect 23688 10332 23694 10782
rect 23684 10308 23694 10332
rect 22710 10260 22726 10306
rect 23682 10260 23694 10308
rect 23728 10782 23740 10836
rect 24696 10836 24756 10984
rect 25206 10926 25266 11094
rect 24994 10920 25482 10926
rect 24994 10886 25006 10920
rect 25470 10886 25482 10920
rect 24994 10880 25482 10886
rect 24696 10794 24712 10836
rect 23728 10332 23734 10782
rect 24706 10336 24712 10794
rect 23728 10260 23744 10332
rect 24696 10260 24712 10336
rect 24746 10794 24756 10836
rect 25720 10836 25780 11226
rect 26220 11160 26280 11166
rect 26220 10926 26280 11100
rect 27256 11160 27316 11166
rect 27256 10926 27316 11100
rect 26012 10920 26500 10926
rect 26012 10886 26024 10920
rect 26488 10886 26500 10920
rect 26012 10880 26500 10886
rect 27030 10920 27518 10926
rect 27030 10886 27042 10920
rect 27506 10886 27518 10920
rect 27030 10880 27518 10886
rect 26742 10836 26788 10848
rect 27750 10836 27810 11226
rect 28262 11160 28322 11166
rect 29270 11100 29276 11160
rect 29336 11100 29342 11160
rect 28262 10926 28322 11100
rect 29276 10926 29336 11100
rect 28048 10920 28536 10926
rect 28048 10886 28060 10920
rect 28524 10886 28536 10920
rect 28048 10880 28536 10886
rect 29066 10920 29554 10926
rect 29066 10886 29078 10920
rect 29542 10886 29554 10920
rect 29066 10880 29554 10886
rect 24746 10336 24752 10794
rect 25720 10762 25730 10836
rect 24746 10320 24756 10336
rect 24746 10260 24760 10320
rect 25724 10316 25730 10762
rect 25716 10260 25730 10316
rect 25764 10762 25780 10836
rect 26736 10786 26748 10836
rect 25764 10316 25770 10762
rect 26742 10324 26748 10786
rect 25764 10260 25776 10316
rect 26736 10296 26748 10324
rect 26734 10260 26748 10296
rect 26782 10786 26796 10836
rect 26782 10324 26788 10786
rect 27750 10768 27766 10836
rect 27760 10336 27766 10768
rect 26782 10260 26796 10324
rect 20922 10210 21410 10216
rect 20922 10176 20934 10210
rect 21398 10176 21410 10210
rect 20922 10170 21410 10176
rect 19608 10062 20686 10122
rect 20626 9906 20686 10062
rect 21136 10012 21196 10170
rect 21644 10122 21704 10260
rect 21940 10210 22428 10216
rect 21940 10176 21952 10210
rect 22416 10176 22428 10210
rect 21940 10170 22428 10176
rect 21638 10062 21644 10122
rect 21704 10062 21710 10122
rect 21130 9952 21136 10012
rect 21196 9952 21202 10012
rect 20620 9846 20626 9906
rect 20686 9846 20692 9906
rect 19606 9740 19612 9800
rect 19672 9740 19678 9800
rect 20104 9740 20110 9800
rect 20170 9740 20176 9800
rect 20616 9740 20622 9800
rect 20682 9740 20688 9800
rect 19612 9604 19672 9740
rect 20110 9694 20170 9740
rect 19904 9688 20392 9694
rect 19904 9654 19916 9688
rect 20380 9654 20392 9688
rect 19904 9648 20392 9654
rect 19612 9564 19622 9604
rect 19616 9028 19622 9564
rect 19656 9564 19672 9604
rect 20622 9604 20682 9740
rect 21136 9694 21196 9952
rect 20922 9688 21410 9694
rect 20922 9654 20934 9688
rect 21398 9654 21410 9688
rect 20922 9648 21410 9654
rect 19656 9028 19662 9564
rect 20622 9558 20640 9604
rect 19616 9016 19662 9028
rect 20634 9028 20640 9558
rect 20674 9558 20682 9604
rect 21644 9604 21704 10062
rect 22158 10012 22218 10170
rect 22152 9952 22158 10012
rect 22218 9952 22224 10012
rect 22158 9694 22218 9952
rect 22666 9906 22726 10260
rect 22958 10210 23446 10216
rect 22958 10176 22970 10210
rect 23434 10176 23446 10210
rect 22958 10170 23446 10176
rect 23172 10012 23232 10170
rect 23684 10122 23744 10260
rect 24706 10248 24752 10260
rect 23976 10210 24464 10216
rect 23976 10176 23988 10210
rect 24452 10176 24464 10210
rect 23976 10170 24464 10176
rect 24994 10210 25482 10216
rect 24994 10176 25006 10210
rect 25470 10176 25482 10210
rect 24994 10170 25482 10176
rect 23678 10062 23684 10122
rect 23744 10062 23750 10122
rect 23166 9952 23172 10012
rect 23232 9952 23238 10012
rect 22660 9846 22666 9906
rect 22726 9846 22732 9906
rect 23172 9694 23232 9952
rect 21940 9688 22428 9694
rect 21940 9654 21952 9688
rect 22416 9654 22428 9688
rect 21940 9648 22428 9654
rect 22958 9688 23446 9694
rect 22958 9654 22970 9688
rect 23434 9654 23446 9688
rect 22958 9648 23446 9654
rect 22670 9604 22716 9616
rect 23684 9604 23744 10062
rect 24186 10012 24246 10170
rect 25204 10012 25264 10170
rect 25716 10122 25776 10260
rect 26012 10210 26500 10216
rect 26012 10176 26024 10210
rect 26488 10176 26500 10210
rect 26012 10170 26500 10176
rect 25710 10062 25716 10122
rect 25776 10062 25782 10122
rect 24180 9952 24186 10012
rect 24246 9952 24252 10012
rect 25198 9952 25204 10012
rect 25264 9952 25270 10012
rect 24186 9694 24246 9952
rect 24690 9846 24696 9906
rect 24756 9846 24762 9906
rect 23976 9688 24464 9694
rect 23976 9654 23988 9688
rect 24452 9654 24464 9688
rect 23976 9648 24464 9654
rect 21644 9566 21658 9604
rect 20674 9028 20680 9558
rect 21652 9086 21658 9566
rect 20634 9016 20680 9028
rect 21638 9028 21658 9086
rect 21692 9566 21704 9604
rect 21692 9028 21698 9566
rect 22664 9552 22676 9604
rect 22670 9048 22676 9552
rect 19904 8978 20392 8984
rect 19904 8944 19916 8978
rect 20380 8944 20392 8978
rect 19904 8938 20392 8944
rect 20922 8978 21410 8984
rect 20922 8944 20934 8978
rect 21398 8944 21410 8978
rect 20922 8938 21410 8944
rect 19476 8850 19482 8910
rect 19542 8850 19548 8910
rect 21638 8806 21698 9028
rect 22660 9028 22676 9048
rect 22710 9552 22724 9604
rect 22710 9048 22716 9552
rect 23682 9540 23694 9604
rect 23688 9092 23694 9540
rect 22710 9028 22720 9048
rect 21940 8978 22428 8984
rect 21940 8944 21952 8978
rect 22416 8944 22428 8978
rect 21940 8938 22428 8944
rect 19600 8746 19606 8806
rect 19666 8746 19672 8806
rect 21120 8746 21126 8806
rect 21186 8746 21192 8806
rect 21632 8746 21638 8806
rect 21698 8746 21704 8806
rect 19370 8624 19376 8684
rect 19436 8624 19442 8684
rect 19258 8510 19264 8570
rect 19324 8510 19330 8570
rect 19376 7442 19436 8624
rect 19606 8370 19666 8746
rect 20106 8510 20112 8570
rect 20172 8510 20178 8570
rect 20112 8460 20172 8510
rect 21126 8460 21186 8746
rect 21638 8512 21644 8572
rect 21704 8512 21710 8572
rect 19902 8454 20390 8460
rect 19902 8420 19914 8454
rect 20378 8420 20390 8454
rect 19902 8414 20390 8420
rect 20920 8454 21408 8460
rect 20920 8420 20932 8454
rect 21396 8420 21408 8454
rect 20920 8414 21408 8420
rect 20632 8370 20678 8382
rect 21644 8370 21704 8512
rect 22142 8460 22202 8938
rect 22660 8910 22720 9028
rect 23674 9028 23694 9092
rect 23728 9570 23744 9604
rect 24696 9604 24756 9846
rect 25204 9694 25264 9952
rect 24994 9688 25482 9694
rect 24994 9654 25006 9688
rect 25470 9654 25482 9688
rect 24994 9648 25482 9654
rect 25716 9604 25776 10062
rect 26230 10012 26290 10170
rect 26736 10052 26796 10260
rect 27748 10260 27766 10336
rect 27800 10768 27810 10836
rect 28778 10836 28824 10848
rect 27800 10336 27806 10768
rect 27800 10260 27808 10336
rect 28778 10322 28784 10836
rect 28772 10320 28784 10322
rect 27030 10210 27518 10216
rect 27030 10176 27042 10210
rect 27506 10176 27518 10210
rect 27030 10170 27518 10176
rect 26224 9952 26230 10012
rect 26290 9952 26296 10012
rect 26736 9992 26962 10052
rect 27250 10012 27310 10170
rect 27748 10122 27808 10260
rect 28770 10260 28784 10320
rect 28818 10322 28824 10836
rect 29790 10836 29850 11226
rect 30292 11160 30352 11166
rect 30292 10926 30352 11100
rect 31300 11160 31360 11166
rect 31360 11100 31362 11106
rect 31300 11094 31362 11100
rect 31302 10926 31362 11094
rect 30084 10920 30572 10926
rect 30084 10886 30096 10920
rect 30560 10886 30572 10920
rect 30084 10880 30572 10886
rect 31102 10920 31590 10926
rect 31102 10886 31114 10920
rect 31578 10886 31590 10920
rect 31102 10880 31590 10886
rect 30814 10836 30860 10848
rect 31822 10836 31882 11226
rect 32316 11160 32376 11166
rect 33340 11160 33400 11166
rect 32376 11100 32378 11106
rect 32316 11094 32378 11100
rect 32318 10926 32378 11094
rect 33340 10926 33400 11100
rect 32120 10920 32608 10926
rect 32120 10886 32132 10920
rect 32596 10886 32608 10920
rect 32120 10880 32608 10886
rect 33138 10920 33626 10926
rect 33138 10886 33150 10920
rect 33614 10886 33626 10920
rect 33138 10880 33626 10886
rect 32850 10836 32896 10848
rect 33862 10836 33922 11226
rect 34362 11160 34422 11166
rect 35384 11160 35444 11166
rect 34362 10926 34422 11100
rect 35382 11100 35384 11106
rect 35382 11094 35444 11100
rect 34878 10984 34884 11044
rect 34944 10984 34950 11044
rect 34156 10920 34644 10926
rect 34156 10886 34168 10920
rect 34632 10886 34644 10920
rect 34156 10880 34644 10886
rect 29790 10768 29802 10836
rect 29796 10326 29802 10768
rect 28818 10260 28832 10322
rect 29784 10260 29802 10326
rect 29836 10768 29850 10836
rect 30804 10802 30820 10836
rect 29836 10326 29842 10768
rect 29836 10260 29844 10326
rect 30814 10308 30820 10802
rect 28048 10210 28536 10216
rect 28048 10176 28060 10210
rect 28524 10176 28536 10210
rect 28048 10170 28536 10176
rect 27742 10062 27748 10122
rect 27808 10062 27814 10122
rect 26230 9694 26290 9952
rect 26730 9846 26736 9906
rect 26796 9846 26802 9906
rect 26012 9688 26500 9694
rect 26012 9654 26024 9688
rect 26488 9654 26500 9688
rect 26012 9648 26500 9654
rect 26736 9604 26796 9846
rect 26902 9800 26962 9992
rect 27244 9952 27250 10012
rect 27310 9952 27316 10012
rect 26896 9740 26902 9800
rect 26962 9740 26968 9800
rect 27250 9694 27310 9952
rect 27030 9688 27518 9694
rect 27030 9654 27042 9688
rect 27506 9654 27518 9688
rect 27030 9648 27518 9654
rect 23728 9540 23742 9570
rect 24696 9560 24712 9604
rect 23728 9028 23734 9540
rect 22958 8978 23446 8984
rect 22958 8944 22970 8978
rect 23434 8944 23446 8978
rect 22958 8938 23446 8944
rect 22654 8850 22660 8910
rect 22720 8850 22726 8910
rect 22656 8746 22662 8806
rect 22722 8746 22728 8806
rect 21938 8454 22426 8460
rect 21938 8420 21950 8454
rect 22414 8420 22426 8454
rect 21938 8414 22426 8420
rect 19606 8314 19620 8370
rect 19614 7794 19620 8314
rect 19654 8314 19666 8370
rect 20626 8338 20638 8370
rect 19654 7794 19660 8314
rect 20632 7838 20638 8338
rect 19614 7782 19660 7794
rect 20626 7794 20638 7838
rect 20672 8338 20686 8370
rect 21644 8344 21656 8370
rect 20672 7838 20678 8338
rect 20672 7794 20686 7838
rect 19902 7744 20390 7750
rect 19902 7710 19914 7744
rect 20378 7710 20390 7744
rect 19902 7704 20390 7710
rect 20626 7642 20686 7794
rect 21650 7794 21656 8344
rect 21690 8344 21704 8370
rect 22662 8370 22722 8746
rect 23162 8460 23222 8938
rect 23674 8806 23734 9028
rect 24706 9028 24712 9560
rect 24746 9570 24758 9604
rect 24746 9560 24756 9570
rect 25716 9562 25730 9604
rect 24746 9028 24752 9560
rect 25724 9070 25730 9562
rect 25716 9028 25730 9070
rect 25764 9562 25776 9604
rect 25764 9070 25770 9562
rect 26732 9542 26748 9604
rect 25764 9028 25776 9070
rect 26742 9028 26748 9542
rect 26782 9564 26796 9604
rect 27748 9604 27808 10062
rect 28270 10012 28330 10170
rect 28264 9952 28270 10012
rect 28330 9952 28336 10012
rect 28270 9694 28330 9952
rect 28770 9906 28830 10260
rect 29066 10210 29554 10216
rect 29066 10176 29078 10210
rect 29542 10176 29554 10210
rect 29066 10170 29554 10176
rect 29272 10012 29332 10170
rect 29784 10122 29844 10260
rect 30806 10260 30820 10308
rect 30854 10802 30864 10836
rect 30854 10308 30860 10802
rect 31822 10782 31838 10836
rect 31832 10320 31838 10782
rect 30854 10260 30866 10308
rect 30084 10210 30572 10216
rect 30084 10176 30096 10210
rect 30560 10176 30572 10210
rect 30084 10170 30572 10176
rect 29778 10062 29784 10122
rect 29844 10062 29850 10122
rect 29266 9952 29272 10012
rect 29332 9952 29338 10012
rect 28764 9846 28770 9906
rect 28830 9846 28836 9906
rect 28764 9740 28770 9800
rect 28830 9740 28836 9800
rect 28048 9688 28536 9694
rect 28048 9654 28060 9688
rect 28524 9654 28536 9688
rect 28048 9648 28536 9654
rect 28770 9604 28830 9740
rect 29272 9694 29332 9952
rect 29066 9688 29554 9694
rect 29066 9654 29078 9688
rect 29542 9654 29554 9688
rect 29066 9648 29554 9654
rect 29784 9604 29844 10062
rect 30298 10012 30358 10170
rect 30292 9952 30298 10012
rect 30358 9952 30364 10012
rect 30298 9694 30358 9952
rect 30806 9906 30866 10260
rect 31820 10260 31838 10320
rect 31872 10782 31882 10836
rect 32842 10796 32856 10836
rect 31872 10320 31878 10782
rect 32850 10326 32856 10796
rect 31872 10260 31880 10320
rect 32846 10300 32856 10326
rect 31102 10210 31590 10216
rect 31102 10176 31114 10210
rect 31578 10176 31590 10210
rect 31102 10170 31590 10176
rect 31316 10012 31376 10170
rect 31820 10122 31880 10260
rect 32844 10260 32856 10300
rect 32890 10796 32902 10836
rect 32890 10326 32896 10796
rect 33862 10782 33874 10836
rect 32890 10260 32906 10326
rect 33868 10310 33874 10782
rect 33858 10260 33874 10310
rect 33908 10782 33922 10836
rect 34884 10836 34944 10984
rect 35382 10926 35442 11094
rect 35174 10920 35662 10926
rect 35174 10886 35186 10920
rect 35650 10886 35662 10920
rect 35174 10880 35662 10886
rect 33908 10310 33914 10782
rect 34884 10772 34892 10836
rect 34886 10316 34892 10772
rect 33908 10260 33918 10310
rect 34878 10260 34892 10316
rect 34926 10772 34944 10836
rect 35898 10836 35958 11226
rect 36402 11160 36462 11166
rect 37416 11160 37476 11166
rect 36462 11100 36464 11106
rect 36402 11094 36464 11100
rect 37476 11100 37478 11106
rect 37416 11094 37478 11100
rect 36404 10926 36464 11094
rect 37418 10926 37478 11094
rect 36192 10920 36680 10926
rect 36192 10886 36204 10920
rect 36668 10886 36680 10920
rect 36192 10880 36680 10886
rect 37210 10920 37698 10926
rect 37210 10886 37222 10920
rect 37686 10886 37698 10920
rect 37210 10880 37698 10886
rect 36922 10836 36968 10848
rect 37932 10836 37992 11226
rect 38440 11160 38500 11166
rect 38438 11100 38440 11106
rect 38438 11094 38500 11100
rect 38438 10926 38498 11094
rect 38950 10984 38956 11044
rect 39016 10984 39022 11044
rect 40082 10984 40088 11044
rect 40148 10984 40154 11044
rect 38228 10920 38716 10926
rect 38228 10886 38240 10920
rect 38704 10886 38716 10920
rect 38228 10880 38716 10886
rect 38956 10836 39016 10984
rect 39246 10920 39734 10926
rect 39246 10886 39258 10920
rect 39722 10886 39734 10920
rect 39246 10880 39734 10886
rect 35898 10776 35910 10836
rect 34926 10316 34932 10772
rect 34926 10314 34938 10316
rect 34926 10260 34940 10314
rect 35904 10296 35910 10776
rect 35896 10260 35910 10296
rect 35944 10776 35958 10836
rect 36914 10796 36928 10836
rect 35944 10296 35950 10776
rect 36922 10316 36928 10796
rect 35944 10260 35956 10296
rect 32120 10210 32608 10216
rect 32120 10176 32132 10210
rect 32596 10176 32608 10210
rect 32120 10170 32608 10176
rect 31814 10062 31820 10122
rect 31880 10062 31886 10122
rect 31310 9952 31316 10012
rect 31376 9952 31382 10012
rect 30800 9846 30806 9906
rect 30866 9846 30872 9906
rect 30802 9740 30808 9800
rect 30868 9740 30874 9800
rect 30084 9688 30572 9694
rect 30084 9654 30096 9688
rect 30560 9654 30572 9688
rect 30084 9648 30572 9654
rect 30808 9604 30868 9740
rect 31316 9694 31376 9952
rect 31102 9688 31590 9694
rect 31102 9654 31114 9688
rect 31578 9654 31590 9688
rect 31102 9648 31590 9654
rect 31820 9604 31880 10062
rect 32324 10012 32384 10170
rect 32844 10044 32904 10260
rect 33336 10216 33396 10218
rect 33138 10210 33626 10216
rect 33138 10176 33150 10210
rect 33614 10176 33626 10210
rect 33138 10170 33626 10176
rect 32318 9952 32324 10012
rect 32384 9952 32390 10012
rect 32688 9984 32904 10044
rect 33336 10012 33396 10170
rect 33858 10122 33918 10260
rect 34886 10248 34932 10260
rect 34368 10216 34428 10218
rect 34156 10210 34644 10216
rect 34156 10176 34168 10210
rect 34632 10176 34644 10210
rect 34156 10170 34644 10176
rect 35174 10210 35662 10216
rect 35174 10176 35186 10210
rect 35650 10176 35662 10210
rect 35174 10170 35662 10176
rect 33852 10062 33858 10122
rect 33918 10062 33924 10122
rect 32324 9694 32384 9952
rect 32688 9800 32748 9984
rect 33330 9952 33336 10012
rect 33396 9952 33402 10012
rect 32836 9846 32842 9906
rect 32902 9846 32908 9906
rect 32682 9740 32688 9800
rect 32748 9740 32754 9800
rect 32120 9688 32608 9694
rect 32120 9654 32132 9688
rect 32596 9654 32608 9688
rect 32120 9648 32608 9654
rect 26782 9542 26792 9564
rect 27748 9548 27766 9604
rect 26782 9028 26788 9542
rect 27760 9070 27766 9548
rect 24706 9016 24752 9028
rect 25724 9016 25770 9028
rect 26742 9016 26788 9028
rect 27752 9028 27766 9070
rect 27800 9548 27808 9604
rect 28768 9552 28784 9604
rect 27800 9070 27806 9548
rect 27800 9028 27812 9070
rect 23976 8978 24464 8984
rect 23976 8944 23988 8978
rect 24452 8944 24464 8978
rect 23976 8938 24464 8944
rect 24994 8978 25482 8984
rect 24994 8944 25006 8978
rect 25470 8944 25482 8978
rect 24994 8938 25482 8944
rect 26012 8978 26500 8984
rect 26012 8944 26024 8978
rect 26488 8944 26500 8978
rect 26012 8938 26500 8944
rect 27030 8978 27518 8984
rect 27030 8944 27042 8978
rect 27506 8944 27518 8978
rect 27030 8938 27518 8944
rect 23668 8746 23674 8806
rect 23734 8746 23740 8806
rect 23674 8512 23680 8572
rect 23740 8512 23746 8572
rect 22956 8454 23444 8460
rect 22956 8420 22968 8454
rect 23432 8420 23444 8454
rect 22956 8414 23444 8420
rect 21690 7794 21696 8344
rect 22662 8338 22674 8370
rect 22668 7834 22674 8338
rect 21650 7782 21696 7794
rect 22660 7794 22674 7834
rect 22708 8338 22722 8370
rect 23680 8370 23740 8512
rect 24174 8460 24234 8938
rect 24688 8746 24694 8806
rect 24754 8746 24760 8806
rect 23974 8454 24462 8460
rect 23974 8420 23986 8454
rect 24450 8420 24462 8454
rect 23974 8414 24462 8420
rect 23680 8340 23692 8370
rect 22708 7834 22714 8338
rect 22708 7794 22720 7834
rect 20920 7744 21408 7750
rect 20920 7710 20932 7744
rect 21396 7710 21408 7744
rect 20920 7704 21408 7710
rect 21938 7744 22426 7750
rect 21938 7710 21950 7744
rect 22414 7710 22426 7744
rect 21938 7704 22426 7710
rect 19482 7582 19488 7642
rect 19548 7582 19554 7642
rect 20620 7582 20626 7642
rect 20686 7582 20692 7642
rect 19370 7382 19376 7442
rect 19436 7382 19442 7442
rect 19264 7280 19270 7340
rect 19330 7280 19336 7340
rect 19154 3828 19160 3888
rect 19220 3828 19226 3888
rect 19270 3850 19330 7280
rect 19376 6206 19436 7382
rect 19370 6146 19376 6206
rect 19436 6146 19442 6206
rect 18922 3678 18928 3738
rect 18988 3678 18994 3738
rect 19160 152 19220 3828
rect 19264 3790 19270 3850
rect 19330 3790 19336 3850
rect 19270 1360 19330 3790
rect 19376 1486 19436 6146
rect 19488 4868 19548 7582
rect 20618 7382 20624 7442
rect 20684 7382 20690 7442
rect 20624 7338 20684 7382
rect 19608 7278 20684 7338
rect 19608 7276 20172 7278
rect 19608 7136 19668 7276
rect 20112 7226 20172 7276
rect 19902 7220 20390 7226
rect 19902 7186 19914 7220
rect 20378 7186 20390 7220
rect 19902 7180 20390 7186
rect 19608 7104 19620 7136
rect 19614 6560 19620 7104
rect 19654 7104 19668 7136
rect 20624 7136 20684 7278
rect 21128 7226 21188 7704
rect 21636 7502 21642 7562
rect 21702 7502 21708 7562
rect 20920 7220 21408 7226
rect 20920 7186 20932 7220
rect 21396 7186 21408 7220
rect 20920 7180 21408 7186
rect 19654 6560 19660 7104
rect 20624 7100 20638 7136
rect 19614 6548 19660 6560
rect 20632 6560 20638 7100
rect 20672 7100 20684 7136
rect 21642 7136 21702 7502
rect 22156 7448 22216 7704
rect 22660 7666 22720 7794
rect 23686 7794 23692 8340
rect 23726 8340 23740 8370
rect 24694 8370 24754 8746
rect 25200 8460 25260 8938
rect 25710 8850 25716 8910
rect 25776 8850 25782 8910
rect 24992 8454 25480 8460
rect 24992 8420 25004 8454
rect 25468 8420 25480 8454
rect 24992 8414 25480 8420
rect 23726 7794 23732 8340
rect 24694 8326 24710 8370
rect 24704 7844 24710 8326
rect 23686 7782 23732 7794
rect 24696 7794 24710 7844
rect 24744 8326 24754 8370
rect 25716 8370 25776 8850
rect 27752 8806 27812 9028
rect 28778 9028 28784 9552
rect 28818 9560 28832 9604
rect 28818 9552 28828 9560
rect 29784 9556 29802 9604
rect 28818 9028 28824 9552
rect 29796 9076 29802 9556
rect 28778 9016 28824 9028
rect 29790 9028 29802 9076
rect 29836 9556 29844 9604
rect 30804 9564 30820 9604
rect 29836 9076 29842 9556
rect 29836 9028 29850 9076
rect 28048 8978 28536 8984
rect 28048 8944 28060 8978
rect 28524 8944 28536 8978
rect 28048 8938 28536 8944
rect 29066 8978 29554 8984
rect 29066 8944 29078 8978
rect 29542 8944 29554 8978
rect 29066 8938 29554 8944
rect 29790 8806 29850 9028
rect 30814 9028 30820 9564
rect 30854 9566 30870 9604
rect 30854 9564 30868 9566
rect 30854 9028 30860 9564
rect 31820 9558 31838 9604
rect 31832 9082 31838 9558
rect 31820 9028 31838 9082
rect 31872 9558 31880 9604
rect 32842 9604 32902 9846
rect 33336 9694 33396 9952
rect 33138 9688 33626 9694
rect 33138 9654 33150 9688
rect 33614 9654 33626 9688
rect 33138 9648 33626 9654
rect 33858 9604 33918 10062
rect 34368 10012 34428 10170
rect 35382 10012 35442 10170
rect 35896 10122 35956 10260
rect 36912 10260 36928 10316
rect 36962 10796 36974 10836
rect 36962 10316 36968 10796
rect 36962 10260 36972 10316
rect 36192 10210 36680 10216
rect 36192 10176 36204 10210
rect 36668 10176 36680 10210
rect 36192 10170 36680 10176
rect 35890 10062 35896 10122
rect 35956 10062 35962 10122
rect 34362 9952 34368 10012
rect 34428 9952 34434 10012
rect 35376 9952 35382 10012
rect 35442 9952 35448 10012
rect 34368 9694 34428 9952
rect 34876 9846 34882 9906
rect 34942 9846 34948 9906
rect 34156 9688 34644 9694
rect 34156 9654 34168 9688
rect 34632 9654 34644 9688
rect 34156 9648 34644 9654
rect 34882 9604 34942 9846
rect 35382 9694 35442 9952
rect 35174 9688 35662 9694
rect 35174 9654 35186 9688
rect 35650 9654 35662 9688
rect 35174 9648 35662 9654
rect 31872 9082 31878 9558
rect 32842 9552 32856 9604
rect 31872 9028 31880 9082
rect 32850 9028 32856 9552
rect 32890 9562 32906 9604
rect 32890 9552 32902 9562
rect 32890 9028 32896 9552
rect 30814 9016 30860 9028
rect 31832 9016 31878 9028
rect 32850 9016 32896 9028
rect 33858 9028 33874 9604
rect 33908 9028 33918 9604
rect 34878 9562 34892 9604
rect 34882 9542 34892 9562
rect 30084 8978 30572 8984
rect 30084 8944 30096 8978
rect 30560 8944 30572 8978
rect 30084 8938 30572 8944
rect 31102 8978 31590 8984
rect 31102 8944 31114 8978
rect 31578 8944 31590 8978
rect 31102 8938 31590 8944
rect 32120 8978 32608 8984
rect 32120 8944 32132 8978
rect 32596 8944 32608 8978
rect 32120 8938 32608 8944
rect 33138 8978 33626 8984
rect 33138 8944 33150 8978
rect 33614 8944 33626 8978
rect 33138 8938 33626 8944
rect 31816 8850 31822 8910
rect 31882 8850 31888 8910
rect 27746 8746 27752 8806
rect 27812 8746 27818 8806
rect 29784 8746 29790 8806
rect 29850 8746 29856 8806
rect 26730 8624 26736 8684
rect 26796 8624 26802 8684
rect 28764 8624 28770 8684
rect 28830 8624 28836 8684
rect 30794 8624 30800 8684
rect 30860 8624 30866 8684
rect 26010 8454 26498 8460
rect 26010 8420 26022 8454
rect 26486 8420 26498 8454
rect 26010 8414 26498 8420
rect 24744 7844 24750 8326
rect 25716 8308 25728 8370
rect 24744 7794 24756 7844
rect 25722 7830 25728 8308
rect 22956 7744 23444 7750
rect 22956 7710 22968 7744
rect 23432 7710 23444 7744
rect 22956 7704 23444 7710
rect 23974 7744 24462 7750
rect 23974 7710 23986 7744
rect 24450 7710 24462 7744
rect 23974 7704 24462 7710
rect 22654 7606 22660 7666
rect 22720 7606 22726 7666
rect 22150 7388 22156 7448
rect 22216 7388 22222 7448
rect 22156 7226 22216 7388
rect 21938 7220 22426 7226
rect 21938 7186 21950 7220
rect 22414 7186 22426 7220
rect 21938 7180 22426 7186
rect 20672 6560 20678 7100
rect 21642 7094 21656 7136
rect 21650 6618 21656 7094
rect 20632 6548 20678 6560
rect 21644 6560 21656 6618
rect 21690 7094 21702 7136
rect 22660 7136 22720 7606
rect 23158 7454 23218 7704
rect 23676 7502 23682 7562
rect 23742 7502 23748 7562
rect 23158 7448 23220 7454
rect 23158 7388 23160 7448
rect 23158 7382 23220 7388
rect 23158 7226 23218 7382
rect 22956 7220 23444 7226
rect 22956 7186 22968 7220
rect 23432 7186 23444 7220
rect 22956 7180 23444 7186
rect 21690 6618 21696 7094
rect 22660 7092 22674 7136
rect 21690 6560 21704 6618
rect 22668 6608 22674 7092
rect 19902 6510 20390 6516
rect 19902 6476 19914 6510
rect 20378 6476 20390 6510
rect 19902 6470 20390 6476
rect 20920 6510 21408 6516
rect 20920 6476 20932 6510
rect 21396 6476 21408 6510
rect 20920 6470 21408 6476
rect 20618 6350 20624 6410
rect 20684 6350 20690 6410
rect 19902 5988 20390 5994
rect 19902 5954 19914 5988
rect 20378 5954 20390 5988
rect 19902 5948 20390 5954
rect 19614 5904 19660 5916
rect 19614 5374 19620 5904
rect 19604 5328 19620 5374
rect 19654 5374 19660 5904
rect 20624 5904 20684 6350
rect 21130 6308 21190 6470
rect 21124 6248 21130 6308
rect 21190 6248 21196 6308
rect 21644 6106 21704 6560
rect 22662 6560 22674 6608
rect 22708 7092 22720 7136
rect 23682 7136 23742 7502
rect 24174 7454 24234 7704
rect 24696 7666 24756 7794
rect 25714 7794 25728 7830
rect 25762 8308 25776 8370
rect 26736 8370 26796 8624
rect 27028 8454 27516 8460
rect 27028 8420 27040 8454
rect 27504 8420 27516 8454
rect 27028 8414 27516 8420
rect 28046 8454 28534 8460
rect 28046 8420 28058 8454
rect 28522 8420 28534 8454
rect 28046 8414 28534 8420
rect 26736 8314 26746 8370
rect 25762 7830 25768 8308
rect 25762 7794 25774 7830
rect 24992 7744 25480 7750
rect 24992 7710 25004 7744
rect 25468 7710 25480 7744
rect 24992 7704 25480 7710
rect 24690 7606 24696 7666
rect 24756 7606 24762 7666
rect 24172 7448 24234 7454
rect 24232 7388 24234 7448
rect 24172 7382 24234 7388
rect 24174 7226 24234 7382
rect 23974 7220 24462 7226
rect 23974 7186 23986 7220
rect 24450 7186 24462 7220
rect 23974 7180 24462 7186
rect 23682 7094 23692 7136
rect 22708 6608 22714 7092
rect 22708 6560 22722 6608
rect 21938 6510 22426 6516
rect 21938 6476 21950 6510
rect 22414 6476 22426 6510
rect 21938 6470 22426 6476
rect 22662 6410 22722 6560
rect 23686 6560 23692 7094
rect 23726 7094 23742 7136
rect 24696 7136 24756 7606
rect 25192 7448 25252 7704
rect 25714 7562 25774 7794
rect 26740 7794 26746 8314
rect 26780 8314 26796 8370
rect 27758 8370 27804 8382
rect 26780 7794 26786 8314
rect 27758 7824 27764 8370
rect 26740 7782 26786 7794
rect 27748 7794 27764 7824
rect 27798 7824 27804 8370
rect 28770 8370 28830 8624
rect 29064 8454 29552 8460
rect 29064 8420 29076 8454
rect 29540 8420 29552 8454
rect 29064 8414 29552 8420
rect 30082 8454 30570 8460
rect 30082 8420 30094 8454
rect 30558 8420 30570 8454
rect 30082 8414 30570 8420
rect 28770 8320 28782 8370
rect 27798 7794 27808 7824
rect 26010 7744 26498 7750
rect 26010 7710 26022 7744
rect 26486 7710 26498 7744
rect 26010 7704 26498 7710
rect 27028 7744 27516 7750
rect 27028 7710 27040 7744
rect 27504 7710 27516 7744
rect 27028 7704 27516 7710
rect 25708 7502 25714 7562
rect 25774 7502 25780 7562
rect 26204 7506 26264 7704
rect 27246 7506 27306 7704
rect 27748 7562 27808 7794
rect 28776 7794 28782 8320
rect 28816 8320 28830 8370
rect 29794 8370 29840 8382
rect 28816 7794 28822 8320
rect 29794 7836 29800 8370
rect 28776 7782 28822 7794
rect 29788 7794 29800 7836
rect 29834 7836 29840 8370
rect 30800 8370 30860 8624
rect 31100 8454 31588 8460
rect 31100 8420 31112 8454
rect 31576 8420 31588 8454
rect 31100 8414 31588 8420
rect 30800 8326 30818 8370
rect 29834 7794 29848 7836
rect 28046 7744 28534 7750
rect 28046 7710 28058 7744
rect 28522 7710 28534 7744
rect 28046 7704 28534 7710
rect 29064 7744 29552 7750
rect 29064 7710 29076 7744
rect 29540 7710 29552 7744
rect 29064 7704 29552 7710
rect 25708 7390 25714 7450
rect 25774 7390 25780 7450
rect 26204 7446 27306 7506
rect 27742 7502 27748 7562
rect 27808 7502 27814 7562
rect 25192 7226 25252 7388
rect 24992 7220 25480 7226
rect 24992 7186 25004 7220
rect 25468 7186 25480 7220
rect 24992 7180 25480 7186
rect 23726 6560 23732 7094
rect 24696 7088 24710 7136
rect 24704 6610 24710 7088
rect 23686 6548 23732 6560
rect 24698 6560 24710 6610
rect 24744 7088 24756 7136
rect 25714 7136 25774 7390
rect 26204 7226 26264 7446
rect 26726 7280 26732 7340
rect 26792 7280 26798 7340
rect 26010 7220 26498 7226
rect 26010 7186 26022 7220
rect 26486 7186 26498 7220
rect 26010 7180 26498 7186
rect 24744 6610 24750 7088
rect 25714 7078 25728 7136
rect 24744 6560 24758 6610
rect 22956 6510 23444 6516
rect 22956 6476 22968 6510
rect 23432 6476 23444 6510
rect 22956 6470 23444 6476
rect 23974 6510 24462 6516
rect 23974 6476 23986 6510
rect 24450 6476 24462 6510
rect 23974 6470 24462 6476
rect 22656 6350 22662 6410
rect 22722 6350 22728 6410
rect 22654 6146 22660 6206
rect 22720 6146 22726 6206
rect 23168 6200 23228 6470
rect 24190 6200 24250 6470
rect 24698 6410 24758 6560
rect 25722 6560 25728 7078
rect 25762 7078 25774 7136
rect 26732 7136 26792 7280
rect 27246 7226 27306 7446
rect 27744 7390 27750 7450
rect 27810 7390 27816 7450
rect 27028 7220 27516 7226
rect 27028 7186 27040 7220
rect 27504 7186 27516 7220
rect 27028 7180 27516 7186
rect 26732 7090 26746 7136
rect 25762 6560 25768 7078
rect 25722 6548 25768 6560
rect 26740 6560 26746 7090
rect 26780 7090 26792 7136
rect 27750 7136 27810 7390
rect 28246 7226 28306 7704
rect 28760 7280 28766 7340
rect 28826 7280 28832 7340
rect 28046 7220 28534 7226
rect 28046 7186 28058 7220
rect 28522 7186 28534 7220
rect 28046 7180 28534 7186
rect 26780 6560 26786 7090
rect 27750 7068 27764 7136
rect 26740 6548 26786 6560
rect 27758 6560 27764 7068
rect 27798 7068 27810 7136
rect 28766 7136 28826 7280
rect 29280 7226 29340 7704
rect 29788 7562 29848 7794
rect 30812 7794 30818 8326
rect 30852 8326 30860 8370
rect 31822 8370 31882 8850
rect 32344 8460 32404 8938
rect 32834 8746 32840 8806
rect 32900 8746 32906 8806
rect 32118 8454 32606 8460
rect 32118 8420 32130 8454
rect 32594 8420 32606 8454
rect 32118 8414 32606 8420
rect 30852 7794 30858 8326
rect 31822 8318 31836 8370
rect 31830 7846 31836 8318
rect 30812 7782 30858 7794
rect 31822 7794 31836 7846
rect 31870 8318 31882 8370
rect 32840 8370 32900 8746
rect 33346 8460 33406 8938
rect 33858 8806 33918 9028
rect 34886 9028 34892 9542
rect 34926 9542 34942 9604
rect 35896 9604 35956 10062
rect 36400 10012 36460 10170
rect 36394 9952 36400 10012
rect 36460 9952 36466 10012
rect 36400 9694 36460 9952
rect 36912 9906 36972 10260
rect 37932 10260 37946 10836
rect 37980 10804 37994 10836
rect 38952 10808 38964 10836
rect 37980 10260 37992 10804
rect 38956 10772 38964 10808
rect 38958 10320 38964 10772
rect 37210 10210 37698 10216
rect 37210 10176 37222 10210
rect 37686 10176 37698 10210
rect 37210 10170 37698 10176
rect 37424 10012 37484 10170
rect 37932 10122 37992 10260
rect 38952 10260 38964 10320
rect 38998 10772 39016 10836
rect 39976 10836 40022 10848
rect 38998 10320 39004 10772
rect 38998 10260 39012 10320
rect 39976 10308 39982 10836
rect 38228 10210 38716 10216
rect 38228 10176 38240 10210
rect 38704 10176 38716 10210
rect 38228 10170 38716 10176
rect 37926 10062 37932 10122
rect 37992 10062 37998 10122
rect 37418 9952 37424 10012
rect 37484 9952 37490 10012
rect 36906 9846 36912 9906
rect 36972 9846 36978 9906
rect 36906 9742 36912 9802
rect 36972 9742 36978 9802
rect 36192 9688 36680 9694
rect 36192 9654 36204 9688
rect 36668 9654 36680 9688
rect 36192 9648 36680 9654
rect 36392 9636 36452 9648
rect 36912 9604 36972 9742
rect 37424 9694 37484 9952
rect 37210 9688 37698 9694
rect 37210 9654 37222 9688
rect 37686 9654 37698 9688
rect 37210 9648 37698 9654
rect 35896 9546 35910 9604
rect 34926 9028 34932 9542
rect 35904 9076 35910 9546
rect 34886 9016 34932 9028
rect 35894 9028 35910 9076
rect 35944 9546 35956 9604
rect 36910 9558 36928 9604
rect 35944 9076 35950 9546
rect 36912 9530 36928 9558
rect 36922 9082 36928 9530
rect 35944 9028 35954 9076
rect 34156 8978 34644 8984
rect 34156 8944 34168 8978
rect 34632 8944 34644 8978
rect 34156 8938 34644 8944
rect 35174 8978 35662 8984
rect 35174 8944 35186 8978
rect 35650 8944 35662 8978
rect 35174 8938 35662 8944
rect 33852 8746 33858 8806
rect 33918 8746 33924 8806
rect 34358 8460 34418 8938
rect 34872 8746 34878 8806
rect 34938 8746 34944 8806
rect 33136 8454 33624 8460
rect 33136 8420 33148 8454
rect 33612 8420 33624 8454
rect 33136 8414 33624 8420
rect 34154 8454 34642 8460
rect 34154 8420 34166 8454
rect 34630 8420 34642 8454
rect 34154 8414 34642 8420
rect 32840 8322 32854 8370
rect 31870 7846 31876 8318
rect 31870 7794 31882 7846
rect 32848 7826 32854 8322
rect 30082 7744 30570 7750
rect 30082 7710 30094 7744
rect 30558 7710 30570 7744
rect 30082 7704 30570 7710
rect 31100 7744 31588 7750
rect 31100 7710 31112 7744
rect 31576 7710 31588 7744
rect 31100 7704 31588 7710
rect 29782 7502 29788 7562
rect 29848 7502 29854 7562
rect 30302 7506 30362 7704
rect 31310 7506 31370 7704
rect 31822 7562 31882 7794
rect 32840 7794 32854 7826
rect 32888 8322 32900 8370
rect 33866 8370 33912 8382
rect 32888 7826 32894 8322
rect 33866 7830 33872 8370
rect 32888 7794 32900 7826
rect 32118 7744 32606 7750
rect 32118 7710 32130 7744
rect 32594 7710 32606 7744
rect 32118 7704 32606 7710
rect 29780 7390 29786 7450
rect 29846 7390 29852 7450
rect 30302 7446 31370 7506
rect 31816 7502 31822 7562
rect 31882 7502 31888 7562
rect 32012 7498 32018 7558
rect 32078 7498 32084 7558
rect 29064 7220 29552 7226
rect 29064 7186 29076 7220
rect 29540 7186 29552 7220
rect 29064 7180 29552 7186
rect 28766 7088 28782 7136
rect 27798 6560 27804 7068
rect 27758 6548 27804 6560
rect 28776 6560 28782 7088
rect 28816 7088 28826 7136
rect 29786 7136 29846 7390
rect 30302 7226 30362 7446
rect 30800 7280 30806 7340
rect 30866 7280 30872 7340
rect 30082 7220 30570 7226
rect 30082 7186 30094 7220
rect 30558 7186 30570 7220
rect 30082 7180 30570 7186
rect 28816 6560 28822 7088
rect 29786 7086 29800 7136
rect 28776 6548 28822 6560
rect 29794 6560 29800 7086
rect 29834 7086 29846 7136
rect 30806 7136 30866 7280
rect 31310 7226 31370 7446
rect 31816 7390 31822 7450
rect 31882 7390 31888 7450
rect 31100 7220 31588 7226
rect 31100 7186 31112 7220
rect 31576 7186 31588 7220
rect 31100 7180 31588 7186
rect 30806 7098 30818 7136
rect 29834 6560 29840 7086
rect 30812 6606 30818 7098
rect 29794 6548 29840 6560
rect 30806 6560 30818 6606
rect 30852 7098 30866 7136
rect 31822 7136 31882 7390
rect 32018 7340 32078 7498
rect 32312 7342 32372 7704
rect 32840 7666 32900 7794
rect 33856 7794 33872 7830
rect 33906 7830 33912 8370
rect 34878 8370 34938 8746
rect 35392 8460 35452 8938
rect 35894 8806 35954 9028
rect 36916 9028 36928 9082
rect 36962 9530 36972 9604
rect 37932 9604 37992 10062
rect 38444 10012 38504 10170
rect 38952 10112 39012 10260
rect 39968 10260 39982 10308
rect 40016 10308 40022 10836
rect 40016 10260 40028 10308
rect 39246 10210 39734 10216
rect 39246 10176 39258 10210
rect 39722 10176 39734 10210
rect 39246 10170 39734 10176
rect 39462 10112 39522 10170
rect 39968 10112 40028 10260
rect 40088 10112 40148 10984
rect 38952 10052 40148 10112
rect 38438 9952 38444 10012
rect 38504 9952 38510 10012
rect 38444 9694 38504 9952
rect 38946 9846 38952 9906
rect 39012 9846 39018 9906
rect 38952 9804 39012 9846
rect 38952 9744 40030 9804
rect 40088 9802 40148 10052
rect 38228 9688 38716 9694
rect 38228 9654 38240 9688
rect 38704 9654 38716 9688
rect 38228 9648 38716 9654
rect 37932 9578 37946 9604
rect 36962 9082 36968 9530
rect 37940 9086 37946 9578
rect 36962 9028 36976 9082
rect 36192 8978 36680 8984
rect 36192 8944 36204 8978
rect 36668 8944 36680 8978
rect 36192 8938 36680 8944
rect 36916 8910 36976 9028
rect 37930 9028 37946 9086
rect 37980 9578 37992 9604
rect 38952 9604 39012 9744
rect 39438 9694 39498 9744
rect 39246 9688 39734 9694
rect 39246 9654 39258 9688
rect 39722 9654 39734 9688
rect 39246 9648 39734 9654
rect 39970 9604 40030 9744
rect 40082 9742 40088 9802
rect 40148 9742 40154 9802
rect 37980 9086 37986 9578
rect 38952 9548 38964 9604
rect 37980 9028 37990 9086
rect 37210 8978 37698 8984
rect 37210 8944 37222 8978
rect 37686 8944 37698 8978
rect 37210 8938 37698 8944
rect 36910 8850 36916 8910
rect 36976 8850 36982 8910
rect 37930 8806 37990 9028
rect 38958 9028 38964 9548
rect 38998 9548 39012 9604
rect 39966 9568 39982 9604
rect 39970 9562 39982 9568
rect 38998 9028 39004 9548
rect 39976 9072 39982 9562
rect 38958 9016 39004 9028
rect 39972 9028 39982 9072
rect 40016 9562 40030 9604
rect 40016 9072 40022 9562
rect 40016 9028 40032 9072
rect 38228 8978 38716 8984
rect 38228 8944 38240 8978
rect 38704 8944 38716 8978
rect 38228 8938 38716 8944
rect 39246 8978 39734 8984
rect 39246 8944 39258 8978
rect 39722 8944 39734 8978
rect 39246 8938 39734 8944
rect 35888 8746 35894 8806
rect 35954 8746 35960 8806
rect 37924 8746 37930 8806
rect 37990 8746 37996 8806
rect 38420 8460 38480 8938
rect 39972 8902 40032 9028
rect 39972 8842 40262 8902
rect 39458 8536 40026 8596
rect 39458 8460 39518 8536
rect 35172 8454 35660 8460
rect 35172 8420 35184 8454
rect 35648 8420 35660 8454
rect 35172 8414 35660 8420
rect 36190 8454 36678 8460
rect 36190 8420 36202 8454
rect 36666 8420 36678 8454
rect 36190 8414 36678 8420
rect 37208 8454 37696 8460
rect 37208 8420 37220 8454
rect 37684 8420 37696 8454
rect 37208 8414 37696 8420
rect 38226 8454 38714 8460
rect 38226 8420 38238 8454
rect 38702 8420 38714 8454
rect 38226 8414 38714 8420
rect 39244 8454 39732 8460
rect 39244 8420 39256 8454
rect 39720 8420 39732 8454
rect 39244 8414 39732 8420
rect 34878 8312 34890 8370
rect 34884 7840 34890 8312
rect 33906 7794 33916 7830
rect 33136 7744 33624 7750
rect 33136 7710 33148 7744
rect 33612 7710 33624 7744
rect 33136 7704 33624 7710
rect 32834 7606 32840 7666
rect 32900 7606 32906 7666
rect 32012 7280 32018 7340
rect 32078 7280 32084 7340
rect 32306 7282 32312 7342
rect 32372 7282 32378 7342
rect 32312 7226 32372 7282
rect 32118 7220 32606 7226
rect 32118 7186 32130 7220
rect 32594 7186 32606 7220
rect 32118 7180 32606 7186
rect 30852 6606 30858 7098
rect 31822 7092 31836 7136
rect 30852 6560 30866 6606
rect 24992 6510 25480 6516
rect 24992 6476 25004 6510
rect 25468 6476 25480 6510
rect 24992 6470 25480 6476
rect 26010 6510 26498 6516
rect 26010 6476 26022 6510
rect 26486 6476 26498 6510
rect 26010 6470 26498 6476
rect 27028 6510 27516 6516
rect 27028 6476 27040 6510
rect 27504 6476 27516 6510
rect 27028 6470 27516 6476
rect 28046 6510 28534 6516
rect 28046 6476 28058 6510
rect 28522 6476 28534 6510
rect 28046 6470 28534 6476
rect 29064 6510 29552 6516
rect 29064 6476 29076 6510
rect 29540 6476 29552 6510
rect 29064 6470 29552 6476
rect 30082 6510 30570 6516
rect 30082 6476 30094 6510
rect 30558 6476 30570 6510
rect 30082 6470 30570 6476
rect 24692 6350 24698 6410
rect 24758 6350 24764 6410
rect 21638 6046 21644 6106
rect 21704 6046 21710 6106
rect 20920 5988 21408 5994
rect 20920 5954 20932 5988
rect 21396 5954 21408 5988
rect 20920 5948 21408 5954
rect 20624 5866 20638 5904
rect 19654 5328 19664 5374
rect 20632 5370 20638 5866
rect 19604 5166 19664 5328
rect 20622 5328 20638 5370
rect 20672 5866 20684 5904
rect 21644 5904 21704 6046
rect 21938 5988 22426 5994
rect 21938 5954 21950 5988
rect 22414 5954 22426 5988
rect 21938 5948 22426 5954
rect 20672 5370 20678 5866
rect 21644 5864 21656 5904
rect 20672 5328 20682 5370
rect 19902 5278 20390 5284
rect 19902 5244 19914 5278
rect 20378 5244 20390 5278
rect 19902 5238 20390 5244
rect 20116 5166 20176 5238
rect 20622 5166 20682 5328
rect 21650 5328 21656 5864
rect 21690 5864 21704 5904
rect 22660 5904 22720 6146
rect 23162 6140 23168 6200
rect 23228 6140 23234 6200
rect 24184 6140 24190 6200
rect 24250 6140 24256 6200
rect 23672 6046 23678 6106
rect 23738 6046 23744 6106
rect 22956 5988 23444 5994
rect 22956 5954 22968 5988
rect 23432 5954 23444 5988
rect 22956 5948 23444 5954
rect 21690 5328 21696 5864
rect 22660 5852 22674 5904
rect 21650 5316 21696 5328
rect 22668 5328 22674 5852
rect 22708 5852 22720 5904
rect 23678 5904 23738 6046
rect 24190 5994 24250 6140
rect 23974 5988 24462 5994
rect 23974 5954 23986 5988
rect 24450 5954 24462 5988
rect 23974 5948 24462 5954
rect 23678 5860 23692 5904
rect 22708 5328 22714 5852
rect 23686 5364 23692 5860
rect 22668 5316 22714 5328
rect 23678 5328 23692 5364
rect 23726 5860 23738 5904
rect 24698 5904 24758 6350
rect 25204 6200 25264 6470
rect 26222 6308 26282 6470
rect 27242 6420 27302 6470
rect 28242 6420 28302 6470
rect 29280 6420 29340 6470
rect 30308 6420 30368 6470
rect 26724 6350 26730 6410
rect 26790 6350 26796 6410
rect 27242 6360 30368 6420
rect 26216 6248 26222 6308
rect 26282 6248 26288 6308
rect 25198 6140 25204 6200
rect 25264 6140 25270 6200
rect 26216 6140 26222 6200
rect 26282 6140 26288 6200
rect 25204 5994 25264 6140
rect 25708 6046 25714 6106
rect 25774 6046 25780 6106
rect 24992 5988 25480 5994
rect 24992 5954 25004 5988
rect 25468 5954 25480 5988
rect 24992 5948 25480 5954
rect 23726 5364 23732 5860
rect 23726 5328 23738 5364
rect 20920 5278 21408 5284
rect 20920 5244 20932 5278
rect 21396 5244 21408 5278
rect 20920 5238 21408 5244
rect 21938 5278 22426 5284
rect 21938 5244 21950 5278
rect 22414 5244 22426 5278
rect 21938 5238 22426 5244
rect 22956 5278 23444 5284
rect 22956 5244 22968 5278
rect 23432 5244 23444 5278
rect 22956 5238 23444 5244
rect 21126 5182 21186 5238
rect 19604 5106 20682 5166
rect 21120 5122 21126 5182
rect 21186 5122 21192 5182
rect 22030 5122 22036 5182
rect 22096 5122 22102 5182
rect 21120 4906 21126 4966
rect 21186 4906 21192 4966
rect 21126 4900 21188 4906
rect 19488 4862 19550 4868
rect 19488 4802 19490 4862
rect 19488 4796 19550 4802
rect 19488 2618 19548 4796
rect 21128 4760 21188 4900
rect 22036 4760 22096 5122
rect 22164 4966 22224 5238
rect 23032 5122 23038 5182
rect 23098 5122 23104 5182
rect 22164 4900 22224 4906
rect 23038 4760 23098 5122
rect 23178 4966 23238 5238
rect 23678 5080 23738 5328
rect 24698 5328 24710 5904
rect 24744 5328 24758 5904
rect 25714 5904 25774 6046
rect 26222 5994 26282 6140
rect 26010 5988 26498 5994
rect 26010 5954 26022 5988
rect 26486 5954 26498 5988
rect 26010 5948 26498 5954
rect 25714 5868 25728 5904
rect 23974 5278 24462 5284
rect 23974 5244 23986 5278
rect 24450 5244 24462 5278
rect 23974 5238 24462 5244
rect 24190 5182 24250 5238
rect 24184 5122 24190 5182
rect 24250 5122 24256 5182
rect 23672 5020 23678 5080
rect 23738 5020 23744 5080
rect 23172 4906 23178 4966
rect 23238 4906 23244 4966
rect 24190 4760 24250 5122
rect 19902 4754 20390 4760
rect 19902 4720 19914 4754
rect 20378 4720 20390 4754
rect 19902 4714 20390 4720
rect 20920 4754 21408 4760
rect 20920 4720 20932 4754
rect 21396 4720 21408 4754
rect 20920 4714 21408 4720
rect 21938 4754 22426 4760
rect 21938 4720 21950 4754
rect 22414 4720 22426 4754
rect 21938 4714 22426 4720
rect 22956 4754 23444 4760
rect 22956 4720 22968 4754
rect 23432 4720 23444 4754
rect 22956 4714 23444 4720
rect 23974 4754 24462 4760
rect 23974 4720 23986 4754
rect 24450 4720 24462 4754
rect 23974 4714 24462 4720
rect 19614 4670 19660 4682
rect 19614 4132 19620 4670
rect 19608 4094 19620 4132
rect 19654 4132 19660 4670
rect 20632 4670 20678 4682
rect 20632 4132 20638 4670
rect 19654 4094 19668 4132
rect 19608 3964 19668 4094
rect 20626 4094 20638 4132
rect 20672 4132 20678 4670
rect 21650 4670 21696 4682
rect 21650 4144 21656 4670
rect 20672 4094 20686 4132
rect 19902 4044 20390 4050
rect 19902 4010 19914 4044
rect 20378 4010 20390 4044
rect 19902 4004 20390 4010
rect 20106 3964 20166 4004
rect 20626 3964 20686 4094
rect 21642 4094 21656 4144
rect 21690 4144 21696 4670
rect 22668 4670 22714 4682
rect 22668 4152 22674 4670
rect 21690 4094 21702 4144
rect 20920 4044 21408 4050
rect 20920 4010 20932 4044
rect 21396 4010 21408 4044
rect 20920 4004 21408 4010
rect 19608 3904 20686 3964
rect 20626 3850 20686 3904
rect 21118 3894 21124 3954
rect 21184 3894 21190 3954
rect 20620 3790 20626 3850
rect 20686 3790 20692 3850
rect 20616 3580 20622 3640
rect 20682 3580 20688 3640
rect 19902 3520 20390 3526
rect 19902 3486 19914 3520
rect 20378 3486 20390 3520
rect 19902 3480 20390 3486
rect 19614 3436 19660 3448
rect 19614 2894 19620 3436
rect 19604 2860 19620 2894
rect 19654 2894 19660 3436
rect 20622 3436 20682 3580
rect 21124 3526 21184 3894
rect 21642 3738 21702 4094
rect 22660 4094 22674 4152
rect 22708 4152 22714 4670
rect 23686 4670 23732 4682
rect 22708 4094 22720 4152
rect 23686 4140 23692 4670
rect 21938 4044 22426 4050
rect 21938 4010 21950 4044
rect 22414 4010 22426 4044
rect 21938 4004 22426 4010
rect 22132 3954 22192 4004
rect 22126 3894 22132 3954
rect 22192 3894 22198 3954
rect 21636 3678 21642 3738
rect 21702 3678 21708 3738
rect 22660 3640 22720 4094
rect 23680 4094 23692 4140
rect 23726 4140 23732 4670
rect 24698 4670 24758 5328
rect 25722 5328 25728 5868
rect 25762 5868 25774 5904
rect 26730 5904 26790 6350
rect 27236 6140 27242 6200
rect 27302 6140 27308 6200
rect 30308 6184 30368 6360
rect 30806 6294 30866 6560
rect 31830 6560 31836 7092
rect 31870 7092 31882 7136
rect 32840 7136 32900 7606
rect 33342 7348 33402 7704
rect 33856 7450 33916 7794
rect 34876 7794 34890 7840
rect 34924 8312 34938 8370
rect 35902 8370 35948 8382
rect 34924 7840 34930 8312
rect 35902 7850 35908 8370
rect 34924 7794 34936 7840
rect 34154 7744 34642 7750
rect 34154 7710 34166 7744
rect 34630 7710 34642 7744
rect 34154 7704 34642 7710
rect 33850 7390 33856 7450
rect 33916 7390 33922 7450
rect 33340 7342 33402 7348
rect 33400 7282 33402 7342
rect 33340 7276 33402 7282
rect 33852 7276 33858 7336
rect 33918 7276 33924 7336
rect 33342 7226 33402 7276
rect 33136 7220 33624 7226
rect 33136 7186 33148 7220
rect 33612 7186 33624 7220
rect 33136 7180 33624 7186
rect 32840 7092 32854 7136
rect 31870 6560 31876 7092
rect 31830 6548 31876 6560
rect 32848 6560 32854 7092
rect 32888 7092 32900 7136
rect 33858 7136 33918 7276
rect 34366 7226 34426 7704
rect 34876 7666 34936 7794
rect 35894 7794 35908 7850
rect 35942 7850 35948 8370
rect 36920 8370 36966 8382
rect 35942 7794 35954 7850
rect 36920 7838 36926 8370
rect 35172 7744 35660 7750
rect 35172 7710 35184 7744
rect 35648 7710 35660 7744
rect 35172 7704 35660 7710
rect 34870 7606 34876 7666
rect 34936 7606 34942 7666
rect 34154 7220 34642 7226
rect 34154 7186 34166 7220
rect 34630 7186 34642 7220
rect 34154 7180 34642 7186
rect 33858 7106 33872 7136
rect 32888 6560 32894 7092
rect 33866 6600 33872 7106
rect 32848 6548 32894 6560
rect 33858 6560 33872 6600
rect 33906 7106 33918 7136
rect 34876 7136 34936 7606
rect 35392 7226 35452 7704
rect 35894 7450 35954 7794
rect 36910 7794 36926 7838
rect 36960 7838 36966 8370
rect 37938 8370 37984 8382
rect 37938 7838 37944 8370
rect 36960 7794 36970 7838
rect 36190 7744 36678 7750
rect 36190 7710 36202 7744
rect 36666 7710 36678 7744
rect 36190 7704 36678 7710
rect 35888 7390 35894 7450
rect 35954 7390 35960 7450
rect 36400 7400 36460 7704
rect 36910 7558 36970 7794
rect 37934 7794 37944 7838
rect 37978 7838 37984 8370
rect 38956 8370 39002 8382
rect 38956 7844 38962 8370
rect 37978 7794 37994 7838
rect 37208 7744 37696 7750
rect 37208 7710 37220 7744
rect 37684 7710 37696 7744
rect 37208 7704 37696 7710
rect 37416 7560 37476 7704
rect 36904 7498 36910 7558
rect 36970 7498 36976 7558
rect 37414 7554 37476 7560
rect 37474 7494 37476 7554
rect 37414 7488 37476 7494
rect 37416 7400 37476 7488
rect 37934 7450 37994 7794
rect 38950 7794 38962 7844
rect 38996 7844 39002 8370
rect 39966 8370 40026 8536
rect 40068 8512 40074 8572
rect 40134 8512 40140 8572
rect 40202 8554 40262 8842
rect 39966 8342 39980 8370
rect 39974 7852 39980 8342
rect 38996 7794 39010 7844
rect 38226 7744 38714 7750
rect 38226 7710 38238 7744
rect 38702 7710 38714 7744
rect 38226 7704 38714 7710
rect 36400 7340 37476 7400
rect 37928 7390 37934 7450
rect 37994 7390 38000 7450
rect 35888 7276 35894 7336
rect 35954 7276 35960 7336
rect 35172 7220 35660 7226
rect 35172 7186 35184 7220
rect 35648 7186 35660 7220
rect 35172 7180 35660 7186
rect 33906 6600 33912 7106
rect 34876 7096 34890 7136
rect 33906 6560 33918 6600
rect 34884 6594 34890 7096
rect 31100 6510 31588 6516
rect 31100 6476 31112 6510
rect 31576 6476 31588 6510
rect 31100 6470 31588 6476
rect 32118 6510 32606 6516
rect 32118 6476 32130 6510
rect 32594 6476 32606 6510
rect 32118 6470 32606 6476
rect 33136 6510 33624 6516
rect 33136 6476 33148 6510
rect 33612 6476 33624 6510
rect 33136 6470 33624 6476
rect 31312 6422 31372 6470
rect 30800 6234 30806 6294
rect 30866 6234 30872 6294
rect 31312 6184 31372 6362
rect 27242 5994 27302 6140
rect 30308 6124 31372 6184
rect 32836 6036 32842 6096
rect 32902 6036 32908 6096
rect 27028 5988 27516 5994
rect 27028 5954 27040 5988
rect 27504 5954 27516 5988
rect 27028 5948 27516 5954
rect 28046 5988 28534 5994
rect 28046 5954 28058 5988
rect 28522 5954 28534 5988
rect 28046 5948 28534 5954
rect 29064 5988 29552 5994
rect 29064 5954 29076 5988
rect 29540 5954 29552 5988
rect 29064 5948 29552 5954
rect 30082 5988 30570 5994
rect 30082 5954 30094 5988
rect 30558 5954 30570 5988
rect 30082 5948 30570 5954
rect 31100 5988 31588 5994
rect 31100 5954 31112 5988
rect 31576 5954 31588 5988
rect 31100 5948 31588 5954
rect 32118 5988 32606 5994
rect 32118 5954 32130 5988
rect 32594 5954 32606 5988
rect 32118 5948 32606 5954
rect 25762 5328 25768 5868
rect 26730 5866 26746 5904
rect 25722 5316 25768 5328
rect 26740 5328 26746 5866
rect 26780 5866 26790 5904
rect 27758 5904 27804 5916
rect 26780 5328 26786 5866
rect 27758 5370 27764 5904
rect 26740 5316 26786 5328
rect 27750 5328 27764 5370
rect 27798 5370 27804 5904
rect 28776 5904 28822 5916
rect 27798 5328 27810 5370
rect 28776 5366 28782 5904
rect 24992 5278 25480 5284
rect 24992 5244 25004 5278
rect 25468 5244 25480 5278
rect 24992 5238 25480 5244
rect 26010 5278 26498 5284
rect 26010 5244 26022 5278
rect 26486 5244 26498 5278
rect 26010 5238 26498 5244
rect 27028 5278 27516 5284
rect 27028 5244 27040 5278
rect 27504 5244 27516 5278
rect 27028 5238 27516 5244
rect 25200 5182 25260 5238
rect 26206 5182 26266 5238
rect 27250 5182 27310 5238
rect 27750 5188 27810 5328
rect 28770 5328 28782 5366
rect 28816 5366 28822 5904
rect 29794 5904 29840 5916
rect 28816 5328 28830 5366
rect 29794 5360 29800 5904
rect 28046 5278 28534 5284
rect 28046 5244 28058 5278
rect 28522 5244 28534 5278
rect 28046 5238 28534 5244
rect 25194 5122 25200 5182
rect 25260 5122 25266 5182
rect 26200 5122 26206 5182
rect 26266 5122 26272 5182
rect 27244 5122 27250 5182
rect 27310 5122 27316 5182
rect 27744 5128 27750 5188
rect 27810 5128 27816 5188
rect 25200 4760 25260 5122
rect 26198 4906 26204 4966
rect 26264 4906 26270 4966
rect 27238 4906 27244 4966
rect 27304 4906 27310 4966
rect 26204 4760 26264 4906
rect 26722 4802 26728 4862
rect 26788 4802 26794 4862
rect 24992 4754 25480 4760
rect 24992 4720 25004 4754
rect 25468 4720 25480 4754
rect 24992 4714 25480 4720
rect 26010 4754 26498 4760
rect 26010 4720 26022 4754
rect 26486 4720 26498 4754
rect 26010 4714 26498 4720
rect 24698 4588 24710 4670
rect 24704 4140 24710 4588
rect 23726 4094 23740 4140
rect 22956 4044 23444 4050
rect 22956 4010 22968 4044
rect 23432 4010 23444 4044
rect 22956 4004 23444 4010
rect 23146 3954 23206 4004
rect 23140 3894 23146 3954
rect 23206 3894 23212 3954
rect 23680 3738 23740 4094
rect 24700 4094 24710 4140
rect 24744 4588 24758 4670
rect 25722 4670 25768 4682
rect 24744 4140 24750 4588
rect 24744 4094 24760 4140
rect 25722 4138 25728 4670
rect 23974 4044 24462 4050
rect 23974 4010 23986 4044
rect 24450 4010 24462 4044
rect 23974 4004 24462 4010
rect 24184 3954 24244 4004
rect 24178 3894 24184 3954
rect 24244 3894 24250 3954
rect 23674 3678 23680 3738
rect 23740 3678 23746 3738
rect 22654 3580 22660 3640
rect 22720 3580 22726 3640
rect 24184 3526 24244 3894
rect 24700 3640 24760 4094
rect 25718 4094 25728 4138
rect 25762 4138 25768 4670
rect 26728 4670 26788 4802
rect 27244 4760 27304 4906
rect 27028 4754 27516 4760
rect 27028 4720 27040 4754
rect 27504 4720 27516 4754
rect 27028 4714 27516 4720
rect 26728 4606 26746 4670
rect 25762 4094 25778 4138
rect 24992 4044 25480 4050
rect 24992 4010 25004 4044
rect 25468 4010 25480 4044
rect 24992 4004 25480 4010
rect 25202 3954 25262 4004
rect 25718 3960 25778 4094
rect 26740 4094 26746 4606
rect 26780 4606 26788 4670
rect 27750 4670 27810 5128
rect 28258 4966 28318 5238
rect 28252 4906 28258 4966
rect 28318 4906 28324 4966
rect 28258 4760 28318 4906
rect 28770 4862 28830 5328
rect 29786 5328 29800 5360
rect 29834 5360 29840 5904
rect 30812 5904 30858 5916
rect 30812 5362 30818 5904
rect 29834 5328 29846 5360
rect 29064 5278 29552 5284
rect 29064 5244 29076 5278
rect 29540 5244 29552 5278
rect 29064 5238 29552 5244
rect 29266 4966 29326 5238
rect 29786 5188 29846 5328
rect 30808 5328 30818 5362
rect 30852 5362 30858 5904
rect 31830 5904 31876 5916
rect 30852 5328 30868 5362
rect 31830 5360 31836 5904
rect 30082 5278 30570 5284
rect 30082 5244 30094 5278
rect 30558 5244 30570 5278
rect 30082 5238 30570 5244
rect 29780 5128 29786 5188
rect 29846 5128 29852 5188
rect 30310 4966 30370 5238
rect 29260 4906 29266 4966
rect 29326 4906 29332 4966
rect 30304 4906 30310 4966
rect 30370 4906 30376 4966
rect 28764 4802 28770 4862
rect 28830 4802 28836 4862
rect 28046 4754 28534 4760
rect 28046 4720 28058 4754
rect 28522 4720 28534 4754
rect 28046 4714 28534 4720
rect 27750 4634 27764 4670
rect 26780 4094 26786 4606
rect 27758 4152 27764 4634
rect 26740 4082 26786 4094
rect 27754 4094 27764 4152
rect 27798 4634 27810 4670
rect 28770 4670 28830 4802
rect 29266 4760 29326 4906
rect 30310 4760 30370 4906
rect 30808 4862 30868 5328
rect 31822 5328 31836 5360
rect 31870 5360 31876 5904
rect 32842 5904 32902 6036
rect 33136 5988 33624 5994
rect 33136 5954 33148 5988
rect 33612 5954 33624 5988
rect 33136 5948 33624 5954
rect 31870 5328 31882 5360
rect 31100 5278 31588 5284
rect 31100 5244 31112 5278
rect 31576 5244 31588 5278
rect 31100 5238 31588 5244
rect 31300 4966 31360 5238
rect 31822 5188 31882 5328
rect 32842 5328 32854 5904
rect 32888 5328 32902 5904
rect 33858 5904 33918 6560
rect 34878 6560 34890 6594
rect 34924 7096 34936 7136
rect 35894 7136 35954 7276
rect 36400 7226 36460 7340
rect 37416 7226 37476 7340
rect 37926 7276 37932 7336
rect 37992 7276 37998 7336
rect 36190 7220 36678 7226
rect 36190 7186 36202 7220
rect 36666 7186 36678 7220
rect 36190 7180 36678 7186
rect 37208 7220 37696 7226
rect 37208 7186 37220 7220
rect 37684 7186 37696 7220
rect 37208 7180 37696 7186
rect 34924 6594 34930 7096
rect 35894 7094 35908 7136
rect 34924 6560 34938 6594
rect 34154 6510 34642 6516
rect 34154 6476 34166 6510
rect 34630 6476 34642 6510
rect 34154 6470 34642 6476
rect 34354 6200 34414 6470
rect 34348 6140 34354 6200
rect 34414 6140 34420 6200
rect 34354 5994 34414 6140
rect 34154 5988 34642 5994
rect 34154 5954 34166 5988
rect 34630 5954 34642 5988
rect 34154 5948 34642 5954
rect 33858 5864 33872 5904
rect 33866 5360 33872 5864
rect 32118 5278 32606 5284
rect 32118 5244 32130 5278
rect 32594 5244 32606 5278
rect 32118 5238 32606 5244
rect 31816 5128 31822 5188
rect 31882 5128 31888 5188
rect 32318 4966 32378 5238
rect 31294 4906 31300 4966
rect 31360 4906 31366 4966
rect 32312 4906 32318 4966
rect 32378 4906 32384 4966
rect 30802 4802 30808 4862
rect 30868 4802 30874 4862
rect 29064 4754 29552 4760
rect 29064 4720 29076 4754
rect 29540 4720 29552 4754
rect 29064 4714 29552 4720
rect 30082 4754 30570 4760
rect 30082 4720 30094 4754
rect 30558 4720 30570 4754
rect 30082 4714 30570 4720
rect 27798 4152 27804 4634
rect 28770 4632 28782 4670
rect 27798 4094 27814 4152
rect 26010 4044 26498 4050
rect 26010 4010 26022 4044
rect 26486 4010 26498 4044
rect 26010 4004 26498 4010
rect 27028 4044 27516 4050
rect 27028 4010 27040 4044
rect 27504 4010 27516 4044
rect 27028 4004 27516 4010
rect 27754 3960 27814 4094
rect 28776 4094 28782 4632
rect 28816 4632 28830 4670
rect 29794 4670 29840 4682
rect 28816 4094 28822 4632
rect 29794 4144 29800 4670
rect 28776 4082 28822 4094
rect 29786 4094 29800 4144
rect 29834 4144 29840 4670
rect 30808 4670 30868 4802
rect 31300 4760 31360 4906
rect 32842 4862 32902 5328
rect 33860 5328 33872 5360
rect 33906 5864 33918 5904
rect 34878 5904 34938 6560
rect 35902 6560 35908 7094
rect 35942 7094 35954 7136
rect 36920 7136 36966 7148
rect 35942 6560 35948 7094
rect 36920 6618 36926 7136
rect 35902 6548 35948 6560
rect 36912 6560 36926 6618
rect 36960 6618 36966 7136
rect 37932 7136 37992 7276
rect 38434 7226 38494 7704
rect 38950 7666 39010 7794
rect 39968 7794 39980 7852
rect 40014 8342 40026 8370
rect 40014 7852 40020 8342
rect 40014 7794 40028 7852
rect 39244 7744 39732 7750
rect 39244 7710 39256 7744
rect 39720 7710 39732 7744
rect 39244 7704 39732 7710
rect 39968 7684 40028 7794
rect 38944 7606 38950 7666
rect 39010 7606 39016 7666
rect 39962 7624 39968 7684
rect 40028 7624 40034 7684
rect 38950 7388 39010 7606
rect 38950 7328 40024 7388
rect 40074 7336 40134 8512
rect 40196 8494 40202 8554
rect 40262 8494 40268 8554
rect 40568 7554 40628 11440
rect 40562 7494 40568 7554
rect 40628 7494 40634 7554
rect 40312 7390 40318 7450
rect 40378 7390 40384 7450
rect 38226 7220 38714 7226
rect 38226 7186 38238 7220
rect 38702 7186 38714 7220
rect 38226 7180 38714 7186
rect 37932 7094 37944 7136
rect 36960 6560 36972 6618
rect 35384 6516 35444 6518
rect 35172 6510 35660 6516
rect 35172 6476 35184 6510
rect 35648 6476 35660 6510
rect 35172 6470 35660 6476
rect 36190 6510 36678 6516
rect 36190 6476 36202 6510
rect 36666 6476 36678 6510
rect 36190 6470 36678 6476
rect 35384 6200 35444 6470
rect 36406 6422 36466 6470
rect 36400 6362 36406 6422
rect 36466 6362 36472 6422
rect 36538 6366 36544 6426
rect 36604 6366 36610 6426
rect 36544 6200 36604 6366
rect 36912 6200 36972 6560
rect 37938 6560 37944 7094
rect 37978 7094 37992 7136
rect 38950 7136 39010 7328
rect 39454 7226 39514 7328
rect 39244 7220 39732 7226
rect 39244 7186 39256 7220
rect 39720 7186 39732 7220
rect 39244 7180 39732 7186
rect 38950 7102 38962 7136
rect 37978 6560 37984 7094
rect 38956 6600 38962 7102
rect 37938 6548 37984 6560
rect 38950 6560 38962 6600
rect 38996 7102 39010 7136
rect 39964 7136 40024 7328
rect 40068 7276 40074 7336
rect 40134 7276 40140 7336
rect 39964 7112 39980 7136
rect 38996 6600 39002 7102
rect 38996 6560 39010 6600
rect 37208 6510 37696 6516
rect 37208 6476 37220 6510
rect 37684 6476 37696 6510
rect 37208 6470 37696 6476
rect 38226 6510 38714 6516
rect 38226 6476 38238 6510
rect 38702 6476 38714 6510
rect 38226 6470 38714 6476
rect 38432 6426 38492 6470
rect 37420 6366 37426 6426
rect 37486 6366 37492 6426
rect 38426 6366 38432 6426
rect 38492 6366 38498 6426
rect 38950 6422 39010 6560
rect 39974 6560 39980 7112
rect 40014 7112 40024 7136
rect 40014 6560 40020 7112
rect 39974 6548 40020 6560
rect 39244 6510 39732 6516
rect 39244 6476 39256 6510
rect 39720 6476 39732 6510
rect 39244 6470 39732 6476
rect 35378 6140 35384 6200
rect 35444 6140 35450 6200
rect 36538 6140 36544 6200
rect 36604 6140 36610 6200
rect 36906 6140 36912 6200
rect 36972 6140 36978 6200
rect 35384 5994 35444 6140
rect 36544 5994 36604 6140
rect 36912 6096 36972 6140
rect 36906 6036 36912 6096
rect 36972 6036 36978 6096
rect 37426 5994 37486 6366
rect 38944 6362 38950 6422
rect 39010 6362 39016 6422
rect 38944 6234 38950 6294
rect 39010 6234 39016 6294
rect 37922 6038 37928 6098
rect 37988 6038 37994 6098
rect 35172 5988 35660 5994
rect 35172 5954 35184 5988
rect 35648 5954 35660 5988
rect 35172 5948 35660 5954
rect 36190 5988 36678 5994
rect 36190 5954 36202 5988
rect 36666 5954 36678 5988
rect 36190 5948 36678 5954
rect 37208 5988 37696 5994
rect 37208 5954 37220 5988
rect 37684 5954 37696 5988
rect 37208 5948 37696 5954
rect 37426 5946 37486 5948
rect 33906 5360 33912 5864
rect 34878 5858 34890 5904
rect 34884 5372 34890 5858
rect 33906 5328 33920 5360
rect 33136 5278 33624 5284
rect 33136 5244 33148 5278
rect 33612 5244 33624 5278
rect 33136 5238 33624 5244
rect 33352 4966 33412 5238
rect 33860 5188 33920 5328
rect 34876 5328 34890 5372
rect 34924 5858 34938 5904
rect 35902 5904 35948 5916
rect 34924 5372 34930 5858
rect 34924 5328 34936 5372
rect 35902 5368 35908 5904
rect 34154 5278 34642 5284
rect 34154 5244 34166 5278
rect 34630 5244 34642 5278
rect 34154 5238 34642 5244
rect 33854 5128 33860 5188
rect 33920 5128 33926 5188
rect 33846 5020 33852 5080
rect 33912 5020 33918 5080
rect 33346 4906 33352 4966
rect 33412 4906 33418 4966
rect 32836 4802 32842 4862
rect 32902 4802 32908 4862
rect 33348 4798 33354 4858
rect 33414 4798 33420 4858
rect 33354 4760 33414 4798
rect 31100 4754 31588 4760
rect 31100 4720 31112 4754
rect 31576 4720 31588 4754
rect 31100 4714 31588 4720
rect 32118 4754 32606 4760
rect 32118 4720 32130 4754
rect 32594 4720 32606 4754
rect 32118 4714 32606 4720
rect 33136 4754 33624 4760
rect 33136 4720 33148 4754
rect 33612 4720 33624 4754
rect 33136 4714 33624 4720
rect 30808 4634 30818 4670
rect 29834 4094 29846 4144
rect 28046 4044 28534 4050
rect 28046 4010 28058 4044
rect 28522 4010 28534 4044
rect 28046 4004 28534 4010
rect 29064 4044 29552 4050
rect 29064 4010 29076 4044
rect 29540 4010 29552 4044
rect 29064 4004 29552 4010
rect 29786 3960 29846 4094
rect 30812 4094 30818 4634
rect 30852 4634 30868 4670
rect 31830 4670 31876 4682
rect 30852 4094 30858 4634
rect 31830 4156 31836 4670
rect 30812 4082 30858 4094
rect 31820 4094 31836 4156
rect 31870 4156 31876 4670
rect 32848 4670 32894 4682
rect 31870 4094 31880 4156
rect 32848 4136 32854 4670
rect 30082 4044 30570 4050
rect 30082 4010 30094 4044
rect 30558 4010 30570 4044
rect 30082 4004 30570 4010
rect 31100 4044 31588 4050
rect 31100 4010 31112 4044
rect 31576 4010 31588 4044
rect 31100 4004 31588 4010
rect 31820 3960 31880 4094
rect 32842 4094 32854 4136
rect 32888 4136 32894 4670
rect 33852 4670 33912 5020
rect 34376 4858 34436 5238
rect 34876 4864 34936 5328
rect 35896 5328 35908 5368
rect 35942 5368 35948 5904
rect 36920 5904 36966 5916
rect 36920 5372 36926 5904
rect 35942 5328 35956 5368
rect 35172 5278 35660 5284
rect 35172 5244 35184 5278
rect 35648 5244 35660 5278
rect 35172 5238 35660 5244
rect 34370 4798 34376 4858
rect 34436 4798 34442 4858
rect 34870 4804 34876 4864
rect 34936 4804 34942 4864
rect 34376 4760 34436 4798
rect 34154 4754 34642 4760
rect 34154 4720 34166 4754
rect 34630 4720 34642 4754
rect 34154 4714 34642 4720
rect 33852 4634 33872 4670
rect 32888 4094 32902 4136
rect 32118 4044 32606 4050
rect 32118 4010 32130 4044
rect 32594 4010 32606 4044
rect 32118 4004 32606 4010
rect 25196 3894 25202 3954
rect 25262 3894 25268 3954
rect 25712 3900 25718 3960
rect 25778 3900 25784 3960
rect 29780 3900 29786 3960
rect 29846 3900 29852 3960
rect 31814 3900 31820 3960
rect 31880 3900 31886 3960
rect 24694 3580 24700 3640
rect 24760 3580 24766 3640
rect 20920 3520 21408 3526
rect 20920 3486 20932 3520
rect 21396 3486 21408 3520
rect 20920 3480 21408 3486
rect 21938 3520 22426 3526
rect 21938 3486 21950 3520
rect 22414 3486 22426 3520
rect 21938 3480 22426 3486
rect 22956 3520 23444 3526
rect 22956 3486 22968 3520
rect 23432 3486 23444 3520
rect 22956 3480 23444 3486
rect 23974 3520 24462 3526
rect 23974 3486 23986 3520
rect 24450 3486 24462 3520
rect 23974 3480 24462 3486
rect 20622 3382 20638 3436
rect 19654 2860 19664 2894
rect 20632 2890 20638 3382
rect 19604 2728 19664 2860
rect 20628 2860 20638 2890
rect 20672 3382 20682 3436
rect 21650 3436 21696 3448
rect 20672 2890 20678 3382
rect 21650 2906 21656 3436
rect 20672 2860 20688 2890
rect 19902 2810 20390 2816
rect 19902 2776 19914 2810
rect 20378 2776 20390 2810
rect 19902 2770 20390 2776
rect 20124 2728 20184 2770
rect 20628 2728 20688 2860
rect 21642 2860 21656 2906
rect 21690 2906 21696 3436
rect 22668 3436 22714 3448
rect 21690 2860 21702 2906
rect 22668 2890 22674 3436
rect 20920 2810 21408 2816
rect 20920 2776 20932 2810
rect 21396 2776 21408 2810
rect 20920 2770 21408 2776
rect 19604 2668 20688 2728
rect 19482 2558 19488 2618
rect 19548 2558 19554 2618
rect 20628 2522 20688 2668
rect 19604 2462 20688 2522
rect 19604 2204 19664 2462
rect 20116 2294 20176 2462
rect 20628 2402 20688 2462
rect 20622 2342 20628 2402
rect 20688 2342 20694 2402
rect 19902 2288 20390 2294
rect 19902 2254 19914 2288
rect 20378 2254 20390 2288
rect 19902 2248 20390 2254
rect 19604 2168 19620 2204
rect 19614 1628 19620 2168
rect 19654 2168 19664 2204
rect 20628 2204 20688 2342
rect 21120 2294 21180 2770
rect 21642 2716 21702 2860
rect 22660 2860 22674 2890
rect 22708 2890 22714 3436
rect 23686 3436 23732 3448
rect 23686 2902 23692 3436
rect 22708 2860 22720 2890
rect 21938 2810 22426 2816
rect 21938 2776 21950 2810
rect 22414 2776 22426 2810
rect 21938 2770 22426 2776
rect 21636 2656 21642 2716
rect 21702 2656 21708 2716
rect 21640 2462 21646 2522
rect 21706 2462 21712 2522
rect 20920 2288 21408 2294
rect 20920 2254 20932 2288
rect 21396 2254 21408 2288
rect 20920 2248 21408 2254
rect 19654 1628 19660 2168
rect 20628 2164 20638 2204
rect 19614 1616 19660 1628
rect 20632 1628 20638 2164
rect 20672 2164 20688 2204
rect 21646 2204 21706 2462
rect 22140 2458 22200 2770
rect 22660 2618 22720 2860
rect 23678 2860 23692 2902
rect 23726 2902 23732 3436
rect 24700 3436 24760 3580
rect 25202 3526 25262 3894
rect 24992 3520 25480 3526
rect 24992 3486 25004 3520
rect 25468 3486 25480 3520
rect 24992 3480 25480 3486
rect 24700 3406 24710 3436
rect 24704 2924 24710 3406
rect 23726 2860 23738 2902
rect 22956 2810 23444 2816
rect 22956 2776 22968 2810
rect 23432 2776 23444 2810
rect 22956 2770 23444 2776
rect 22654 2558 22660 2618
rect 22720 2558 22726 2618
rect 23174 2458 23234 2770
rect 23678 2716 23738 2860
rect 24696 2860 24710 2924
rect 24744 3406 24760 3436
rect 25718 3436 25778 3900
rect 27754 3894 27814 3900
rect 28764 3790 28770 3850
rect 28830 3790 28836 3850
rect 30800 3790 30806 3850
rect 30866 3790 30872 3850
rect 27746 3678 27752 3738
rect 27812 3678 27818 3738
rect 26730 3580 26736 3640
rect 26796 3580 26802 3640
rect 26010 3520 26498 3526
rect 26010 3486 26022 3520
rect 26486 3486 26498 3520
rect 26010 3480 26498 3486
rect 24744 2924 24750 3406
rect 25718 3394 25728 3436
rect 24744 2860 24756 2924
rect 25722 2900 25728 3394
rect 23974 2810 24462 2816
rect 23974 2776 23986 2810
rect 24450 2776 24462 2810
rect 23974 2770 24462 2776
rect 23672 2656 23678 2716
rect 23738 2656 23744 2716
rect 24184 2618 24244 2770
rect 24178 2558 24184 2618
rect 24244 2558 24250 2618
rect 23676 2462 23682 2522
rect 23742 2462 23748 2522
rect 22140 2398 23234 2458
rect 22140 2294 22200 2398
rect 23174 2294 23234 2398
rect 21938 2288 22426 2294
rect 21938 2254 21950 2288
rect 22414 2254 22426 2288
rect 21938 2248 22426 2254
rect 22956 2288 23444 2294
rect 22956 2254 22968 2288
rect 23432 2254 23444 2288
rect 22956 2248 23444 2254
rect 20672 1628 20678 2164
rect 21646 2160 21656 2204
rect 20632 1616 20678 1628
rect 21650 1628 21656 2160
rect 21690 2160 21706 2204
rect 22668 2204 22714 2216
rect 21690 1628 21696 2160
rect 22668 1670 22674 2204
rect 21650 1616 21696 1628
rect 22660 1628 22674 1670
rect 22708 1670 22714 2204
rect 23682 2204 23742 2462
rect 24184 2294 24244 2558
rect 24696 2402 24756 2860
rect 25716 2860 25728 2900
rect 25762 3394 25778 3436
rect 26736 3436 26796 3580
rect 27028 3520 27516 3526
rect 27028 3486 27040 3520
rect 27504 3486 27516 3520
rect 27028 3480 27516 3486
rect 26736 3400 26746 3436
rect 25762 2900 25768 3394
rect 25762 2860 25776 2900
rect 26740 2894 26746 3400
rect 24992 2810 25480 2816
rect 24992 2776 25004 2810
rect 25468 2776 25480 2810
rect 24992 2770 25480 2776
rect 25206 2618 25266 2770
rect 25716 2716 25776 2860
rect 26730 2860 26746 2894
rect 26780 3400 26796 3436
rect 27752 3436 27812 3678
rect 28046 3520 28534 3526
rect 28046 3486 28058 3520
rect 28522 3486 28534 3520
rect 28046 3480 28534 3486
rect 27752 3410 27764 3436
rect 26780 2894 26786 3400
rect 27758 2916 27764 3410
rect 26780 2860 26790 2894
rect 26010 2810 26498 2816
rect 26010 2776 26022 2810
rect 26486 2776 26498 2810
rect 26010 2770 26498 2776
rect 25710 2656 25716 2716
rect 25776 2656 25782 2716
rect 26230 2624 26290 2770
rect 24690 2342 24696 2402
rect 24756 2342 24762 2402
rect 23974 2288 24462 2294
rect 23974 2254 23986 2288
rect 24450 2254 24462 2288
rect 23974 2248 24462 2254
rect 23682 2152 23692 2204
rect 22708 1628 22720 1670
rect 19902 1578 20390 1584
rect 19902 1544 19914 1578
rect 20378 1544 20390 1578
rect 19902 1538 20390 1544
rect 20920 1578 21408 1584
rect 20920 1544 20932 1578
rect 21396 1544 21408 1578
rect 20920 1538 21408 1544
rect 21938 1578 22426 1584
rect 21938 1544 21950 1578
rect 22414 1544 22426 1578
rect 21938 1538 22426 1544
rect 19370 1426 19376 1486
rect 19436 1426 19442 1486
rect 19264 1300 19270 1360
rect 19330 1300 19336 1360
rect 19604 1120 20684 1180
rect 19604 970 19664 1120
rect 20112 1060 20172 1120
rect 19902 1054 20390 1060
rect 19902 1020 19914 1054
rect 20378 1020 20390 1054
rect 19902 1014 20390 1020
rect 19604 914 19620 970
rect 19614 394 19620 914
rect 19654 914 19664 970
rect 20624 970 20684 1120
rect 21122 1060 21182 1538
rect 22660 1360 22720 1628
rect 23686 1628 23692 2152
rect 23726 2152 23742 2204
rect 24696 2204 24756 2342
rect 25206 2294 25266 2558
rect 26228 2618 26290 2624
rect 26288 2558 26290 2618
rect 26228 2552 26290 2558
rect 25704 2462 25710 2522
rect 25770 2462 25776 2522
rect 24992 2288 25480 2294
rect 24992 2254 25004 2288
rect 25468 2254 25480 2288
rect 24992 2248 25480 2254
rect 24696 2164 24710 2204
rect 23726 1628 23732 2152
rect 24704 1682 24710 2164
rect 23686 1616 23732 1628
rect 24698 1628 24710 1682
rect 24744 2164 24756 2204
rect 25710 2204 25770 2462
rect 26230 2294 26290 2552
rect 26730 2402 26790 2860
rect 27748 2860 27764 2916
rect 27798 3410 27812 3436
rect 28770 3436 28830 3790
rect 29064 3520 29552 3526
rect 29064 3486 29076 3520
rect 29540 3486 29552 3520
rect 29064 3480 29552 3486
rect 30082 3520 30570 3526
rect 30082 3486 30094 3520
rect 30558 3486 30570 3520
rect 30082 3480 30570 3486
rect 27798 2916 27804 3410
rect 28770 3404 28782 3436
rect 27798 2860 27808 2916
rect 27028 2810 27516 2816
rect 27028 2776 27040 2810
rect 27504 2776 27516 2810
rect 27028 2770 27516 2776
rect 27232 2618 27292 2770
rect 27578 2736 27638 2742
rect 27748 2736 27808 2860
rect 28776 2860 28782 3404
rect 28816 3404 28830 3436
rect 29794 3436 29840 3448
rect 28816 2860 28822 3404
rect 29794 2930 29800 3436
rect 28776 2848 28822 2860
rect 29790 2860 29800 2930
rect 29834 2930 29840 3436
rect 30806 3436 30866 3790
rect 32348 3752 32408 4004
rect 32842 3962 32902 4094
rect 33866 4094 33872 4634
rect 33906 4094 33912 4670
rect 34876 4670 34936 4804
rect 35354 4760 35414 5238
rect 35896 5188 35956 5328
rect 36910 5328 36926 5372
rect 36960 5372 36966 5904
rect 37928 5904 37988 6038
rect 38226 5988 38714 5994
rect 38226 5954 38238 5988
rect 38702 5954 38714 5988
rect 38226 5948 38714 5954
rect 37928 5854 37944 5904
rect 36960 5328 36970 5372
rect 37938 5356 37944 5854
rect 36190 5278 36678 5284
rect 36190 5244 36202 5278
rect 36666 5244 36678 5278
rect 36190 5238 36678 5244
rect 35890 5128 35896 5188
rect 35956 5128 35962 5188
rect 35886 5020 35892 5080
rect 35952 5020 35958 5080
rect 35172 4754 35660 4760
rect 35172 4720 35184 4754
rect 35648 4720 35660 4754
rect 35172 4714 35660 4720
rect 34876 4576 34890 4670
rect 34884 4136 34890 4576
rect 33866 4082 33912 4094
rect 34876 4094 34890 4136
rect 34924 4576 34936 4670
rect 35892 4670 35952 5020
rect 36378 4906 36384 4966
rect 36444 4906 36450 4966
rect 36384 4760 36444 4906
rect 36910 4864 36970 5328
rect 37934 5328 37944 5356
rect 37978 5854 37988 5904
rect 38950 5904 39010 6234
rect 39244 5988 39732 5994
rect 39244 5954 39256 5988
rect 39720 5954 39732 5988
rect 39244 5948 39732 5954
rect 37978 5356 37984 5854
rect 38950 5852 38962 5904
rect 38956 5356 38962 5852
rect 37978 5328 37994 5356
rect 37208 5278 37696 5284
rect 37208 5244 37220 5278
rect 37684 5244 37696 5278
rect 37208 5238 37696 5244
rect 37934 5188 37994 5328
rect 38950 5328 38962 5356
rect 38996 5852 39010 5904
rect 39974 5904 40020 5916
rect 38996 5356 39002 5852
rect 39974 5362 39980 5904
rect 38996 5328 39010 5356
rect 38226 5278 38714 5284
rect 38226 5244 38238 5278
rect 38702 5244 38714 5278
rect 38226 5238 38714 5244
rect 37928 5128 37934 5188
rect 37994 5128 38000 5188
rect 37924 5020 37930 5080
rect 37990 5020 37996 5080
rect 37416 4906 37422 4966
rect 37482 4906 37488 4966
rect 36904 4804 36910 4864
rect 36970 4804 36976 4864
rect 37422 4760 37482 4906
rect 36190 4754 36678 4760
rect 36190 4720 36202 4754
rect 36666 4720 36678 4754
rect 36190 4714 36678 4720
rect 37208 4754 37696 4760
rect 37208 4720 37220 4754
rect 37684 4720 37696 4754
rect 37208 4714 37696 4720
rect 35892 4604 35908 4670
rect 34924 4136 34930 4576
rect 34924 4094 34936 4136
rect 33136 4044 33624 4050
rect 33136 4010 33148 4044
rect 33612 4010 33624 4044
rect 33136 4004 33624 4010
rect 34154 4044 34642 4050
rect 34154 4010 34166 4044
rect 34630 4010 34642 4044
rect 34154 4004 34642 4010
rect 32836 3902 32842 3962
rect 32902 3902 32908 3962
rect 33190 3902 33196 3962
rect 33256 3902 33262 3962
rect 32832 3790 32838 3850
rect 32898 3790 32904 3850
rect 32342 3692 32348 3752
rect 32408 3692 32414 3752
rect 31100 3520 31588 3526
rect 31100 3486 31112 3520
rect 31576 3486 31588 3520
rect 31100 3480 31588 3486
rect 32118 3520 32606 3526
rect 32118 3486 32130 3520
rect 32594 3486 32606 3520
rect 32118 3480 32606 3486
rect 30806 3398 30818 3436
rect 29834 2860 29850 2930
rect 28046 2810 28534 2816
rect 28046 2776 28058 2810
rect 28522 2776 28534 2810
rect 28046 2770 28534 2776
rect 29064 2810 29552 2816
rect 29064 2776 29076 2810
rect 29540 2776 29552 2810
rect 29064 2770 29552 2776
rect 27742 2676 27748 2736
rect 27808 2676 27814 2736
rect 27226 2558 27232 2618
rect 27292 2558 27298 2618
rect 26724 2342 26730 2402
rect 26790 2342 26796 2402
rect 26010 2288 26498 2294
rect 26010 2254 26022 2288
rect 26486 2254 26498 2288
rect 26010 2248 26498 2254
rect 24744 1682 24750 2164
rect 25710 2144 25728 2204
rect 24744 1628 24758 1682
rect 22956 1578 23444 1584
rect 22956 1544 22968 1578
rect 23432 1544 23444 1578
rect 22956 1538 23444 1544
rect 23974 1578 24462 1584
rect 23974 1544 23986 1578
rect 24450 1544 24462 1578
rect 23974 1538 24462 1544
rect 23180 1372 23240 1538
rect 22654 1300 22660 1360
rect 22720 1300 22726 1360
rect 23174 1312 23180 1372
rect 23240 1312 23246 1372
rect 21636 1198 21642 1258
rect 21702 1198 21708 1258
rect 23672 1198 23678 1258
rect 23738 1198 23744 1258
rect 20920 1054 21408 1060
rect 20920 1020 20932 1054
rect 21396 1020 21408 1054
rect 20920 1014 21408 1020
rect 19654 394 19660 914
rect 19614 382 19660 394
rect 20624 394 20638 970
rect 20672 394 20684 970
rect 21642 970 21702 1198
rect 22654 1094 22660 1154
rect 22720 1094 22726 1154
rect 21938 1054 22426 1060
rect 21938 1020 21950 1054
rect 22414 1020 22426 1054
rect 21938 1014 22426 1020
rect 21642 910 21656 970
rect 21650 430 21656 910
rect 19902 344 20390 350
rect 19902 310 19914 344
rect 20378 310 20390 344
rect 19902 304 20390 310
rect 19482 196 19488 256
rect 19548 196 19554 256
rect 19154 92 19160 152
rect 19220 92 19226 152
rect 19488 -74 19548 196
rect 20624 152 20684 394
rect 21644 394 21656 430
rect 21690 910 21702 970
rect 22660 970 22720 1094
rect 22956 1054 23444 1060
rect 22956 1020 22968 1054
rect 23432 1020 23444 1054
rect 22956 1014 23444 1020
rect 22660 916 22674 970
rect 21690 430 21696 910
rect 22668 434 22674 916
rect 21690 394 21704 430
rect 20920 344 21408 350
rect 20920 310 20932 344
rect 21396 310 21408 344
rect 20920 304 21408 310
rect 20618 92 20624 152
rect 20684 92 20690 152
rect 21132 46 21192 304
rect 21126 -14 21132 46
rect 21192 -14 21198 46
rect 19488 -134 20688 -74
rect 18104 -968 18110 -908
rect 18170 -968 18176 -908
rect 19488 -986 19548 -134
rect 19608 -262 19668 -134
rect 20094 -172 20154 -134
rect 19902 -178 20390 -172
rect 19902 -212 19914 -178
rect 20378 -212 20390 -178
rect 19902 -218 20390 -212
rect 19608 -334 19620 -262
rect 19614 -838 19620 -334
rect 19654 -334 19668 -262
rect 20628 -262 20688 -134
rect 21132 -172 21192 -14
rect 21644 -64 21704 394
rect 22658 394 22674 434
rect 22708 916 22720 970
rect 23678 970 23738 1198
rect 24180 1060 24240 1538
rect 24698 1258 24758 1628
rect 25722 1628 25728 2144
rect 25762 2144 25770 2204
rect 26730 2204 26790 2342
rect 27232 2294 27292 2558
rect 27578 2522 27638 2676
rect 27572 2462 27578 2522
rect 27638 2462 27644 2522
rect 27748 2468 27754 2528
rect 27814 2468 27820 2528
rect 27028 2288 27516 2294
rect 27028 2254 27040 2288
rect 27504 2254 27516 2288
rect 27028 2248 27516 2254
rect 26730 2164 26746 2204
rect 25762 1628 25768 2144
rect 26740 1694 26746 2164
rect 25722 1616 25768 1628
rect 26734 1628 26746 1694
rect 26780 2164 26790 2204
rect 27754 2204 27814 2468
rect 28270 2466 28330 2770
rect 29284 2630 29344 2770
rect 29790 2736 29850 2860
rect 30812 2860 30818 3398
rect 30852 3398 30866 3436
rect 31830 3436 31876 3448
rect 30852 2860 30858 3398
rect 31830 2930 31836 3436
rect 30812 2848 30858 2860
rect 31822 2860 31836 2930
rect 31870 2930 31876 3436
rect 32838 3436 32898 3790
rect 33196 3644 33256 3902
rect 33386 3752 33446 4004
rect 34362 3752 34422 4004
rect 33380 3692 33386 3752
rect 33446 3692 33452 3752
rect 34356 3692 34362 3752
rect 34422 3692 34428 3752
rect 34876 3640 34936 4094
rect 35902 4094 35908 4604
rect 35942 4604 35952 4670
rect 36920 4670 36966 4682
rect 35942 4094 35948 4604
rect 36920 4138 36926 4670
rect 35902 4082 35948 4094
rect 36914 4094 36926 4138
rect 36960 4138 36966 4670
rect 37930 4670 37990 5020
rect 38448 4966 38508 5238
rect 38950 5146 39010 5328
rect 39964 5328 39980 5362
rect 40014 5362 40020 5904
rect 40014 5328 40024 5362
rect 39244 5278 39732 5284
rect 39244 5244 39256 5278
rect 39720 5244 39732 5278
rect 39244 5238 39732 5244
rect 39458 5146 39518 5238
rect 39964 5146 40024 5328
rect 38950 5086 40024 5146
rect 38442 4906 38448 4966
rect 38508 4906 38514 4966
rect 38946 4804 38952 4864
rect 39012 4804 39018 4864
rect 38226 4754 38714 4760
rect 38226 4720 38238 4754
rect 38702 4720 38714 4754
rect 38226 4714 38714 4720
rect 37930 4618 37944 4670
rect 37938 4144 37944 4618
rect 36960 4094 36974 4138
rect 35172 4044 35660 4050
rect 35172 4010 35184 4044
rect 35648 4010 35660 4044
rect 35172 4004 35660 4010
rect 36190 4044 36678 4050
rect 36190 4010 36202 4044
rect 36666 4010 36678 4044
rect 36190 4004 36678 4010
rect 35378 3752 35438 4004
rect 36914 3962 36974 4094
rect 37932 4094 37944 4144
rect 37978 4618 37990 4670
rect 38952 4670 39012 4804
rect 39244 4754 39732 4760
rect 39244 4720 39256 4754
rect 39720 4720 39732 4754
rect 39244 4714 39732 4720
rect 38952 4636 38962 4670
rect 37978 4144 37984 4618
rect 37978 4094 37992 4144
rect 38956 4138 38962 4636
rect 37208 4044 37696 4050
rect 37208 4010 37220 4044
rect 37684 4010 37696 4044
rect 37208 4004 37696 4010
rect 36908 3902 36914 3962
rect 36974 3902 36980 3962
rect 35372 3692 35378 3752
rect 35438 3692 35444 3752
rect 37398 3692 37404 3752
rect 37464 3692 37470 3752
rect 33196 3578 33256 3584
rect 34870 3580 34876 3640
rect 34936 3580 34942 3640
rect 36906 3580 36912 3640
rect 36972 3580 36978 3640
rect 33136 3520 33624 3526
rect 33136 3486 33148 3520
rect 33612 3486 33624 3520
rect 33136 3480 33624 3486
rect 34154 3520 34642 3526
rect 34154 3486 34166 3520
rect 34630 3486 34642 3520
rect 34154 3480 34642 3486
rect 32838 3394 32854 3436
rect 31870 2860 31882 2930
rect 30082 2810 30570 2816
rect 30082 2776 30094 2810
rect 30558 2776 30570 2810
rect 30082 2770 30570 2776
rect 31100 2810 31588 2816
rect 31100 2776 31112 2810
rect 31576 2776 31588 2810
rect 31100 2770 31588 2776
rect 29784 2676 29790 2736
rect 29850 2676 29856 2736
rect 30306 2630 30366 2770
rect 31320 2630 31380 2770
rect 31822 2736 31882 2860
rect 32848 2860 32854 3394
rect 32888 3394 32898 3436
rect 33866 3436 33912 3448
rect 32888 2860 32894 3394
rect 33866 2896 33872 3436
rect 32848 2848 32894 2860
rect 33862 2860 33872 2896
rect 33906 2896 33912 3436
rect 34876 3436 34936 3580
rect 35172 3520 35660 3526
rect 35172 3486 35184 3520
rect 35648 3486 35660 3520
rect 35172 3480 35660 3486
rect 36190 3520 36678 3526
rect 36190 3486 36202 3520
rect 36666 3486 36678 3520
rect 36190 3480 36678 3486
rect 34876 3398 34890 3436
rect 34884 2912 34890 3398
rect 33906 2860 33922 2896
rect 32118 2810 32606 2816
rect 32118 2776 32130 2810
rect 32594 2776 32606 2810
rect 32118 2770 32606 2776
rect 33136 2810 33624 2816
rect 33136 2776 33148 2810
rect 33612 2776 33624 2810
rect 33136 2770 33624 2776
rect 31816 2676 31822 2736
rect 31882 2676 31888 2736
rect 32322 2730 32382 2770
rect 33348 2730 33408 2770
rect 33862 2736 33922 2860
rect 34880 2860 34890 2912
rect 34924 3398 34936 3436
rect 35902 3436 35948 3448
rect 34924 2912 34930 3398
rect 34924 2860 34940 2912
rect 35902 2904 35908 3436
rect 34154 2810 34642 2816
rect 34154 2776 34166 2810
rect 34630 2776 34642 2810
rect 34154 2770 34642 2776
rect 32322 2670 33408 2730
rect 33856 2676 33862 2736
rect 33922 2676 33928 2736
rect 32322 2630 32382 2670
rect 29284 2570 32382 2630
rect 32834 2578 32840 2638
rect 32900 2578 32906 2638
rect 29284 2466 29344 2570
rect 29776 2468 29782 2528
rect 29842 2468 29848 2528
rect 28270 2406 29344 2466
rect 28270 2294 28330 2406
rect 29284 2294 29344 2406
rect 28046 2288 28534 2294
rect 28046 2254 28058 2288
rect 28522 2254 28534 2288
rect 28046 2248 28534 2254
rect 29064 2288 29552 2294
rect 29064 2254 29076 2288
rect 29540 2254 29552 2288
rect 29064 2248 29552 2254
rect 26780 1694 26786 2164
rect 27754 2160 27764 2204
rect 26780 1628 26794 1694
rect 27758 1686 27764 2160
rect 24992 1578 25480 1584
rect 24992 1544 25004 1578
rect 25468 1544 25480 1578
rect 24992 1538 25480 1544
rect 26010 1578 26498 1584
rect 26010 1544 26022 1578
rect 26486 1544 26498 1578
rect 26010 1538 26498 1544
rect 24692 1198 24698 1258
rect 24758 1198 24764 1258
rect 25202 1060 25262 1538
rect 25708 1198 25714 1258
rect 25774 1198 25780 1258
rect 23974 1054 24462 1060
rect 23974 1020 23986 1054
rect 24450 1020 24462 1054
rect 23974 1014 24462 1020
rect 24992 1054 25480 1060
rect 24992 1020 25004 1054
rect 25468 1020 25480 1054
rect 24992 1014 25480 1020
rect 23678 920 23692 970
rect 22708 434 22714 916
rect 22708 394 22718 434
rect 23686 418 23692 920
rect 21938 344 22426 350
rect 21938 310 21950 344
rect 22414 310 22426 344
rect 21938 304 22426 310
rect 22152 46 22212 304
rect 22658 256 22718 394
rect 23680 394 23692 418
rect 23726 920 23738 970
rect 24704 970 24750 982
rect 23726 418 23732 920
rect 23726 394 23740 418
rect 24704 408 24710 970
rect 22956 344 23444 350
rect 22956 310 22968 344
rect 23432 310 23444 344
rect 22956 304 23444 310
rect 22652 196 22658 256
rect 22718 196 22724 256
rect 22658 92 22664 152
rect 22724 92 22730 152
rect 22146 -14 22152 46
rect 22212 -14 22218 46
rect 21638 -124 21644 -64
rect 21704 -124 21710 -64
rect 20920 -178 21408 -172
rect 20920 -212 20932 -178
rect 21396 -212 21408 -178
rect 20920 -218 21408 -212
rect 19654 -838 19660 -334
rect 20628 -338 20638 -262
rect 20632 -790 20638 -338
rect 19614 -850 19660 -838
rect 20624 -838 20638 -790
rect 20672 -338 20688 -262
rect 21644 -262 21704 -124
rect 22152 -172 22212 -14
rect 21938 -178 22426 -172
rect 21938 -212 21950 -178
rect 22414 -212 22426 -178
rect 21938 -218 22426 -212
rect 20672 -790 20678 -338
rect 20672 -838 20684 -790
rect 19902 -888 20390 -882
rect 19902 -922 19914 -888
rect 20378 -922 20390 -888
rect 19902 -928 20390 -922
rect 20624 -986 20684 -838
rect 21644 -838 21656 -262
rect 21690 -838 21704 -262
rect 22664 -262 22724 92
rect 23176 46 23236 304
rect 23170 -14 23176 46
rect 23236 -14 23242 46
rect 23176 -172 23236 -14
rect 23680 -64 23740 394
rect 24694 394 24710 408
rect 24744 408 24750 970
rect 25714 970 25774 1198
rect 26214 1060 26274 1538
rect 26734 1258 26794 1628
rect 27746 1628 27764 1686
rect 27798 2160 27814 2204
rect 28776 2204 28822 2216
rect 27798 1686 27804 2160
rect 27798 1628 27806 1686
rect 28776 1680 28782 2204
rect 27028 1578 27516 1584
rect 27028 1544 27040 1578
rect 27504 1544 27516 1578
rect 27028 1538 27516 1544
rect 26728 1198 26734 1258
rect 26794 1198 26800 1258
rect 27244 1060 27304 1538
rect 27746 1426 27806 1628
rect 28764 1628 28782 1680
rect 28816 1680 28822 2204
rect 29782 2204 29842 2468
rect 30306 2294 30366 2570
rect 31320 2294 31380 2570
rect 31820 2468 31826 2528
rect 31886 2468 31892 2528
rect 30082 2288 30570 2294
rect 30082 2254 30094 2288
rect 30558 2254 30570 2288
rect 30082 2248 30570 2254
rect 31100 2288 31588 2294
rect 31100 2254 31112 2288
rect 31576 2254 31588 2288
rect 31100 2248 31588 2254
rect 29782 2160 29800 2204
rect 28816 1628 28824 1680
rect 28046 1578 28534 1584
rect 28046 1544 28058 1578
rect 28522 1544 28534 1578
rect 28046 1538 28534 1544
rect 27596 1366 27806 1426
rect 28260 1372 28320 1538
rect 28764 1486 28824 1628
rect 29794 1628 29800 2160
rect 29834 2160 29842 2204
rect 30812 2204 30858 2216
rect 29834 1628 29840 2160
rect 30812 1680 30818 2204
rect 29794 1616 29840 1628
rect 30806 1628 30818 1680
rect 30852 1680 30858 2204
rect 31826 2204 31886 2468
rect 32322 2294 32382 2570
rect 32118 2288 32606 2294
rect 32118 2254 32130 2288
rect 32594 2254 32606 2288
rect 32118 2248 32606 2254
rect 31826 2156 31836 2204
rect 30852 1628 30866 1680
rect 29064 1578 29552 1584
rect 29064 1544 29076 1578
rect 29540 1544 29552 1578
rect 29064 1538 29552 1544
rect 30082 1578 30570 1584
rect 30082 1544 30094 1578
rect 30558 1544 30570 1578
rect 30082 1538 30570 1544
rect 30806 1486 30866 1628
rect 31830 1628 31836 2156
rect 31870 2156 31886 2204
rect 32840 2204 32900 2578
rect 33348 2294 33408 2670
rect 33848 2468 33854 2528
rect 33914 2468 33920 2528
rect 33136 2288 33624 2294
rect 33136 2254 33148 2288
rect 33612 2254 33624 2288
rect 33136 2248 33624 2254
rect 32840 2168 32854 2204
rect 31870 1628 31876 2156
rect 32848 1672 32854 2168
rect 31830 1616 31876 1628
rect 32842 1628 32854 1672
rect 32888 2168 32900 2204
rect 33854 2204 33914 2468
rect 34368 2294 34428 2770
rect 34880 2402 34940 2860
rect 35892 2860 35908 2904
rect 35942 2904 35948 3436
rect 36912 3436 36972 3580
rect 37404 3526 37464 3692
rect 37208 3520 37696 3526
rect 37208 3486 37220 3520
rect 37684 3486 37696 3520
rect 37208 3480 37696 3486
rect 36912 3378 36926 3436
rect 35942 2860 35952 2904
rect 36920 2900 36926 3378
rect 35172 2810 35660 2816
rect 35172 2776 35184 2810
rect 35648 2776 35660 2810
rect 35172 2770 35660 2776
rect 34874 2342 34880 2402
rect 34940 2342 34946 2402
rect 34154 2288 34642 2294
rect 34154 2254 34166 2288
rect 34630 2254 34642 2288
rect 34154 2248 34642 2254
rect 32888 1672 32894 2168
rect 33854 2156 33872 2204
rect 32888 1628 32902 1672
rect 33866 1668 33872 2156
rect 31100 1578 31588 1584
rect 31100 1544 31112 1578
rect 31576 1544 31588 1578
rect 31100 1538 31588 1544
rect 32118 1578 32606 1584
rect 32118 1544 32130 1578
rect 32594 1544 32606 1578
rect 32118 1538 32606 1544
rect 32842 1486 32902 1628
rect 33856 1628 33872 1668
rect 33906 2156 33914 2204
rect 34880 2204 34940 2342
rect 35384 2294 35444 2770
rect 35892 2528 35952 2860
rect 36910 2860 36926 2900
rect 36960 3378 36972 3436
rect 37932 3436 37992 4094
rect 38948 4094 38962 4138
rect 38996 4636 39012 4670
rect 39974 4670 40020 4682
rect 38996 4138 39002 4636
rect 38996 4094 39008 4138
rect 39974 4124 39980 4670
rect 38226 4044 38714 4050
rect 38226 4010 38238 4044
rect 38702 4010 38714 4044
rect 38226 4004 38714 4010
rect 38434 3752 38494 4004
rect 38948 3912 39008 4094
rect 39964 4094 39980 4124
rect 40014 4124 40020 4670
rect 40014 4094 40024 4124
rect 39244 4044 39732 4050
rect 39244 4010 39256 4044
rect 39720 4010 39732 4044
rect 39244 4004 39732 4010
rect 39454 3912 39514 4004
rect 39964 3912 40024 4094
rect 38948 3852 40024 3912
rect 38428 3692 38434 3752
rect 38494 3692 38500 3752
rect 38948 3640 39008 3852
rect 38942 3580 38948 3640
rect 39008 3580 39014 3640
rect 38226 3520 38714 3526
rect 38226 3486 38238 3520
rect 38702 3486 38714 3520
rect 38226 3480 38714 3486
rect 39244 3520 39732 3526
rect 39244 3486 39256 3520
rect 39720 3486 39732 3520
rect 39244 3480 39732 3486
rect 37932 3394 37944 3436
rect 36960 2900 36966 3378
rect 37938 2914 37944 3394
rect 36960 2860 36970 2900
rect 36190 2810 36678 2816
rect 36190 2776 36202 2810
rect 36666 2776 36678 2810
rect 36190 2770 36678 2776
rect 35886 2468 35892 2528
rect 35952 2468 35958 2528
rect 36418 2294 36478 2770
rect 36910 2402 36970 2860
rect 37932 2860 37944 2914
rect 37978 3394 37992 3436
rect 38956 3436 39002 3448
rect 37978 2914 37984 3394
rect 37978 2860 37992 2914
rect 38956 2906 38962 3436
rect 37208 2810 37696 2816
rect 37208 2776 37220 2810
rect 37684 2776 37696 2810
rect 37208 2770 37696 2776
rect 37436 2404 37496 2770
rect 37932 2528 37992 2860
rect 38946 2860 38962 2906
rect 38996 2906 39002 3436
rect 39974 3436 40020 3448
rect 38996 2860 39006 2906
rect 39974 2888 39980 3436
rect 38226 2810 38714 2816
rect 38226 2776 38238 2810
rect 38702 2776 38714 2810
rect 38226 2770 38714 2776
rect 38450 2532 38510 2770
rect 38946 2734 39006 2860
rect 39966 2860 39980 2888
rect 40014 2888 40020 3436
rect 40014 2860 40026 2888
rect 39244 2810 39732 2816
rect 39244 2776 39256 2810
rect 39720 2776 39732 2810
rect 39244 2770 39732 2776
rect 39452 2736 39512 2770
rect 39966 2736 40026 2860
rect 39452 2734 40026 2736
rect 38946 2674 40026 2734
rect 38946 2638 39006 2674
rect 38940 2578 38946 2638
rect 39006 2578 39012 2638
rect 37926 2468 37932 2528
rect 37992 2468 37998 2528
rect 38444 2472 38450 2532
rect 38510 2472 38516 2532
rect 39956 2472 39962 2532
rect 40022 2472 40028 2532
rect 36904 2342 36910 2402
rect 36970 2342 36976 2402
rect 35172 2288 35660 2294
rect 35172 2254 35184 2288
rect 35648 2254 35660 2288
rect 35172 2248 35660 2254
rect 36190 2288 36678 2294
rect 36190 2254 36202 2288
rect 36666 2254 36678 2288
rect 36190 2248 36678 2254
rect 34880 2158 34890 2204
rect 33906 1668 33912 2156
rect 34884 1688 34890 2158
rect 33906 1628 33916 1668
rect 33136 1578 33624 1584
rect 33136 1544 33148 1578
rect 33612 1544 33624 1578
rect 33136 1538 33624 1544
rect 28758 1426 28764 1486
rect 28824 1426 28830 1486
rect 30800 1426 30806 1486
rect 30866 1426 30872 1486
rect 32836 1426 32842 1486
rect 32902 1426 32908 1486
rect 33348 1376 33408 1538
rect 33856 1478 33916 1628
rect 34878 1628 34890 1688
rect 34924 2158 34940 2204
rect 35902 2204 35948 2216
rect 34924 1688 34930 2158
rect 34924 1628 34938 1688
rect 35902 1672 35908 2204
rect 34154 1578 34642 1584
rect 34154 1544 34166 1578
rect 34630 1544 34642 1578
rect 34154 1538 34642 1544
rect 33856 1418 34062 1478
rect 27596 1154 27656 1366
rect 28254 1312 28260 1372
rect 28320 1312 28326 1372
rect 33342 1316 33348 1376
rect 33408 1316 33414 1376
rect 27746 1198 27752 1258
rect 27812 1198 27818 1258
rect 29776 1198 29782 1258
rect 29842 1198 29848 1258
rect 31814 1198 31820 1258
rect 31880 1198 31886 1258
rect 33850 1198 33856 1258
rect 33916 1198 33922 1258
rect 27590 1094 27596 1154
rect 27656 1094 27662 1154
rect 26010 1054 26498 1060
rect 26010 1020 26022 1054
rect 26486 1020 26498 1054
rect 26010 1014 26498 1020
rect 27028 1054 27516 1060
rect 27028 1020 27040 1054
rect 27504 1020 27516 1054
rect 27028 1014 27516 1020
rect 25714 488 25728 970
rect 25722 414 25728 488
rect 24744 394 24754 408
rect 23974 344 24462 350
rect 23974 310 23986 344
rect 24450 310 24462 344
rect 23974 304 24462 310
rect 24194 46 24254 304
rect 24694 152 24754 394
rect 25718 394 25728 414
rect 25762 488 25774 970
rect 26740 970 26786 982
rect 25762 414 25768 488
rect 26740 420 26746 970
rect 25762 394 25778 414
rect 24992 344 25480 350
rect 24992 310 25004 344
rect 25468 310 25480 344
rect 24992 304 25480 310
rect 24688 92 24694 152
rect 24754 92 24760 152
rect 25208 46 25268 304
rect 24188 -14 24194 46
rect 24254 -14 24260 46
rect 25202 -14 25208 46
rect 25268 -14 25274 46
rect 23674 -124 23680 -64
rect 23740 -124 23746 -64
rect 22956 -178 23444 -172
rect 22956 -212 22968 -178
rect 23432 -212 23444 -178
rect 22956 -218 23444 -212
rect 22664 -276 22674 -262
rect 20920 -888 21408 -882
rect 20920 -922 20932 -888
rect 21396 -922 21408 -888
rect 20920 -928 21408 -922
rect 19482 -1046 19488 -986
rect 19548 -1046 19554 -986
rect 20618 -1046 20624 -986
rect 20684 -1046 20690 -986
rect 21136 -1094 21196 -928
rect 21130 -1154 21136 -1094
rect 21196 -1154 21202 -1094
rect 21644 -1350 21704 -838
rect 22668 -838 22674 -276
rect 22708 -276 22724 -262
rect 23680 -262 23740 -124
rect 24194 -172 24254 -14
rect 25208 -172 25268 -14
rect 25718 -64 25778 394
rect 26734 394 26746 420
rect 26780 420 26786 970
rect 27752 970 27812 1198
rect 28046 1054 28534 1060
rect 28046 1020 28058 1054
rect 28522 1020 28534 1054
rect 28046 1014 28534 1020
rect 29064 1054 29552 1060
rect 29064 1020 29076 1054
rect 29540 1020 29552 1054
rect 29064 1014 29552 1020
rect 28776 970 28822 982
rect 29782 970 29842 1198
rect 30082 1054 30570 1060
rect 30082 1020 30094 1054
rect 30558 1020 30570 1054
rect 30082 1014 30570 1020
rect 31100 1054 31588 1060
rect 31100 1020 31112 1054
rect 31576 1020 31588 1054
rect 31100 1014 31588 1020
rect 30812 970 30858 982
rect 31820 970 31880 1198
rect 32118 1054 32606 1060
rect 32118 1020 32130 1054
rect 32594 1020 32606 1054
rect 32118 1014 32606 1020
rect 33136 1054 33624 1060
rect 33136 1020 33148 1054
rect 33612 1020 33624 1054
rect 33136 1014 33624 1020
rect 27752 914 27764 970
rect 26780 394 26794 420
rect 27758 418 27764 914
rect 26010 344 26498 350
rect 26010 310 26022 344
rect 26486 310 26498 344
rect 26010 304 26498 310
rect 26240 46 26300 304
rect 26734 152 26794 394
rect 27756 394 27764 418
rect 27798 914 27812 970
rect 28770 934 28782 970
rect 27798 418 27804 914
rect 28776 446 28782 934
rect 27798 394 27816 418
rect 27028 344 27516 350
rect 27028 310 27040 344
rect 27504 310 27516 344
rect 27028 304 27516 310
rect 26882 198 26888 258
rect 26948 198 26954 258
rect 26728 92 26734 152
rect 26794 92 26800 152
rect 26234 -14 26240 46
rect 26300 -14 26306 46
rect 26888 14 26948 198
rect 27252 46 27312 304
rect 25712 -124 25718 -64
rect 25778 -124 25784 -64
rect 23974 -178 24462 -172
rect 23974 -212 23986 -178
rect 24450 -212 24462 -178
rect 23974 -218 24462 -212
rect 24992 -178 25480 -172
rect 24992 -212 25004 -178
rect 25468 -212 25480 -178
rect 24992 -218 25480 -212
rect 22708 -838 22714 -276
rect 22668 -850 22714 -838
rect 23680 -838 23692 -262
rect 23726 -838 23740 -262
rect 24704 -262 24750 -250
rect 24704 -796 24710 -262
rect 21938 -888 22426 -882
rect 21938 -922 21950 -888
rect 22414 -922 22426 -888
rect 21938 -928 22426 -922
rect 22956 -888 23444 -882
rect 22956 -922 22968 -888
rect 23432 -922 23444 -888
rect 22956 -928 23444 -922
rect 22150 -1094 22210 -928
rect 22150 -1160 22210 -1154
rect 23172 -1094 23232 -928
rect 23172 -1160 23232 -1154
rect 23680 -1350 23740 -838
rect 24694 -838 24710 -796
rect 24744 -796 24750 -262
rect 25718 -262 25778 -124
rect 26240 -172 26300 -14
rect 26732 -46 26948 14
rect 27246 -14 27252 46
rect 27312 -14 27318 46
rect 26010 -178 26498 -172
rect 26010 -212 26022 -178
rect 26486 -212 26498 -178
rect 26010 -218 26498 -212
rect 24744 -838 24754 -796
rect 23974 -888 24462 -882
rect 23974 -922 23986 -888
rect 24450 -922 24462 -888
rect 23974 -928 24462 -922
rect 24184 -1088 24244 -928
rect 24694 -986 24754 -838
rect 25718 -838 25728 -262
rect 25762 -838 25778 -262
rect 26732 -262 26792 -46
rect 27252 -172 27312 -14
rect 27756 -64 27816 394
rect 28766 394 28782 446
rect 28816 934 28830 970
rect 28816 446 28822 934
rect 29782 920 29800 970
rect 28816 394 28826 446
rect 29794 424 29800 920
rect 28046 344 28534 350
rect 28046 310 28058 344
rect 28522 310 28534 344
rect 28046 304 28534 310
rect 28260 46 28320 304
rect 28766 258 28826 394
rect 29792 394 29800 424
rect 29834 920 29842 970
rect 30806 938 30818 970
rect 29834 424 29840 920
rect 30812 434 30818 938
rect 29834 394 29852 424
rect 29064 344 29552 350
rect 29064 310 29076 344
rect 29540 310 29552 344
rect 29064 304 29552 310
rect 28760 198 28766 258
rect 28826 198 28832 258
rect 28764 92 28770 152
rect 28830 92 28836 152
rect 28254 -14 28260 46
rect 28320 -14 28326 46
rect 27750 -124 27756 -64
rect 27816 -124 27822 -64
rect 27028 -178 27516 -172
rect 27028 -212 27040 -178
rect 27504 -212 27516 -178
rect 27028 -218 27516 -212
rect 26732 -288 26746 -262
rect 24992 -888 25480 -882
rect 24992 -922 25004 -888
rect 25468 -922 25480 -888
rect 24992 -928 25480 -922
rect 24688 -1046 24694 -986
rect 24754 -1046 24760 -986
rect 25210 -1088 25270 -928
rect 24184 -1094 24246 -1088
rect 24184 -1100 24186 -1094
rect 25210 -1094 25272 -1088
rect 25210 -1100 25212 -1094
rect 24186 -1160 24246 -1154
rect 25212 -1160 25272 -1154
rect 25718 -1350 25778 -838
rect 26740 -838 26746 -288
rect 26780 -288 26792 -262
rect 27756 -262 27816 -124
rect 28260 -172 28320 -14
rect 28046 -178 28534 -172
rect 28046 -212 28058 -178
rect 28522 -212 28534 -178
rect 28046 -218 28534 -212
rect 26780 -838 26786 -288
rect 26740 -850 26786 -838
rect 27756 -838 27764 -262
rect 27798 -838 27816 -262
rect 28770 -262 28830 92
rect 29278 46 29338 304
rect 29272 -14 29278 46
rect 29338 -14 29344 46
rect 29278 -172 29338 -14
rect 29792 -64 29852 394
rect 30804 394 30818 434
rect 30852 938 30866 970
rect 30852 434 30858 938
rect 31820 926 31836 970
rect 30852 394 30864 434
rect 31830 418 31836 926
rect 30082 344 30570 350
rect 30082 310 30094 344
rect 30558 310 30570 344
rect 30082 304 30570 310
rect 30304 46 30364 304
rect 30804 258 30864 394
rect 31828 394 31836 418
rect 31870 926 31880 970
rect 32848 970 32894 982
rect 31870 418 31876 926
rect 32848 440 32854 970
rect 31870 394 31888 418
rect 31100 344 31588 350
rect 31100 310 31112 344
rect 31576 310 31588 344
rect 31100 304 31588 310
rect 30798 198 30804 258
rect 30864 198 30870 258
rect 30800 92 30806 152
rect 30866 92 30872 152
rect 30298 -14 30304 46
rect 30364 -14 30370 46
rect 29786 -124 29792 -64
rect 29852 -124 29858 -64
rect 29064 -178 29552 -172
rect 29064 -212 29076 -178
rect 29540 -212 29552 -178
rect 29064 -218 29552 -212
rect 28770 -288 28782 -262
rect 26010 -888 26498 -882
rect 26010 -922 26022 -888
rect 26486 -922 26498 -888
rect 26010 -928 26498 -922
rect 27028 -888 27516 -882
rect 27028 -922 27040 -888
rect 27504 -922 27516 -888
rect 27028 -928 27516 -922
rect 26224 -1094 26284 -928
rect 26224 -1160 26284 -1154
rect 27260 -1094 27320 -928
rect 27260 -1160 27320 -1154
rect 27756 -1350 27816 -838
rect 28776 -838 28782 -288
rect 28816 -288 28830 -262
rect 29792 -262 29852 -124
rect 30304 -172 30364 -14
rect 30082 -178 30570 -172
rect 30082 -212 30094 -178
rect 30558 -212 30570 -178
rect 30082 -218 30570 -212
rect 28816 -838 28822 -288
rect 28776 -850 28822 -838
rect 29792 -838 29800 -262
rect 29834 -838 29852 -262
rect 30806 -262 30866 92
rect 31306 46 31366 304
rect 31300 -14 31306 46
rect 31366 -14 31372 46
rect 31306 -172 31366 -14
rect 31828 -64 31888 394
rect 32840 394 32854 440
rect 32888 440 32894 970
rect 33856 970 33916 1198
rect 34002 1154 34062 1418
rect 33996 1094 34002 1154
rect 34062 1094 34068 1154
rect 34366 1060 34426 1538
rect 34878 1258 34938 1628
rect 35896 1628 35908 1672
rect 35942 1672 35948 2204
rect 36910 2204 36970 2342
rect 37436 2294 37496 2344
rect 38450 2294 38510 2472
rect 38944 2344 38950 2404
rect 39010 2344 39016 2404
rect 37208 2288 37696 2294
rect 37208 2254 37220 2288
rect 37684 2254 37696 2288
rect 37208 2248 37696 2254
rect 38226 2288 38714 2294
rect 38226 2254 38238 2288
rect 38702 2254 38714 2288
rect 38226 2248 38714 2254
rect 36910 2158 36926 2204
rect 36920 1676 36926 2158
rect 35942 1628 35956 1672
rect 35172 1578 35660 1584
rect 35172 1544 35184 1578
rect 35648 1544 35660 1578
rect 35172 1538 35660 1544
rect 34872 1198 34878 1258
rect 34938 1198 34944 1258
rect 35386 1060 35446 1538
rect 35896 1486 35956 1628
rect 36912 1628 36926 1676
rect 36960 2158 36970 2204
rect 37938 2204 37984 2216
rect 38950 2204 39010 2344
rect 39244 2288 39732 2294
rect 39244 2254 39256 2288
rect 39720 2254 39732 2288
rect 39244 2248 39732 2254
rect 36960 1676 36966 2158
rect 36960 1628 36972 1676
rect 37938 1672 37944 2204
rect 36190 1578 36678 1584
rect 36190 1544 36202 1578
rect 36666 1544 36678 1578
rect 36190 1538 36678 1544
rect 35890 1426 35896 1486
rect 35956 1426 35962 1486
rect 35892 1198 35898 1258
rect 35958 1198 35964 1258
rect 34154 1054 34642 1060
rect 34154 1020 34166 1054
rect 34630 1020 34642 1054
rect 34154 1014 34642 1020
rect 35172 1054 35660 1060
rect 35172 1020 35184 1054
rect 35648 1020 35660 1054
rect 35172 1014 35660 1020
rect 33856 926 33872 970
rect 32888 394 32900 440
rect 33866 420 33872 926
rect 32118 344 32606 350
rect 32118 310 32130 344
rect 32594 310 32606 344
rect 32118 304 32606 310
rect 32326 46 32386 304
rect 32668 198 32674 258
rect 32734 198 32740 258
rect 32320 -14 32326 46
rect 32386 -14 32392 46
rect 32674 6 32734 198
rect 32840 152 32900 394
rect 33860 394 33872 420
rect 33906 926 33916 970
rect 34884 970 34930 982
rect 33906 420 33912 926
rect 34884 434 34890 970
rect 33906 394 33920 420
rect 33136 344 33624 350
rect 33136 310 33148 344
rect 33612 310 33624 344
rect 33136 304 33624 310
rect 32834 92 32840 152
rect 32900 92 32906 152
rect 33346 46 33406 304
rect 31822 -124 31828 -64
rect 31888 -124 31894 -64
rect 31100 -178 31588 -172
rect 31100 -212 31112 -178
rect 31576 -212 31588 -178
rect 31100 -218 31588 -212
rect 30806 -298 30818 -262
rect 28046 -888 28534 -882
rect 28046 -922 28058 -888
rect 28522 -922 28534 -888
rect 28046 -928 28534 -922
rect 29064 -888 29552 -882
rect 29064 -922 29076 -888
rect 29540 -922 29552 -888
rect 29064 -928 29552 -922
rect 28266 -1094 28326 -928
rect 29280 -1094 29340 -928
rect 29274 -1154 29280 -1094
rect 29340 -1154 29346 -1094
rect 28266 -1160 28326 -1154
rect 29792 -1350 29852 -838
rect 30812 -838 30818 -298
rect 30852 -298 30866 -262
rect 31828 -262 31888 -124
rect 32326 -172 32386 -14
rect 32674 -54 32900 6
rect 33340 -14 33346 46
rect 33406 -14 33412 46
rect 32118 -178 32606 -172
rect 32118 -212 32130 -178
rect 32594 -212 32606 -178
rect 32118 -218 32606 -212
rect 30852 -838 30858 -298
rect 30812 -850 30858 -838
rect 31828 -838 31836 -262
rect 31870 -838 31888 -262
rect 32840 -262 32900 -54
rect 33346 -172 33406 -14
rect 33860 -64 33920 394
rect 34880 394 34890 434
rect 34924 434 34930 970
rect 35898 970 35958 1198
rect 36400 1060 36460 1538
rect 36912 1258 36972 1628
rect 37928 1628 37944 1672
rect 37978 1672 37984 2204
rect 38948 2170 38962 2204
rect 38950 2160 38962 2170
rect 37978 1628 37988 1672
rect 37208 1578 37696 1584
rect 37208 1544 37220 1578
rect 37684 1544 37696 1578
rect 37208 1538 37696 1544
rect 36906 1198 36912 1258
rect 36972 1198 36978 1258
rect 36906 1094 36912 1154
rect 36972 1094 36978 1154
rect 36190 1054 36678 1060
rect 36190 1020 36202 1054
rect 36666 1020 36678 1054
rect 36190 1014 36678 1020
rect 36408 1010 36468 1014
rect 35898 904 35908 970
rect 35902 440 35908 904
rect 34924 394 34940 434
rect 34154 344 34642 350
rect 34154 310 34166 344
rect 34630 310 34642 344
rect 34154 304 34642 310
rect 34372 46 34432 304
rect 34880 152 34940 394
rect 35892 394 35908 440
rect 35942 904 35958 970
rect 36912 970 36972 1094
rect 37436 1060 37496 1538
rect 37928 1486 37988 1628
rect 38956 1628 38962 2160
rect 38996 2160 39010 2204
rect 39962 2204 40022 2472
rect 38996 1628 39002 2160
rect 39962 2150 39980 2204
rect 38956 1616 39002 1628
rect 39974 1628 39980 2150
rect 40014 2166 40026 2204
rect 40014 2150 40022 2166
rect 40014 1628 40020 2150
rect 39974 1616 40020 1628
rect 38226 1578 38714 1584
rect 38226 1544 38238 1578
rect 38702 1544 38714 1578
rect 38226 1538 38714 1544
rect 39244 1578 39732 1584
rect 39244 1544 39256 1578
rect 39720 1544 39732 1578
rect 39244 1538 39732 1544
rect 37922 1426 37928 1486
rect 37988 1426 37994 1486
rect 38448 1376 38508 1538
rect 39456 1376 39516 1538
rect 40074 1486 40134 7276
rect 40196 6362 40202 6422
rect 40262 6362 40268 6422
rect 40202 4864 40262 6362
rect 40318 6098 40378 7390
rect 40434 6140 40440 6200
rect 40500 6140 40506 6200
rect 40312 6038 40318 6098
rect 40378 6038 40384 6098
rect 40196 4804 40202 4864
rect 40262 4804 40268 4864
rect 40192 3902 40198 3962
rect 40258 3902 40264 3962
rect 40198 2638 40258 3902
rect 40318 2736 40378 6038
rect 40312 2676 40318 2736
rect 40378 2676 40384 2736
rect 40192 2578 40198 2638
rect 40258 2578 40264 2638
rect 40068 1426 40074 1486
rect 40134 1426 40140 1486
rect 38442 1316 38448 1376
rect 38508 1316 38514 1376
rect 39450 1316 39456 1376
rect 39516 1316 39522 1376
rect 40318 1260 40378 2676
rect 40440 2404 40500 6140
rect 40568 4972 40628 7494
rect 40566 4966 40628 4972
rect 40626 4906 40628 4966
rect 40566 4900 40628 4906
rect 40568 2532 40628 4900
rect 40562 2472 40568 2532
rect 40628 2472 40634 2532
rect 40434 2344 40440 2404
rect 40500 2344 40506 2404
rect 40690 1376 40750 12304
rect 40796 8494 40802 8554
rect 40862 8494 40868 8554
rect 40684 1316 40690 1376
rect 40750 1316 40756 1376
rect 37928 1198 37934 1258
rect 37994 1198 38000 1258
rect 38950 1200 40378 1260
rect 37208 1054 37696 1060
rect 37208 1020 37220 1054
rect 37684 1020 37696 1054
rect 37208 1014 37696 1020
rect 36912 924 36926 970
rect 35942 440 35948 904
rect 35942 394 35952 440
rect 35172 344 35660 350
rect 35172 310 35184 344
rect 35648 310 35660 344
rect 35172 304 35660 310
rect 34874 92 34880 152
rect 34940 92 34946 152
rect 35390 46 35450 304
rect 34366 -14 34372 46
rect 34432 -14 34438 46
rect 35384 -14 35390 46
rect 35450 -14 35456 46
rect 33854 -124 33860 -64
rect 33920 -124 33926 -64
rect 33136 -178 33624 -172
rect 33136 -212 33148 -178
rect 33612 -212 33624 -178
rect 33136 -218 33624 -212
rect 32840 -298 32854 -262
rect 30082 -888 30570 -882
rect 30082 -922 30094 -888
rect 30558 -922 30570 -888
rect 30082 -928 30570 -922
rect 31100 -888 31588 -882
rect 31100 -922 31112 -888
rect 31576 -922 31588 -888
rect 31100 -928 31588 -922
rect 30296 -1094 30356 -928
rect 31306 -1088 31366 -928
rect 30296 -1160 30356 -1154
rect 31304 -1094 31366 -1088
rect 31364 -1100 31366 -1094
rect 31304 -1160 31364 -1154
rect 31828 -1350 31888 -838
rect 32848 -838 32854 -298
rect 32888 -298 32900 -262
rect 33860 -262 33920 -124
rect 34372 -172 34432 -14
rect 35390 -172 35450 -14
rect 35892 -64 35952 394
rect 36920 394 36926 924
rect 36960 924 36972 970
rect 37934 970 37994 1198
rect 38226 1054 38714 1060
rect 38226 1020 38238 1054
rect 38702 1020 38714 1054
rect 38226 1014 38714 1020
rect 36960 394 36966 924
rect 37934 910 37944 970
rect 37938 418 37944 910
rect 36920 382 36966 394
rect 37932 394 37944 418
rect 37978 910 37994 970
rect 38950 970 39010 1200
rect 39448 1060 39508 1200
rect 39244 1054 39732 1060
rect 39244 1020 39256 1054
rect 39720 1020 39732 1054
rect 39244 1014 39732 1020
rect 37978 418 37984 910
rect 37978 394 37992 418
rect 36190 344 36678 350
rect 36190 310 36202 344
rect 36666 310 36678 344
rect 36190 304 36678 310
rect 37208 344 37696 350
rect 37208 310 37220 344
rect 37684 310 37696 344
rect 37208 304 37696 310
rect 36404 46 36464 304
rect 36904 92 36910 152
rect 36970 92 36976 152
rect 36398 -14 36404 46
rect 36464 -14 36470 46
rect 35886 -124 35892 -64
rect 35952 -124 35958 -64
rect 34154 -178 34642 -172
rect 34154 -212 34166 -178
rect 34630 -212 34642 -178
rect 34154 -218 34642 -212
rect 35172 -178 35660 -172
rect 35172 -212 35184 -178
rect 35648 -212 35660 -178
rect 35172 -218 35660 -212
rect 32888 -838 32894 -298
rect 32848 -850 32894 -838
rect 33860 -838 33872 -262
rect 33906 -838 33920 -262
rect 34884 -262 34930 -250
rect 34884 -786 34890 -262
rect 33344 -882 33404 -880
rect 32118 -888 32606 -882
rect 32118 -922 32130 -888
rect 32594 -922 32606 -888
rect 32118 -928 32606 -922
rect 33136 -888 33624 -882
rect 33136 -922 33148 -888
rect 33612 -922 33624 -888
rect 33136 -928 33624 -922
rect 32322 -1088 32382 -928
rect 32320 -1094 32382 -1088
rect 32380 -1100 32382 -1094
rect 33344 -1094 33404 -928
rect 32320 -1160 32380 -1154
rect 33344 -1160 33404 -1154
rect 33860 -1350 33920 -838
rect 34874 -838 34890 -786
rect 34924 -786 34930 -262
rect 35892 -262 35952 -124
rect 36404 -172 36464 -14
rect 36190 -178 36678 -172
rect 36190 -212 36202 -178
rect 36666 -212 36678 -178
rect 36190 -218 36678 -212
rect 34924 -838 34934 -786
rect 34154 -888 34642 -882
rect 34154 -922 34166 -888
rect 34630 -922 34642 -888
rect 34154 -928 34642 -922
rect 34366 -1094 34426 -928
rect 34874 -986 34934 -838
rect 35892 -838 35908 -262
rect 35942 -838 35952 -262
rect 36910 -262 36970 92
rect 37418 46 37478 304
rect 37412 -14 37418 46
rect 37478 -14 37484 46
rect 37418 -172 37478 -14
rect 37932 -64 37992 394
rect 38950 394 38962 970
rect 38996 394 39010 970
rect 39964 970 40024 1200
rect 40088 1094 40094 1154
rect 40154 1094 40160 1154
rect 39964 916 39980 970
rect 38226 344 38714 350
rect 38226 310 38238 344
rect 38702 310 38714 344
rect 38226 304 38714 310
rect 38440 46 38500 304
rect 38950 258 39010 394
rect 39974 394 39980 916
rect 40014 916 40024 970
rect 40014 394 40020 916
rect 39974 382 40020 394
rect 39244 344 39732 350
rect 39244 310 39256 344
rect 39720 310 39732 344
rect 39244 304 39732 310
rect 38944 198 38950 258
rect 39010 198 39016 258
rect 38944 92 38950 152
rect 39010 92 39016 152
rect 38434 -14 38440 46
rect 38500 -14 38506 46
rect 37926 -124 37932 -64
rect 37992 -124 37998 -64
rect 37208 -178 37696 -172
rect 37208 -212 37220 -178
rect 37684 -212 37696 -178
rect 37208 -218 37696 -212
rect 36910 -306 36926 -262
rect 35172 -888 35660 -882
rect 35172 -922 35184 -888
rect 35648 -922 35660 -888
rect 35172 -928 35660 -922
rect 34868 -1046 34874 -986
rect 34934 -1046 34940 -986
rect 35386 -1088 35446 -928
rect 35386 -1094 35448 -1088
rect 35386 -1100 35388 -1094
rect 34366 -1160 34426 -1154
rect 35388 -1160 35448 -1154
rect 35892 -1350 35952 -838
rect 36920 -838 36926 -306
rect 36960 -306 36970 -262
rect 37932 -262 37992 -124
rect 38440 -172 38500 -14
rect 38950 -64 39010 92
rect 38950 -124 40028 -64
rect 38226 -178 38714 -172
rect 38226 -212 38238 -178
rect 38702 -212 38714 -178
rect 38226 -218 38714 -212
rect 36960 -838 36966 -306
rect 36920 -850 36966 -838
rect 37932 -838 37944 -262
rect 37978 -838 37992 -262
rect 38950 -262 39010 -124
rect 39466 -172 39526 -124
rect 39244 -178 39732 -172
rect 39244 -212 39256 -178
rect 39720 -212 39732 -178
rect 39244 -218 39732 -212
rect 38950 -270 38962 -262
rect 36408 -882 36468 -880
rect 36190 -888 36678 -882
rect 36190 -922 36202 -888
rect 36666 -922 36678 -888
rect 36190 -928 36678 -922
rect 37208 -888 37696 -882
rect 37208 -922 37220 -888
rect 37684 -922 37696 -888
rect 37208 -928 37696 -922
rect 36408 -1088 36468 -928
rect 37422 -1088 37482 -928
rect 36406 -1094 36468 -1088
rect 36466 -1100 36468 -1094
rect 37420 -1094 37482 -1088
rect 36406 -1160 36466 -1154
rect 37480 -1100 37482 -1094
rect 37420 -1160 37480 -1154
rect 37932 -1350 37992 -838
rect 38956 -838 38962 -270
rect 38996 -270 39010 -262
rect 39968 -262 40028 -124
rect 38996 -838 39002 -270
rect 39968 -280 39980 -262
rect 38956 -850 39002 -838
rect 39974 -838 39980 -280
rect 40014 -280 40028 -262
rect 40014 -838 40020 -280
rect 39974 -850 40020 -838
rect 38442 -882 38502 -880
rect 38226 -888 38714 -882
rect 38226 -922 38238 -888
rect 38702 -922 38714 -888
rect 38226 -928 38714 -922
rect 39244 -888 39732 -882
rect 39244 -922 39256 -888
rect 39720 -922 39732 -888
rect 39244 -928 39732 -922
rect 38442 -1088 38502 -928
rect 40094 -986 40154 1094
rect 40802 152 40862 8494
rect 40796 92 40802 152
rect 40862 92 40868 152
rect 40088 -1046 40094 -986
rect 40154 -1046 40160 -986
rect 38442 -1094 38504 -1088
rect 38442 -1100 38444 -1094
rect 38444 -1160 38504 -1154
rect 41856 -1250 41862 13010
rect 41962 -1250 41968 13010
rect 8922 -1396 9072 -1350
rect 9118 -1396 12292 -1350
rect 12352 -1396 18744 -1350
rect 18804 -1396 40846 -1350
rect 40906 -1396 41008 -1350
rect 8922 -1550 8968 -1396
rect 40968 -1550 41008 -1396
rect 8922 -1596 41008 -1550
rect 5424 -2036 5434 -1736
rect 41246 -2036 41256 -1736
rect 41856 -2036 41968 -1250
rect 4712 -2042 41968 -2036
rect 4712 -2142 4818 -2042
rect 41862 -2142 41968 -2042
rect 4712 -2148 41968 -2142
<< via1 >>
rect 17524 28996 18124 29296
rect 41156 28996 41756 29296
rect 21101 28700 37886 28914
rect 25026 26938 25086 26998
rect 26108 26938 26168 26998
rect 27066 26938 27126 26998
rect 25552 26692 25612 26752
rect 27588 26692 27648 26752
rect 23370 25760 23430 25820
rect 24534 25760 24594 25820
rect 23240 25556 23300 25616
rect 21232 23372 21292 23432
rect 24534 25556 24594 25616
rect 30130 26938 30190 26998
rect 31148 26938 31208 26998
rect 29626 26694 29686 26754
rect 26570 25656 26630 25716
rect 25020 24406 25080 24466
rect 32172 26938 32232 26998
rect 33184 26938 33244 26998
rect 31656 26694 31716 26754
rect 28606 25656 28666 25716
rect 33698 26696 33758 26756
rect 30644 25760 30704 25820
rect 30640 25556 30700 25616
rect 27076 24622 27136 24682
rect 27586 24622 27646 24682
rect 26568 24520 26632 24584
rect 26058 24406 26118 24466
rect 27070 24406 27130 24466
rect 23370 23086 23430 23146
rect 23726 20678 23786 20738
rect 23600 20068 23660 20128
rect 20716 19114 20776 19174
rect 20824 19002 20884 19062
rect 19054 18080 19114 18140
rect 21738 19114 21798 19174
rect 21608 19002 21668 19062
rect 20214 17970 20274 18030
rect 22248 18080 22308 18140
rect 18928 16992 18988 17052
rect 20730 17046 20790 17106
rect 20836 16946 20896 17006
rect 23400 17970 23460 18030
rect 21740 17046 21800 17106
rect 23592 17842 23652 17902
rect 21622 16946 21682 17006
rect 18442 15936 18502 15996
rect 18582 15760 18642 15820
rect 19482 15586 19542 15646
rect 23842 20068 23902 20128
rect 24528 23232 24592 23296
rect 24352 23086 24412 23146
rect 28444 24520 28508 24584
rect 34708 26696 34768 26756
rect 36242 26938 36302 26998
rect 37254 26938 37314 26998
rect 35730 26696 35790 26756
rect 32678 25760 32738 25820
rect 32676 25556 32736 25616
rect 33178 25556 33238 25616
rect 29620 24622 29680 24682
rect 28080 24414 28140 24474
rect 29104 24414 29164 24474
rect 25550 23484 25610 23544
rect 26566 23370 26630 23434
rect 30132 24414 30192 24474
rect 38272 26938 38332 26998
rect 37766 26696 37826 26756
rect 34712 25656 34772 25716
rect 34198 25556 34258 25616
rect 31658 24620 31718 24680
rect 27586 23484 27646 23544
rect 28108 23484 28168 23544
rect 28606 23484 28666 23544
rect 35224 25556 35284 25616
rect 36746 25656 36806 25716
rect 35730 25552 35790 25612
rect 36244 25552 36304 25612
rect 36748 25552 36808 25612
rect 37254 25552 37314 25612
rect 37774 25552 37834 25612
rect 32678 24522 32738 24582
rect 38786 25760 38846 25820
rect 40036 25760 40096 25820
rect 33694 24620 33754 24680
rect 34194 24620 34254 24680
rect 34708 24620 34768 24680
rect 35232 24620 35292 24680
rect 35730 24620 35790 24680
rect 36232 24620 36292 24680
rect 29080 23480 29140 23540
rect 24468 22980 24528 23040
rect 25030 22980 25090 23040
rect 26072 22980 26132 23040
rect 27072 22980 27132 23040
rect 29620 23542 29680 23544
rect 29588 23484 29680 23542
rect 30080 23484 30140 23544
rect 29588 23482 29648 23484
rect 30638 23228 30702 23292
rect 31124 23486 31184 23546
rect 30234 22980 30294 23040
rect 31656 23484 31716 23544
rect 36746 24618 36806 24678
rect 37254 24618 37314 24678
rect 37764 24618 37824 24678
rect 36236 24406 36296 24466
rect 37248 24406 37308 24466
rect 33168 23486 33228 23546
rect 32674 23086 32738 23150
rect 31244 22980 31304 23040
rect 32186 22980 32246 23040
rect 33694 23540 33754 23542
rect 33662 23482 33754 23540
rect 33662 23480 33722 23482
rect 34190 23476 34250 23536
rect 34678 23538 34738 23540
rect 34678 23480 34772 23538
rect 34712 23478 34772 23480
rect 38786 24522 38846 24582
rect 38250 24406 38310 24466
rect 35190 23476 35250 23536
rect 35730 23480 35790 23540
rect 37764 23480 37824 23540
rect 36746 23370 36810 23434
rect 40032 23232 40096 23296
rect 38780 23086 38840 23146
rect 24582 22778 24642 22838
rect 27760 22778 27820 22838
rect 25726 21842 25786 21902
rect 26230 21734 26290 21794
rect 27760 21842 27820 21902
rect 27252 21734 27312 21794
rect 28270 21734 28330 21794
rect 25722 20810 25782 20870
rect 26228 20676 26288 20736
rect 31828 22778 31888 22838
rect 29802 21842 29862 21902
rect 29294 21734 29354 21794
rect 30308 21734 30368 21794
rect 27242 20672 27302 20732
rect 28274 20680 28334 20740
rect 31828 21842 31888 21902
rect 31326 21734 31386 21794
rect 32336 21734 32396 21794
rect 29802 20810 29862 20870
rect 29272 20680 29332 20740
rect 30316 20680 30376 20740
rect 35904 22778 35964 22838
rect 33870 21842 33930 21902
rect 33358 21734 33418 21794
rect 34372 21734 34432 21794
rect 31320 20676 31380 20736
rect 32336 20676 32396 20736
rect 31120 20468 31180 20528
rect 24352 20150 24412 20210
rect 25518 20150 25578 20210
rect 24084 19104 24144 19164
rect 23842 17946 23902 18006
rect 23838 17732 23898 17792
rect 23726 16690 23786 16750
rect 18322 15436 18382 15496
rect 24220 19006 24280 19066
rect 24084 15432 24144 15492
rect 27554 20150 27614 20210
rect 28062 20146 28126 20210
rect 26536 19202 26596 19262
rect 39100 22778 39160 22838
rect 35906 21842 35966 21902
rect 35404 21734 35464 21794
rect 36414 21734 36474 21794
rect 33870 20810 33930 20870
rect 33340 20676 33400 20736
rect 34372 20680 34432 20740
rect 32856 20468 32916 20528
rect 32136 20268 32200 20332
rect 37942 21842 38002 21902
rect 37436 21734 37496 21794
rect 35388 20676 35448 20736
rect 36416 20676 36476 20736
rect 37938 20810 37998 20870
rect 37436 20676 37496 20736
rect 39894 20678 39954 20738
rect 38754 20452 38814 20512
rect 36200 20268 36264 20332
rect 37224 20268 37288 20332
rect 38236 20268 38300 20332
rect 32138 20146 32202 20210
rect 28572 19202 28632 19262
rect 28914 19204 28974 19264
rect 26536 19006 26596 19066
rect 27556 19008 27616 19068
rect 25522 18896 25582 18956
rect 27556 18896 27616 18956
rect 24504 17732 24564 17792
rect 31628 19204 31688 19264
rect 35700 20150 35760 20210
rect 37734 20150 37794 20210
rect 32646 19008 32706 19068
rect 30612 18894 30672 18954
rect 32646 18894 32706 18954
rect 26538 17842 26598 17902
rect 26538 17638 26598 17698
rect 28574 17842 28634 17902
rect 28572 17740 28632 17800
rect 28572 17638 28632 17698
rect 25520 16690 25580 16750
rect 24352 16482 24412 16542
rect 26534 16380 26594 16440
rect 30608 17946 30668 18006
rect 27556 16690 27616 16750
rect 27556 16582 27616 16642
rect 31628 17946 31688 18006
rect 31628 17640 31688 17700
rect 35702 18894 35762 18954
rect 32646 17640 32706 17700
rect 36716 19202 36776 19262
rect 37736 18894 37796 18954
rect 38752 19202 38812 19262
rect 33664 17946 33724 18006
rect 33662 17640 33722 17700
rect 28574 16698 28634 16758
rect 30376 16698 30436 16758
rect 28568 16380 28628 16440
rect 28772 16368 28832 16428
rect 25516 15432 25576 15492
rect 30610 16692 30670 16752
rect 35698 17842 35758 17902
rect 36566 17960 36626 18020
rect 36714 17850 36774 17910
rect 36566 17640 36626 17700
rect 36718 17642 36778 17702
rect 32646 16692 32706 16752
rect 32644 16582 32704 16642
rect 27552 15432 27612 15492
rect 24220 15302 24280 15362
rect 19376 15174 19436 15234
rect 19256 15056 19316 15116
rect 32134 16368 32194 16428
rect 37734 17740 37794 17800
rect 40330 20810 40390 20870
rect 40036 20450 40096 20510
rect 40178 20150 40238 20210
rect 40018 19008 40078 19068
rect 38754 17850 38814 17910
rect 39894 17850 39954 17910
rect 38752 17642 38812 17702
rect 33150 16368 33210 16428
rect 35700 16694 35760 16754
rect 36210 16368 36270 16428
rect 36722 16380 36782 16440
rect 37736 16694 37796 16754
rect 40018 17642 40078 17702
rect 39894 16582 39954 16642
rect 38756 16380 38816 16440
rect 35704 15432 35764 15492
rect 37740 15432 37800 15492
rect 28574 15162 28634 15222
rect 40330 18894 40390 18954
rect 40178 15162 40238 15222
rect 18810 14938 18870 14998
rect 3410 14410 14174 14702
rect 18928 13662 18988 13722
rect 19256 13672 19316 13732
rect 18322 13526 18382 13586
rect 18442 13528 18502 13588
rect 18582 13546 18642 13606
rect 18810 13562 18870 13622
rect 18190 13398 18250 13458
rect 15478 12800 15538 12860
rect 4704 1198 4718 12790
rect 4718 1198 4818 12790
rect 4818 1198 4962 12790
rect 17004 12666 17064 12726
rect 18190 6198 18250 6258
rect 13642 5272 13702 5332
rect 7532 5126 7592 5186
rect 11612 5126 11672 5186
rect 6378 4998 6438 5058
rect 9056 4998 9116 5058
rect 10088 4998 10148 5058
rect 8036 4036 8096 4096
rect 7536 3932 7596 3992
rect 9060 4036 9120 4096
rect 8554 3828 8614 3888
rect 6378 2766 6438 2826
rect -156 942 4718 986
rect -156 896 -102 942
rect -102 896 4302 942
rect 4302 896 4718 942
rect 4718 896 4818 986
rect 4818 896 4924 986
rect -2 688 58 748
rect 142 564 202 624
rect 790 688 850 748
rect 1818 564 1878 624
rect 2338 564 2398 624
rect 3366 688 3426 748
rect 662 -170 722 -110
rect 920 -168 980 -108
rect 532 -418 592 -358
rect 790 -300 850 -240
rect 1692 -170 1752 -110
rect 1952 -170 2012 -110
rect 1564 -300 1624 -240
rect 1050 -418 1110 -358
rect 142 -1152 202 -1092
rect 1822 -418 1882 -358
rect 2208 -170 2268 -110
rect 2466 -170 2526 -110
rect 2080 -300 2140 -240
rect 2336 -418 2396 -358
rect -2 -1278 58 -1218
rect 532 -1152 592 -1092
rect 1048 -1152 1108 -1092
rect 2598 -300 2658 -240
rect 4134 688 4194 748
rect 3998 564 4058 624
rect 3242 -170 3302 -110
rect 3502 -170 3562 -110
rect 3112 -418 3172 -358
rect 3368 -300 3428 -240
rect 3626 -418 3686 -358
rect 3112 -1152 3172 -1092
rect 3626 -1152 3686 -1092
rect 3998 -1152 4058 -1092
rect 1560 -1278 1620 -1218
rect 2082 -1278 2142 -1218
rect 2596 -1278 2656 -1218
rect 4134 -1278 4194 -1218
rect 258 -1506 3950 -1402
rect -96 -1936 504 -1636
rect 3696 -1936 4296 -1636
rect 13148 4998 13208 5058
rect 10092 4036 10152 4096
rect 9572 3932 9632 3992
rect 15672 5126 15732 5186
rect 17856 5126 17916 5186
rect 14144 4998 14204 5058
rect 11092 4036 11152 4096
rect 12112 4036 12172 4096
rect 11608 3932 11668 3992
rect 10590 3828 10650 3888
rect 8028 2766 8088 2826
rect 9566 2886 9626 2946
rect 13132 4036 13192 4096
rect 12622 3828 12682 3888
rect 11098 2766 11158 2826
rect 14142 4036 14202 4096
rect 13642 3932 13702 3992
rect 15156 4036 15216 4096
rect 16174 4036 16234 4096
rect 15678 3932 15738 3992
rect 14656 3828 14716 3888
rect 12106 2766 12166 2826
rect 8554 1822 8614 1882
rect 7540 1714 7600 1774
rect 8034 1602 8094 1662
rect 9576 1714 9636 1774
rect 9058 1602 9118 1662
rect 13642 2886 13702 2946
rect 10590 1822 10650 1882
rect 10090 1602 10150 1662
rect 16700 3828 16760 3888
rect 15168 2766 15228 2826
rect 17976 4036 18036 4096
rect 17856 2886 17916 2946
rect 16194 2766 16254 2826
rect 12622 1822 12682 1882
rect 11612 1714 11672 1774
rect 11090 1602 11150 1662
rect 12110 1602 12170 1662
rect 13646 1714 13706 1774
rect 13130 1602 13190 1662
rect 6378 640 6438 700
rect 9048 640 9108 700
rect 10080 640 10140 700
rect 14140 1602 14200 1662
rect 14656 1822 14716 1882
rect 16700 1822 16760 1882
rect 15682 1714 15742 1774
rect 15154 1602 15214 1662
rect 16172 1602 16232 1662
rect 13140 640 13200 700
rect 14136 640 14196 700
rect 17976 1602 18036 1662
rect 7534 510 7594 570
rect 11614 510 11674 570
rect 15674 510 15734 570
rect 17856 510 17916 570
rect 9012 -856 9072 -796
rect 11050 -856 11110 -796
rect 13086 -856 13146 -796
rect 10030 -968 10090 -908
rect 15122 -856 15182 -796
rect 14104 -968 14164 -908
rect 18322 5126 18382 5186
rect 18442 4998 18502 5058
rect 18700 13408 18760 13468
rect 18810 12666 18870 12726
rect 19376 13664 19436 13724
rect 19256 12800 19316 12860
rect 19052 11442 19112 11502
rect 18926 9740 18986 9800
rect 18700 7280 18760 7340
rect 18582 4036 18642 4096
rect 19264 11106 19324 11166
rect 19160 9846 19220 9906
rect 19052 8746 19112 8806
rect 19482 13528 19542 13588
rect 30294 13178 30354 13238
rect 35398 13178 35458 13238
rect 39458 13172 39518 13232
rect 20626 11442 20686 11502
rect 21640 11226 21700 11286
rect 23680 11226 23740 11286
rect 25720 11226 25780 11286
rect 27750 11226 27810 11286
rect 29790 11226 29850 11286
rect 31822 11226 31882 11286
rect 33862 11226 33922 11286
rect 35898 11226 35958 11286
rect 37932 11226 37992 11286
rect 19608 11106 19668 11166
rect 21132 11100 21192 11160
rect 19482 10984 19542 11044
rect 22146 11100 22206 11160
rect 23168 11100 23228 11160
rect 24182 11100 24242 11160
rect 25208 11100 25268 11160
rect 24696 10984 24756 11044
rect 26220 11100 26280 11160
rect 27256 11100 27316 11160
rect 28262 11100 28322 11160
rect 29276 11100 29336 11160
rect 21644 10062 21704 10122
rect 21136 9952 21196 10012
rect 20626 9846 20686 9906
rect 19612 9740 19672 9800
rect 20110 9740 20170 9800
rect 20622 9740 20682 9800
rect 22158 9952 22218 10012
rect 23684 10062 23744 10122
rect 23172 9952 23232 10012
rect 22666 9846 22726 9906
rect 25716 10062 25776 10122
rect 24186 9952 24246 10012
rect 25204 9952 25264 10012
rect 24696 9846 24756 9906
rect 19482 8850 19542 8910
rect 19606 8746 19666 8806
rect 21126 8746 21186 8806
rect 21638 8746 21698 8806
rect 19376 8624 19436 8684
rect 19264 8510 19324 8570
rect 20112 8510 20172 8570
rect 21644 8512 21704 8572
rect 26230 9952 26290 10012
rect 30292 11100 30352 11160
rect 31300 11100 31360 11160
rect 32316 11100 32376 11160
rect 33340 11100 33400 11160
rect 34362 11100 34422 11160
rect 35384 11100 35444 11160
rect 34884 10984 34944 11044
rect 27748 10062 27808 10122
rect 26736 9846 26796 9906
rect 27250 9952 27310 10012
rect 26902 9740 26962 9800
rect 22660 8850 22720 8910
rect 22662 8746 22722 8806
rect 28270 9952 28330 10012
rect 29784 10062 29844 10122
rect 29272 9952 29332 10012
rect 28770 9846 28830 9906
rect 28770 9740 28830 9800
rect 30298 9952 30358 10012
rect 36402 11100 36462 11160
rect 37416 11100 37476 11160
rect 38440 11100 38500 11160
rect 38956 10984 39016 11044
rect 40088 10984 40148 11044
rect 31820 10062 31880 10122
rect 31316 9952 31376 10012
rect 30806 9846 30866 9906
rect 30808 9740 30868 9800
rect 32324 9952 32384 10012
rect 33858 10062 33918 10122
rect 33336 9952 33396 10012
rect 32842 9846 32902 9906
rect 32688 9740 32748 9800
rect 23674 8746 23734 8806
rect 23680 8512 23740 8572
rect 24694 8746 24754 8806
rect 19488 7582 19548 7642
rect 20626 7582 20686 7642
rect 19376 7382 19436 7442
rect 19270 7280 19330 7340
rect 19160 3828 19220 3888
rect 19376 6146 19436 6206
rect 18928 3678 18988 3738
rect 19270 3790 19330 3850
rect 20624 7382 20684 7442
rect 21642 7502 21702 7562
rect 25716 8850 25776 8910
rect 35896 10062 35956 10122
rect 34368 9952 34428 10012
rect 35382 9952 35442 10012
rect 34882 9846 34942 9906
rect 31822 8850 31882 8910
rect 27752 8746 27812 8806
rect 29790 8746 29850 8806
rect 26736 8624 26796 8684
rect 28770 8624 28830 8684
rect 30800 8624 30860 8684
rect 22660 7606 22720 7666
rect 22156 7388 22216 7448
rect 23682 7502 23742 7562
rect 23160 7388 23220 7448
rect 20624 6350 20684 6410
rect 21130 6248 21190 6308
rect 24696 7606 24756 7666
rect 24172 7388 24232 7448
rect 25714 7502 25774 7562
rect 25192 7388 25252 7448
rect 25714 7390 25774 7450
rect 27748 7502 27808 7562
rect 26732 7280 26792 7340
rect 22662 6350 22722 6410
rect 22660 6146 22720 6206
rect 27750 7390 27810 7450
rect 28766 7280 28826 7340
rect 32840 8746 32900 8806
rect 36400 9952 36460 10012
rect 37932 10062 37992 10122
rect 37424 9952 37484 10012
rect 36912 9846 36972 9906
rect 36912 9742 36972 9802
rect 33858 8746 33918 8806
rect 34878 8746 34938 8806
rect 29788 7502 29848 7562
rect 29786 7390 29846 7450
rect 31822 7502 31882 7562
rect 32018 7498 32078 7558
rect 30806 7280 30866 7340
rect 31822 7390 31882 7450
rect 38444 9952 38504 10012
rect 38952 9846 39012 9906
rect 40088 9742 40148 9802
rect 36916 8850 36976 8910
rect 35894 8746 35954 8806
rect 37930 8746 37990 8806
rect 32840 7606 32900 7666
rect 32018 7280 32078 7340
rect 32312 7282 32372 7342
rect 24698 6350 24758 6410
rect 21644 6046 21704 6106
rect 23168 6140 23228 6200
rect 24190 6140 24250 6200
rect 23678 6046 23738 6106
rect 26730 6350 26790 6410
rect 26222 6248 26282 6308
rect 25204 6140 25264 6200
rect 26222 6140 26282 6200
rect 25714 6046 25774 6106
rect 21126 5122 21186 5182
rect 22036 5122 22096 5182
rect 21126 4906 21186 4966
rect 19490 4802 19550 4862
rect 23038 5122 23098 5182
rect 22164 4906 22224 4966
rect 24190 5122 24250 5182
rect 23678 5020 23738 5080
rect 23178 4906 23238 4966
rect 21124 3894 21184 3954
rect 20626 3790 20686 3850
rect 20622 3580 20682 3640
rect 22132 3894 22192 3954
rect 21642 3678 21702 3738
rect 27242 6140 27302 6200
rect 33856 7390 33916 7450
rect 33340 7282 33400 7342
rect 33858 7276 33918 7336
rect 34876 7606 34936 7666
rect 35894 7390 35954 7450
rect 36910 7498 36970 7558
rect 37414 7494 37474 7554
rect 40074 8512 40134 8572
rect 37934 7390 37994 7450
rect 35894 7276 35954 7336
rect 31312 6362 31372 6422
rect 30806 6234 30866 6294
rect 32842 6036 32902 6096
rect 25200 5122 25260 5182
rect 26206 5122 26266 5182
rect 27250 5122 27310 5182
rect 27750 5128 27810 5188
rect 26204 4906 26264 4966
rect 27244 4906 27304 4966
rect 26728 4802 26788 4862
rect 23146 3894 23206 3954
rect 24184 3894 24244 3954
rect 23680 3678 23740 3738
rect 22660 3580 22720 3640
rect 28258 4906 28318 4966
rect 29786 5128 29846 5188
rect 29266 4906 29326 4966
rect 30310 4906 30370 4966
rect 28770 4802 28830 4862
rect 37932 7276 37992 7336
rect 34354 6140 34414 6200
rect 31822 5128 31882 5188
rect 31300 4906 31360 4966
rect 32318 4906 32378 4966
rect 30808 4802 30868 4862
rect 38950 7606 39010 7666
rect 39968 7624 40028 7684
rect 40202 8494 40262 8554
rect 40568 7494 40628 7554
rect 40318 7390 40378 7450
rect 36406 6362 36466 6422
rect 36544 6366 36604 6426
rect 40074 7276 40134 7336
rect 37426 6366 37486 6426
rect 38432 6366 38492 6426
rect 35384 6140 35444 6200
rect 36544 6140 36604 6200
rect 36912 6140 36972 6200
rect 36912 6036 36972 6096
rect 38950 6362 39010 6422
rect 38950 6234 39010 6294
rect 37928 6038 37988 6098
rect 33860 5128 33920 5188
rect 33852 5020 33912 5080
rect 33352 4906 33412 4966
rect 32842 4802 32902 4862
rect 33354 4798 33414 4858
rect 34376 4798 34436 4858
rect 34876 4804 34936 4864
rect 25202 3894 25262 3954
rect 25718 3900 25778 3960
rect 27754 3900 27814 3960
rect 29786 3900 29846 3960
rect 31820 3900 31880 3960
rect 24700 3580 24760 3640
rect 19488 2558 19548 2618
rect 20628 2342 20688 2402
rect 21642 2656 21702 2716
rect 21646 2462 21706 2522
rect 22660 2558 22720 2618
rect 28770 3790 28830 3850
rect 30806 3790 30866 3850
rect 27752 3678 27812 3738
rect 26736 3580 26796 3640
rect 23678 2656 23738 2716
rect 24184 2558 24244 2618
rect 23682 2462 23742 2522
rect 25716 2656 25776 2716
rect 25206 2558 25266 2618
rect 24696 2342 24756 2402
rect 19376 1426 19436 1486
rect 19270 1300 19330 1360
rect 26228 2558 26288 2618
rect 25710 2462 25770 2522
rect 35896 5128 35956 5188
rect 35892 5020 35952 5080
rect 36384 4906 36444 4966
rect 37934 5128 37994 5188
rect 37930 5020 37990 5080
rect 37422 4906 37482 4966
rect 36910 4804 36970 4864
rect 32842 3902 32902 3962
rect 33196 3902 33256 3962
rect 32838 3790 32898 3850
rect 32348 3692 32408 3752
rect 27578 2676 27638 2736
rect 27748 2676 27808 2736
rect 27232 2558 27292 2618
rect 26730 2342 26790 2402
rect 22660 1300 22720 1360
rect 23180 1312 23240 1372
rect 21642 1198 21702 1258
rect 23678 1198 23738 1258
rect 22660 1094 22720 1154
rect 19488 196 19548 256
rect 19160 92 19220 152
rect 20624 92 20684 152
rect 21132 -14 21192 46
rect 18110 -968 18170 -908
rect 27578 2462 27638 2522
rect 27754 2468 27814 2528
rect 33386 3692 33446 3752
rect 34362 3692 34422 3752
rect 33196 3584 33256 3644
rect 38448 4906 38508 4966
rect 38952 4804 39012 4864
rect 36914 3902 36974 3962
rect 35378 3692 35438 3752
rect 37404 3692 37464 3752
rect 34876 3580 34936 3640
rect 36912 3580 36972 3640
rect 29790 2676 29850 2736
rect 31822 2676 31882 2736
rect 33862 2676 33922 2736
rect 32840 2578 32900 2638
rect 29782 2468 29842 2528
rect 24698 1198 24758 1258
rect 25714 1198 25774 1258
rect 22658 196 22718 256
rect 22664 92 22724 152
rect 22152 -14 22212 46
rect 21644 -124 21704 -64
rect 23176 -14 23236 46
rect 26734 1198 26794 1258
rect 31826 2468 31886 2528
rect 33854 2468 33914 2528
rect 34880 2342 34940 2402
rect 38434 3692 38494 3752
rect 38948 3580 39008 3640
rect 35892 2468 35952 2528
rect 38946 2578 39006 2638
rect 37932 2468 37992 2528
rect 38450 2472 38510 2532
rect 39962 2472 40022 2532
rect 36910 2342 36970 2402
rect 37436 2344 37496 2404
rect 28764 1426 28824 1486
rect 30806 1426 30866 1486
rect 32842 1426 32902 1486
rect 28260 1312 28320 1372
rect 33348 1316 33408 1376
rect 27752 1198 27812 1258
rect 29782 1198 29842 1258
rect 31820 1198 31880 1258
rect 33856 1198 33916 1258
rect 27596 1094 27656 1154
rect 24694 92 24754 152
rect 24194 -14 24254 46
rect 25208 -14 25268 46
rect 23680 -124 23740 -64
rect 19488 -1046 19548 -986
rect 20624 -1046 20684 -986
rect 21136 -1154 21196 -1094
rect 26888 198 26948 258
rect 26734 92 26794 152
rect 26240 -14 26300 46
rect 25718 -124 25778 -64
rect 22150 -1154 22210 -1094
rect 23172 -1154 23232 -1094
rect 27252 -14 27312 46
rect 28766 198 28826 258
rect 28770 92 28830 152
rect 28260 -14 28320 46
rect 27756 -124 27816 -64
rect 24694 -1046 24754 -986
rect 24186 -1154 24246 -1094
rect 25212 -1154 25272 -1094
rect 29278 -14 29338 46
rect 30804 198 30864 258
rect 30806 92 30866 152
rect 30304 -14 30364 46
rect 29792 -124 29852 -64
rect 26224 -1154 26284 -1094
rect 27260 -1154 27320 -1094
rect 31306 -14 31366 46
rect 34002 1094 34062 1154
rect 38950 2344 39010 2404
rect 34878 1198 34938 1258
rect 35896 1426 35956 1486
rect 35898 1198 35958 1258
rect 32674 198 32734 258
rect 32326 -14 32386 46
rect 32840 92 32900 152
rect 31828 -124 31888 -64
rect 28266 -1154 28326 -1094
rect 29280 -1154 29340 -1094
rect 33346 -14 33406 46
rect 36912 1198 36972 1258
rect 36912 1094 36972 1154
rect 37928 1426 37988 1486
rect 40202 6362 40262 6422
rect 40440 6140 40500 6200
rect 40318 6038 40378 6098
rect 40202 4804 40262 4864
rect 40198 3902 40258 3962
rect 40318 2676 40378 2736
rect 40198 2578 40258 2638
rect 40074 1426 40134 1486
rect 38448 1316 38508 1376
rect 39456 1316 39516 1376
rect 40566 4906 40626 4966
rect 40568 2472 40628 2532
rect 40440 2344 40500 2404
rect 40802 8494 40862 8554
rect 40690 1316 40750 1376
rect 37934 1198 37994 1258
rect 34880 92 34940 152
rect 34372 -14 34432 46
rect 35390 -14 35450 46
rect 33860 -124 33920 -64
rect 30296 -1154 30356 -1094
rect 31304 -1154 31364 -1094
rect 36910 92 36970 152
rect 36404 -14 36464 46
rect 35892 -124 35952 -64
rect 32320 -1154 32380 -1094
rect 33344 -1154 33404 -1094
rect 37418 -14 37478 46
rect 40094 1094 40154 1154
rect 38950 198 39010 258
rect 38950 92 39010 152
rect 38440 -14 38500 46
rect 37932 -124 37992 -64
rect 34874 -1046 34934 -986
rect 34366 -1154 34426 -1094
rect 35388 -1154 35448 -1094
rect 36406 -1154 36466 -1094
rect 37420 -1154 37480 -1094
rect 40802 92 40862 152
rect 40094 -1046 40154 -986
rect 38444 -1154 38504 -1094
rect 8968 -1550 40968 -1396
rect 4824 -2036 5424 -1736
rect 41256 -2036 41856 -1736
<< metal2 >>
rect 17524 29296 18124 29306
rect 17524 28986 18124 28996
rect 41156 29296 41756 29306
rect 41156 28986 41756 28996
rect 21038 28914 37918 28946
rect 21038 28700 21101 28914
rect 37886 28700 37918 28914
rect 21038 28680 37918 28700
rect 21038 28678 25392 28680
rect 25026 26998 25086 27004
rect 26108 26998 26168 27004
rect 27066 26998 27126 27004
rect 30130 26998 30190 27004
rect 31148 26998 31208 27004
rect 32172 26998 32232 27004
rect 33184 26998 33244 27004
rect 36242 26998 36302 27004
rect 37254 26998 37314 27004
rect 38272 26998 38332 27004
rect 25086 26938 26108 26998
rect 26168 26938 27066 26998
rect 27126 26938 30130 26998
rect 30190 26938 31148 26998
rect 31208 26938 32172 26998
rect 32232 26938 33184 26998
rect 33244 26938 36242 26998
rect 36302 26938 37254 26998
rect 37314 26938 38272 26998
rect 25026 26932 25086 26938
rect 26108 26932 26168 26938
rect 27066 26932 27126 26938
rect 30130 26932 30190 26938
rect 31148 26932 31208 26938
rect 32172 26932 32232 26938
rect 33184 26932 33244 26938
rect 36242 26932 36302 26938
rect 37254 26932 37314 26938
rect 38272 26932 38332 26938
rect 25552 26752 25612 26758
rect 27588 26752 27648 26758
rect 29626 26754 29686 26760
rect 31656 26754 31716 26760
rect 33698 26756 33758 26762
rect 34708 26756 34768 26762
rect 35730 26756 35790 26762
rect 37766 26756 37826 26762
rect 25612 26692 27588 26752
rect 27648 26694 29626 26752
rect 29686 26694 31656 26754
rect 31716 26696 33698 26754
rect 33758 26696 34708 26756
rect 34768 26696 35730 26756
rect 35790 26696 37766 26756
rect 31716 26694 33896 26696
rect 27648 26692 29808 26694
rect 25552 26686 25612 26692
rect 27588 26686 27648 26692
rect 29626 26688 29686 26692
rect 31656 26688 31716 26694
rect 33698 26690 33758 26694
rect 34708 26690 34768 26696
rect 35730 26690 35790 26696
rect 37766 26690 37826 26696
rect 23370 25820 23430 25826
rect 24534 25820 24594 25826
rect 30644 25820 30704 25826
rect 23430 25760 24534 25820
rect 24594 25760 30644 25820
rect 23370 25754 23430 25760
rect 24534 25754 24594 25760
rect 30644 25754 30704 25760
rect 32678 25820 32738 25826
rect 38786 25820 38846 25826
rect 40036 25820 40096 25826
rect 32738 25760 38786 25820
rect 38846 25760 40036 25820
rect 32678 25754 32738 25760
rect 38786 25754 38846 25760
rect 40036 25754 40096 25760
rect 26570 25716 26630 25722
rect 28606 25716 28666 25722
rect 34712 25716 34772 25722
rect 36746 25716 36806 25722
rect 26630 25656 28606 25716
rect 28666 25708 29084 25716
rect 29300 25708 34712 25716
rect 28666 25662 34712 25708
rect 28666 25658 31100 25662
rect 28666 25656 30074 25658
rect 30312 25656 31100 25658
rect 31316 25656 34712 25662
rect 34772 25656 36746 25716
rect 26570 25650 26630 25656
rect 28606 25650 28666 25656
rect 34712 25650 34772 25656
rect 36746 25650 36806 25656
rect 23240 25616 23300 25622
rect 24534 25616 24594 25622
rect 30640 25616 30700 25622
rect 32676 25616 32736 25622
rect 23300 25556 24534 25616
rect 24594 25556 30640 25616
rect 30700 25556 32676 25616
rect 23240 25550 23300 25556
rect 24534 25550 24594 25556
rect 30640 25550 30700 25556
rect 32676 25550 32736 25556
rect 33178 25616 33238 25622
rect 34198 25616 34258 25622
rect 35224 25616 35284 25622
rect 33238 25556 34198 25616
rect 34258 25556 35224 25616
rect 33178 25550 33238 25556
rect 34198 25550 34258 25556
rect 35224 25550 35284 25556
rect 35730 25612 35790 25618
rect 36244 25612 36304 25618
rect 36748 25612 36808 25618
rect 37254 25612 37314 25618
rect 35790 25552 36244 25612
rect 36304 25552 36748 25612
rect 36808 25552 37254 25612
rect 37314 25552 37774 25612
rect 37834 25552 37840 25612
rect 35730 25546 35790 25552
rect 36244 25546 36304 25552
rect 36748 25546 36808 25552
rect 37254 25546 37314 25552
rect 27586 24682 27646 24688
rect 29620 24682 29680 24688
rect 31658 24682 31718 24686
rect 27070 24622 27076 24682
rect 27136 24622 27586 24682
rect 27646 24622 29620 24682
rect 29680 24680 31862 24682
rect 33694 24680 33754 24686
rect 34194 24680 34254 24686
rect 34708 24680 34768 24686
rect 35232 24680 35292 24686
rect 35730 24680 35790 24686
rect 36232 24680 36292 24686
rect 29680 24622 31658 24680
rect 27586 24616 27646 24622
rect 29620 24616 29680 24622
rect 31718 24620 33694 24680
rect 33754 24620 34194 24680
rect 34254 24620 34708 24680
rect 34768 24620 35232 24680
rect 35292 24620 35730 24680
rect 35790 24620 36232 24680
rect 36292 24678 36600 24680
rect 36746 24678 36806 24684
rect 37254 24678 37314 24684
rect 37764 24678 37824 24684
rect 36292 24620 36746 24678
rect 31658 24614 31718 24620
rect 33694 24614 33754 24620
rect 34194 24614 34254 24620
rect 34708 24614 34768 24620
rect 35232 24614 35292 24620
rect 35629 24618 36144 24620
rect 35730 24614 35790 24618
rect 36232 24614 36292 24620
rect 36394 24618 36746 24620
rect 36806 24618 37254 24678
rect 37314 24618 37764 24678
rect 36746 24612 36806 24618
rect 37254 24612 37314 24618
rect 37764 24612 37824 24618
rect 26568 24584 26632 24590
rect 28444 24584 28508 24590
rect 26632 24520 28444 24584
rect 26568 24514 26632 24520
rect 28444 24514 28508 24520
rect 32678 24582 32738 24588
rect 38786 24582 38846 24588
rect 32738 24522 38786 24582
rect 32678 24516 32738 24522
rect 38786 24516 38846 24522
rect 28080 24474 28140 24480
rect 29104 24474 29164 24480
rect 30132 24474 30192 24480
rect 26058 24466 26118 24472
rect 27070 24466 27130 24472
rect 25014 24406 25020 24466
rect 25080 24406 26058 24466
rect 26118 24406 27070 24466
rect 28140 24414 29104 24474
rect 29164 24414 30132 24474
rect 28080 24408 28140 24414
rect 29104 24408 29164 24414
rect 30132 24408 30192 24414
rect 36236 24466 36296 24472
rect 37248 24466 37308 24472
rect 38250 24466 38310 24472
rect 26058 24400 26118 24406
rect 27070 24400 27130 24406
rect 36296 24406 37248 24466
rect 37308 24406 38250 24466
rect 36236 24400 36296 24406
rect 37248 24400 37308 24406
rect 38250 24400 38310 24406
rect 25550 23544 25610 23550
rect 27586 23544 27646 23550
rect 28108 23544 28168 23550
rect 28606 23544 28666 23550
rect 29620 23544 29680 23550
rect 30080 23544 30140 23550
rect 31118 23544 31124 23546
rect 25610 23484 27586 23544
rect 27646 23484 28108 23544
rect 28168 23484 28606 23544
rect 28666 23542 29620 23544
rect 28666 23540 29588 23542
rect 28666 23484 29080 23540
rect 25550 23478 25610 23484
rect 27586 23478 27646 23484
rect 28108 23478 28168 23484
rect 28606 23478 28666 23484
rect 29074 23480 29080 23484
rect 29140 23484 29588 23540
rect 29680 23484 30080 23544
rect 30140 23486 31124 23544
rect 31184 23544 31190 23546
rect 31656 23544 31716 23550
rect 33162 23544 33168 23546
rect 31184 23486 31656 23544
rect 30140 23484 31656 23486
rect 31716 23486 33168 23544
rect 33228 23544 33234 23546
rect 33228 23542 33540 23544
rect 33694 23542 33754 23548
rect 35730 23542 35790 23546
rect 33228 23540 33694 23542
rect 33754 23540 35918 23542
rect 37764 23540 37824 23546
rect 33228 23486 33662 23540
rect 31716 23484 33662 23486
rect 29140 23480 29146 23484
rect 29582 23482 29588 23484
rect 29648 23482 29680 23484
rect 29620 23478 29680 23482
rect 30080 23478 30140 23484
rect 31656 23478 31716 23484
rect 31800 23482 33126 23484
rect 33332 23482 33662 23484
rect 33754 23536 34678 23540
rect 34738 23538 35730 23540
rect 33754 23482 34190 23536
rect 33656 23480 33662 23482
rect 33722 23480 33754 23482
rect 33694 23476 33754 23480
rect 34184 23476 34190 23482
rect 34250 23482 34678 23536
rect 34250 23476 34256 23482
rect 34672 23480 34678 23482
rect 34772 23536 35730 23538
rect 34772 23482 35190 23536
rect 34706 23478 34712 23480
rect 34772 23478 34778 23482
rect 35184 23476 35190 23482
rect 35250 23482 35730 23536
rect 35250 23476 35256 23482
rect 35790 23480 37764 23540
rect 35730 23474 35790 23480
rect 37764 23474 37824 23480
rect 21232 23434 21292 23438
rect 26566 23434 26630 23440
rect 36746 23434 36810 23440
rect 21230 23432 26566 23434
rect 21230 23372 21232 23432
rect 21292 23372 26566 23432
rect 21230 23370 26566 23372
rect 26630 23370 36746 23434
rect 21232 23366 21292 23370
rect 26566 23364 26630 23370
rect 36746 23364 36810 23370
rect 24528 23296 24592 23302
rect 24592 23292 40032 23296
rect 24592 23232 30638 23292
rect 24528 23226 24592 23232
rect 30632 23228 30638 23232
rect 30702 23232 40032 23292
rect 40096 23232 40102 23296
rect 30702 23228 30708 23232
rect 23370 23146 23430 23152
rect 32674 23150 32738 23156
rect 23430 23086 24352 23146
rect 24412 23086 32674 23146
rect 38780 23146 38840 23152
rect 32738 23086 38780 23146
rect 23370 23080 23430 23086
rect 32674 23080 32738 23086
rect 38780 23080 38840 23086
rect 24468 23040 24528 23046
rect 25030 23040 25090 23046
rect 26072 23040 26132 23046
rect 27072 23040 27132 23046
rect 30234 23040 30294 23046
rect 31244 23040 31304 23046
rect 32186 23040 32246 23046
rect 24528 22980 25030 23040
rect 25090 22980 26072 23040
rect 26132 22980 27072 23040
rect 27132 22980 30234 23040
rect 30294 22980 31244 23040
rect 31304 22980 32186 23040
rect 24468 22974 24528 22980
rect 25030 22974 25090 22980
rect 26072 22974 26132 22980
rect 27072 22974 27132 22980
rect 30234 22974 30294 22980
rect 31244 22974 31304 22980
rect 32186 22974 32246 22980
rect 24582 22838 24642 22844
rect 27760 22838 27820 22844
rect 31828 22838 31888 22844
rect 35904 22838 35964 22844
rect 39100 22838 39160 22844
rect 24642 22778 27760 22838
rect 27820 22778 31828 22838
rect 31888 22778 35904 22838
rect 35964 22778 39100 22838
rect 24582 22772 24642 22778
rect 27760 22772 27820 22778
rect 31828 22772 31888 22778
rect 35904 22772 35964 22778
rect 39100 22772 39160 22778
rect 25726 21902 25786 21908
rect 27760 21902 27820 21908
rect 29802 21902 29862 21908
rect 31828 21902 31888 21908
rect 33870 21902 33930 21908
rect 35906 21902 35966 21908
rect 37942 21902 38002 21908
rect 25786 21842 27760 21902
rect 27820 21842 29802 21902
rect 29862 21842 31828 21902
rect 31888 21842 33870 21902
rect 33930 21842 35906 21902
rect 35966 21842 37942 21902
rect 25726 21836 25786 21842
rect 27760 21836 27820 21842
rect 29802 21836 29862 21842
rect 31828 21836 31888 21842
rect 33870 21836 33930 21842
rect 35906 21836 35966 21842
rect 37942 21836 38002 21842
rect 26230 21794 26290 21800
rect 26290 21734 27252 21794
rect 27312 21734 28270 21794
rect 28330 21734 29294 21794
rect 29354 21734 30308 21794
rect 30368 21734 31326 21794
rect 31386 21734 32336 21794
rect 32396 21734 33358 21794
rect 33418 21734 34372 21794
rect 34432 21734 35404 21794
rect 35464 21734 36414 21794
rect 36474 21734 37436 21794
rect 37496 21734 37502 21794
rect 26230 21728 26290 21734
rect 25722 20870 25782 20876
rect 29802 20870 29862 20876
rect 33870 20870 33930 20876
rect 37938 20870 37998 20876
rect 40330 20870 40390 20876
rect 18190 20810 25722 20870
rect 25782 20810 29802 20870
rect 29862 20810 33870 20870
rect 33930 20810 37938 20870
rect 37998 20810 40330 20870
rect 3048 14702 14318 14958
rect 3048 14410 3410 14702
rect 14262 14410 14318 14702
rect 3048 14102 14318 14410
rect 3048 13780 15400 14102
rect 18190 13458 18250 20810
rect 25722 20804 25782 20810
rect 29802 20804 29862 20810
rect 33870 20804 33930 20810
rect 37938 20804 37998 20810
rect 40330 20804 40390 20810
rect 23726 20738 23786 20744
rect 28268 20738 28274 20740
rect 23786 20736 28274 20738
rect 23786 20678 26228 20736
rect 23726 20672 23786 20678
rect 26222 20676 26228 20678
rect 26288 20732 28274 20736
rect 26288 20678 27242 20732
rect 26288 20676 26294 20678
rect 27236 20672 27242 20678
rect 27302 20680 28274 20732
rect 28334 20738 28340 20740
rect 29266 20738 29272 20740
rect 28334 20680 29272 20738
rect 29332 20738 29338 20740
rect 30310 20738 30316 20740
rect 29332 20680 30316 20738
rect 30376 20738 30382 20740
rect 34366 20738 34372 20740
rect 30376 20736 34372 20738
rect 30376 20680 31320 20736
rect 27302 20678 31320 20680
rect 27302 20672 27308 20678
rect 31314 20676 31320 20678
rect 31380 20678 32336 20736
rect 31380 20676 31386 20678
rect 32330 20676 32336 20678
rect 32396 20678 33340 20736
rect 32396 20676 32402 20678
rect 33334 20676 33340 20678
rect 33400 20680 34372 20736
rect 34432 20738 34438 20740
rect 39894 20738 39954 20744
rect 34432 20736 39894 20738
rect 34432 20680 35388 20736
rect 33400 20678 35388 20680
rect 33400 20676 33406 20678
rect 35382 20676 35388 20678
rect 35448 20678 36416 20736
rect 35448 20676 35454 20678
rect 36410 20676 36416 20678
rect 36476 20678 37436 20736
rect 36476 20676 36482 20678
rect 37430 20676 37436 20678
rect 37496 20678 39894 20736
rect 37496 20676 37502 20678
rect 39894 20672 39954 20678
rect 31120 20528 31180 20534
rect 31180 20468 32856 20528
rect 32916 20468 32922 20528
rect 38754 20514 38814 20518
rect 38752 20512 40096 20514
rect 31120 20462 31180 20468
rect 38752 20452 38754 20512
rect 38814 20510 40096 20512
rect 38814 20452 40036 20510
rect 38752 20450 40036 20452
rect 40096 20450 40102 20510
rect 38754 20446 38814 20450
rect 32136 20332 32200 20338
rect 36200 20332 36264 20338
rect 37224 20332 37288 20338
rect 38236 20332 38300 20338
rect 32200 20268 36200 20332
rect 36264 20268 37224 20332
rect 37288 20268 38236 20332
rect 32136 20262 32200 20268
rect 36200 20262 36264 20268
rect 37224 20262 37288 20268
rect 38236 20262 38300 20268
rect 24352 20210 24412 20216
rect 25518 20210 25578 20216
rect 27554 20210 27614 20216
rect 24412 20150 25518 20210
rect 25578 20150 27554 20210
rect 24352 20144 24412 20150
rect 25518 20144 25578 20150
rect 27554 20144 27614 20150
rect 28062 20210 28126 20216
rect 32138 20210 32202 20216
rect 28126 20146 32138 20210
rect 28062 20140 28126 20146
rect 32138 20140 32202 20146
rect 35700 20210 35760 20216
rect 37734 20210 37794 20216
rect 40178 20210 40238 20216
rect 35760 20150 37734 20210
rect 37794 20150 40178 20210
rect 35700 20144 35760 20150
rect 37734 20144 37794 20150
rect 40178 20144 40238 20150
rect 23600 20128 23660 20134
rect 23842 20128 23902 20134
rect 23660 20068 23842 20128
rect 23600 20062 23660 20068
rect 23842 20062 23902 20068
rect 26536 19262 26596 19268
rect 28572 19262 28632 19268
rect 26596 19202 28572 19262
rect 26536 19196 26596 19202
rect 28572 19196 28632 19202
rect 28914 19264 28974 19270
rect 31628 19264 31688 19270
rect 28974 19204 31628 19264
rect 28914 19198 28974 19204
rect 31628 19198 31688 19204
rect 36716 19262 36776 19268
rect 38752 19262 38812 19268
rect 36776 19202 38752 19262
rect 36716 19196 36776 19202
rect 20716 19174 20776 19180
rect 21738 19174 21798 19180
rect 20776 19114 21738 19174
rect 20716 19108 20776 19114
rect 21738 19108 21798 19114
rect 24084 19164 24144 19170
rect 36824 19164 36884 19202
rect 38752 19196 38812 19202
rect 24144 19104 36884 19164
rect 24084 19098 24144 19104
rect 20824 19062 20884 19068
rect 21608 19062 21668 19068
rect 20884 19002 21608 19062
rect 20824 18996 20884 19002
rect 21608 18996 21668 19002
rect 24220 19066 24280 19072
rect 26536 19066 26596 19072
rect 24280 19006 26536 19066
rect 24220 19000 24280 19006
rect 26536 19000 26596 19006
rect 27556 19068 27616 19074
rect 32646 19068 32706 19074
rect 40018 19068 40078 19074
rect 27616 19008 32646 19068
rect 32706 19008 40018 19068
rect 27556 19002 27616 19008
rect 32646 19002 32706 19008
rect 40018 19002 40078 19008
rect 25522 18956 25582 18962
rect 27556 18956 27616 18962
rect 25582 18896 27556 18956
rect 25522 18890 25582 18896
rect 27556 18890 27616 18896
rect 30612 18954 30672 18960
rect 32646 18954 32706 18960
rect 30672 18894 32646 18954
rect 30612 18888 30672 18894
rect 32646 18888 32706 18894
rect 35702 18954 35762 18960
rect 37736 18956 37796 18960
rect 37668 18954 37796 18956
rect 40330 18954 40390 18960
rect 35762 18894 37736 18954
rect 37796 18894 40330 18954
rect 35702 18888 35762 18894
rect 37668 18892 37796 18894
rect 37736 18888 37796 18892
rect 40330 18888 40390 18894
rect 19054 18140 19114 18146
rect 22248 18140 22308 18146
rect 19114 18080 22248 18140
rect 19054 18074 19114 18080
rect 22248 18074 22308 18080
rect 20214 18030 20274 18036
rect 23400 18030 23460 18036
rect 20274 17970 23400 18030
rect 36566 18020 36626 18026
rect 20214 17964 20274 17970
rect 23400 17964 23460 17970
rect 23842 18006 23902 18012
rect 30608 18006 30668 18012
rect 31628 18006 31688 18012
rect 33664 18006 33724 18012
rect 23902 17946 30608 18006
rect 30668 17946 31628 18006
rect 31688 17946 33664 18006
rect 36626 17960 40988 18020
rect 36566 17954 36626 17960
rect 23842 17940 23902 17946
rect 30608 17940 30668 17946
rect 31628 17940 31688 17946
rect 33664 17940 33724 17946
rect 36714 17910 36774 17916
rect 38754 17910 38814 17916
rect 39894 17910 39954 17916
rect 23592 17902 23652 17908
rect 28574 17902 28634 17908
rect 35698 17902 35758 17908
rect 23652 17842 26538 17902
rect 26598 17842 28574 17902
rect 28634 17842 35698 17902
rect 36774 17850 38754 17910
rect 38814 17850 39894 17910
rect 36714 17844 36774 17850
rect 38754 17844 38814 17850
rect 39894 17844 39954 17850
rect 23592 17836 23652 17842
rect 28574 17836 28634 17842
rect 35698 17836 35758 17842
rect 28572 17800 28632 17806
rect 37734 17800 37794 17806
rect 23838 17792 23898 17798
rect 24504 17792 24564 17798
rect 23898 17732 24504 17792
rect 28632 17740 37734 17800
rect 28572 17734 28632 17740
rect 37734 17734 37794 17740
rect 23838 17726 23898 17732
rect 24504 17726 24564 17732
rect 26538 17698 26598 17704
rect 28572 17698 28632 17704
rect 26598 17638 28572 17698
rect 26538 17632 26598 17638
rect 28572 17632 28632 17638
rect 31628 17700 31688 17706
rect 32646 17700 32706 17706
rect 33662 17700 33722 17706
rect 36566 17700 36626 17706
rect 31688 17640 32646 17700
rect 32706 17640 33662 17700
rect 33722 17640 36566 17700
rect 31628 17634 31688 17640
rect 32646 17634 32706 17640
rect 33662 17634 33722 17640
rect 36566 17634 36626 17640
rect 36718 17702 36778 17708
rect 38752 17702 38812 17708
rect 40018 17702 40078 17708
rect 36778 17642 38752 17702
rect 38812 17642 40018 17702
rect 40078 17642 40860 17702
rect 36718 17636 36778 17642
rect 38752 17636 38812 17642
rect 40018 17636 40078 17642
rect 20730 17106 20790 17112
rect 21740 17106 21800 17112
rect 18922 16992 18928 17052
rect 18988 16992 18994 17052
rect 20790 17046 21740 17106
rect 20730 17040 20790 17046
rect 21740 17040 21800 17046
rect 20836 17006 20896 17012
rect 21622 17006 21682 17012
rect 18436 15936 18442 15996
rect 18502 15936 18508 15996
rect 18316 15436 18322 15496
rect 18382 15436 18388 15496
rect 18322 13586 18382 15436
rect 18322 13520 18382 13526
rect 18442 13588 18502 15936
rect 18576 15760 18582 15820
rect 18642 15760 18648 15820
rect 18582 13606 18642 15760
rect 18804 14938 18810 14998
rect 18870 14938 18876 14998
rect 18810 13622 18870 14938
rect 18928 13722 18988 16992
rect 20896 16946 21622 17006
rect 20836 16940 20896 16946
rect 21622 16940 21682 16946
rect 28574 16758 28634 16764
rect 30376 16758 30436 16764
rect 23726 16750 23786 16756
rect 25520 16750 25580 16756
rect 27556 16750 27616 16756
rect 23786 16690 25520 16750
rect 25580 16690 27556 16750
rect 28634 16698 30376 16758
rect 28574 16692 28634 16698
rect 30376 16692 30436 16698
rect 30610 16752 30670 16758
rect 32646 16752 32706 16758
rect 30670 16692 32646 16752
rect 23726 16684 23786 16690
rect 19476 15586 19482 15646
rect 19542 15586 19548 15646
rect 19370 15174 19376 15234
rect 19436 15174 19442 15234
rect 19250 15056 19256 15116
rect 19316 15056 19322 15116
rect 19256 13732 19316 15056
rect 19376 14140 19436 15174
rect 19359 14131 19449 14140
rect 19359 14032 19449 14041
rect 18922 13662 18928 13722
rect 18988 13662 18994 13722
rect 19376 13724 19436 14032
rect 19256 13666 19316 13672
rect 19370 13664 19376 13724
rect 19436 13664 19442 13724
rect 19482 13588 19542 15586
rect 18810 13556 18870 13562
rect 18582 13540 18642 13546
rect 19476 13528 19482 13588
rect 19542 13528 19548 13588
rect 18442 13522 18502 13528
rect 18700 13468 18760 13474
rect 23954 13468 24014 16690
rect 25520 16684 25580 16690
rect 27556 16684 27616 16690
rect 30610 16686 30670 16692
rect 32646 16686 32706 16692
rect 35700 16754 35760 16760
rect 37736 16754 37796 16760
rect 35760 16694 37736 16754
rect 35700 16688 35760 16694
rect 37736 16688 37796 16694
rect 27556 16642 27616 16648
rect 32644 16642 32704 16648
rect 39894 16642 39954 16648
rect 27616 16582 32644 16642
rect 32704 16582 39894 16642
rect 27556 16576 27616 16582
rect 32644 16576 32704 16582
rect 39894 16576 39954 16582
rect 24352 16542 24412 16548
rect 24412 16482 36936 16542
rect 24352 16476 24412 16482
rect 26534 16440 26594 16446
rect 28568 16440 28628 16446
rect 26594 16380 28568 16440
rect 36722 16440 36782 16446
rect 36876 16440 36936 16482
rect 38756 16440 38816 16446
rect 26534 16374 26594 16380
rect 28568 16374 28628 16380
rect 28772 16428 28832 16434
rect 28832 16368 32134 16428
rect 32194 16368 33150 16428
rect 33210 16368 36210 16428
rect 36270 16368 36276 16428
rect 36782 16380 38756 16440
rect 36722 16374 36782 16380
rect 38756 16374 38816 16380
rect 28772 16362 28832 16368
rect 24084 15492 24144 15498
rect 25516 15492 25576 15498
rect 27552 15492 27612 15498
rect 24144 15432 25516 15492
rect 25576 15432 27552 15492
rect 24084 15426 24144 15432
rect 25516 15426 25576 15432
rect 27552 15426 27612 15432
rect 35704 15492 35764 15498
rect 37740 15492 37800 15498
rect 35764 15432 37740 15492
rect 35704 15426 35764 15432
rect 24220 15362 24280 15368
rect 35834 15362 35894 15432
rect 37740 15426 37800 15432
rect 24280 15302 35894 15362
rect 24220 15296 24280 15302
rect 28574 15222 28634 15228
rect 40178 15222 40238 15228
rect 28634 15162 40178 15222
rect 28574 15156 28634 15162
rect 18760 13408 24014 13468
rect 18700 13402 18760 13408
rect 18190 13392 18250 13398
rect 30294 13238 30354 15162
rect 30294 13172 30354 13178
rect 35398 13238 35458 15162
rect 39458 13232 39518 15162
rect 40178 15156 40238 15162
rect 35398 13172 35458 13178
rect 39452 13172 39458 13232
rect 39518 13172 39524 13232
rect 4216 12972 5348 13072
rect 1875 12090 1965 12094
rect 4216 12090 4316 12972
rect 1870 12085 4316 12090
rect 1870 11995 1875 12085
rect 1965 11995 4316 12085
rect 1870 11990 4316 11995
rect 4636 12790 5024 12860
rect 1875 11986 1965 11990
rect 1574 9681 1676 9686
rect 1570 9589 1579 9681
rect 1671 9589 1680 9681
rect 1574 9539 1676 9589
rect 919 9437 1676 9539
rect 919 9387 1021 9437
rect 919 9276 1021 9285
rect 1286 4681 1390 4686
rect 1282 4587 1291 4681
rect 1385 4587 1394 4681
rect 1286 4532 1390 4587
rect 1286 4428 1746 4532
rect 1642 4366 1746 4428
rect 1642 4253 1746 4262
rect 4636 1198 4704 12790
rect 4962 1198 5024 12790
rect 5248 12784 5348 12972
rect 15478 12860 15538 12866
rect 19256 12860 19316 12866
rect 15538 12800 19256 12860
rect 15478 12794 15538 12800
rect 19256 12794 19316 12800
rect 5248 12675 5348 12684
rect 17004 12726 17064 12732
rect 18810 12726 18870 12732
rect 17064 12666 18810 12726
rect 17004 12660 17064 12666
rect 18810 12660 18870 12666
rect 19052 11502 19112 11508
rect 19112 11442 20626 11502
rect 20686 11442 20692 11502
rect 19052 11436 19112 11442
rect 21640 11286 21700 11292
rect 23680 11286 23740 11292
rect 25720 11286 25780 11292
rect 27750 11286 27810 11292
rect 29790 11286 29850 11292
rect 31822 11286 31882 11292
rect 33862 11286 33922 11292
rect 35898 11286 35958 11292
rect 37932 11286 37992 11292
rect 21700 11226 23680 11286
rect 23740 11226 25720 11286
rect 25780 11226 27750 11286
rect 27810 11226 29790 11286
rect 29850 11226 31822 11286
rect 31882 11226 33862 11286
rect 33922 11226 35898 11286
rect 35958 11226 37932 11286
rect 21640 11220 21700 11226
rect 23680 11220 23740 11226
rect 25720 11220 25780 11226
rect 27750 11220 27810 11226
rect 29790 11220 29850 11226
rect 31822 11220 31882 11226
rect 33862 11220 33922 11226
rect 35898 11220 35958 11226
rect 37932 11220 37992 11226
rect 19264 11166 19324 11172
rect 19608 11166 19668 11172
rect 19324 11106 19608 11166
rect 19264 11100 19324 11106
rect 19608 11100 19668 11106
rect 21132 11160 21192 11166
rect 29276 11160 29336 11166
rect 21192 11100 22146 11160
rect 22206 11100 23168 11160
rect 23228 11100 24182 11160
rect 24242 11100 25208 11160
rect 25268 11100 26220 11160
rect 26280 11100 27256 11160
rect 27316 11100 28262 11160
rect 28322 11100 29276 11160
rect 29336 11100 30292 11160
rect 30352 11100 31300 11160
rect 31360 11100 32316 11160
rect 32376 11100 33340 11160
rect 33400 11100 34362 11160
rect 34422 11100 35384 11160
rect 35444 11100 36402 11160
rect 36462 11100 37416 11160
rect 37476 11100 38440 11160
rect 38500 11100 38506 11160
rect 21132 11094 21192 11100
rect 29276 11094 29336 11100
rect 19482 11044 19542 11050
rect 24696 11044 24756 11050
rect 34884 11044 34944 11050
rect 38956 11044 39016 11050
rect 40088 11044 40148 11050
rect 19542 10984 24696 11044
rect 24756 10984 34884 11044
rect 34944 10984 38956 11044
rect 39016 10984 40088 11044
rect 19482 10978 19542 10984
rect 24696 10978 24756 10984
rect 34884 10978 34944 10984
rect 38956 10978 39016 10984
rect 40088 10978 40148 10984
rect 21644 10122 21704 10128
rect 23684 10122 23744 10128
rect 25716 10122 25776 10128
rect 27748 10122 27808 10128
rect 29784 10122 29844 10128
rect 31820 10122 31880 10128
rect 33858 10122 33918 10128
rect 35896 10122 35956 10128
rect 37932 10122 37992 10128
rect 21704 10062 23684 10122
rect 23744 10062 25716 10122
rect 25776 10062 27748 10122
rect 27808 10062 29784 10122
rect 29844 10062 31820 10122
rect 31880 10062 33858 10122
rect 33918 10062 35896 10122
rect 35956 10062 37932 10122
rect 21644 10056 21704 10062
rect 23684 10056 23744 10062
rect 25716 10056 25776 10062
rect 27748 10056 27808 10062
rect 29784 10056 29844 10062
rect 31820 10056 31880 10062
rect 33858 10056 33918 10062
rect 35896 10056 35956 10062
rect 37932 10056 37992 10062
rect 21136 10012 21196 10018
rect 22158 10012 22218 10018
rect 23172 10012 23232 10018
rect 24186 10012 24246 10018
rect 25204 10012 25264 10018
rect 26230 10012 26290 10018
rect 27250 10012 27310 10018
rect 28270 10012 28330 10018
rect 29272 10012 29332 10018
rect 30298 10012 30358 10018
rect 31316 10012 31376 10018
rect 32324 10012 32384 10018
rect 33336 10012 33396 10018
rect 34368 10012 34428 10018
rect 35382 10012 35442 10018
rect 36400 10012 36460 10018
rect 37424 10012 37484 10018
rect 38444 10012 38504 10018
rect 21196 9952 22158 10012
rect 22218 9952 23172 10012
rect 23232 9952 24186 10012
rect 24246 9952 25204 10012
rect 25264 9952 26230 10012
rect 26290 9952 27250 10012
rect 27310 9952 28270 10012
rect 28330 9952 29272 10012
rect 29332 9952 30298 10012
rect 30358 9952 31316 10012
rect 31376 9952 32324 10012
rect 32384 9952 33336 10012
rect 33396 9952 34368 10012
rect 34428 9952 35382 10012
rect 35442 9952 36400 10012
rect 36460 9952 37424 10012
rect 37484 9952 38444 10012
rect 21136 9946 21196 9952
rect 22158 9946 22218 9952
rect 23172 9946 23232 9952
rect 24186 9946 24246 9952
rect 25204 9946 25264 9952
rect 26230 9946 26290 9952
rect 27250 9946 27310 9952
rect 28270 9946 28330 9952
rect 29272 9946 29332 9952
rect 30298 9946 30358 9952
rect 31316 9946 31376 9952
rect 32324 9946 32384 9952
rect 33336 9946 33396 9952
rect 34368 9946 34428 9952
rect 35382 9946 35442 9952
rect 36400 9946 36460 9952
rect 37424 9946 37484 9952
rect 38444 9946 38504 9952
rect 19160 9906 19220 9912
rect 20626 9906 20686 9912
rect 22666 9906 22726 9912
rect 24696 9906 24756 9912
rect 26736 9906 26796 9912
rect 28770 9906 28830 9912
rect 30806 9906 30866 9912
rect 32842 9906 32902 9912
rect 34882 9906 34942 9912
rect 36912 9906 36972 9912
rect 38952 9906 39012 9912
rect 19220 9846 20626 9906
rect 20686 9846 22666 9906
rect 22726 9846 24696 9906
rect 24756 9846 26736 9906
rect 26796 9846 28770 9906
rect 28830 9846 30806 9906
rect 30866 9846 32842 9906
rect 32902 9846 34882 9906
rect 34942 9846 36912 9906
rect 36972 9846 38952 9906
rect 19160 9840 19220 9846
rect 20626 9840 20686 9846
rect 22666 9840 22726 9846
rect 24696 9840 24756 9846
rect 26736 9840 26796 9846
rect 28770 9840 28830 9846
rect 30806 9840 30866 9846
rect 32842 9840 32902 9846
rect 34882 9840 34942 9846
rect 36912 9840 36972 9846
rect 38952 9840 39012 9846
rect 19612 9800 19672 9806
rect 20110 9800 20170 9806
rect 20622 9800 20682 9806
rect 26902 9800 26962 9806
rect 28770 9800 28830 9806
rect 30808 9800 30868 9806
rect 32688 9800 32748 9806
rect 18920 9740 18926 9800
rect 18986 9740 19612 9800
rect 19672 9740 20110 9800
rect 20170 9740 20622 9800
rect 20682 9740 26902 9800
rect 26962 9740 28770 9800
rect 28830 9740 30808 9800
rect 30868 9740 32688 9800
rect 19612 9734 19672 9740
rect 20110 9734 20170 9740
rect 20622 9734 20682 9740
rect 26902 9734 26962 9740
rect 28770 9734 28830 9740
rect 30808 9734 30868 9740
rect 32688 9734 32748 9740
rect 36912 9802 36972 9808
rect 40088 9802 40148 9808
rect 36972 9742 40088 9802
rect 36912 9736 36972 9742
rect 40088 9736 40148 9742
rect 19482 8910 19542 8916
rect 22660 8910 22720 8916
rect 25716 8910 25776 8916
rect 31822 8910 31882 8916
rect 36916 8910 36976 8916
rect 19542 8850 22660 8910
rect 22720 8850 25716 8910
rect 25776 8850 31822 8910
rect 31882 8850 36916 8910
rect 19482 8844 19542 8850
rect 22660 8844 22720 8850
rect 25716 8844 25776 8850
rect 31822 8844 31882 8850
rect 36916 8844 36976 8850
rect 19052 8806 19112 8812
rect 19606 8806 19666 8812
rect 21126 8806 21186 8812
rect 19112 8746 19606 8806
rect 19666 8746 21126 8806
rect 19052 8740 19112 8746
rect 19606 8740 19666 8746
rect 21126 8740 21186 8746
rect 21638 8806 21698 8812
rect 22662 8806 22722 8812
rect 23674 8806 23734 8812
rect 24694 8806 24754 8812
rect 27752 8806 27812 8812
rect 29790 8806 29850 8812
rect 32840 8806 32900 8812
rect 33858 8806 33918 8812
rect 34878 8806 34938 8812
rect 35894 8806 35954 8812
rect 37930 8806 37990 8812
rect 21698 8746 22662 8806
rect 22722 8746 23674 8806
rect 23734 8746 24694 8806
rect 24754 8746 27752 8806
rect 27812 8746 29790 8806
rect 29850 8746 32840 8806
rect 32900 8746 33858 8806
rect 33918 8746 34878 8806
rect 34938 8746 35894 8806
rect 35954 8746 37930 8806
rect 21638 8740 21698 8746
rect 22662 8740 22722 8746
rect 23674 8740 23734 8746
rect 24694 8740 24754 8746
rect 27752 8740 27812 8746
rect 29790 8740 29850 8746
rect 32840 8740 32900 8746
rect 33858 8740 33918 8746
rect 34878 8740 34938 8746
rect 35894 8740 35954 8746
rect 37930 8740 37990 8746
rect 19376 8684 19436 8690
rect 26736 8684 26796 8690
rect 28770 8684 28830 8690
rect 30800 8684 30860 8690
rect 40800 8684 40860 17642
rect 19436 8624 26736 8684
rect 26796 8624 28770 8684
rect 28830 8624 30800 8684
rect 30860 8624 40860 8684
rect 19376 8618 19436 8624
rect 26736 8618 26796 8624
rect 28770 8618 28830 8624
rect 30800 8618 30860 8624
rect 19264 8570 19324 8576
rect 20112 8570 20172 8576
rect 19324 8510 20112 8570
rect 19264 8504 19324 8510
rect 20112 8504 20172 8510
rect 21644 8572 21704 8578
rect 23680 8572 23740 8578
rect 40074 8572 40134 8578
rect 21704 8512 23680 8572
rect 23740 8512 40074 8572
rect 21644 8506 21704 8512
rect 23680 8506 23740 8512
rect 40074 8506 40134 8512
rect 40202 8554 40262 8560
rect 40802 8554 40862 8560
rect 40262 8494 40802 8554
rect 40202 8488 40262 8494
rect 40802 8488 40862 8494
rect 39968 7684 40028 7690
rect 40928 7684 40988 17960
rect 22660 7666 22720 7672
rect 24696 7666 24756 7672
rect 32840 7666 32900 7672
rect 34876 7666 34936 7672
rect 38950 7666 39010 7672
rect 19488 7642 19548 7648
rect 20626 7642 20686 7648
rect 19548 7582 20626 7642
rect 20686 7582 21508 7642
rect 22720 7606 24696 7666
rect 24756 7606 32840 7666
rect 32900 7606 34876 7666
rect 34936 7606 38950 7666
rect 40028 7624 40988 7684
rect 39968 7618 40028 7624
rect 22660 7600 22720 7606
rect 24696 7600 24756 7606
rect 32840 7600 32900 7606
rect 34876 7600 34936 7606
rect 38950 7600 39010 7606
rect 19488 7576 19548 7582
rect 20626 7576 20686 7582
rect 19376 7442 19436 7448
rect 20624 7442 20684 7448
rect 19436 7382 20624 7442
rect 21448 7446 21508 7582
rect 21642 7562 21702 7568
rect 23682 7562 23742 7568
rect 25714 7562 25774 7568
rect 27748 7562 27808 7568
rect 29788 7562 29848 7568
rect 31822 7562 31882 7568
rect 21702 7502 23682 7562
rect 23742 7502 25714 7562
rect 25774 7502 27748 7562
rect 27808 7502 29788 7562
rect 29848 7502 31822 7562
rect 21642 7496 21702 7502
rect 23682 7496 23742 7502
rect 25714 7496 25774 7502
rect 27748 7496 27808 7502
rect 29788 7496 29848 7502
rect 31822 7496 31882 7502
rect 32018 7558 32078 7564
rect 36910 7558 36970 7564
rect 32078 7498 36910 7558
rect 40568 7554 40628 7560
rect 32018 7492 32078 7498
rect 36910 7492 36970 7498
rect 37408 7494 37414 7554
rect 37474 7494 40568 7554
rect 40568 7488 40628 7494
rect 22156 7448 22216 7454
rect 25714 7450 25774 7456
rect 27750 7450 27810 7456
rect 29786 7450 29846 7456
rect 31822 7450 31882 7456
rect 33856 7450 33916 7456
rect 35894 7450 35954 7456
rect 37934 7450 37994 7456
rect 40318 7450 40378 7456
rect 21448 7388 22156 7446
rect 22216 7388 23160 7448
rect 23220 7388 24172 7448
rect 24232 7388 25192 7448
rect 25252 7388 25258 7448
rect 25774 7390 27750 7450
rect 27810 7390 29786 7450
rect 29846 7390 31822 7450
rect 31882 7390 33856 7450
rect 33916 7390 35894 7450
rect 35954 7390 37934 7450
rect 37994 7390 40318 7450
rect 21448 7386 22498 7388
rect 22156 7382 22216 7386
rect 25714 7384 25774 7390
rect 27750 7384 27810 7390
rect 29786 7384 29846 7390
rect 31822 7384 31882 7390
rect 33856 7384 33916 7390
rect 35894 7384 35954 7390
rect 37934 7384 37994 7390
rect 40318 7384 40378 7390
rect 19376 7376 19436 7382
rect 20624 7376 20684 7382
rect 18700 7340 18760 7346
rect 19270 7340 19330 7346
rect 26732 7340 26792 7346
rect 28766 7340 28826 7346
rect 30806 7340 30866 7346
rect 32018 7340 32078 7346
rect 18760 7280 19270 7340
rect 19330 7280 26732 7340
rect 26792 7280 28766 7340
rect 28826 7280 30806 7340
rect 30866 7280 32018 7340
rect 18700 7274 18760 7280
rect 19270 7274 19330 7280
rect 26732 7274 26792 7280
rect 28766 7274 28826 7280
rect 30806 7274 30866 7280
rect 32018 7274 32078 7280
rect 32312 7342 32372 7348
rect 32372 7282 33340 7342
rect 33400 7282 33406 7342
rect 33858 7336 33918 7342
rect 35894 7336 35954 7342
rect 37932 7336 37992 7342
rect 40074 7336 40134 7342
rect 32312 7276 32372 7282
rect 33918 7276 35894 7336
rect 35954 7276 37932 7336
rect 37992 7276 40074 7336
rect 33858 7270 33918 7276
rect 35894 7270 35954 7276
rect 37932 7270 37992 7276
rect 40074 7270 40134 7276
rect 36406 6422 36466 6428
rect 20624 6410 20684 6416
rect 22662 6410 22722 6416
rect 24698 6410 24758 6416
rect 26730 6410 26790 6416
rect 20684 6350 22662 6410
rect 22722 6350 24698 6410
rect 24758 6350 26730 6410
rect 31306 6362 31312 6422
rect 31372 6362 36406 6422
rect 36406 6356 36466 6362
rect 36544 6426 36604 6432
rect 37426 6426 37486 6432
rect 38432 6426 38492 6432
rect 36604 6366 37426 6426
rect 37486 6366 38432 6426
rect 36544 6360 36604 6366
rect 37426 6360 37486 6366
rect 38432 6360 38492 6366
rect 38950 6422 39010 6428
rect 40202 6422 40262 6428
rect 39010 6362 40202 6422
rect 38950 6356 39010 6362
rect 40202 6356 40262 6362
rect 20624 6344 20684 6350
rect 22662 6344 22722 6350
rect 24698 6344 24758 6350
rect 26730 6344 26790 6350
rect 21130 6308 21190 6314
rect 26222 6308 26282 6314
rect 18190 6258 18250 6264
rect 21190 6248 26222 6308
rect 21130 6242 21190 6248
rect 26222 6242 26282 6248
rect 30806 6294 30866 6300
rect 38950 6294 39010 6300
rect 30866 6234 38950 6294
rect 30806 6228 30866 6234
rect 38950 6228 39010 6234
rect 13642 5332 13702 5338
rect 18190 5332 18250 6198
rect 19376 6206 19436 6212
rect 22660 6206 22720 6212
rect 19436 6146 22660 6206
rect 19376 6140 19436 6146
rect 22660 6140 22720 6146
rect 23168 6200 23228 6206
rect 24190 6200 24250 6206
rect 25204 6200 25264 6206
rect 26222 6200 26282 6206
rect 27242 6200 27302 6206
rect 34354 6200 34414 6206
rect 35384 6200 35444 6206
rect 36544 6200 36604 6206
rect 23228 6140 24190 6200
rect 24250 6140 25204 6200
rect 25264 6140 26222 6200
rect 26282 6140 27242 6200
rect 27302 6140 34354 6200
rect 34414 6140 35384 6200
rect 35444 6140 36544 6200
rect 23168 6134 23228 6140
rect 24190 6134 24250 6140
rect 25204 6134 25264 6140
rect 26222 6134 26282 6140
rect 27242 6134 27302 6140
rect 34354 6134 34414 6140
rect 35384 6134 35444 6140
rect 36544 6134 36604 6140
rect 36912 6200 36972 6206
rect 40440 6200 40500 6206
rect 36972 6140 40440 6200
rect 36912 6134 36972 6140
rect 40440 6134 40500 6140
rect 21644 6106 21704 6112
rect 23678 6106 23738 6112
rect 25714 6106 25774 6112
rect 21704 6046 23678 6106
rect 23738 6046 25714 6106
rect 21644 6040 21704 6046
rect 23678 6040 23738 6046
rect 25714 6040 25774 6046
rect 32842 6096 32902 6102
rect 36912 6096 36972 6102
rect 32902 6036 36912 6096
rect 32842 6030 32902 6036
rect 36912 6030 36972 6036
rect 37928 6098 37988 6104
rect 40318 6098 40378 6104
rect 37988 6038 40318 6098
rect 37928 6032 37988 6038
rect 40318 6032 40378 6038
rect 13702 5272 18250 5332
rect 13642 5266 13702 5272
rect 11612 5186 11672 5192
rect 15672 5186 15732 5192
rect 17856 5186 17916 5192
rect 18322 5186 18382 5192
rect 27750 5188 27810 5194
rect 29786 5188 29846 5194
rect 31822 5188 31882 5194
rect 33860 5188 33920 5194
rect 7526 5126 7532 5186
rect 7592 5126 11612 5186
rect 11672 5126 15672 5186
rect 15732 5126 17856 5186
rect 17916 5126 18322 5186
rect 11612 5120 11672 5126
rect 15672 5120 15732 5126
rect 17856 5120 17916 5126
rect 18322 5120 18382 5126
rect 21126 5182 21186 5188
rect 22036 5182 22096 5188
rect 23038 5182 23098 5188
rect 24190 5182 24250 5188
rect 25200 5182 25260 5188
rect 26206 5182 26266 5188
rect 27250 5182 27310 5188
rect 21186 5122 22036 5182
rect 22096 5122 23038 5182
rect 23098 5122 24190 5182
rect 24250 5122 25200 5182
rect 25260 5122 26206 5182
rect 26266 5122 27250 5182
rect 27810 5128 29786 5188
rect 29846 5128 31822 5188
rect 31882 5128 33860 5188
rect 27750 5122 27810 5128
rect 29786 5122 29846 5128
rect 31822 5122 31882 5128
rect 33860 5122 33920 5128
rect 35896 5188 35956 5194
rect 37934 5188 37994 5194
rect 35956 5128 37934 5188
rect 35896 5122 35956 5128
rect 37934 5122 37994 5128
rect 21126 5116 21186 5122
rect 22036 5116 22096 5122
rect 23038 5116 23098 5122
rect 24190 5116 24250 5122
rect 25200 5116 25260 5122
rect 26206 5116 26266 5122
rect 27250 5116 27310 5122
rect 23678 5080 23738 5086
rect 33852 5080 33912 5086
rect 35892 5080 35952 5086
rect 37930 5080 37990 5086
rect 6378 5058 6438 5064
rect 9056 5058 9116 5064
rect 10088 5058 10148 5064
rect 13148 5058 13208 5064
rect 14144 5058 14204 5064
rect 18442 5058 18502 5064
rect 6438 4998 9056 5058
rect 9116 4998 10088 5058
rect 10148 4998 13148 5058
rect 13208 4998 14144 5058
rect 14204 4998 18442 5058
rect 23738 5020 33852 5080
rect 33912 5020 35892 5080
rect 35952 5020 37930 5080
rect 23678 5014 23738 5020
rect 33852 5014 33912 5020
rect 35892 5014 35952 5020
rect 37930 5014 37990 5020
rect 6378 4992 6438 4998
rect 9056 4992 9116 4998
rect 10088 4992 10148 4998
rect 13148 4992 13208 4998
rect 14144 4992 14204 4998
rect 18442 4992 18502 4998
rect 21126 4966 21186 4972
rect 23178 4966 23238 4972
rect 26204 4966 26264 4972
rect 27244 4966 27304 4972
rect 28258 4966 28318 4972
rect 29266 4966 29326 4972
rect 30310 4966 30370 4972
rect 31300 4966 31360 4972
rect 32318 4966 32378 4972
rect 33352 4966 33412 4972
rect 36384 4966 36444 4972
rect 37422 4966 37482 4972
rect 38448 4966 38508 4972
rect 21186 4906 22164 4966
rect 22224 4906 23178 4966
rect 23238 4906 26204 4966
rect 26264 4906 27244 4966
rect 27304 4906 28258 4966
rect 28318 4906 29266 4966
rect 29326 4906 30310 4966
rect 30370 4906 31300 4966
rect 31360 4906 32318 4966
rect 32378 4906 33352 4966
rect 33412 4906 36384 4966
rect 36444 4906 37422 4966
rect 37482 4906 38448 4966
rect 38508 4906 40566 4966
rect 40626 4906 40632 4966
rect 21126 4900 21186 4906
rect 23178 4900 23238 4906
rect 26204 4900 26264 4906
rect 27244 4900 27304 4906
rect 28258 4900 28318 4906
rect 29266 4900 29326 4906
rect 30310 4900 30370 4906
rect 31300 4900 31360 4906
rect 32318 4900 32378 4906
rect 33352 4900 33412 4906
rect 36384 4900 36444 4906
rect 37422 4900 37482 4906
rect 38448 4900 38508 4906
rect 26728 4862 26788 4868
rect 28770 4862 28830 4868
rect 30808 4862 30868 4868
rect 32842 4862 32902 4868
rect 34876 4864 34936 4870
rect 36910 4864 36970 4870
rect 38952 4864 39012 4870
rect 40202 4864 40262 4870
rect 19484 4802 19490 4862
rect 19550 4802 26728 4862
rect 26788 4802 28770 4862
rect 28830 4802 30808 4862
rect 30868 4802 32842 4862
rect 26728 4796 26788 4802
rect 28770 4796 28830 4802
rect 30808 4796 30868 4802
rect 32842 4796 32902 4802
rect 33354 4858 33414 4864
rect 34376 4858 34436 4864
rect 33414 4798 34376 4858
rect 34936 4804 36910 4864
rect 36970 4804 38952 4864
rect 39012 4804 40202 4864
rect 34876 4798 34936 4804
rect 36910 4798 36970 4804
rect 38952 4798 39012 4804
rect 40202 4798 40262 4804
rect 33354 4792 33414 4798
rect 34376 4792 34436 4798
rect 8036 4096 8096 4102
rect 9060 4096 9120 4102
rect 10092 4096 10152 4102
rect 11092 4096 11152 4102
rect 12112 4096 12172 4102
rect 13132 4096 13192 4102
rect 15156 4096 15216 4102
rect 17976 4096 18036 4102
rect 18582 4096 18642 4102
rect 8096 4036 9060 4096
rect 9120 4036 10092 4096
rect 10152 4036 11092 4096
rect 11152 4036 12112 4096
rect 12172 4036 13132 4096
rect 13192 4036 14142 4096
rect 14202 4036 15156 4096
rect 15216 4036 16174 4096
rect 16234 4036 17976 4096
rect 18036 4036 18582 4096
rect 8036 4030 8096 4036
rect 9060 4030 9120 4036
rect 10092 4030 10152 4036
rect 11092 4030 11152 4036
rect 12112 4030 12172 4036
rect 13132 4030 13192 4036
rect 15156 4030 15216 4036
rect 17976 4030 18036 4036
rect 18582 4030 18642 4036
rect 7536 3992 7596 3998
rect 9572 3992 9632 3998
rect 11608 3992 11668 3998
rect 13642 3992 13702 3998
rect 15678 3992 15738 3998
rect 7596 3932 9572 3992
rect 9632 3932 11608 3992
rect 11668 3932 13642 3992
rect 13702 3932 15678 3992
rect 25718 3960 25778 3966
rect 29786 3960 29846 3966
rect 31820 3960 31880 3966
rect 7536 3926 7596 3932
rect 9572 3926 9632 3932
rect 11608 3926 11668 3932
rect 13642 3926 13702 3932
rect 15678 3926 15738 3932
rect 21124 3954 21184 3960
rect 22132 3954 22192 3960
rect 23146 3954 23206 3960
rect 24184 3954 24244 3960
rect 25202 3954 25262 3960
rect 21184 3894 22132 3954
rect 22192 3894 23146 3954
rect 23206 3894 24184 3954
rect 24244 3894 25202 3954
rect 25778 3900 27754 3960
rect 27814 3900 29786 3960
rect 29846 3900 31820 3960
rect 25718 3894 25778 3900
rect 29786 3894 29846 3900
rect 31820 3894 31880 3900
rect 32842 3962 32902 3968
rect 33196 3962 33256 3968
rect 32902 3902 33196 3962
rect 32842 3896 32902 3902
rect 33196 3896 33256 3902
rect 36914 3962 36974 3968
rect 40198 3962 40258 3968
rect 36974 3902 40198 3962
rect 36914 3896 36974 3902
rect 40198 3896 40258 3902
rect 12622 3888 12682 3894
rect 19160 3888 19220 3894
rect 21124 3888 21184 3894
rect 22132 3888 22192 3894
rect 23146 3888 23206 3894
rect 24184 3888 24244 3894
rect 25202 3888 25262 3894
rect 8548 3828 8554 3888
rect 8614 3828 10590 3888
rect 10650 3828 12622 3888
rect 12682 3828 14656 3888
rect 14716 3828 16700 3888
rect 16760 3828 19160 3888
rect 12622 3822 12682 3828
rect 19160 3822 19220 3828
rect 19270 3850 19330 3856
rect 20626 3850 20686 3856
rect 28770 3850 28830 3856
rect 30806 3850 30866 3856
rect 32838 3850 32898 3856
rect 19330 3790 20626 3850
rect 20686 3790 28770 3850
rect 28830 3790 30806 3850
rect 30866 3790 32838 3850
rect 19270 3784 19330 3790
rect 20626 3784 20686 3790
rect 28770 3784 28830 3790
rect 30806 3784 30866 3790
rect 32838 3784 32898 3790
rect 32348 3752 32408 3758
rect 33386 3752 33446 3758
rect 34362 3752 34422 3758
rect 35378 3752 35438 3758
rect 37404 3752 37464 3758
rect 38434 3752 38494 3758
rect 18928 3738 18988 3744
rect 21642 3738 21702 3744
rect 23680 3738 23740 3744
rect 27752 3738 27812 3744
rect 18988 3678 21642 3738
rect 21702 3678 23680 3738
rect 23740 3678 27752 3738
rect 32408 3692 33386 3752
rect 33446 3692 34362 3752
rect 34422 3692 35378 3752
rect 35438 3692 37404 3752
rect 37464 3692 38434 3752
rect 32348 3686 32408 3692
rect 33386 3686 33446 3692
rect 34362 3686 34422 3692
rect 35378 3686 35438 3692
rect 37404 3686 37464 3692
rect 38434 3686 38494 3692
rect 18928 3672 18988 3678
rect 21642 3672 21702 3678
rect 23680 3672 23740 3678
rect 27752 3672 27812 3678
rect 20622 3640 20682 3646
rect 22660 3640 22720 3646
rect 24700 3640 24760 3646
rect 26736 3640 26796 3646
rect 32840 3640 32900 3646
rect 33190 3640 33196 3644
rect 20682 3580 22660 3640
rect 22720 3580 24700 3640
rect 24760 3580 26736 3640
rect 26796 3584 33196 3640
rect 33256 3640 33262 3644
rect 34876 3640 34936 3646
rect 36912 3640 36972 3646
rect 38948 3640 39008 3646
rect 33256 3584 34876 3640
rect 26796 3580 34876 3584
rect 34936 3580 36912 3640
rect 36972 3580 38948 3640
rect 20622 3574 20682 3580
rect 22660 3574 22720 3580
rect 24700 3574 24760 3580
rect 26736 3574 26796 3580
rect 32840 3574 32900 3580
rect 34876 3574 34936 3580
rect 36912 3574 36972 3580
rect 38948 3574 39008 3580
rect 9566 2946 9626 2952
rect 13642 2946 13702 2952
rect 17856 2946 17916 2952
rect 9626 2886 13642 2946
rect 13702 2886 17856 2946
rect 9566 2880 9626 2886
rect 13642 2880 13702 2886
rect 17856 2880 17916 2886
rect 6378 2826 6438 2832
rect 8028 2826 8088 2832
rect 11098 2826 11158 2832
rect 12106 2826 12166 2832
rect 15168 2826 15228 2832
rect 16194 2826 16254 2832
rect 6438 2766 8028 2826
rect 8088 2766 11098 2826
rect 11158 2766 12106 2826
rect 12166 2766 15168 2826
rect 15228 2766 16194 2826
rect 6378 2760 6438 2766
rect 8028 2760 8088 2766
rect 11098 2760 11158 2766
rect 12106 2760 12166 2766
rect 15168 2760 15228 2766
rect 16194 2760 16254 2766
rect 27748 2736 27808 2742
rect 29790 2736 29850 2742
rect 31822 2736 31882 2742
rect 33862 2736 33922 2742
rect 40318 2736 40378 2742
rect 21642 2716 21702 2722
rect 23678 2716 23738 2722
rect 25716 2716 25776 2722
rect 21702 2656 23678 2716
rect 23738 2656 25716 2716
rect 27572 2676 27578 2736
rect 27638 2676 27748 2736
rect 27808 2676 29790 2736
rect 29850 2676 31822 2736
rect 31882 2676 33862 2736
rect 33922 2676 40318 2736
rect 27748 2670 27808 2676
rect 29790 2670 29850 2676
rect 31822 2670 31882 2676
rect 33862 2670 33922 2676
rect 40318 2670 40378 2676
rect 21642 2650 21702 2656
rect 23678 2650 23738 2656
rect 25716 2650 25776 2656
rect 32840 2638 32900 2644
rect 38946 2638 39006 2644
rect 40198 2638 40258 2644
rect 19488 2618 19548 2624
rect 22660 2618 22720 2624
rect 19548 2558 22660 2618
rect 19488 2552 19548 2558
rect 22660 2552 22720 2558
rect 24184 2618 24244 2624
rect 27232 2618 27292 2624
rect 24244 2558 25206 2618
rect 25266 2558 26228 2618
rect 26288 2558 27232 2618
rect 32900 2578 38946 2638
rect 39006 2578 40198 2638
rect 32840 2572 32900 2578
rect 38946 2572 39006 2578
rect 40198 2572 40258 2578
rect 24184 2552 24244 2558
rect 27232 2552 27292 2558
rect 27754 2528 27814 2534
rect 29782 2528 29842 2534
rect 31826 2528 31886 2534
rect 33854 2528 33914 2534
rect 35892 2528 35952 2534
rect 37932 2528 37992 2534
rect 21646 2522 21706 2528
rect 23682 2522 23742 2528
rect 25710 2522 25770 2528
rect 27578 2522 27638 2528
rect 21706 2462 23682 2522
rect 23742 2462 25710 2522
rect 25770 2462 27578 2522
rect 27814 2468 29782 2528
rect 29842 2468 31826 2528
rect 31886 2468 33854 2528
rect 33914 2468 35892 2528
rect 35952 2468 37932 2528
rect 27754 2462 27814 2468
rect 29782 2462 29842 2468
rect 31826 2462 31886 2468
rect 33854 2462 33914 2468
rect 35892 2462 35952 2468
rect 37932 2462 37992 2468
rect 38450 2532 38510 2538
rect 39962 2532 40022 2538
rect 40568 2532 40628 2538
rect 38510 2472 39962 2532
rect 40022 2472 40568 2532
rect 38450 2466 38510 2472
rect 39962 2466 40022 2472
rect 40568 2466 40628 2472
rect 21646 2456 21706 2462
rect 23682 2456 23742 2462
rect 25710 2456 25770 2462
rect 27578 2456 27638 2462
rect 20628 2402 20688 2408
rect 24696 2402 24756 2408
rect 26730 2402 26790 2408
rect 34880 2402 34940 2408
rect 36910 2402 36970 2408
rect 38950 2404 39010 2410
rect 40440 2404 40500 2410
rect 20688 2342 24696 2402
rect 24756 2342 26730 2402
rect 26790 2342 34880 2402
rect 34940 2342 36910 2402
rect 37430 2344 37436 2404
rect 37496 2344 38950 2404
rect 39010 2344 40440 2404
rect 20628 2336 20688 2342
rect 24696 2336 24756 2342
rect 26730 2336 26790 2342
rect 34880 2336 34940 2342
rect 36910 2336 36970 2342
rect 38950 2338 39010 2344
rect 40440 2338 40500 2344
rect 16700 1882 16760 1888
rect 8548 1822 8554 1882
rect 8614 1822 10590 1882
rect 10650 1822 12622 1882
rect 12682 1822 14656 1882
rect 14716 1822 16700 1882
rect 16700 1816 16760 1822
rect 7540 1774 7600 1780
rect 9576 1774 9636 1780
rect 11612 1774 11672 1780
rect 13646 1774 13706 1780
rect 15682 1774 15742 1780
rect 7600 1714 9576 1774
rect 9636 1714 11612 1774
rect 11672 1714 13646 1774
rect 13706 1714 15682 1774
rect 7540 1708 7600 1714
rect 9576 1708 9636 1714
rect 11612 1708 11672 1714
rect 13646 1708 13706 1714
rect 15682 1708 15742 1714
rect 8034 1662 8094 1668
rect 9058 1662 9118 1668
rect 10090 1662 10150 1668
rect 11090 1662 11150 1668
rect 12110 1662 12170 1668
rect 13130 1662 13190 1668
rect 15154 1662 15214 1668
rect 17976 1662 18036 1668
rect 4636 1148 5024 1198
rect 5564 1602 8034 1662
rect 8094 1602 9058 1662
rect 9118 1602 10090 1662
rect 10150 1602 11090 1662
rect 11150 1602 12110 1662
rect 12170 1602 13130 1662
rect 13190 1602 14140 1662
rect 14200 1602 15154 1662
rect 15214 1602 16172 1662
rect 16232 1602 17976 1662
rect -202 986 4964 1026
rect -202 896 -156 986
rect 4924 896 4964 986
rect -202 846 4964 896
rect -2 748 58 754
rect 790 748 850 754
rect 3366 748 3426 754
rect 4134 748 4194 754
rect 58 688 790 748
rect 850 688 3366 748
rect 3426 688 4134 748
rect -2 682 58 688
rect 790 682 850 688
rect 3366 682 3426 688
rect 4134 682 4194 688
rect 1033 639 1123 648
rect 142 624 202 630
rect 202 564 1033 624
rect 142 558 202 564
rect 1818 624 1878 630
rect 2338 624 2398 630
rect 3998 624 4058 630
rect 5564 624 5624 1602
rect 8034 1596 8094 1602
rect 9058 1596 9118 1602
rect 10090 1596 10150 1602
rect 11090 1596 11150 1602
rect 12110 1596 12170 1602
rect 13130 1596 13190 1602
rect 15154 1596 15214 1602
rect 17976 1596 18036 1602
rect 19376 1486 19436 1492
rect 28764 1486 28824 1492
rect 30806 1486 30866 1492
rect 32842 1486 32902 1492
rect 19436 1426 28764 1486
rect 28824 1426 30806 1486
rect 30866 1426 32842 1486
rect 19376 1420 19436 1426
rect 28764 1420 28824 1426
rect 30806 1420 30866 1426
rect 32842 1420 32902 1426
rect 35896 1486 35956 1492
rect 37928 1486 37988 1492
rect 40074 1486 40134 1492
rect 35956 1426 37928 1486
rect 37988 1426 40074 1486
rect 35896 1420 35956 1426
rect 37928 1420 37988 1426
rect 40074 1420 40134 1426
rect 23180 1372 23240 1378
rect 28260 1372 28320 1378
rect 19270 1360 19330 1366
rect 22660 1360 22720 1366
rect 19330 1300 22660 1360
rect 23240 1312 28260 1372
rect 23180 1306 23240 1312
rect 28260 1306 28320 1312
rect 33348 1376 33408 1382
rect 38448 1376 38508 1382
rect 33408 1316 38448 1376
rect 33348 1310 33408 1316
rect 38448 1310 38508 1316
rect 39456 1376 39516 1382
rect 40690 1376 40750 1382
rect 39516 1316 40690 1376
rect 39456 1310 39516 1316
rect 40690 1310 40750 1316
rect 19270 1294 19330 1300
rect 22660 1294 22720 1300
rect 21642 1258 21702 1264
rect 23678 1258 23738 1264
rect 24698 1258 24758 1264
rect 25714 1258 25774 1264
rect 26734 1258 26794 1264
rect 27752 1258 27812 1264
rect 29782 1258 29842 1264
rect 31820 1258 31880 1264
rect 33856 1258 33916 1264
rect 34878 1258 34938 1264
rect 35898 1258 35958 1264
rect 36912 1258 36972 1264
rect 37934 1258 37994 1264
rect 21702 1198 23678 1258
rect 23738 1198 24698 1258
rect 24758 1198 25714 1258
rect 25774 1198 26734 1258
rect 26794 1198 27752 1258
rect 27812 1198 29782 1258
rect 29842 1198 31820 1258
rect 31880 1198 33856 1258
rect 33916 1198 34878 1258
rect 34938 1198 35898 1258
rect 35958 1198 36912 1258
rect 36972 1198 37934 1258
rect 21642 1192 21702 1198
rect 23678 1192 23738 1198
rect 24698 1192 24758 1198
rect 25714 1192 25774 1198
rect 26734 1192 26794 1198
rect 27752 1192 27812 1198
rect 29782 1192 29842 1198
rect 31820 1192 31880 1198
rect 33856 1192 33916 1198
rect 34878 1192 34938 1198
rect 35898 1192 35958 1198
rect 36912 1192 36972 1198
rect 37934 1192 37994 1198
rect 22660 1154 22720 1160
rect 27596 1154 27656 1160
rect 34002 1154 34062 1160
rect 36912 1154 36972 1160
rect 40094 1154 40154 1160
rect 22720 1094 27596 1154
rect 27656 1094 34002 1154
rect 34062 1094 36912 1154
rect 36972 1094 40094 1154
rect 22660 1088 22720 1094
rect 27596 1088 27656 1094
rect 34002 1088 34062 1094
rect 36912 1088 36972 1094
rect 40094 1088 40154 1094
rect 6378 700 6438 706
rect 9048 700 9108 706
rect 10080 700 10140 706
rect 13140 700 13200 706
rect 14136 700 14196 706
rect 6438 640 9048 700
rect 9108 640 10080 700
rect 10140 640 13140 700
rect 13200 640 14136 700
rect 6378 634 6508 640
rect 9048 634 9108 640
rect 10080 634 10140 640
rect 13140 634 13200 640
rect 14136 634 14196 640
rect 1123 564 1818 624
rect 1878 564 2338 624
rect 2398 564 3998 624
rect 4058 564 5624 624
rect 1818 558 1878 564
rect 2338 558 2398 564
rect 3998 558 4058 564
rect 1033 540 1123 549
rect 662 -110 722 -104
rect 920 -108 980 -102
rect 722 -168 920 -110
rect 1692 -110 1752 -104
rect 1952 -110 2012 -104
rect 2208 -110 2268 -104
rect 2466 -110 2526 -104
rect 3242 -110 3302 -104
rect 3502 -110 3562 -104
rect 980 -168 1692 -110
rect 722 -170 1692 -168
rect 1752 -170 1952 -110
rect 2012 -170 2208 -110
rect 2268 -170 2466 -110
rect 2526 -170 3242 -110
rect 3302 -170 3502 -110
rect 662 -176 722 -170
rect 920 -174 980 -170
rect 1692 -176 1752 -170
rect 1952 -176 2012 -170
rect 2208 -176 2268 -170
rect 2466 -176 2526 -170
rect 3242 -176 3302 -170
rect 3502 -176 3562 -170
rect 790 -240 850 -234
rect 1564 -240 1624 -234
rect 2080 -240 2140 -234
rect 2598 -240 2658 -234
rect 3368 -240 3428 -234
rect 850 -300 1564 -240
rect 1624 -300 2080 -240
rect 2140 -300 2598 -240
rect 2658 -300 3368 -240
rect 3428 -300 5112 -240
rect 5172 -300 5181 -240
rect 790 -306 850 -300
rect 1564 -306 1624 -300
rect 2080 -306 2140 -300
rect 2598 -306 2658 -300
rect 3368 -306 3428 -300
rect 3607 -341 3697 -332
rect 532 -358 592 -352
rect 1050 -358 1110 -352
rect 1822 -358 1882 -352
rect 2336 -358 2396 -352
rect 3112 -358 3172 -352
rect 6448 -358 6508 634
rect 11614 570 11674 576
rect 15674 570 15734 576
rect 17856 570 17916 576
rect 7528 510 7534 570
rect 7594 510 11614 570
rect 11674 510 15674 570
rect 15734 510 17856 570
rect 11614 504 11674 510
rect 15674 504 15734 510
rect 17856 504 17916 510
rect 19488 256 19548 262
rect 22658 256 22718 262
rect 19548 196 22658 256
rect 19488 190 19548 196
rect 22658 190 22718 196
rect 26888 258 26948 264
rect 28766 258 28826 264
rect 30804 258 30864 264
rect 32674 258 32734 264
rect 38950 258 39010 264
rect 26948 198 28766 258
rect 28826 198 30804 258
rect 30864 198 32674 258
rect 32734 198 38950 258
rect 26888 192 26948 198
rect 28766 192 28826 198
rect 30804 192 30864 198
rect 32674 192 32734 198
rect 38950 192 39010 198
rect 19160 152 19220 158
rect 20624 152 20684 158
rect 22664 152 22724 158
rect 24694 152 24754 158
rect 26734 152 26794 158
rect 28770 152 28830 158
rect 30806 152 30866 158
rect 32840 152 32900 158
rect 34880 152 34940 158
rect 36910 152 36970 158
rect 38950 152 39010 158
rect 40802 152 40862 158
rect 19220 92 20624 152
rect 20684 92 22664 152
rect 22724 92 24694 152
rect 24754 92 26734 152
rect 26794 92 28770 152
rect 28830 92 30806 152
rect 30866 92 32840 152
rect 32900 92 34880 152
rect 34940 92 36910 152
rect 36970 92 38950 152
rect 39010 92 40802 152
rect 19160 86 19220 92
rect 20624 86 20684 92
rect 22664 86 22724 92
rect 24694 86 24754 92
rect 26734 86 26794 92
rect 28770 86 28830 92
rect 30806 86 30866 92
rect 32840 86 32900 92
rect 34880 86 34940 92
rect 36910 86 36970 92
rect 38950 86 39010 92
rect 40802 86 40862 92
rect 21132 46 21192 52
rect 22152 46 22212 52
rect 23176 46 23236 52
rect 24194 46 24254 52
rect 25208 46 25268 52
rect 26240 46 26300 52
rect 27252 46 27312 52
rect 28260 46 28320 52
rect 29278 46 29338 52
rect 30304 46 30364 52
rect 31306 46 31366 52
rect 32326 46 32386 52
rect 33346 46 33406 52
rect 34372 46 34432 52
rect 35390 46 35450 52
rect 36404 46 36464 52
rect 37418 46 37478 52
rect 38440 46 38500 52
rect 21192 -14 22152 46
rect 22212 -14 23176 46
rect 23236 -14 24194 46
rect 24254 -14 25208 46
rect 25268 -14 26240 46
rect 26300 -14 27252 46
rect 27312 -14 28260 46
rect 28320 -14 29278 46
rect 29338 -14 30304 46
rect 30364 -14 31306 46
rect 31366 -14 32326 46
rect 32386 -14 33346 46
rect 33406 -14 34372 46
rect 34432 -14 35390 46
rect 35450 -14 36404 46
rect 36464 -14 37418 46
rect 37478 -14 38440 46
rect 21132 -20 21192 -14
rect 22152 -20 22212 -14
rect 23176 -20 23236 -14
rect 24194 -20 24254 -14
rect 25208 -20 25268 -14
rect 26240 -20 26300 -14
rect 27252 -20 27312 -14
rect 28260 -20 28320 -14
rect 29278 -20 29338 -14
rect 30304 -20 30364 -14
rect 31306 -20 31366 -14
rect 32326 -20 32386 -14
rect 33346 -20 33406 -14
rect 34372 -20 34432 -14
rect 35390 -20 35450 -14
rect 36404 -20 36464 -14
rect 37418 -20 37478 -14
rect 38440 -20 38500 -14
rect 21644 -64 21704 -58
rect 23680 -64 23740 -58
rect 25718 -64 25778 -58
rect 27756 -64 27816 -58
rect 29792 -64 29852 -58
rect 31828 -64 31888 -58
rect 33860 -64 33920 -58
rect 35892 -64 35952 -58
rect 37932 -64 37992 -58
rect 21704 -124 23680 -64
rect 23740 -124 25718 -64
rect 25778 -124 27756 -64
rect 27816 -124 29792 -64
rect 29852 -124 31828 -64
rect 31888 -124 33860 -64
rect 33920 -124 35892 -64
rect 35952 -124 37932 -64
rect 21644 -130 21704 -124
rect 23680 -130 23740 -124
rect 25718 -130 25778 -124
rect 27756 -130 27816 -124
rect 29792 -130 29852 -124
rect 31828 -130 31888 -124
rect 33860 -130 33920 -124
rect 35892 -130 35952 -124
rect 37932 -130 37992 -124
rect 592 -418 1050 -358
rect 1110 -418 1822 -358
rect 1882 -418 2336 -358
rect 2396 -418 3112 -358
rect 3172 -418 3607 -358
rect 3697 -418 6508 -358
rect 532 -424 592 -418
rect 1050 -424 1110 -418
rect 1822 -424 1882 -418
rect 2336 -424 2396 -418
rect 3112 -424 3172 -418
rect 3607 -440 3697 -431
rect 9012 -796 9072 -790
rect 11050 -796 11110 -790
rect 13086 -796 13146 -790
rect 15122 -796 15182 -790
rect 9072 -856 11050 -796
rect 11110 -856 13086 -796
rect 13146 -856 15122 -796
rect 9012 -862 9072 -856
rect 11050 -862 11110 -856
rect 13086 -862 13146 -856
rect 15122 -862 15182 -856
rect 10030 -908 10090 -902
rect 14104 -908 14164 -902
rect 18110 -908 18170 -902
rect 10090 -968 14104 -908
rect 14164 -968 18110 -908
rect 10030 -974 10090 -968
rect 14104 -974 14164 -968
rect 18110 -974 18170 -968
rect 19488 -986 19548 -980
rect 20624 -986 20684 -980
rect 24694 -986 24754 -980
rect 34874 -986 34934 -980
rect 40094 -986 40154 -980
rect 19548 -1046 20624 -986
rect 20684 -1046 24694 -986
rect 24754 -1046 34874 -986
rect 34934 -1046 40094 -986
rect 19488 -1052 19548 -1046
rect 20624 -1052 20684 -1046
rect 24694 -1052 24754 -1046
rect 34874 -1052 34934 -1046
rect 40094 -1052 40154 -1046
rect 142 -1092 202 -1086
rect 532 -1092 592 -1086
rect 1048 -1092 1108 -1086
rect 3112 -1092 3172 -1086
rect 3626 -1092 3686 -1086
rect 3998 -1092 4058 -1086
rect 202 -1152 532 -1092
rect 592 -1152 1048 -1092
rect 1108 -1152 3112 -1092
rect 3172 -1152 3626 -1092
rect 3686 -1152 3998 -1092
rect 142 -1158 202 -1152
rect 532 -1158 592 -1152
rect 1048 -1158 1108 -1152
rect 3112 -1158 3172 -1152
rect 3626 -1158 3686 -1152
rect 3998 -1158 4058 -1152
rect 21136 -1094 21196 -1088
rect 29280 -1094 29340 -1088
rect 21196 -1154 22150 -1094
rect 22210 -1154 23172 -1094
rect 23232 -1154 24186 -1094
rect 24246 -1154 25212 -1094
rect 25272 -1154 26224 -1094
rect 26284 -1154 27260 -1094
rect 27320 -1154 28266 -1094
rect 28326 -1154 29280 -1094
rect 29340 -1154 30296 -1094
rect 30356 -1154 31304 -1094
rect 31364 -1154 32320 -1094
rect 32380 -1154 33344 -1094
rect 33404 -1154 34366 -1094
rect 34426 -1154 35388 -1094
rect 35448 -1154 36406 -1094
rect 36466 -1154 37420 -1094
rect 37480 -1154 38444 -1094
rect 38504 -1154 38510 -1094
rect 21136 -1160 21196 -1154
rect 29280 -1160 29340 -1154
rect -2 -1218 58 -1212
rect 1560 -1218 1620 -1212
rect 2082 -1218 2142 -1212
rect 2596 -1218 2656 -1212
rect 4134 -1218 4194 -1212
rect 58 -1278 1560 -1218
rect 1620 -1278 2082 -1218
rect 2142 -1278 2596 -1218
rect 2656 -1278 4134 -1218
rect -2 -1284 58 -1278
rect 1560 -1284 1620 -1278
rect 2082 -1284 2142 -1278
rect 2596 -1284 2656 -1278
rect 4134 -1284 4194 -1278
rect 204 -1402 3996 -1352
rect 204 -1506 258 -1402
rect 3950 -1506 3996 -1402
rect 204 -1550 3996 -1506
rect 8922 -1396 41008 -1350
rect 8922 -1550 8968 -1396
rect 40968 -1550 41008 -1396
rect 8922 -1596 41008 -1550
rect -96 -1636 504 -1626
rect -96 -1946 504 -1936
rect 3696 -1636 4296 -1626
rect 3696 -1946 4296 -1936
rect 4824 -1736 5424 -1726
rect 4824 -2046 5424 -2036
rect 41256 -1736 41856 -1726
rect 41256 -2046 41856 -2036
<< via2 >>
rect 17524 28996 18124 29296
rect 41156 28996 41756 29296
rect 21101 28700 37886 28914
rect 3410 14410 14174 14702
rect 14174 14410 14262 14702
rect 19359 14041 19449 14131
rect 1875 11995 1965 12085
rect 1579 9589 1671 9681
rect 919 9285 1021 9387
rect 1291 4587 1385 4681
rect 1642 4262 1746 4366
rect 4704 1198 4962 12790
rect 5248 12684 5348 12784
rect -156 896 4924 986
rect 1033 549 1123 639
rect 5112 -300 5172 -240
rect 3607 -358 3697 -341
rect 3607 -418 3626 -358
rect 3626 -418 3686 -358
rect 3686 -418 3697 -358
rect 3607 -431 3697 -418
rect 258 -1506 3950 -1402
rect 8968 -1550 40968 -1396
rect -96 -1936 504 -1636
rect 3696 -1936 4296 -1636
rect 4824 -2036 5424 -1736
rect 41256 -2036 41856 -1736
<< metal3 >>
rect 17514 29296 18134 29301
rect 17514 28996 17524 29296
rect 18124 28996 18134 29296
rect 17514 28991 18134 28996
rect 41146 29296 41766 29301
rect 41146 28996 41156 29296
rect 41756 28996 41766 29296
rect 41146 28991 41766 28996
rect 21038 28914 37918 28946
rect 21038 28700 21101 28914
rect 37886 28700 37918 28914
rect 21038 28680 37918 28700
rect 21038 28678 25392 28680
rect 1872 28020 16912 28166
rect 1872 28010 16066 28020
rect 1872 27320 2024 28010
rect 2720 27322 16066 28010
rect 16756 27322 16912 28020
rect 2720 27320 16912 27322
rect 1872 26990 16912 27320
rect 1872 14328 3054 26990
rect 3342 15790 15248 26730
rect 15612 15790 16912 26990
rect 3342 14702 16912 15790
rect 14262 14410 16912 14702
rect 14174 14328 16912 14410
rect 1872 14102 16912 14328
rect 19355 14136 19453 14141
rect 19354 14135 19454 14136
rect 1872 14002 15414 14102
rect 19354 14037 19355 14135
rect 19453 14037 19454 14135
rect 19354 14036 19454 14037
rect 19355 14031 19453 14036
rect 1872 13320 2026 14002
rect 2360 13320 15414 14002
rect 1872 13164 15414 13320
rect 1872 12944 5056 13164
rect -1766 12834 5056 12944
rect -1766 12368 -1732 12834
rect -1668 12368 4533 12834
rect 4597 12790 5056 12834
rect 4597 12368 4704 12790
rect -1766 12340 4704 12368
rect -1766 12172 -1052 12340
rect -1766 9628 -1736 12172
rect -1672 11834 -1052 12172
rect 3922 12172 4704 12340
rect 1870 12085 1970 12090
rect -841 12038 -743 12043
rect 1627 12038 1725 12043
rect -844 12037 1726 12038
rect -844 11939 -841 12037
rect -743 11939 1627 12037
rect 1725 11939 1726 12037
rect -844 11938 1726 11939
rect 1870 11995 1875 12085
rect 1965 11995 1970 12085
rect -841 11933 -743 11938
rect 1627 11933 1725 11938
rect 1870 11834 1970 11995
rect -1672 9691 1166 11834
rect -1672 9634 523 9691
rect -1672 9628 -1052 9634
rect -1766 9322 -1052 9628
rect 517 9581 523 9634
rect 633 9634 1166 9691
rect 1476 9681 3676 11834
rect 1476 9634 1579 9681
rect 633 9581 639 9634
rect 1574 9589 1579 9634
rect 1671 9634 3676 9681
rect 1671 9589 1676 9634
rect 3922 9628 4537 12172
rect 4601 9628 4704 12172
rect 3922 9600 4704 9628
rect 1574 9584 1676 9589
rect 522 9580 634 9581
rect 914 9387 1026 9392
rect 2088 9387 2200 9388
rect 914 9334 919 9387
rect -1766 7178 -1736 9322
rect -1672 7178 -1052 9322
rect -1766 6828 -1052 7178
rect -1766 4684 -1736 6828
rect -1672 4684 -1052 6828
rect -1766 4378 -1052 4684
rect -804 9285 919 9334
rect 1021 9336 1026 9387
rect 1021 9334 1298 9336
rect 2083 9334 2089 9387
rect 1021 9285 1396 9334
rect -804 4681 1396 9285
rect -804 4634 1291 4681
rect 1286 4587 1291 4634
rect 1385 4634 1396 4681
rect 1734 9277 2089 9334
rect 2199 9334 2205 9387
rect 3928 9350 4704 9600
rect 3922 9334 4704 9350
rect 2199 9322 4704 9334
rect 2199 9277 4537 9322
rect 1734 7178 4537 9277
rect 4601 7178 4704 9322
rect 1734 6828 4704 7178
rect 1734 4684 4537 6828
rect 4601 4684 4704 6828
rect 1734 4665 4704 4684
rect 1734 4634 2113 4665
rect 1385 4587 1390 4634
rect 1286 4582 1390 4587
rect 2107 4575 2113 4634
rect 2203 4634 4704 4665
rect 2203 4575 2209 4634
rect 2112 4574 2204 4575
rect -1766 1834 -1736 4378
rect -1672 4336 -1052 4378
rect -1672 4334 -478 4336
rect 834 4334 840 4380
rect -1672 4288 840 4334
rect 932 4334 938 4380
rect 3922 4378 4704 4634
rect 1637 4366 1751 4371
rect 1637 4334 1642 4366
rect 932 4288 1156 4334
rect -1672 2134 1156 4288
rect 1478 4262 1642 4334
rect 1746 4334 1751 4366
rect 1746 4262 3678 4334
rect 1478 2134 3678 4262
rect -1672 1834 -1052 2134
rect 1291 2030 1389 2035
rect 1290 2029 1796 2030
rect 1290 1931 1291 2029
rect 1389 1931 1697 2029
rect 1795 1931 1801 2029
rect 1290 1930 1796 1931
rect 1291 1925 1389 1930
rect -1766 1726 -1052 1834
rect 3922 1834 4537 4378
rect 4601 1834 4704 4378
rect 3922 1726 4704 1834
rect -1766 1698 4704 1726
rect -1766 1232 -1732 1698
rect -1668 1232 4533 1698
rect 4597 1232 4704 1698
rect -1766 1198 4704 1232
rect 4962 1198 5056 12790
rect 5243 12784 5353 12789
rect 5243 12779 5248 12784
rect 5348 12779 5353 12784
rect 5243 12673 5353 12679
rect -1766 1126 5056 1198
rect -242 1124 5056 1126
rect -242 986 5054 1124
rect -242 896 -156 986
rect 4924 896 5054 986
rect -242 818 5054 896
rect 1291 644 1389 649
rect 1028 643 1390 644
rect 1028 639 1291 643
rect 1028 549 1033 639
rect 1123 549 1291 639
rect 1028 545 1291 549
rect 1389 545 1390 643
rect 1028 544 1390 545
rect 1291 539 1389 544
rect 5247 -220 5345 -215
rect 5094 -221 5346 -220
rect 5094 -240 5247 -221
rect 5094 -300 5112 -240
rect 5172 -300 5247 -240
rect 5094 -319 5247 -300
rect 5345 -319 5346 -221
rect 5094 -320 5346 -319
rect 5247 -325 5345 -320
rect 4043 -336 4141 -331
rect 3602 -337 4142 -336
rect 3602 -341 4043 -337
rect 3602 -431 3607 -341
rect 3697 -431 4043 -341
rect 3602 -435 4043 -431
rect 4141 -435 4142 -337
rect 3602 -436 4142 -435
rect 4043 -441 4141 -436
rect 204 -1402 3996 -1352
rect 204 -1506 258 -1402
rect 3950 -1506 3996 -1402
rect 204 -1550 3996 -1506
rect 8922 -1396 41008 -1350
rect 8922 -1550 8968 -1396
rect 40968 -1550 41008 -1396
rect 8922 -1596 41008 -1550
rect -106 -1636 514 -1631
rect -106 -1936 -96 -1636
rect 504 -1936 514 -1636
rect -106 -1941 514 -1936
rect 3686 -1636 4306 -1631
rect 3686 -1936 3696 -1636
rect 4296 -1936 4306 -1636
rect 3686 -1941 4306 -1936
rect 4814 -1736 5434 -1731
rect 4814 -2036 4824 -1736
rect 5424 -2036 5434 -1736
rect 4814 -2041 5434 -2036
rect 41246 -1736 41866 -1731
rect 41246 -2036 41256 -1736
rect 41856 -2036 41866 -1736
rect 41246 -2041 41866 -2036
<< via3 >>
rect 17524 28996 18124 29296
rect 41156 28996 41756 29296
rect 21101 28700 37886 28914
rect 2024 27320 2720 28010
rect 16066 27322 16756 28020
rect 3054 26730 15612 26990
rect 3054 14702 3342 26730
rect 15248 15790 15612 26730
rect 3054 14410 3410 14702
rect 3410 14410 14174 14702
rect 3054 14328 14174 14410
rect 19355 14131 19453 14135
rect 19355 14041 19359 14131
rect 19359 14041 19449 14131
rect 19449 14041 19453 14131
rect 19355 14037 19453 14041
rect 2026 13320 2360 14002
rect -1732 12368 -1668 12834
rect 4533 12368 4597 12834
rect -1736 9628 -1672 12172
rect -841 11939 -743 12037
rect 1627 11939 1725 12037
rect 523 9581 633 9691
rect 4537 9628 4601 12172
rect -1736 7178 -1672 9322
rect -1736 4684 -1672 6828
rect 2089 9277 2199 9387
rect 4537 7178 4601 9322
rect 4537 4684 4601 6828
rect 2113 4575 2203 4665
rect -1736 1834 -1672 4378
rect 840 4288 932 4380
rect 1291 1931 1389 2029
rect 1697 1931 1795 2029
rect 4537 1834 4601 4378
rect -1732 1232 -1668 1698
rect 4533 1232 4597 1698
rect 5243 12684 5248 12779
rect 5248 12684 5348 12779
rect 5348 12684 5353 12779
rect 5243 12679 5353 12684
rect 1291 545 1389 643
rect 5247 -319 5345 -221
rect 4043 -435 4141 -337
rect 258 -1506 3950 -1402
rect 8968 -1550 40968 -1396
rect -96 -1936 504 -1636
rect 3696 -1936 4296 -1636
rect 4824 -2036 5424 -1736
rect 41256 -2036 41856 -1736
<< mimcap >>
rect 3058 28016 9258 28066
rect 3058 27716 8908 28016
rect 9208 27716 9258 28016
rect 3058 27666 9258 27716
rect 9458 28016 15658 28066
rect 9458 27716 15308 28016
rect 15608 27716 15658 28016
rect 9458 27666 15658 27716
rect 1972 26934 2772 26984
rect 1972 21234 2422 26934
rect 2722 21234 2772 26934
rect 16016 26934 16816 26984
rect 3912 26016 9112 26066
rect 3912 21316 8762 26016
rect 9062 21316 9112 26016
rect 3912 21266 9112 21316
rect 9512 26016 14712 26066
rect 9512 21316 14362 26016
rect 14662 21316 14712 26016
rect 9512 21266 14712 21316
rect 1972 21184 2772 21234
rect 16016 21234 16466 26934
rect 16766 21234 16816 26934
rect 16016 21184 16816 21234
rect 1972 20442 2772 20492
rect 1972 14742 2422 20442
rect 2722 14742 2772 20442
rect 3912 20416 9112 20466
rect 3912 15716 8762 20416
rect 9062 15716 9112 20416
rect 3912 15666 9112 15716
rect 9512 20416 14712 20466
rect 9512 15716 14362 20416
rect 14662 15716 14712 20416
rect 9512 15666 14712 15716
rect 16016 20442 16816 20492
rect 1972 14692 2772 14742
rect 16016 14742 16466 20442
rect 16766 14742 16816 20442
rect 16016 14692 16816 14742
rect 2558 14016 8758 14066
rect 2558 13716 8408 14016
rect 8708 13716 8758 14016
rect 2558 13666 8758 13716
rect 8958 14016 15158 14066
rect 8958 13716 14808 14016
rect 15108 13716 15158 14016
rect 8958 13666 15158 13716
rect -1553 12800 1247 12840
rect -1553 12480 -1513 12800
rect 1207 12480 1247 12800
rect -1553 12440 1247 12480
rect 1618 12800 4418 12840
rect 1618 12480 1658 12800
rect 4378 12480 4418 12800
rect 1618 12440 4418 12480
rect -1557 12060 -1157 12100
rect -1557 9740 -1517 12060
rect -1197 9740 -1157 12060
rect 4022 12060 4422 12100
rect -1557 9700 -1157 9740
rect -934 11694 1066 11734
rect -934 9774 -894 11694
rect 1026 9774 1066 11694
rect -934 9734 1066 9774
rect 1576 11694 3576 11734
rect 1576 9774 1616 11694
rect 3536 9774 3576 11694
rect 1576 9734 3576 9774
rect 4022 9740 4062 12060
rect 4382 9740 4422 12060
rect 4022 9700 4422 9740
rect -1557 9210 -1157 9250
rect -1557 7290 -1517 9210
rect -1197 7290 -1157 9210
rect -1557 7250 -1157 7290
rect -704 9194 1296 9234
rect -704 7274 -664 9194
rect 1256 7274 1296 9194
rect -704 7234 1296 7274
rect 1834 9194 3834 9234
rect 1834 7274 1874 9194
rect 3794 7274 3834 9194
rect 1834 7234 3834 7274
rect 4022 9210 4422 9250
rect 4022 7290 4062 9210
rect 4382 7290 4422 9210
rect 4022 7250 4422 7290
rect -1557 6716 -1157 6756
rect -1557 4796 -1517 6716
rect -1197 4796 -1157 6716
rect -1557 4756 -1157 4796
rect -704 6694 1296 6734
rect -704 4774 -664 6694
rect 1256 4774 1296 6694
rect -704 4734 1296 4774
rect 1834 6694 3834 6734
rect 1834 4774 1874 6694
rect 3794 4774 3834 6694
rect 1834 4734 3834 4774
rect 4022 6716 4422 6756
rect 4022 4796 4062 6716
rect 4382 4796 4422 6716
rect 4022 4756 4422 4796
rect -1557 4266 -1157 4306
rect -1557 1946 -1517 4266
rect -1197 1946 -1157 4266
rect 4022 4266 4422 4306
rect -944 4194 1056 4234
rect -944 2274 -904 4194
rect 1016 2274 1056 4194
rect -944 2234 1056 2274
rect 1578 4194 3578 4234
rect 1578 2274 1618 4194
rect 3538 2274 3578 4194
rect 1578 2234 3578 2274
rect -1557 1906 -1157 1946
rect 4022 1946 4062 4266
rect 4382 1946 4422 4266
rect 4022 1906 4422 1946
rect -1553 1586 1247 1626
rect -1553 1266 -1513 1586
rect 1207 1266 1247 1586
rect -1553 1226 1247 1266
rect 1618 1586 4418 1626
rect 1618 1266 1658 1586
rect 4378 1266 4418 1586
rect 1618 1226 4418 1266
<< mimcapcontact >>
rect 8908 27716 9208 28016
rect 15308 27716 15608 28016
rect 2422 21234 2722 26934
rect 8762 21316 9062 26016
rect 14362 21316 14662 26016
rect 16466 21234 16766 26934
rect 2422 14742 2722 20442
rect 8762 15716 9062 20416
rect 14362 15716 14662 20416
rect 16466 14742 16766 20442
rect 8408 13716 8708 14016
rect 14808 13716 15108 14016
rect -1513 12480 1207 12800
rect 1658 12480 4378 12800
rect -1517 9740 -1197 12060
rect -894 9774 1026 11694
rect 1616 9774 3536 11694
rect 4062 9740 4382 12060
rect -1517 7290 -1197 9210
rect -664 7274 1256 9194
rect 1874 7274 3794 9194
rect 4062 7290 4382 9210
rect -1517 4796 -1197 6716
rect -664 4774 1256 6694
rect 1874 4774 3794 6694
rect 4062 4796 4382 6716
rect -1517 1946 -1197 4266
rect -904 2274 1016 4194
rect 1618 2274 3538 4194
rect 4062 1946 4382 4266
rect -1513 1266 1207 1586
rect 1658 1266 4378 1586
<< metal4 >>
rect 1872 29296 42040 29480
rect 1872 28996 17524 29296
rect 18124 28996 41156 29296
rect 41756 28996 42040 29296
rect 1872 28914 42040 28996
rect 1872 28700 21101 28914
rect 37886 28700 42040 28914
rect 1872 28680 42040 28700
rect 1872 28020 16912 28166
rect 1872 28016 16066 28020
rect 1872 28010 8908 28016
rect 1872 27320 2024 28010
rect 2720 27716 8908 28010
rect 9208 27716 15308 28016
rect 15608 27716 16066 28016
rect 2720 27322 16066 27716
rect 16756 27322 16912 28020
rect 2720 27320 16912 27322
rect 1872 26990 16912 27320
rect 1872 26934 3054 26990
rect 1872 21234 2422 26934
rect 2722 21234 3054 26934
rect 15612 26934 16912 26990
rect 1872 20442 3054 21234
rect 1872 14742 2422 20442
rect 2722 14742 3054 20442
rect 1872 14328 3054 14742
rect 3812 26016 14812 26166
rect 3812 21316 8762 26016
rect 9062 21316 14362 26016
rect 14662 21316 14812 26016
rect 3812 20416 14812 21316
rect 3812 15716 8762 20416
rect 9062 15716 14362 20416
rect 14662 15716 14812 20416
rect 3812 15264 14812 15716
rect 15612 21234 16466 26934
rect 16766 21234 16912 26934
rect 15612 20442 16912 21234
rect 15612 15644 16466 20442
rect 3812 15167 15713 15264
rect 3812 15166 14812 15167
rect 3542 14702 14318 14784
rect 14206 14328 14318 14702
rect 1872 14242 14318 14328
rect 1874 14102 14318 14242
rect 1874 14016 15318 14102
rect 1874 14002 8408 14016
rect 1874 13320 2026 14002
rect 2360 13716 8408 14002
rect 8708 13716 14808 14016
rect 15108 13716 15318 14016
rect 2360 13320 15318 13716
rect 15616 13680 15713 15167
rect 15982 14742 16466 15644
rect 16766 14742 16912 20442
rect 15982 14232 16912 14742
rect 17266 14135 19454 14136
rect 17266 14037 19355 14135
rect 19453 14037 19454 14135
rect 17266 14036 19454 14037
rect 17266 13680 17366 14036
rect 15616 13580 17366 13680
rect 1874 13164 15318 13320
rect 17174 13068 17274 13580
rect 15670 12968 17274 13068
rect -1748 12834 -1652 12874
rect -1748 12706 -1732 12834
rect -1750 12606 -1732 12706
rect -1748 12368 -1732 12606
rect -1668 12734 -1652 12834
rect 4517 12834 4613 12874
rect -1514 12800 1208 12801
rect -1668 12706 -1644 12734
rect -1514 12706 -1513 12800
rect -1668 12606 -1513 12706
rect -1668 12368 -1644 12606
rect -1514 12480 -1513 12606
rect 1207 12706 1208 12800
rect 1657 12800 4379 12801
rect 1657 12706 1658 12800
rect 1207 12606 1212 12706
rect 1654 12606 1658 12706
rect 1207 12480 1208 12606
rect -1514 12479 1208 12480
rect 1657 12480 1658 12606
rect 4378 12706 4379 12800
rect 4517 12706 4533 12834
rect 4378 12606 4533 12706
rect 4378 12480 4379 12606
rect 1657 12479 4379 12480
rect -1748 12352 -1644 12368
rect 4517 12368 4533 12606
rect 4597 12706 4613 12834
rect 15670 12784 15770 12968
rect 5246 12780 15770 12784
rect 5242 12779 15770 12780
rect 4597 12368 4620 12706
rect 5242 12679 5243 12779
rect 5353 12684 15770 12779
rect 5353 12679 5354 12684
rect 5242 12678 5354 12679
rect 4517 12352 4620 12368
rect -1744 12188 -1644 12352
rect -1752 12172 -1644 12188
rect -1752 9628 -1736 12172
rect -1672 10950 -1644 12172
rect 1238 12182 3888 12282
rect -1518 12060 -1196 12061
rect -1518 10950 -1517 12060
rect -1672 10850 -1517 10950
rect -1672 9628 -1644 10850
rect -1518 9740 -1517 10850
rect -1197 9740 -1196 12060
rect -1518 9739 -1196 9740
rect -1110 12037 -742 12038
rect -1110 11939 -841 12037
rect -743 11939 -742 12037
rect -1110 11938 -742 11939
rect -1752 9612 -1644 9628
rect -1744 9338 -1644 9612
rect -1752 9322 -1644 9338
rect -1752 7178 -1736 9322
rect -1672 8336 -1644 9322
rect -1518 9210 -1196 9211
rect -1518 8336 -1517 9210
rect -1672 8228 -1517 8336
rect -1672 7178 -1644 8228
rect -1518 7290 -1517 8228
rect -1197 7290 -1196 9210
rect -1110 9134 -1010 11938
rect -895 11694 1027 11695
rect -895 9774 -894 11694
rect 1026 11660 1027 11694
rect 1238 11660 1338 12182
rect 1626 12037 1726 12038
rect 1626 11939 1627 12037
rect 1725 11939 1726 12037
rect 1626 11695 1726 11939
rect 1026 11560 1338 11660
rect 1615 11694 3537 11695
rect 1026 9774 1027 11560
rect -895 9773 1027 9774
rect 1615 9774 1616 11694
rect 3536 9774 3537 11694
rect 1615 9773 3537 9774
rect 522 9691 2200 9692
rect 522 9581 523 9691
rect 633 9581 2200 9691
rect 522 9580 2200 9581
rect 2088 9387 2200 9580
rect 2088 9277 2089 9387
rect 2199 9277 2200 9387
rect 2088 9276 2200 9277
rect 3788 9195 3888 12182
rect 4520 12172 4620 12352
rect 4061 12060 4383 12061
rect 4061 9740 4062 12060
rect 4382 10936 4383 12060
rect 4520 10936 4537 12172
rect 4382 10828 4537 10936
rect 4382 9740 4383 10828
rect 4061 9739 4383 9740
rect 4520 9628 4537 10828
rect 4601 9628 4620 12172
rect 4520 9322 4620 9628
rect -665 9194 1257 9195
rect -665 9134 -664 9194
rect -1110 9034 -664 9134
rect -1518 7289 -1196 7290
rect -665 7274 -664 9034
rect 1256 7274 1257 9194
rect -665 7273 1257 7274
rect 1873 9194 3888 9195
rect 1873 7274 1874 9194
rect 3794 9034 3888 9194
rect 4061 9210 4383 9211
rect 3794 7274 3795 9034
rect 4061 7290 4062 9210
rect 4382 8336 4383 9210
rect 4520 8336 4537 9322
rect 4382 8228 4537 8336
rect 4382 7290 4383 8228
rect 4061 7289 4383 7290
rect 1873 7273 3795 7274
rect -1752 7162 -1644 7178
rect -1744 6844 -1644 7162
rect -1752 6828 -1644 6844
rect -1752 4684 -1736 6828
rect -1672 5836 -1644 6828
rect -1518 6716 -1196 6717
rect -1518 5836 -1517 6716
rect -1672 5728 -1517 5836
rect -1672 4684 -1644 5728
rect -1518 4796 -1517 5728
rect -1197 4796 -1196 6716
rect 246 6695 346 7273
rect 2522 6695 2622 7273
rect 4520 7178 4537 8228
rect 4601 7178 4620 9322
rect 4520 6828 4620 7178
rect 4061 6716 4383 6717
rect -665 6694 1257 6695
rect -665 4882 -664 6694
rect -1518 4795 -1196 4796
rect -1752 4668 -1644 4684
rect -1744 4394 -1644 4668
rect -1752 4378 -1644 4394
rect -1752 1834 -1736 4378
rect -1672 3236 -1644 4378
rect -1108 4782 -664 4882
rect -1518 4266 -1196 4267
rect -1518 3236 -1517 4266
rect -1672 3128 -1517 3236
rect -1672 1834 -1644 3128
rect -1518 1946 -1517 3128
rect -1197 1946 -1196 4266
rect -1518 1945 -1196 1946
rect -1108 2030 -1008 4782
rect -665 4774 -664 4782
rect 1256 4774 1257 6694
rect -665 4773 1257 4774
rect 1873 6694 3795 6695
rect 1873 4774 1874 6694
rect 3794 4886 3795 6694
rect 3794 4774 3891 4886
rect 4061 4796 4062 6716
rect 4382 5736 4383 6716
rect 4520 5736 4537 6828
rect 4382 5628 4537 5736
rect 4382 4796 4383 5628
rect 4061 4795 4383 4796
rect 1873 4773 3891 4774
rect 2112 4665 2204 4666
rect 2112 4575 2113 4665
rect 2203 4575 2204 4665
rect 839 4380 933 4381
rect 2112 4380 2204 4575
rect 839 4288 840 4380
rect 932 4288 2204 4380
rect 839 4287 933 4288
rect -905 4194 1017 4195
rect -905 2274 -904 4194
rect 1016 2414 1017 4194
rect 1617 4194 3539 4195
rect 1016 2274 1018 2414
rect -905 2273 1018 2274
rect 1617 2274 1618 4194
rect 3538 2274 3539 4194
rect 1617 2273 3539 2274
rect 890 2196 1018 2273
rect 890 2096 1590 2196
rect -1108 2029 1390 2030
rect -1108 1931 1291 2029
rect 1389 1931 1390 2029
rect -1108 1930 1390 1931
rect -1752 1818 -1644 1834
rect -1744 1714 -1644 1818
rect -1748 1698 -1644 1714
rect -1748 1232 -1732 1698
rect -1668 1478 -1644 1698
rect -1514 1586 1208 1587
rect -1514 1478 -1513 1586
rect -1668 1378 -1513 1478
rect -1668 1232 -1652 1378
rect -1514 1266 -1513 1378
rect 1207 1266 1208 1586
rect -1514 1265 1208 1266
rect -1748 1192 -1652 1232
rect 1290 643 1390 1930
rect 1490 1840 1590 2096
rect 1696 2029 1796 2273
rect 1696 1931 1697 2029
rect 1795 1931 1796 2029
rect 1696 1930 1796 1931
rect 3791 1840 3891 4773
rect 4520 4684 4537 5628
rect 4601 4684 4620 6828
rect 4520 4378 4620 4684
rect 4061 4266 4383 4267
rect 4061 1946 4062 4266
rect 4382 3236 4383 4266
rect 4520 3236 4537 4378
rect 4382 3128 4537 3236
rect 4382 1946 4383 3128
rect 4061 1945 4383 1946
rect 1490 1740 3891 1840
rect 4520 1834 4537 3128
rect 4601 1834 4620 4378
rect 1490 1140 1590 1740
rect 4520 1714 4620 1834
rect 4517 1698 4620 1714
rect 1657 1586 4379 1587
rect 1657 1266 1658 1586
rect 4378 1478 4379 1586
rect 4517 1478 4533 1698
rect 4378 1378 4533 1478
rect 4378 1266 4379 1378
rect 1657 1265 4379 1266
rect 4517 1232 4533 1378
rect 4597 1378 4620 1698
rect 4597 1232 4613 1378
rect 4517 1192 4613 1232
rect 1490 1040 4142 1140
rect 1290 545 1291 643
rect 1389 545 1390 643
rect 1290 544 1390 545
rect 4042 -337 4142 1040
rect 5246 -221 5346 12678
rect 5246 -319 5247 -221
rect 5345 -319 5346 -221
rect 5246 -320 5346 -319
rect 4042 -435 4043 -337
rect 4141 -435 4142 -337
rect 4042 -436 4142 -435
rect -280 -1396 42040 -1320
rect -280 -1402 8968 -1396
rect -280 -1506 258 -1402
rect 3950 -1506 8968 -1402
rect -280 -1550 8968 -1506
rect 40968 -1550 42040 -1396
rect -280 -1636 42040 -1550
rect -280 -1936 -96 -1636
rect 504 -1936 3696 -1636
rect 4296 -1736 42040 -1636
rect 4296 -1936 4824 -1736
rect -280 -2036 4824 -1936
rect 5424 -2036 41256 -1736
rect 41856 -2036 42040 -1736
rect -280 -2120 42040 -2036
<< via4 >>
rect 2024 27320 2720 28010
rect 16066 27322 16756 28020
rect 3054 26730 15612 26990
rect 3054 14702 3342 26730
rect 3342 26526 15248 26730
rect 3342 14702 3542 26526
rect 15156 15790 15248 26526
rect 15248 15790 15612 26730
rect 15156 15644 15612 15790
rect 3054 14328 14174 14702
rect 14174 14328 14206 14702
rect 2026 13320 2360 14002
<< mimcap2 >>
rect 3058 27616 8858 28066
rect 3058 27316 3108 27616
rect 8808 27316 8858 27616
rect 3058 27266 8858 27316
rect 9458 27616 15258 28066
rect 9458 27316 9508 27616
rect 15208 27316 15258 27616
rect 9458 27266 15258 27316
rect 1972 21134 2372 26984
rect 1972 20834 2022 21134
rect 2322 20834 2372 21134
rect 3912 21216 8712 26066
rect 3912 20916 3962 21216
rect 8662 20916 8712 21216
rect 3912 20866 8712 20916
rect 9512 21216 14312 26066
rect 9512 20916 9562 21216
rect 14262 20916 14312 21216
rect 9512 20866 14312 20916
rect 16016 21134 16416 26984
rect 1972 20784 2372 20834
rect 16016 20834 16066 21134
rect 16366 20834 16416 21134
rect 16016 20784 16416 20834
rect 1972 14642 2372 20492
rect 3912 15616 8712 20466
rect 3912 15316 3962 15616
rect 8662 15316 8712 15616
rect 3912 15266 8712 15316
rect 9512 15616 14312 20466
rect 9512 15316 9562 15616
rect 14262 15316 14312 15616
rect 9512 15266 14312 15316
rect 1972 14342 2022 14642
rect 2322 14342 2372 14642
rect 1972 14292 2372 14342
rect 16016 14642 16416 20492
rect 16016 14356 16066 14642
rect 16366 14356 16416 14642
rect 16016 14292 16416 14356
rect 2558 13616 8358 14066
rect 2558 13316 2608 13616
rect 8308 13316 8358 13616
rect 2558 13266 8358 13316
rect 8958 13616 14758 14066
rect 8958 13316 9008 13616
rect 14708 13316 14758 13616
rect 8958 13266 14758 13316
<< mimcap2contact >>
rect 3108 27316 8808 27616
rect 9508 27316 15208 27616
rect 2022 20834 2322 21134
rect 3962 20916 8662 21216
rect 9562 20916 14262 21216
rect 16066 20834 16366 21134
rect 3962 15316 8662 15616
rect 9562 15316 14262 15616
rect 2022 14342 2322 14642
rect 16066 14356 16366 14642
rect 2608 13316 8308 13616
rect 9008 13316 14708 13616
<< metal5 >>
rect 1872 28020 16912 28166
rect 1872 28010 16066 28020
rect 1872 27320 2024 28010
rect 2720 27616 16066 28010
rect 2720 27320 3108 27616
rect 1872 27316 3108 27320
rect 8808 27316 9508 27616
rect 15208 27322 16066 27616
rect 16756 27322 16912 28020
rect 15208 27316 16912 27322
rect 1872 26990 16912 27316
rect 1872 21134 3054 26990
rect 1872 20834 2022 21134
rect 2322 20834 3054 21134
rect 1872 14642 3054 20834
rect 3542 21216 15156 26526
rect 3542 20916 3962 21216
rect 8662 20916 9562 21216
rect 14262 20916 15156 21216
rect 3542 15644 15156 20916
rect 15612 21134 16912 26990
rect 15612 20834 16066 21134
rect 16366 20834 16912 21134
rect 15612 15644 16912 20834
rect 3542 15616 16912 15644
rect 3542 15316 3962 15616
rect 8662 15316 9562 15616
rect 14262 15562 16912 15616
rect 14262 15316 14314 15562
rect 3542 14702 14314 15316
rect 1872 14342 2022 14642
rect 2322 14342 3054 14642
rect 1872 14328 3054 14342
rect 14206 14328 14314 14702
rect 1872 14098 14314 14328
rect 15968 14642 16912 15562
rect 15968 14356 16066 14642
rect 16366 14356 16912 14642
rect 15968 14316 16912 14356
rect 1872 14002 15212 14098
rect 1872 13320 2026 14002
rect 2360 13616 15212 14002
rect 2360 13320 2608 13616
rect 1872 13316 2608 13320
rect 8308 13316 9008 13616
rect 14708 13316 15212 13616
rect 1872 13164 15212 13316
<< labels >>
flabel metal2 2362 -152 2380 -136 1 FreeSans 480 0 0 0 clk
port 2 n
flabel metal2 2348 -280 2366 -264 1 FreeSans 480 0 0 0 vout
port 6 n
flabel metal1 18 -178 30 -162 1 FreeSans 480 0 0 0 vin
port 1 n
flabel metal2 1848 -1132 1870 -1116 1 FreeSans 480 0 0 0 vholdm
flabel metal2 2620 -404 2638 -386 1 FreeSans 480 0 0 0 vhold
port 7 n
flabel metal4 3836 11340 3852 11354 1 FreeSans 480 0 0 0 vhold
flabel metal1 6974 124 6984 136 1 FreeSans 480 0 0 0 ibiasn
port 5 n
flabel metal4 2134 29128 2186 29174 1 FreeSans 480 0 0 0 VDD
port 3 n power bidirectional
flabel metal4 -1076 11268 -1050 11288 1 FreeSans 480 0 0 0 vholdm
flabel metal3 1324 6968 1358 6998 1 FreeSans 480 0 0 0 vout
flabel metal4 -266 -1346 -260 -1342 1 FreeSans 480 0 0 0 VSS
port 4 n ground bidirectional
flabel metal1 8962 12728 8962 12728 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias1
flabel metal1 10834 6054 10834 6054 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias2
flabel metal1 40220 5762 40244 5792 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/VSS
flabel metal1 40596 6610 40596 6610 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias3
flabel metal1 40340 6816 40340 6816 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascnm
flabel metal1 40476 2584 40476 2584 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias4
flabel metal1 19178 6978 19206 7008 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vtail_cascn
flabel metal1 19496 10320 19528 10360 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascnp
flabel metal1 20362 13182 20452 13212 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M8d
flabel metal1 19284 6718 19322 6754 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vmirror
flabel metal1 39978 8450 40014 8480 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M16d
flabel metal1 6394 3540 6422 3584 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vip
flabel metal1 17994 3544 18026 3582 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vim
flabel metal1 11838 114 11934 150 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/ibiasn
flabel metal1 16988 2840 17036 2864 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vtail_cascn
flabel metal4 6120 -1664 6146 -1642 1 FreeSans 3200 0 0 0 se_fold_casc_wide_swing_ota_0/VSS
flabel metal2 10476 5146 10524 5162 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpp
flabel metal1 7552 2912 7584 2940 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpm
flabel metal4 5336 28990 5362 29084 1 FreeSans 3200 0 0 0 se_fold_casc_wide_swing_ota_0/VDD
flabel metal4 17634 14078 17654 14098 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vo
flabel metal1 39648 16708 39654 16726 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vo
flabel metal1 24538 23530 24570 23562 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M9d
flabel metal1 19972 20072 20044 20102 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascnm
flabel metal1 22696 20080 22738 20102 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascnp
flabel metal1 21250 20042 21276 20080 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vtail_cascp
flabel metal1 20738 16034 20768 16060 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vip
flabel metal1 21746 16030 21776 16064 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vim
flabel metal2 37212 20690 37274 20718 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vmirror
flabel metal1 33250 22894 33302 22920 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/VDD
flabel metal2 27486 21852 27554 21882 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpp
flabel metal2 27710 20820 27762 20854 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpm
flabel metal2 25364 26964 25364 26964 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias1
flabel metal2 26342 26702 26372 26730 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/VDD
flabel metal1 23386 25690 23420 25712 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M7d
flabel metal2 24774 25566 24832 25602 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M13d
flabel metal2 26800 23386 26878 23420 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vtail_cascp
flabel metal1 34550 19220 34586 19248 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/VDD
flabel metal2 28906 15172 28960 15206 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M8d
flabel metal2 29330 20160 29412 20192 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias2
flabel metal2 33880 17650 33942 17680 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M16d
flabel metal2 33472 17962 33536 17994 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M13d
flabel metal1 24364 20000 24404 20034 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M7d
flabel metal2 39434 17862 39496 17894 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vmirror
flabel metal2 37548 17752 37598 17788 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpm
flabel metal2 37600 16704 37692 16736 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpp
flabel metal2 24658 19032 24658 19032 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias1
flabel metal2 24528 15446 24584 15480 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M9d
<< end >>
