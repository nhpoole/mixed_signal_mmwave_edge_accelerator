magic
tech sky130A
timestamp 1626065694
<< checkpaint >>
rect -720 -863 720 863
<< metal4 >>
rect -90 219 90 233
rect -90 101 -59 219
rect 59 101 90 219
rect -90 59 90 101
rect -90 -59 -59 59
rect 59 -59 90 59
rect -90 -101 90 -59
rect -90 -219 -59 -101
rect 59 -219 90 -101
rect -90 -233 90 -219
<< via4 >>
rect -59 101 59 219
rect -59 -59 59 59
rect -59 -219 59 -101
<< metal5 >>
rect -90 219 90 233
rect -90 101 -59 219
rect 59 101 90 219
rect -90 59 90 101
rect -90 -59 -59 59
rect 59 -59 90 59
rect -90 -101 90 -59
rect -90 -219 -59 -101
rect 59 -219 90 -101
rect -90 -233 90 -219
<< end >>
