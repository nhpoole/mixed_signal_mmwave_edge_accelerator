magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -1660 -4360 12360 3740
<< nwell >>
rect -358 582 11058 2438
<< pwell >>
rect -348 256 11048 408
rect -348 -2896 -196 256
rect 10896 -2896 11048 256
rect -348 -3048 11048 -2896
<< psubdiff >>
rect -322 349 11022 382
rect -322 315 -141 349
rect -107 315 -73 349
rect -39 315 -5 349
rect 29 315 63 349
rect 97 315 131 349
rect 165 315 199 349
rect 233 315 267 349
rect 301 315 335 349
rect 369 315 403 349
rect 437 315 471 349
rect 505 315 539 349
rect 573 315 607 349
rect 641 315 675 349
rect 709 315 743 349
rect 777 315 811 349
rect 845 315 879 349
rect 913 315 947 349
rect 981 315 1015 349
rect 1049 315 1083 349
rect 1117 315 1151 349
rect 1185 315 1219 349
rect 1253 315 1287 349
rect 1321 315 1355 349
rect 1389 315 1423 349
rect 1457 315 1491 349
rect 1525 315 1559 349
rect 1593 315 1627 349
rect 1661 315 1695 349
rect 1729 315 1763 349
rect 1797 315 1831 349
rect 1865 315 1899 349
rect 1933 315 1967 349
rect 2001 315 2035 349
rect 2069 315 2103 349
rect 2137 315 2171 349
rect 2205 315 2239 349
rect 2273 315 2307 349
rect 2341 315 2375 349
rect 2409 315 2443 349
rect 2477 315 2511 349
rect 2545 315 2579 349
rect 2613 315 2647 349
rect 2681 315 2715 349
rect 2749 315 2783 349
rect 2817 315 2851 349
rect 2885 315 2919 349
rect 2953 315 2987 349
rect 3021 315 3055 349
rect 3089 315 3123 349
rect 3157 315 3191 349
rect 3225 315 3259 349
rect 3293 315 3327 349
rect 3361 315 3395 349
rect 3429 315 3463 349
rect 3497 315 3531 349
rect 3565 315 3599 349
rect 3633 315 3667 349
rect 3701 315 3735 349
rect 3769 315 3803 349
rect 3837 315 3871 349
rect 3905 315 3939 349
rect 3973 315 4007 349
rect 4041 315 4075 349
rect 4109 315 4143 349
rect 4177 315 4211 349
rect 4245 315 4279 349
rect 4313 315 4347 349
rect 4381 315 4415 349
rect 4449 315 4483 349
rect 4517 315 4551 349
rect 4585 315 4619 349
rect 4653 315 4687 349
rect 4721 315 4755 349
rect 4789 315 4823 349
rect 4857 315 4891 349
rect 4925 315 4959 349
rect 4993 315 5027 349
rect 5061 315 5095 349
rect 5129 315 5163 349
rect 5197 315 5231 349
rect 5265 315 5299 349
rect 5333 315 5367 349
rect 5401 315 5435 349
rect 5469 315 5503 349
rect 5537 315 5571 349
rect 5605 315 5639 349
rect 5673 315 5707 349
rect 5741 315 5775 349
rect 5809 315 5843 349
rect 5877 315 5911 349
rect 5945 315 5979 349
rect 6013 315 6047 349
rect 6081 315 6115 349
rect 6149 315 6183 349
rect 6217 315 6251 349
rect 6285 315 6319 349
rect 6353 315 6387 349
rect 6421 315 6455 349
rect 6489 315 6523 349
rect 6557 315 6591 349
rect 6625 315 6659 349
rect 6693 315 6727 349
rect 6761 315 6795 349
rect 6829 315 6863 349
rect 6897 315 6931 349
rect 6965 315 6999 349
rect 7033 315 7067 349
rect 7101 315 7135 349
rect 7169 315 7203 349
rect 7237 315 7271 349
rect 7305 315 7339 349
rect 7373 315 7407 349
rect 7441 315 7475 349
rect 7509 315 7543 349
rect 7577 315 7611 349
rect 7645 315 7679 349
rect 7713 315 7747 349
rect 7781 315 7815 349
rect 7849 315 7883 349
rect 7917 315 7951 349
rect 7985 315 8019 349
rect 8053 315 8087 349
rect 8121 315 8155 349
rect 8189 315 8223 349
rect 8257 315 8291 349
rect 8325 315 8359 349
rect 8393 315 8427 349
rect 8461 315 8495 349
rect 8529 315 8563 349
rect 8597 315 8631 349
rect 8665 315 8699 349
rect 8733 315 8767 349
rect 8801 315 8835 349
rect 8869 315 8903 349
rect 8937 315 8971 349
rect 9005 315 9039 349
rect 9073 315 9107 349
rect 9141 315 9175 349
rect 9209 315 9243 349
rect 9277 315 9311 349
rect 9345 315 9379 349
rect 9413 315 9447 349
rect 9481 315 9515 349
rect 9549 315 9583 349
rect 9617 315 9651 349
rect 9685 315 9719 349
rect 9753 315 9787 349
rect 9821 315 9855 349
rect 9889 315 9923 349
rect 9957 315 9991 349
rect 10025 315 10059 349
rect 10093 315 10127 349
rect 10161 315 10195 349
rect 10229 315 10263 349
rect 10297 315 10331 349
rect 10365 315 10399 349
rect 10433 315 10467 349
rect 10501 315 10535 349
rect 10569 315 10603 349
rect 10637 315 10671 349
rect 10705 315 10739 349
rect 10773 315 10807 349
rect 10841 315 11022 349
rect -322 282 11022 315
rect -322 193 -222 282
rect -322 159 -289 193
rect -255 159 -222 193
rect -322 125 -222 159
rect -322 91 -289 125
rect -255 91 -222 125
rect -322 57 -222 91
rect -322 23 -289 57
rect -255 23 -222 57
rect -322 -11 -222 23
rect -322 -45 -289 -11
rect -255 -45 -222 -11
rect -322 -79 -222 -45
rect -322 -113 -289 -79
rect -255 -113 -222 -79
rect -322 -147 -222 -113
rect -322 -181 -289 -147
rect -255 -181 -222 -147
rect -322 -215 -222 -181
rect -322 -249 -289 -215
rect -255 -249 -222 -215
rect -322 -283 -222 -249
rect -322 -317 -289 -283
rect -255 -317 -222 -283
rect -322 -351 -222 -317
rect -322 -385 -289 -351
rect -255 -385 -222 -351
rect -322 -419 -222 -385
rect -322 -453 -289 -419
rect -255 -453 -222 -419
rect -322 -487 -222 -453
rect -322 -521 -289 -487
rect -255 -521 -222 -487
rect -322 -555 -222 -521
rect -322 -589 -289 -555
rect -255 -589 -222 -555
rect -322 -623 -222 -589
rect -322 -657 -289 -623
rect -255 -657 -222 -623
rect -322 -691 -222 -657
rect -322 -725 -289 -691
rect -255 -725 -222 -691
rect -322 -759 -222 -725
rect -322 -793 -289 -759
rect -255 -793 -222 -759
rect -322 -827 -222 -793
rect -322 -861 -289 -827
rect -255 -861 -222 -827
rect -322 -895 -222 -861
rect -322 -929 -289 -895
rect -255 -929 -222 -895
rect -322 -963 -222 -929
rect -322 -997 -289 -963
rect -255 -997 -222 -963
rect -322 -1031 -222 -997
rect -322 -1065 -289 -1031
rect -255 -1065 -222 -1031
rect -322 -1099 -222 -1065
rect -322 -1133 -289 -1099
rect -255 -1133 -222 -1099
rect -322 -1167 -222 -1133
rect -322 -1201 -289 -1167
rect -255 -1201 -222 -1167
rect -322 -1235 -222 -1201
rect -322 -1269 -289 -1235
rect -255 -1269 -222 -1235
rect -322 -1303 -222 -1269
rect -322 -1337 -289 -1303
rect -255 -1337 -222 -1303
rect -322 -1371 -222 -1337
rect -322 -1405 -289 -1371
rect -255 -1405 -222 -1371
rect -322 -1439 -222 -1405
rect -322 -1473 -289 -1439
rect -255 -1473 -222 -1439
rect -322 -1507 -222 -1473
rect -322 -1541 -289 -1507
rect -255 -1541 -222 -1507
rect -322 -1575 -222 -1541
rect -322 -1609 -289 -1575
rect -255 -1609 -222 -1575
rect -322 -1643 -222 -1609
rect -322 -1677 -289 -1643
rect -255 -1677 -222 -1643
rect -322 -1711 -222 -1677
rect -322 -1745 -289 -1711
rect -255 -1745 -222 -1711
rect -322 -1779 -222 -1745
rect -322 -1813 -289 -1779
rect -255 -1813 -222 -1779
rect -322 -1847 -222 -1813
rect -322 -1881 -289 -1847
rect -255 -1881 -222 -1847
rect -322 -1915 -222 -1881
rect -322 -1949 -289 -1915
rect -255 -1949 -222 -1915
rect -322 -1983 -222 -1949
rect -322 -2017 -289 -1983
rect -255 -2017 -222 -1983
rect -322 -2051 -222 -2017
rect -322 -2085 -289 -2051
rect -255 -2085 -222 -2051
rect -322 -2119 -222 -2085
rect -322 -2153 -289 -2119
rect -255 -2153 -222 -2119
rect -322 -2187 -222 -2153
rect -322 -2221 -289 -2187
rect -255 -2221 -222 -2187
rect -322 -2255 -222 -2221
rect -322 -2289 -289 -2255
rect -255 -2289 -222 -2255
rect -322 -2323 -222 -2289
rect -322 -2357 -289 -2323
rect -255 -2357 -222 -2323
rect -322 -2391 -222 -2357
rect -322 -2425 -289 -2391
rect -255 -2425 -222 -2391
rect -322 -2459 -222 -2425
rect -322 -2493 -289 -2459
rect -255 -2493 -222 -2459
rect -322 -2527 -222 -2493
rect -322 -2561 -289 -2527
rect -255 -2561 -222 -2527
rect -322 -2595 -222 -2561
rect -322 -2629 -289 -2595
rect -255 -2629 -222 -2595
rect -322 -2663 -222 -2629
rect -322 -2697 -289 -2663
rect -255 -2697 -222 -2663
rect -322 -2731 -222 -2697
rect -322 -2765 -289 -2731
rect -255 -2765 -222 -2731
rect -322 -2799 -222 -2765
rect -322 -2833 -289 -2799
rect -255 -2833 -222 -2799
rect -322 -2922 -222 -2833
rect 10922 193 11022 282
rect 10922 159 10955 193
rect 10989 159 11022 193
rect 10922 125 11022 159
rect 10922 91 10955 125
rect 10989 91 11022 125
rect 10922 57 11022 91
rect 10922 23 10955 57
rect 10989 23 11022 57
rect 10922 -11 11022 23
rect 10922 -45 10955 -11
rect 10989 -45 11022 -11
rect 10922 -79 11022 -45
rect 10922 -113 10955 -79
rect 10989 -113 11022 -79
rect 10922 -147 11022 -113
rect 10922 -181 10955 -147
rect 10989 -181 11022 -147
rect 10922 -215 11022 -181
rect 10922 -249 10955 -215
rect 10989 -249 11022 -215
rect 10922 -283 11022 -249
rect 10922 -317 10955 -283
rect 10989 -317 11022 -283
rect 10922 -351 11022 -317
rect 10922 -385 10955 -351
rect 10989 -385 11022 -351
rect 10922 -419 11022 -385
rect 10922 -453 10955 -419
rect 10989 -453 11022 -419
rect 10922 -487 11022 -453
rect 10922 -521 10955 -487
rect 10989 -521 11022 -487
rect 10922 -555 11022 -521
rect 10922 -589 10955 -555
rect 10989 -589 11022 -555
rect 10922 -623 11022 -589
rect 10922 -657 10955 -623
rect 10989 -657 11022 -623
rect 10922 -691 11022 -657
rect 10922 -725 10955 -691
rect 10989 -725 11022 -691
rect 10922 -759 11022 -725
rect 10922 -793 10955 -759
rect 10989 -793 11022 -759
rect 10922 -827 11022 -793
rect 10922 -861 10955 -827
rect 10989 -861 11022 -827
rect 10922 -895 11022 -861
rect 10922 -929 10955 -895
rect 10989 -929 11022 -895
rect 10922 -963 11022 -929
rect 10922 -997 10955 -963
rect 10989 -997 11022 -963
rect 10922 -1031 11022 -997
rect 10922 -1065 10955 -1031
rect 10989 -1065 11022 -1031
rect 10922 -1099 11022 -1065
rect 10922 -1133 10955 -1099
rect 10989 -1133 11022 -1099
rect 10922 -1167 11022 -1133
rect 10922 -1201 10955 -1167
rect 10989 -1201 11022 -1167
rect 10922 -1235 11022 -1201
rect 10922 -1269 10955 -1235
rect 10989 -1269 11022 -1235
rect 10922 -1303 11022 -1269
rect 10922 -1337 10955 -1303
rect 10989 -1337 11022 -1303
rect 10922 -1371 11022 -1337
rect 10922 -1405 10955 -1371
rect 10989 -1405 11022 -1371
rect 10922 -1439 11022 -1405
rect 10922 -1473 10955 -1439
rect 10989 -1473 11022 -1439
rect 10922 -1507 11022 -1473
rect 10922 -1541 10955 -1507
rect 10989 -1541 11022 -1507
rect 10922 -1575 11022 -1541
rect 10922 -1609 10955 -1575
rect 10989 -1609 11022 -1575
rect 10922 -1643 11022 -1609
rect 10922 -1677 10955 -1643
rect 10989 -1677 11022 -1643
rect 10922 -1711 11022 -1677
rect 10922 -1745 10955 -1711
rect 10989 -1745 11022 -1711
rect 10922 -1779 11022 -1745
rect 10922 -1813 10955 -1779
rect 10989 -1813 11022 -1779
rect 10922 -1847 11022 -1813
rect 10922 -1881 10955 -1847
rect 10989 -1881 11022 -1847
rect 10922 -1915 11022 -1881
rect 10922 -1949 10955 -1915
rect 10989 -1949 11022 -1915
rect 10922 -1983 11022 -1949
rect 10922 -2017 10955 -1983
rect 10989 -2017 11022 -1983
rect 10922 -2051 11022 -2017
rect 10922 -2085 10955 -2051
rect 10989 -2085 11022 -2051
rect 10922 -2119 11022 -2085
rect 10922 -2153 10955 -2119
rect 10989 -2153 11022 -2119
rect 10922 -2187 11022 -2153
rect 10922 -2221 10955 -2187
rect 10989 -2221 11022 -2187
rect 10922 -2255 11022 -2221
rect 10922 -2289 10955 -2255
rect 10989 -2289 11022 -2255
rect 10922 -2323 11022 -2289
rect 10922 -2357 10955 -2323
rect 10989 -2357 11022 -2323
rect 10922 -2391 11022 -2357
rect 10922 -2425 10955 -2391
rect 10989 -2425 11022 -2391
rect 10922 -2459 11022 -2425
rect 10922 -2493 10955 -2459
rect 10989 -2493 11022 -2459
rect 10922 -2527 11022 -2493
rect 10922 -2561 10955 -2527
rect 10989 -2561 11022 -2527
rect 10922 -2595 11022 -2561
rect 10922 -2629 10955 -2595
rect 10989 -2629 11022 -2595
rect 10922 -2663 11022 -2629
rect 10922 -2697 10955 -2663
rect 10989 -2697 11022 -2663
rect 10922 -2731 11022 -2697
rect 10922 -2765 10955 -2731
rect 10989 -2765 11022 -2731
rect 10922 -2799 11022 -2765
rect 10922 -2833 10955 -2799
rect 10989 -2833 11022 -2799
rect 10922 -2922 11022 -2833
rect -322 -2955 11022 -2922
rect -322 -2989 -141 -2955
rect -107 -2989 -73 -2955
rect -39 -2989 -5 -2955
rect 29 -2989 63 -2955
rect 97 -2989 131 -2955
rect 165 -2989 199 -2955
rect 233 -2989 267 -2955
rect 301 -2989 335 -2955
rect 369 -2989 403 -2955
rect 437 -2989 471 -2955
rect 505 -2989 539 -2955
rect 573 -2989 607 -2955
rect 641 -2989 675 -2955
rect 709 -2989 743 -2955
rect 777 -2989 811 -2955
rect 845 -2989 879 -2955
rect 913 -2989 947 -2955
rect 981 -2989 1015 -2955
rect 1049 -2989 1083 -2955
rect 1117 -2989 1151 -2955
rect 1185 -2989 1219 -2955
rect 1253 -2989 1287 -2955
rect 1321 -2989 1355 -2955
rect 1389 -2989 1423 -2955
rect 1457 -2989 1491 -2955
rect 1525 -2989 1559 -2955
rect 1593 -2989 1627 -2955
rect 1661 -2989 1695 -2955
rect 1729 -2989 1763 -2955
rect 1797 -2989 1831 -2955
rect 1865 -2989 1899 -2955
rect 1933 -2989 1967 -2955
rect 2001 -2989 2035 -2955
rect 2069 -2989 2103 -2955
rect 2137 -2989 2171 -2955
rect 2205 -2989 2239 -2955
rect 2273 -2989 2307 -2955
rect 2341 -2989 2375 -2955
rect 2409 -2989 2443 -2955
rect 2477 -2989 2511 -2955
rect 2545 -2989 2579 -2955
rect 2613 -2989 2647 -2955
rect 2681 -2989 2715 -2955
rect 2749 -2989 2783 -2955
rect 2817 -2989 2851 -2955
rect 2885 -2989 2919 -2955
rect 2953 -2989 2987 -2955
rect 3021 -2989 3055 -2955
rect 3089 -2989 3123 -2955
rect 3157 -2989 3191 -2955
rect 3225 -2989 3259 -2955
rect 3293 -2989 3327 -2955
rect 3361 -2989 3395 -2955
rect 3429 -2989 3463 -2955
rect 3497 -2989 3531 -2955
rect 3565 -2989 3599 -2955
rect 3633 -2989 3667 -2955
rect 3701 -2989 3735 -2955
rect 3769 -2989 3803 -2955
rect 3837 -2989 3871 -2955
rect 3905 -2989 3939 -2955
rect 3973 -2989 4007 -2955
rect 4041 -2989 4075 -2955
rect 4109 -2989 4143 -2955
rect 4177 -2989 4211 -2955
rect 4245 -2989 4279 -2955
rect 4313 -2989 4347 -2955
rect 4381 -2989 4415 -2955
rect 4449 -2989 4483 -2955
rect 4517 -2989 4551 -2955
rect 4585 -2989 4619 -2955
rect 4653 -2989 4687 -2955
rect 4721 -2989 4755 -2955
rect 4789 -2989 4823 -2955
rect 4857 -2989 4891 -2955
rect 4925 -2989 4959 -2955
rect 4993 -2989 5027 -2955
rect 5061 -2989 5095 -2955
rect 5129 -2989 5163 -2955
rect 5197 -2989 5231 -2955
rect 5265 -2989 5299 -2955
rect 5333 -2989 5367 -2955
rect 5401 -2989 5435 -2955
rect 5469 -2989 5503 -2955
rect 5537 -2989 5571 -2955
rect 5605 -2989 5639 -2955
rect 5673 -2989 5707 -2955
rect 5741 -2989 5775 -2955
rect 5809 -2989 5843 -2955
rect 5877 -2989 5911 -2955
rect 5945 -2989 5979 -2955
rect 6013 -2989 6047 -2955
rect 6081 -2989 6115 -2955
rect 6149 -2989 6183 -2955
rect 6217 -2989 6251 -2955
rect 6285 -2989 6319 -2955
rect 6353 -2989 6387 -2955
rect 6421 -2989 6455 -2955
rect 6489 -2989 6523 -2955
rect 6557 -2989 6591 -2955
rect 6625 -2989 6659 -2955
rect 6693 -2989 6727 -2955
rect 6761 -2989 6795 -2955
rect 6829 -2989 6863 -2955
rect 6897 -2989 6931 -2955
rect 6965 -2989 6999 -2955
rect 7033 -2989 7067 -2955
rect 7101 -2989 7135 -2955
rect 7169 -2989 7203 -2955
rect 7237 -2989 7271 -2955
rect 7305 -2989 7339 -2955
rect 7373 -2989 7407 -2955
rect 7441 -2989 7475 -2955
rect 7509 -2989 7543 -2955
rect 7577 -2989 7611 -2955
rect 7645 -2989 7679 -2955
rect 7713 -2989 7747 -2955
rect 7781 -2989 7815 -2955
rect 7849 -2989 7883 -2955
rect 7917 -2989 7951 -2955
rect 7985 -2989 8019 -2955
rect 8053 -2989 8087 -2955
rect 8121 -2989 8155 -2955
rect 8189 -2989 8223 -2955
rect 8257 -2989 8291 -2955
rect 8325 -2989 8359 -2955
rect 8393 -2989 8427 -2955
rect 8461 -2989 8495 -2955
rect 8529 -2989 8563 -2955
rect 8597 -2989 8631 -2955
rect 8665 -2989 8699 -2955
rect 8733 -2989 8767 -2955
rect 8801 -2989 8835 -2955
rect 8869 -2989 8903 -2955
rect 8937 -2989 8971 -2955
rect 9005 -2989 9039 -2955
rect 9073 -2989 9107 -2955
rect 9141 -2989 9175 -2955
rect 9209 -2989 9243 -2955
rect 9277 -2989 9311 -2955
rect 9345 -2989 9379 -2955
rect 9413 -2989 9447 -2955
rect 9481 -2989 9515 -2955
rect 9549 -2989 9583 -2955
rect 9617 -2989 9651 -2955
rect 9685 -2989 9719 -2955
rect 9753 -2989 9787 -2955
rect 9821 -2989 9855 -2955
rect 9889 -2989 9923 -2955
rect 9957 -2989 9991 -2955
rect 10025 -2989 10059 -2955
rect 10093 -2989 10127 -2955
rect 10161 -2989 10195 -2955
rect 10229 -2989 10263 -2955
rect 10297 -2989 10331 -2955
rect 10365 -2989 10399 -2955
rect 10433 -2989 10467 -2955
rect 10501 -2989 10535 -2955
rect 10569 -2989 10603 -2955
rect 10637 -2989 10671 -2955
rect 10705 -2989 10739 -2955
rect 10773 -2989 10807 -2955
rect 10841 -2989 11022 -2955
rect -322 -3022 11022 -2989
<< nsubdiff >>
rect -322 2369 11022 2402
rect -322 2335 -141 2369
rect -107 2335 -73 2369
rect -39 2335 -5 2369
rect 29 2335 63 2369
rect 97 2335 131 2369
rect 165 2335 199 2369
rect 233 2335 267 2369
rect 301 2335 335 2369
rect 369 2335 403 2369
rect 437 2335 471 2369
rect 505 2335 539 2369
rect 573 2335 607 2369
rect 641 2335 675 2369
rect 709 2335 743 2369
rect 777 2335 811 2369
rect 845 2335 879 2369
rect 913 2335 947 2369
rect 981 2335 1015 2369
rect 1049 2335 1083 2369
rect 1117 2335 1151 2369
rect 1185 2335 1219 2369
rect 1253 2335 1287 2369
rect 1321 2335 1355 2369
rect 1389 2335 1423 2369
rect 1457 2335 1491 2369
rect 1525 2335 1559 2369
rect 1593 2335 1627 2369
rect 1661 2335 1695 2369
rect 1729 2335 1763 2369
rect 1797 2335 1831 2369
rect 1865 2335 1899 2369
rect 1933 2335 1967 2369
rect 2001 2335 2035 2369
rect 2069 2335 2103 2369
rect 2137 2335 2171 2369
rect 2205 2335 2239 2369
rect 2273 2335 2307 2369
rect 2341 2335 2375 2369
rect 2409 2335 2443 2369
rect 2477 2335 2511 2369
rect 2545 2335 2579 2369
rect 2613 2335 2647 2369
rect 2681 2335 2715 2369
rect 2749 2335 2783 2369
rect 2817 2335 2851 2369
rect 2885 2335 2919 2369
rect 2953 2335 2987 2369
rect 3021 2335 3055 2369
rect 3089 2335 3123 2369
rect 3157 2335 3191 2369
rect 3225 2335 3259 2369
rect 3293 2335 3327 2369
rect 3361 2335 3395 2369
rect 3429 2335 3463 2369
rect 3497 2335 3531 2369
rect 3565 2335 3599 2369
rect 3633 2335 3667 2369
rect 3701 2335 3735 2369
rect 3769 2335 3803 2369
rect 3837 2335 3871 2369
rect 3905 2335 3939 2369
rect 3973 2335 4007 2369
rect 4041 2335 4075 2369
rect 4109 2335 4143 2369
rect 4177 2335 4211 2369
rect 4245 2335 4279 2369
rect 4313 2335 4347 2369
rect 4381 2335 4415 2369
rect 4449 2335 4483 2369
rect 4517 2335 4551 2369
rect 4585 2335 4619 2369
rect 4653 2335 4687 2369
rect 4721 2335 4755 2369
rect 4789 2335 4823 2369
rect 4857 2335 4891 2369
rect 4925 2335 4959 2369
rect 4993 2335 5027 2369
rect 5061 2335 5095 2369
rect 5129 2335 5163 2369
rect 5197 2335 5231 2369
rect 5265 2335 5299 2369
rect 5333 2335 5367 2369
rect 5401 2335 5435 2369
rect 5469 2335 5503 2369
rect 5537 2335 5571 2369
rect 5605 2335 5639 2369
rect 5673 2335 5707 2369
rect 5741 2335 5775 2369
rect 5809 2335 5843 2369
rect 5877 2335 5911 2369
rect 5945 2335 5979 2369
rect 6013 2335 6047 2369
rect 6081 2335 6115 2369
rect 6149 2335 6183 2369
rect 6217 2335 6251 2369
rect 6285 2335 6319 2369
rect 6353 2335 6387 2369
rect 6421 2335 6455 2369
rect 6489 2335 6523 2369
rect 6557 2335 6591 2369
rect 6625 2335 6659 2369
rect 6693 2335 6727 2369
rect 6761 2335 6795 2369
rect 6829 2335 6863 2369
rect 6897 2335 6931 2369
rect 6965 2335 6999 2369
rect 7033 2335 7067 2369
rect 7101 2335 7135 2369
rect 7169 2335 7203 2369
rect 7237 2335 7271 2369
rect 7305 2335 7339 2369
rect 7373 2335 7407 2369
rect 7441 2335 7475 2369
rect 7509 2335 7543 2369
rect 7577 2335 7611 2369
rect 7645 2335 7679 2369
rect 7713 2335 7747 2369
rect 7781 2335 7815 2369
rect 7849 2335 7883 2369
rect 7917 2335 7951 2369
rect 7985 2335 8019 2369
rect 8053 2335 8087 2369
rect 8121 2335 8155 2369
rect 8189 2335 8223 2369
rect 8257 2335 8291 2369
rect 8325 2335 8359 2369
rect 8393 2335 8427 2369
rect 8461 2335 8495 2369
rect 8529 2335 8563 2369
rect 8597 2335 8631 2369
rect 8665 2335 8699 2369
rect 8733 2335 8767 2369
rect 8801 2335 8835 2369
rect 8869 2335 8903 2369
rect 8937 2335 8971 2369
rect 9005 2335 9039 2369
rect 9073 2335 9107 2369
rect 9141 2335 9175 2369
rect 9209 2335 9243 2369
rect 9277 2335 9311 2369
rect 9345 2335 9379 2369
rect 9413 2335 9447 2369
rect 9481 2335 9515 2369
rect 9549 2335 9583 2369
rect 9617 2335 9651 2369
rect 9685 2335 9719 2369
rect 9753 2335 9787 2369
rect 9821 2335 9855 2369
rect 9889 2335 9923 2369
rect 9957 2335 9991 2369
rect 10025 2335 10059 2369
rect 10093 2335 10127 2369
rect 10161 2335 10195 2369
rect 10229 2335 10263 2369
rect 10297 2335 10331 2369
rect 10365 2335 10399 2369
rect 10433 2335 10467 2369
rect 10501 2335 10535 2369
rect 10569 2335 10603 2369
rect 10637 2335 10671 2369
rect 10705 2335 10739 2369
rect 10773 2335 10807 2369
rect 10841 2335 11022 2369
rect -322 2302 11022 2335
rect -322 2207 -222 2302
rect -322 2173 -289 2207
rect -255 2173 -222 2207
rect -322 2139 -222 2173
rect -322 2105 -289 2139
rect -255 2105 -222 2139
rect -322 2071 -222 2105
rect -322 2037 -289 2071
rect -255 2037 -222 2071
rect -322 2003 -222 2037
rect -322 1969 -289 2003
rect -255 1969 -222 2003
rect -322 1935 -222 1969
rect -322 1901 -289 1935
rect -255 1901 -222 1935
rect -322 1867 -222 1901
rect -322 1833 -289 1867
rect -255 1833 -222 1867
rect -322 1799 -222 1833
rect -322 1765 -289 1799
rect -255 1765 -222 1799
rect -322 1731 -222 1765
rect -322 1697 -289 1731
rect -255 1697 -222 1731
rect -322 1663 -222 1697
rect -322 1629 -289 1663
rect -255 1629 -222 1663
rect -322 1595 -222 1629
rect -322 1561 -289 1595
rect -255 1561 -222 1595
rect -322 1527 -222 1561
rect -322 1493 -289 1527
rect -255 1493 -222 1527
rect -322 1459 -222 1493
rect -322 1425 -289 1459
rect -255 1425 -222 1459
rect -322 1391 -222 1425
rect -322 1357 -289 1391
rect -255 1357 -222 1391
rect -322 1323 -222 1357
rect -322 1289 -289 1323
rect -255 1289 -222 1323
rect -322 1255 -222 1289
rect -322 1221 -289 1255
rect -255 1221 -222 1255
rect -322 1187 -222 1221
rect -322 1153 -289 1187
rect -255 1153 -222 1187
rect -322 1119 -222 1153
rect -322 1085 -289 1119
rect -255 1085 -222 1119
rect -322 1051 -222 1085
rect -322 1017 -289 1051
rect -255 1017 -222 1051
rect -322 983 -222 1017
rect -322 949 -289 983
rect -255 949 -222 983
rect -322 915 -222 949
rect -322 881 -289 915
rect -255 881 -222 915
rect -322 847 -222 881
rect -322 813 -289 847
rect -255 813 -222 847
rect -322 718 -222 813
rect 10922 2207 11022 2302
rect 10922 2173 10955 2207
rect 10989 2173 11022 2207
rect 10922 2139 11022 2173
rect 10922 2105 10955 2139
rect 10989 2105 11022 2139
rect 10922 2071 11022 2105
rect 10922 2037 10955 2071
rect 10989 2037 11022 2071
rect 10922 2003 11022 2037
rect 10922 1969 10955 2003
rect 10989 1969 11022 2003
rect 10922 1935 11022 1969
rect 10922 1901 10955 1935
rect 10989 1901 11022 1935
rect 10922 1867 11022 1901
rect 10922 1833 10955 1867
rect 10989 1833 11022 1867
rect 10922 1799 11022 1833
rect 10922 1765 10955 1799
rect 10989 1765 11022 1799
rect 10922 1731 11022 1765
rect 10922 1697 10955 1731
rect 10989 1697 11022 1731
rect 10922 1663 11022 1697
rect 10922 1629 10955 1663
rect 10989 1629 11022 1663
rect 10922 1595 11022 1629
rect 10922 1561 10955 1595
rect 10989 1561 11022 1595
rect 10922 1527 11022 1561
rect 10922 1493 10955 1527
rect 10989 1493 11022 1527
rect 10922 1459 11022 1493
rect 10922 1425 10955 1459
rect 10989 1425 11022 1459
rect 10922 1391 11022 1425
rect 10922 1357 10955 1391
rect 10989 1357 11022 1391
rect 10922 1323 11022 1357
rect 10922 1289 10955 1323
rect 10989 1289 11022 1323
rect 10922 1255 11022 1289
rect 10922 1221 10955 1255
rect 10989 1221 11022 1255
rect 10922 1187 11022 1221
rect 10922 1153 10955 1187
rect 10989 1153 11022 1187
rect 10922 1119 11022 1153
rect 10922 1085 10955 1119
rect 10989 1085 11022 1119
rect 10922 1051 11022 1085
rect 10922 1017 10955 1051
rect 10989 1017 11022 1051
rect 10922 983 11022 1017
rect 10922 949 10955 983
rect 10989 949 11022 983
rect 10922 915 11022 949
rect 10922 881 10955 915
rect 10989 881 11022 915
rect 10922 847 11022 881
rect 10922 813 10955 847
rect 10989 813 11022 847
rect 10922 718 11022 813
rect -322 685 11022 718
rect -322 651 -141 685
rect -107 651 -73 685
rect -39 651 -5 685
rect 29 651 63 685
rect 97 651 131 685
rect 165 651 199 685
rect 233 651 267 685
rect 301 651 335 685
rect 369 651 403 685
rect 437 651 471 685
rect 505 651 539 685
rect 573 651 607 685
rect 641 651 675 685
rect 709 651 743 685
rect 777 651 811 685
rect 845 651 879 685
rect 913 651 947 685
rect 981 651 1015 685
rect 1049 651 1083 685
rect 1117 651 1151 685
rect 1185 651 1219 685
rect 1253 651 1287 685
rect 1321 651 1355 685
rect 1389 651 1423 685
rect 1457 651 1491 685
rect 1525 651 1559 685
rect 1593 651 1627 685
rect 1661 651 1695 685
rect 1729 651 1763 685
rect 1797 651 1831 685
rect 1865 651 1899 685
rect 1933 651 1967 685
rect 2001 651 2035 685
rect 2069 651 2103 685
rect 2137 651 2171 685
rect 2205 651 2239 685
rect 2273 651 2307 685
rect 2341 651 2375 685
rect 2409 651 2443 685
rect 2477 651 2511 685
rect 2545 651 2579 685
rect 2613 651 2647 685
rect 2681 651 2715 685
rect 2749 651 2783 685
rect 2817 651 2851 685
rect 2885 651 2919 685
rect 2953 651 2987 685
rect 3021 651 3055 685
rect 3089 651 3123 685
rect 3157 651 3191 685
rect 3225 651 3259 685
rect 3293 651 3327 685
rect 3361 651 3395 685
rect 3429 651 3463 685
rect 3497 651 3531 685
rect 3565 651 3599 685
rect 3633 651 3667 685
rect 3701 651 3735 685
rect 3769 651 3803 685
rect 3837 651 3871 685
rect 3905 651 3939 685
rect 3973 651 4007 685
rect 4041 651 4075 685
rect 4109 651 4143 685
rect 4177 651 4211 685
rect 4245 651 4279 685
rect 4313 651 4347 685
rect 4381 651 4415 685
rect 4449 651 4483 685
rect 4517 651 4551 685
rect 4585 651 4619 685
rect 4653 651 4687 685
rect 4721 651 4755 685
rect 4789 651 4823 685
rect 4857 651 4891 685
rect 4925 651 4959 685
rect 4993 651 5027 685
rect 5061 651 5095 685
rect 5129 651 5163 685
rect 5197 651 5231 685
rect 5265 651 5299 685
rect 5333 651 5367 685
rect 5401 651 5435 685
rect 5469 651 5503 685
rect 5537 651 5571 685
rect 5605 651 5639 685
rect 5673 651 5707 685
rect 5741 651 5775 685
rect 5809 651 5843 685
rect 5877 651 5911 685
rect 5945 651 5979 685
rect 6013 651 6047 685
rect 6081 651 6115 685
rect 6149 651 6183 685
rect 6217 651 6251 685
rect 6285 651 6319 685
rect 6353 651 6387 685
rect 6421 651 6455 685
rect 6489 651 6523 685
rect 6557 651 6591 685
rect 6625 651 6659 685
rect 6693 651 6727 685
rect 6761 651 6795 685
rect 6829 651 6863 685
rect 6897 651 6931 685
rect 6965 651 6999 685
rect 7033 651 7067 685
rect 7101 651 7135 685
rect 7169 651 7203 685
rect 7237 651 7271 685
rect 7305 651 7339 685
rect 7373 651 7407 685
rect 7441 651 7475 685
rect 7509 651 7543 685
rect 7577 651 7611 685
rect 7645 651 7679 685
rect 7713 651 7747 685
rect 7781 651 7815 685
rect 7849 651 7883 685
rect 7917 651 7951 685
rect 7985 651 8019 685
rect 8053 651 8087 685
rect 8121 651 8155 685
rect 8189 651 8223 685
rect 8257 651 8291 685
rect 8325 651 8359 685
rect 8393 651 8427 685
rect 8461 651 8495 685
rect 8529 651 8563 685
rect 8597 651 8631 685
rect 8665 651 8699 685
rect 8733 651 8767 685
rect 8801 651 8835 685
rect 8869 651 8903 685
rect 8937 651 8971 685
rect 9005 651 9039 685
rect 9073 651 9107 685
rect 9141 651 9175 685
rect 9209 651 9243 685
rect 9277 651 9311 685
rect 9345 651 9379 685
rect 9413 651 9447 685
rect 9481 651 9515 685
rect 9549 651 9583 685
rect 9617 651 9651 685
rect 9685 651 9719 685
rect 9753 651 9787 685
rect 9821 651 9855 685
rect 9889 651 9923 685
rect 9957 651 9991 685
rect 10025 651 10059 685
rect 10093 651 10127 685
rect 10161 651 10195 685
rect 10229 651 10263 685
rect 10297 651 10331 685
rect 10365 651 10399 685
rect 10433 651 10467 685
rect 10501 651 10535 685
rect 10569 651 10603 685
rect 10637 651 10671 685
rect 10705 651 10739 685
rect 10773 651 10807 685
rect 10841 651 11022 685
rect -322 618 11022 651
<< psubdiffcont >>
rect -141 315 -107 349
rect -73 315 -39 349
rect -5 315 29 349
rect 63 315 97 349
rect 131 315 165 349
rect 199 315 233 349
rect 267 315 301 349
rect 335 315 369 349
rect 403 315 437 349
rect 471 315 505 349
rect 539 315 573 349
rect 607 315 641 349
rect 675 315 709 349
rect 743 315 777 349
rect 811 315 845 349
rect 879 315 913 349
rect 947 315 981 349
rect 1015 315 1049 349
rect 1083 315 1117 349
rect 1151 315 1185 349
rect 1219 315 1253 349
rect 1287 315 1321 349
rect 1355 315 1389 349
rect 1423 315 1457 349
rect 1491 315 1525 349
rect 1559 315 1593 349
rect 1627 315 1661 349
rect 1695 315 1729 349
rect 1763 315 1797 349
rect 1831 315 1865 349
rect 1899 315 1933 349
rect 1967 315 2001 349
rect 2035 315 2069 349
rect 2103 315 2137 349
rect 2171 315 2205 349
rect 2239 315 2273 349
rect 2307 315 2341 349
rect 2375 315 2409 349
rect 2443 315 2477 349
rect 2511 315 2545 349
rect 2579 315 2613 349
rect 2647 315 2681 349
rect 2715 315 2749 349
rect 2783 315 2817 349
rect 2851 315 2885 349
rect 2919 315 2953 349
rect 2987 315 3021 349
rect 3055 315 3089 349
rect 3123 315 3157 349
rect 3191 315 3225 349
rect 3259 315 3293 349
rect 3327 315 3361 349
rect 3395 315 3429 349
rect 3463 315 3497 349
rect 3531 315 3565 349
rect 3599 315 3633 349
rect 3667 315 3701 349
rect 3735 315 3769 349
rect 3803 315 3837 349
rect 3871 315 3905 349
rect 3939 315 3973 349
rect 4007 315 4041 349
rect 4075 315 4109 349
rect 4143 315 4177 349
rect 4211 315 4245 349
rect 4279 315 4313 349
rect 4347 315 4381 349
rect 4415 315 4449 349
rect 4483 315 4517 349
rect 4551 315 4585 349
rect 4619 315 4653 349
rect 4687 315 4721 349
rect 4755 315 4789 349
rect 4823 315 4857 349
rect 4891 315 4925 349
rect 4959 315 4993 349
rect 5027 315 5061 349
rect 5095 315 5129 349
rect 5163 315 5197 349
rect 5231 315 5265 349
rect 5299 315 5333 349
rect 5367 315 5401 349
rect 5435 315 5469 349
rect 5503 315 5537 349
rect 5571 315 5605 349
rect 5639 315 5673 349
rect 5707 315 5741 349
rect 5775 315 5809 349
rect 5843 315 5877 349
rect 5911 315 5945 349
rect 5979 315 6013 349
rect 6047 315 6081 349
rect 6115 315 6149 349
rect 6183 315 6217 349
rect 6251 315 6285 349
rect 6319 315 6353 349
rect 6387 315 6421 349
rect 6455 315 6489 349
rect 6523 315 6557 349
rect 6591 315 6625 349
rect 6659 315 6693 349
rect 6727 315 6761 349
rect 6795 315 6829 349
rect 6863 315 6897 349
rect 6931 315 6965 349
rect 6999 315 7033 349
rect 7067 315 7101 349
rect 7135 315 7169 349
rect 7203 315 7237 349
rect 7271 315 7305 349
rect 7339 315 7373 349
rect 7407 315 7441 349
rect 7475 315 7509 349
rect 7543 315 7577 349
rect 7611 315 7645 349
rect 7679 315 7713 349
rect 7747 315 7781 349
rect 7815 315 7849 349
rect 7883 315 7917 349
rect 7951 315 7985 349
rect 8019 315 8053 349
rect 8087 315 8121 349
rect 8155 315 8189 349
rect 8223 315 8257 349
rect 8291 315 8325 349
rect 8359 315 8393 349
rect 8427 315 8461 349
rect 8495 315 8529 349
rect 8563 315 8597 349
rect 8631 315 8665 349
rect 8699 315 8733 349
rect 8767 315 8801 349
rect 8835 315 8869 349
rect 8903 315 8937 349
rect 8971 315 9005 349
rect 9039 315 9073 349
rect 9107 315 9141 349
rect 9175 315 9209 349
rect 9243 315 9277 349
rect 9311 315 9345 349
rect 9379 315 9413 349
rect 9447 315 9481 349
rect 9515 315 9549 349
rect 9583 315 9617 349
rect 9651 315 9685 349
rect 9719 315 9753 349
rect 9787 315 9821 349
rect 9855 315 9889 349
rect 9923 315 9957 349
rect 9991 315 10025 349
rect 10059 315 10093 349
rect 10127 315 10161 349
rect 10195 315 10229 349
rect 10263 315 10297 349
rect 10331 315 10365 349
rect 10399 315 10433 349
rect 10467 315 10501 349
rect 10535 315 10569 349
rect 10603 315 10637 349
rect 10671 315 10705 349
rect 10739 315 10773 349
rect 10807 315 10841 349
rect -289 159 -255 193
rect -289 91 -255 125
rect -289 23 -255 57
rect -289 -45 -255 -11
rect -289 -113 -255 -79
rect -289 -181 -255 -147
rect -289 -249 -255 -215
rect -289 -317 -255 -283
rect -289 -385 -255 -351
rect -289 -453 -255 -419
rect -289 -521 -255 -487
rect -289 -589 -255 -555
rect -289 -657 -255 -623
rect -289 -725 -255 -691
rect -289 -793 -255 -759
rect -289 -861 -255 -827
rect -289 -929 -255 -895
rect -289 -997 -255 -963
rect -289 -1065 -255 -1031
rect -289 -1133 -255 -1099
rect -289 -1201 -255 -1167
rect -289 -1269 -255 -1235
rect -289 -1337 -255 -1303
rect -289 -1405 -255 -1371
rect -289 -1473 -255 -1439
rect -289 -1541 -255 -1507
rect -289 -1609 -255 -1575
rect -289 -1677 -255 -1643
rect -289 -1745 -255 -1711
rect -289 -1813 -255 -1779
rect -289 -1881 -255 -1847
rect -289 -1949 -255 -1915
rect -289 -2017 -255 -1983
rect -289 -2085 -255 -2051
rect -289 -2153 -255 -2119
rect -289 -2221 -255 -2187
rect -289 -2289 -255 -2255
rect -289 -2357 -255 -2323
rect -289 -2425 -255 -2391
rect -289 -2493 -255 -2459
rect -289 -2561 -255 -2527
rect -289 -2629 -255 -2595
rect -289 -2697 -255 -2663
rect -289 -2765 -255 -2731
rect -289 -2833 -255 -2799
rect 10955 159 10989 193
rect 10955 91 10989 125
rect 10955 23 10989 57
rect 10955 -45 10989 -11
rect 10955 -113 10989 -79
rect 10955 -181 10989 -147
rect 10955 -249 10989 -215
rect 10955 -317 10989 -283
rect 10955 -385 10989 -351
rect 10955 -453 10989 -419
rect 10955 -521 10989 -487
rect 10955 -589 10989 -555
rect 10955 -657 10989 -623
rect 10955 -725 10989 -691
rect 10955 -793 10989 -759
rect 10955 -861 10989 -827
rect 10955 -929 10989 -895
rect 10955 -997 10989 -963
rect 10955 -1065 10989 -1031
rect 10955 -1133 10989 -1099
rect 10955 -1201 10989 -1167
rect 10955 -1269 10989 -1235
rect 10955 -1337 10989 -1303
rect 10955 -1405 10989 -1371
rect 10955 -1473 10989 -1439
rect 10955 -1541 10989 -1507
rect 10955 -1609 10989 -1575
rect 10955 -1677 10989 -1643
rect 10955 -1745 10989 -1711
rect 10955 -1813 10989 -1779
rect 10955 -1881 10989 -1847
rect 10955 -1949 10989 -1915
rect 10955 -2017 10989 -1983
rect 10955 -2085 10989 -2051
rect 10955 -2153 10989 -2119
rect 10955 -2221 10989 -2187
rect 10955 -2289 10989 -2255
rect 10955 -2357 10989 -2323
rect 10955 -2425 10989 -2391
rect 10955 -2493 10989 -2459
rect 10955 -2561 10989 -2527
rect 10955 -2629 10989 -2595
rect 10955 -2697 10989 -2663
rect 10955 -2765 10989 -2731
rect 10955 -2833 10989 -2799
rect -141 -2989 -107 -2955
rect -73 -2989 -39 -2955
rect -5 -2989 29 -2955
rect 63 -2989 97 -2955
rect 131 -2989 165 -2955
rect 199 -2989 233 -2955
rect 267 -2989 301 -2955
rect 335 -2989 369 -2955
rect 403 -2989 437 -2955
rect 471 -2989 505 -2955
rect 539 -2989 573 -2955
rect 607 -2989 641 -2955
rect 675 -2989 709 -2955
rect 743 -2989 777 -2955
rect 811 -2989 845 -2955
rect 879 -2989 913 -2955
rect 947 -2989 981 -2955
rect 1015 -2989 1049 -2955
rect 1083 -2989 1117 -2955
rect 1151 -2989 1185 -2955
rect 1219 -2989 1253 -2955
rect 1287 -2989 1321 -2955
rect 1355 -2989 1389 -2955
rect 1423 -2989 1457 -2955
rect 1491 -2989 1525 -2955
rect 1559 -2989 1593 -2955
rect 1627 -2989 1661 -2955
rect 1695 -2989 1729 -2955
rect 1763 -2989 1797 -2955
rect 1831 -2989 1865 -2955
rect 1899 -2989 1933 -2955
rect 1967 -2989 2001 -2955
rect 2035 -2989 2069 -2955
rect 2103 -2989 2137 -2955
rect 2171 -2989 2205 -2955
rect 2239 -2989 2273 -2955
rect 2307 -2989 2341 -2955
rect 2375 -2989 2409 -2955
rect 2443 -2989 2477 -2955
rect 2511 -2989 2545 -2955
rect 2579 -2989 2613 -2955
rect 2647 -2989 2681 -2955
rect 2715 -2989 2749 -2955
rect 2783 -2989 2817 -2955
rect 2851 -2989 2885 -2955
rect 2919 -2989 2953 -2955
rect 2987 -2989 3021 -2955
rect 3055 -2989 3089 -2955
rect 3123 -2989 3157 -2955
rect 3191 -2989 3225 -2955
rect 3259 -2989 3293 -2955
rect 3327 -2989 3361 -2955
rect 3395 -2989 3429 -2955
rect 3463 -2989 3497 -2955
rect 3531 -2989 3565 -2955
rect 3599 -2989 3633 -2955
rect 3667 -2989 3701 -2955
rect 3735 -2989 3769 -2955
rect 3803 -2989 3837 -2955
rect 3871 -2989 3905 -2955
rect 3939 -2989 3973 -2955
rect 4007 -2989 4041 -2955
rect 4075 -2989 4109 -2955
rect 4143 -2989 4177 -2955
rect 4211 -2989 4245 -2955
rect 4279 -2989 4313 -2955
rect 4347 -2989 4381 -2955
rect 4415 -2989 4449 -2955
rect 4483 -2989 4517 -2955
rect 4551 -2989 4585 -2955
rect 4619 -2989 4653 -2955
rect 4687 -2989 4721 -2955
rect 4755 -2989 4789 -2955
rect 4823 -2989 4857 -2955
rect 4891 -2989 4925 -2955
rect 4959 -2989 4993 -2955
rect 5027 -2989 5061 -2955
rect 5095 -2989 5129 -2955
rect 5163 -2989 5197 -2955
rect 5231 -2989 5265 -2955
rect 5299 -2989 5333 -2955
rect 5367 -2989 5401 -2955
rect 5435 -2989 5469 -2955
rect 5503 -2989 5537 -2955
rect 5571 -2989 5605 -2955
rect 5639 -2989 5673 -2955
rect 5707 -2989 5741 -2955
rect 5775 -2989 5809 -2955
rect 5843 -2989 5877 -2955
rect 5911 -2989 5945 -2955
rect 5979 -2989 6013 -2955
rect 6047 -2989 6081 -2955
rect 6115 -2989 6149 -2955
rect 6183 -2989 6217 -2955
rect 6251 -2989 6285 -2955
rect 6319 -2989 6353 -2955
rect 6387 -2989 6421 -2955
rect 6455 -2989 6489 -2955
rect 6523 -2989 6557 -2955
rect 6591 -2989 6625 -2955
rect 6659 -2989 6693 -2955
rect 6727 -2989 6761 -2955
rect 6795 -2989 6829 -2955
rect 6863 -2989 6897 -2955
rect 6931 -2989 6965 -2955
rect 6999 -2989 7033 -2955
rect 7067 -2989 7101 -2955
rect 7135 -2989 7169 -2955
rect 7203 -2989 7237 -2955
rect 7271 -2989 7305 -2955
rect 7339 -2989 7373 -2955
rect 7407 -2989 7441 -2955
rect 7475 -2989 7509 -2955
rect 7543 -2989 7577 -2955
rect 7611 -2989 7645 -2955
rect 7679 -2989 7713 -2955
rect 7747 -2989 7781 -2955
rect 7815 -2989 7849 -2955
rect 7883 -2989 7917 -2955
rect 7951 -2989 7985 -2955
rect 8019 -2989 8053 -2955
rect 8087 -2989 8121 -2955
rect 8155 -2989 8189 -2955
rect 8223 -2989 8257 -2955
rect 8291 -2989 8325 -2955
rect 8359 -2989 8393 -2955
rect 8427 -2989 8461 -2955
rect 8495 -2989 8529 -2955
rect 8563 -2989 8597 -2955
rect 8631 -2989 8665 -2955
rect 8699 -2989 8733 -2955
rect 8767 -2989 8801 -2955
rect 8835 -2989 8869 -2955
rect 8903 -2989 8937 -2955
rect 8971 -2989 9005 -2955
rect 9039 -2989 9073 -2955
rect 9107 -2989 9141 -2955
rect 9175 -2989 9209 -2955
rect 9243 -2989 9277 -2955
rect 9311 -2989 9345 -2955
rect 9379 -2989 9413 -2955
rect 9447 -2989 9481 -2955
rect 9515 -2989 9549 -2955
rect 9583 -2989 9617 -2955
rect 9651 -2989 9685 -2955
rect 9719 -2989 9753 -2955
rect 9787 -2989 9821 -2955
rect 9855 -2989 9889 -2955
rect 9923 -2989 9957 -2955
rect 9991 -2989 10025 -2955
rect 10059 -2989 10093 -2955
rect 10127 -2989 10161 -2955
rect 10195 -2989 10229 -2955
rect 10263 -2989 10297 -2955
rect 10331 -2989 10365 -2955
rect 10399 -2989 10433 -2955
rect 10467 -2989 10501 -2955
rect 10535 -2989 10569 -2955
rect 10603 -2989 10637 -2955
rect 10671 -2989 10705 -2955
rect 10739 -2989 10773 -2955
rect 10807 -2989 10841 -2955
<< nsubdiffcont >>
rect -141 2335 -107 2369
rect -73 2335 -39 2369
rect -5 2335 29 2369
rect 63 2335 97 2369
rect 131 2335 165 2369
rect 199 2335 233 2369
rect 267 2335 301 2369
rect 335 2335 369 2369
rect 403 2335 437 2369
rect 471 2335 505 2369
rect 539 2335 573 2369
rect 607 2335 641 2369
rect 675 2335 709 2369
rect 743 2335 777 2369
rect 811 2335 845 2369
rect 879 2335 913 2369
rect 947 2335 981 2369
rect 1015 2335 1049 2369
rect 1083 2335 1117 2369
rect 1151 2335 1185 2369
rect 1219 2335 1253 2369
rect 1287 2335 1321 2369
rect 1355 2335 1389 2369
rect 1423 2335 1457 2369
rect 1491 2335 1525 2369
rect 1559 2335 1593 2369
rect 1627 2335 1661 2369
rect 1695 2335 1729 2369
rect 1763 2335 1797 2369
rect 1831 2335 1865 2369
rect 1899 2335 1933 2369
rect 1967 2335 2001 2369
rect 2035 2335 2069 2369
rect 2103 2335 2137 2369
rect 2171 2335 2205 2369
rect 2239 2335 2273 2369
rect 2307 2335 2341 2369
rect 2375 2335 2409 2369
rect 2443 2335 2477 2369
rect 2511 2335 2545 2369
rect 2579 2335 2613 2369
rect 2647 2335 2681 2369
rect 2715 2335 2749 2369
rect 2783 2335 2817 2369
rect 2851 2335 2885 2369
rect 2919 2335 2953 2369
rect 2987 2335 3021 2369
rect 3055 2335 3089 2369
rect 3123 2335 3157 2369
rect 3191 2335 3225 2369
rect 3259 2335 3293 2369
rect 3327 2335 3361 2369
rect 3395 2335 3429 2369
rect 3463 2335 3497 2369
rect 3531 2335 3565 2369
rect 3599 2335 3633 2369
rect 3667 2335 3701 2369
rect 3735 2335 3769 2369
rect 3803 2335 3837 2369
rect 3871 2335 3905 2369
rect 3939 2335 3973 2369
rect 4007 2335 4041 2369
rect 4075 2335 4109 2369
rect 4143 2335 4177 2369
rect 4211 2335 4245 2369
rect 4279 2335 4313 2369
rect 4347 2335 4381 2369
rect 4415 2335 4449 2369
rect 4483 2335 4517 2369
rect 4551 2335 4585 2369
rect 4619 2335 4653 2369
rect 4687 2335 4721 2369
rect 4755 2335 4789 2369
rect 4823 2335 4857 2369
rect 4891 2335 4925 2369
rect 4959 2335 4993 2369
rect 5027 2335 5061 2369
rect 5095 2335 5129 2369
rect 5163 2335 5197 2369
rect 5231 2335 5265 2369
rect 5299 2335 5333 2369
rect 5367 2335 5401 2369
rect 5435 2335 5469 2369
rect 5503 2335 5537 2369
rect 5571 2335 5605 2369
rect 5639 2335 5673 2369
rect 5707 2335 5741 2369
rect 5775 2335 5809 2369
rect 5843 2335 5877 2369
rect 5911 2335 5945 2369
rect 5979 2335 6013 2369
rect 6047 2335 6081 2369
rect 6115 2335 6149 2369
rect 6183 2335 6217 2369
rect 6251 2335 6285 2369
rect 6319 2335 6353 2369
rect 6387 2335 6421 2369
rect 6455 2335 6489 2369
rect 6523 2335 6557 2369
rect 6591 2335 6625 2369
rect 6659 2335 6693 2369
rect 6727 2335 6761 2369
rect 6795 2335 6829 2369
rect 6863 2335 6897 2369
rect 6931 2335 6965 2369
rect 6999 2335 7033 2369
rect 7067 2335 7101 2369
rect 7135 2335 7169 2369
rect 7203 2335 7237 2369
rect 7271 2335 7305 2369
rect 7339 2335 7373 2369
rect 7407 2335 7441 2369
rect 7475 2335 7509 2369
rect 7543 2335 7577 2369
rect 7611 2335 7645 2369
rect 7679 2335 7713 2369
rect 7747 2335 7781 2369
rect 7815 2335 7849 2369
rect 7883 2335 7917 2369
rect 7951 2335 7985 2369
rect 8019 2335 8053 2369
rect 8087 2335 8121 2369
rect 8155 2335 8189 2369
rect 8223 2335 8257 2369
rect 8291 2335 8325 2369
rect 8359 2335 8393 2369
rect 8427 2335 8461 2369
rect 8495 2335 8529 2369
rect 8563 2335 8597 2369
rect 8631 2335 8665 2369
rect 8699 2335 8733 2369
rect 8767 2335 8801 2369
rect 8835 2335 8869 2369
rect 8903 2335 8937 2369
rect 8971 2335 9005 2369
rect 9039 2335 9073 2369
rect 9107 2335 9141 2369
rect 9175 2335 9209 2369
rect 9243 2335 9277 2369
rect 9311 2335 9345 2369
rect 9379 2335 9413 2369
rect 9447 2335 9481 2369
rect 9515 2335 9549 2369
rect 9583 2335 9617 2369
rect 9651 2335 9685 2369
rect 9719 2335 9753 2369
rect 9787 2335 9821 2369
rect 9855 2335 9889 2369
rect 9923 2335 9957 2369
rect 9991 2335 10025 2369
rect 10059 2335 10093 2369
rect 10127 2335 10161 2369
rect 10195 2335 10229 2369
rect 10263 2335 10297 2369
rect 10331 2335 10365 2369
rect 10399 2335 10433 2369
rect 10467 2335 10501 2369
rect 10535 2335 10569 2369
rect 10603 2335 10637 2369
rect 10671 2335 10705 2369
rect 10739 2335 10773 2369
rect 10807 2335 10841 2369
rect -289 2173 -255 2207
rect -289 2105 -255 2139
rect -289 2037 -255 2071
rect -289 1969 -255 2003
rect -289 1901 -255 1935
rect -289 1833 -255 1867
rect -289 1765 -255 1799
rect -289 1697 -255 1731
rect -289 1629 -255 1663
rect -289 1561 -255 1595
rect -289 1493 -255 1527
rect -289 1425 -255 1459
rect -289 1357 -255 1391
rect -289 1289 -255 1323
rect -289 1221 -255 1255
rect -289 1153 -255 1187
rect -289 1085 -255 1119
rect -289 1017 -255 1051
rect -289 949 -255 983
rect -289 881 -255 915
rect -289 813 -255 847
rect 10955 2173 10989 2207
rect 10955 2105 10989 2139
rect 10955 2037 10989 2071
rect 10955 1969 10989 2003
rect 10955 1901 10989 1935
rect 10955 1833 10989 1867
rect 10955 1765 10989 1799
rect 10955 1697 10989 1731
rect 10955 1629 10989 1663
rect 10955 1561 10989 1595
rect 10955 1493 10989 1527
rect 10955 1425 10989 1459
rect 10955 1357 10989 1391
rect 10955 1289 10989 1323
rect 10955 1221 10989 1255
rect 10955 1153 10989 1187
rect 10955 1085 10989 1119
rect 10955 1017 10989 1051
rect 10955 949 10989 983
rect 10955 881 10989 915
rect 10955 813 10989 847
rect -141 651 -107 685
rect -73 651 -39 685
rect -5 651 29 685
rect 63 651 97 685
rect 131 651 165 685
rect 199 651 233 685
rect 267 651 301 685
rect 335 651 369 685
rect 403 651 437 685
rect 471 651 505 685
rect 539 651 573 685
rect 607 651 641 685
rect 675 651 709 685
rect 743 651 777 685
rect 811 651 845 685
rect 879 651 913 685
rect 947 651 981 685
rect 1015 651 1049 685
rect 1083 651 1117 685
rect 1151 651 1185 685
rect 1219 651 1253 685
rect 1287 651 1321 685
rect 1355 651 1389 685
rect 1423 651 1457 685
rect 1491 651 1525 685
rect 1559 651 1593 685
rect 1627 651 1661 685
rect 1695 651 1729 685
rect 1763 651 1797 685
rect 1831 651 1865 685
rect 1899 651 1933 685
rect 1967 651 2001 685
rect 2035 651 2069 685
rect 2103 651 2137 685
rect 2171 651 2205 685
rect 2239 651 2273 685
rect 2307 651 2341 685
rect 2375 651 2409 685
rect 2443 651 2477 685
rect 2511 651 2545 685
rect 2579 651 2613 685
rect 2647 651 2681 685
rect 2715 651 2749 685
rect 2783 651 2817 685
rect 2851 651 2885 685
rect 2919 651 2953 685
rect 2987 651 3021 685
rect 3055 651 3089 685
rect 3123 651 3157 685
rect 3191 651 3225 685
rect 3259 651 3293 685
rect 3327 651 3361 685
rect 3395 651 3429 685
rect 3463 651 3497 685
rect 3531 651 3565 685
rect 3599 651 3633 685
rect 3667 651 3701 685
rect 3735 651 3769 685
rect 3803 651 3837 685
rect 3871 651 3905 685
rect 3939 651 3973 685
rect 4007 651 4041 685
rect 4075 651 4109 685
rect 4143 651 4177 685
rect 4211 651 4245 685
rect 4279 651 4313 685
rect 4347 651 4381 685
rect 4415 651 4449 685
rect 4483 651 4517 685
rect 4551 651 4585 685
rect 4619 651 4653 685
rect 4687 651 4721 685
rect 4755 651 4789 685
rect 4823 651 4857 685
rect 4891 651 4925 685
rect 4959 651 4993 685
rect 5027 651 5061 685
rect 5095 651 5129 685
rect 5163 651 5197 685
rect 5231 651 5265 685
rect 5299 651 5333 685
rect 5367 651 5401 685
rect 5435 651 5469 685
rect 5503 651 5537 685
rect 5571 651 5605 685
rect 5639 651 5673 685
rect 5707 651 5741 685
rect 5775 651 5809 685
rect 5843 651 5877 685
rect 5911 651 5945 685
rect 5979 651 6013 685
rect 6047 651 6081 685
rect 6115 651 6149 685
rect 6183 651 6217 685
rect 6251 651 6285 685
rect 6319 651 6353 685
rect 6387 651 6421 685
rect 6455 651 6489 685
rect 6523 651 6557 685
rect 6591 651 6625 685
rect 6659 651 6693 685
rect 6727 651 6761 685
rect 6795 651 6829 685
rect 6863 651 6897 685
rect 6931 651 6965 685
rect 6999 651 7033 685
rect 7067 651 7101 685
rect 7135 651 7169 685
rect 7203 651 7237 685
rect 7271 651 7305 685
rect 7339 651 7373 685
rect 7407 651 7441 685
rect 7475 651 7509 685
rect 7543 651 7577 685
rect 7611 651 7645 685
rect 7679 651 7713 685
rect 7747 651 7781 685
rect 7815 651 7849 685
rect 7883 651 7917 685
rect 7951 651 7985 685
rect 8019 651 8053 685
rect 8087 651 8121 685
rect 8155 651 8189 685
rect 8223 651 8257 685
rect 8291 651 8325 685
rect 8359 651 8393 685
rect 8427 651 8461 685
rect 8495 651 8529 685
rect 8563 651 8597 685
rect 8631 651 8665 685
rect 8699 651 8733 685
rect 8767 651 8801 685
rect 8835 651 8869 685
rect 8903 651 8937 685
rect 8971 651 9005 685
rect 9039 651 9073 685
rect 9107 651 9141 685
rect 9175 651 9209 685
rect 9243 651 9277 685
rect 9311 651 9345 685
rect 9379 651 9413 685
rect 9447 651 9481 685
rect 9515 651 9549 685
rect 9583 651 9617 685
rect 9651 651 9685 685
rect 9719 651 9753 685
rect 9787 651 9821 685
rect 9855 651 9889 685
rect 9923 651 9957 685
rect 9991 651 10025 685
rect 10059 651 10093 685
rect 10127 651 10161 685
rect 10195 651 10229 685
rect 10263 651 10297 685
rect 10331 651 10365 685
rect 10399 651 10433 685
rect 10467 651 10501 685
rect 10535 651 10569 685
rect 10603 651 10637 685
rect 10671 651 10705 685
rect 10739 651 10773 685
rect 10807 651 10841 685
<< locali >>
rect -322 2369 11022 2402
rect -322 2335 -211 2369
rect -177 2335 -141 2369
rect -105 2335 -73 2369
rect -33 2335 -5 2369
rect 39 2335 63 2369
rect 111 2335 131 2369
rect 183 2335 199 2369
rect 255 2335 267 2369
rect 327 2335 335 2369
rect 399 2335 403 2369
rect 505 2335 509 2369
rect 573 2335 581 2369
rect 641 2335 653 2369
rect 709 2335 725 2369
rect 777 2335 797 2369
rect 845 2335 869 2369
rect 913 2335 941 2369
rect 981 2335 1013 2369
rect 1049 2335 1083 2369
rect 1119 2335 1151 2369
rect 1191 2335 1219 2369
rect 1263 2335 1287 2369
rect 1335 2335 1355 2369
rect 1407 2335 1423 2369
rect 1479 2335 1491 2369
rect 1551 2335 1559 2369
rect 1623 2335 1627 2369
rect 1729 2335 1733 2369
rect 1797 2335 1805 2369
rect 1865 2335 1877 2369
rect 1933 2335 1949 2369
rect 2001 2335 2021 2369
rect 2069 2335 2093 2369
rect 2137 2335 2165 2369
rect 2205 2335 2237 2369
rect 2273 2335 2307 2369
rect 2343 2335 2375 2369
rect 2415 2335 2443 2369
rect 2487 2335 2511 2369
rect 2559 2335 2579 2369
rect 2631 2335 2647 2369
rect 2703 2335 2715 2369
rect 2775 2335 2783 2369
rect 2847 2335 2851 2369
rect 2953 2335 2957 2369
rect 3021 2335 3029 2369
rect 3089 2335 3101 2369
rect 3157 2335 3173 2369
rect 3225 2335 3245 2369
rect 3293 2335 3317 2369
rect 3361 2335 3389 2369
rect 3429 2335 3461 2369
rect 3497 2335 3531 2369
rect 3567 2335 3599 2369
rect 3639 2335 3667 2369
rect 3711 2335 3735 2369
rect 3783 2335 3803 2369
rect 3855 2335 3871 2369
rect 3927 2335 3939 2369
rect 3999 2335 4007 2369
rect 4071 2335 4075 2369
rect 4177 2335 4181 2369
rect 4245 2335 4253 2369
rect 4313 2335 4325 2369
rect 4381 2335 4397 2369
rect 4449 2335 4469 2369
rect 4517 2335 4541 2369
rect 4585 2335 4613 2369
rect 4653 2335 4685 2369
rect 4721 2335 4755 2369
rect 4791 2335 4823 2369
rect 4863 2335 4891 2369
rect 4935 2335 4959 2369
rect 5007 2335 5027 2369
rect 5079 2335 5095 2369
rect 5151 2335 5163 2369
rect 5223 2335 5231 2369
rect 5295 2335 5299 2369
rect 5401 2335 5405 2369
rect 5469 2335 5477 2369
rect 5537 2335 5549 2369
rect 5605 2335 5621 2369
rect 5673 2335 5693 2369
rect 5741 2335 5765 2369
rect 5809 2335 5837 2369
rect 5877 2335 5909 2369
rect 5945 2335 5979 2369
rect 6015 2335 6047 2369
rect 6087 2335 6115 2369
rect 6159 2335 6183 2369
rect 6231 2335 6251 2369
rect 6303 2335 6319 2369
rect 6375 2335 6387 2369
rect 6447 2335 6455 2369
rect 6519 2335 6523 2369
rect 6625 2335 6629 2369
rect 6693 2335 6701 2369
rect 6761 2335 6773 2369
rect 6829 2335 6845 2369
rect 6897 2335 6917 2369
rect 6965 2335 6989 2369
rect 7033 2335 7061 2369
rect 7101 2335 7133 2369
rect 7169 2335 7203 2369
rect 7239 2335 7271 2369
rect 7311 2335 7339 2369
rect 7383 2335 7407 2369
rect 7455 2335 7475 2369
rect 7527 2335 7543 2369
rect 7599 2335 7611 2369
rect 7671 2335 7679 2369
rect 7743 2335 7747 2369
rect 7849 2335 7853 2369
rect 7917 2335 7925 2369
rect 7985 2335 7997 2369
rect 8053 2335 8069 2369
rect 8121 2335 8141 2369
rect 8189 2335 8213 2369
rect 8257 2335 8285 2369
rect 8325 2335 8357 2369
rect 8393 2335 8427 2369
rect 8463 2335 8495 2369
rect 8535 2335 8563 2369
rect 8607 2335 8631 2369
rect 8679 2335 8699 2369
rect 8751 2335 8767 2369
rect 8823 2335 8835 2369
rect 8895 2335 8903 2369
rect 8967 2335 8971 2369
rect 9073 2335 9077 2369
rect 9141 2335 9149 2369
rect 9209 2335 9221 2369
rect 9277 2335 9293 2369
rect 9345 2335 9365 2369
rect 9413 2335 9437 2369
rect 9481 2335 9509 2369
rect 9549 2335 9581 2369
rect 9617 2335 9651 2369
rect 9687 2335 9719 2369
rect 9759 2335 9787 2369
rect 9831 2335 9855 2369
rect 9903 2335 9923 2369
rect 9975 2335 9991 2369
rect 10047 2335 10059 2369
rect 10119 2335 10127 2369
rect 10191 2335 10195 2369
rect 10297 2335 10301 2369
rect 10365 2335 10373 2369
rect 10433 2335 10445 2369
rect 10501 2335 10517 2369
rect 10569 2335 10589 2369
rect 10637 2335 10661 2369
rect 10705 2335 10733 2369
rect 10773 2335 10805 2369
rect 10841 2335 10877 2369
rect 10911 2335 11022 2369
rect -322 2302 11022 2335
rect -322 2211 -222 2302
rect -322 2173 -289 2211
rect -255 2173 -222 2211
rect -322 2139 -222 2173
rect -322 2105 -289 2139
rect -255 2105 -222 2139
rect -322 2071 -222 2105
rect -322 2033 -289 2071
rect -255 2033 -222 2071
rect -322 2003 -222 2033
rect -322 1961 -289 2003
rect -255 1961 -222 2003
rect -322 1935 -222 1961
rect -322 1889 -289 1935
rect -255 1889 -222 1935
rect -322 1867 -222 1889
rect -322 1817 -289 1867
rect -255 1817 -222 1867
rect -322 1799 -222 1817
rect -322 1745 -289 1799
rect -255 1745 -222 1799
rect -322 1731 -222 1745
rect -322 1673 -289 1731
rect -255 1673 -222 1731
rect -322 1663 -222 1673
rect -322 1601 -289 1663
rect -255 1601 -222 1663
rect -322 1595 -222 1601
rect -322 1529 -289 1595
rect -255 1529 -222 1595
rect -322 1527 -222 1529
rect -322 1493 -289 1527
rect -255 1493 -222 1527
rect -322 1491 -222 1493
rect -322 1425 -289 1491
rect -255 1425 -222 1491
rect -322 1419 -222 1425
rect -322 1357 -289 1419
rect -255 1357 -222 1419
rect -322 1347 -222 1357
rect -322 1289 -289 1347
rect -255 1289 -222 1347
rect -322 1275 -222 1289
rect -322 1221 -289 1275
rect -255 1221 -222 1275
rect -322 1203 -222 1221
rect -322 1153 -289 1203
rect -255 1153 -222 1203
rect -322 1131 -222 1153
rect -322 1085 -289 1131
rect -255 1085 -222 1131
rect -322 1059 -222 1085
rect -322 1017 -289 1059
rect -255 1017 -222 1059
rect -322 987 -222 1017
rect -322 949 -289 987
rect -255 949 -222 987
rect -322 915 -222 949
rect -322 881 -289 915
rect -255 881 -222 915
rect -322 847 -222 881
rect -322 809 -289 847
rect -255 809 -222 847
rect -322 718 -222 809
rect 10922 2211 11022 2302
rect 10922 2173 10955 2211
rect 10989 2173 11022 2211
rect 10922 2139 11022 2173
rect 10922 2105 10955 2139
rect 10989 2105 11022 2139
rect 10922 2071 11022 2105
rect 10922 2033 10955 2071
rect 10989 2033 11022 2071
rect 10922 2003 11022 2033
rect 10922 1961 10955 2003
rect 10989 1961 11022 2003
rect 10922 1935 11022 1961
rect 10922 1889 10955 1935
rect 10989 1889 11022 1935
rect 10922 1867 11022 1889
rect 10922 1817 10955 1867
rect 10989 1817 11022 1867
rect 10922 1799 11022 1817
rect 10922 1745 10955 1799
rect 10989 1745 11022 1799
rect 10922 1731 11022 1745
rect 10922 1673 10955 1731
rect 10989 1673 11022 1731
rect 10922 1663 11022 1673
rect 10922 1601 10955 1663
rect 10989 1601 11022 1663
rect 10922 1595 11022 1601
rect 10922 1529 10955 1595
rect 10989 1529 11022 1595
rect 10922 1527 11022 1529
rect 10922 1493 10955 1527
rect 10989 1493 11022 1527
rect 10922 1491 11022 1493
rect 10922 1425 10955 1491
rect 10989 1425 11022 1491
rect 10922 1419 11022 1425
rect 10922 1357 10955 1419
rect 10989 1357 11022 1419
rect 10922 1347 11022 1357
rect 10922 1289 10955 1347
rect 10989 1289 11022 1347
rect 10922 1275 11022 1289
rect 10922 1221 10955 1275
rect 10989 1221 11022 1275
rect 10922 1203 11022 1221
rect 10922 1153 10955 1203
rect 10989 1153 11022 1203
rect 10922 1131 11022 1153
rect 10922 1085 10955 1131
rect 10989 1085 11022 1131
rect 10922 1059 11022 1085
rect 10922 1017 10955 1059
rect 10989 1017 11022 1059
rect 10922 987 11022 1017
rect 10922 949 10955 987
rect 10989 949 11022 987
rect 10922 915 11022 949
rect 10922 881 10955 915
rect 10989 881 11022 915
rect 10922 847 11022 881
rect 10922 809 10955 847
rect 10989 809 11022 847
rect 10922 718 11022 809
rect -322 685 11022 718
rect -322 651 -211 685
rect -177 651 -141 685
rect -105 651 -73 685
rect -33 651 -5 685
rect 39 651 63 685
rect 111 651 131 685
rect 183 651 199 685
rect 255 651 267 685
rect 327 651 335 685
rect 399 651 403 685
rect 505 651 509 685
rect 573 651 581 685
rect 641 651 653 685
rect 709 651 725 685
rect 777 651 797 685
rect 845 651 869 685
rect 913 651 941 685
rect 981 651 1013 685
rect 1049 651 1083 685
rect 1119 651 1151 685
rect 1191 651 1219 685
rect 1263 651 1287 685
rect 1335 651 1355 685
rect 1407 651 1423 685
rect 1479 651 1491 685
rect 1551 651 1559 685
rect 1623 651 1627 685
rect 1729 651 1733 685
rect 1797 651 1805 685
rect 1865 651 1877 685
rect 1933 651 1949 685
rect 2001 651 2021 685
rect 2069 651 2093 685
rect 2137 651 2165 685
rect 2205 651 2237 685
rect 2273 651 2307 685
rect 2343 651 2375 685
rect 2415 651 2443 685
rect 2487 651 2511 685
rect 2559 651 2579 685
rect 2631 651 2647 685
rect 2703 651 2715 685
rect 2775 651 2783 685
rect 2847 651 2851 685
rect 2953 651 2957 685
rect 3021 651 3029 685
rect 3089 651 3101 685
rect 3157 651 3173 685
rect 3225 651 3245 685
rect 3293 651 3317 685
rect 3361 651 3389 685
rect 3429 651 3461 685
rect 3497 651 3531 685
rect 3567 651 3599 685
rect 3639 651 3667 685
rect 3711 651 3735 685
rect 3783 651 3803 685
rect 3855 651 3871 685
rect 3927 651 3939 685
rect 3999 651 4007 685
rect 4071 651 4075 685
rect 4177 651 4181 685
rect 4245 651 4253 685
rect 4313 651 4325 685
rect 4381 651 4397 685
rect 4449 651 4469 685
rect 4517 651 4541 685
rect 4585 651 4613 685
rect 4653 651 4685 685
rect 4721 651 4755 685
rect 4791 651 4823 685
rect 4863 651 4891 685
rect 4935 651 4959 685
rect 5007 651 5027 685
rect 5079 651 5095 685
rect 5151 651 5163 685
rect 5223 651 5231 685
rect 5295 651 5299 685
rect 5401 651 5405 685
rect 5469 651 5477 685
rect 5537 651 5549 685
rect 5605 651 5621 685
rect 5673 651 5693 685
rect 5741 651 5765 685
rect 5809 651 5837 685
rect 5877 651 5909 685
rect 5945 651 5979 685
rect 6015 651 6047 685
rect 6087 651 6115 685
rect 6159 651 6183 685
rect 6231 651 6251 685
rect 6303 651 6319 685
rect 6375 651 6387 685
rect 6447 651 6455 685
rect 6519 651 6523 685
rect 6625 651 6629 685
rect 6693 651 6701 685
rect 6761 651 6773 685
rect 6829 651 6845 685
rect 6897 651 6917 685
rect 6965 651 6989 685
rect 7033 651 7061 685
rect 7101 651 7133 685
rect 7169 651 7203 685
rect 7239 651 7271 685
rect 7311 651 7339 685
rect 7383 651 7407 685
rect 7455 651 7475 685
rect 7527 651 7543 685
rect 7599 651 7611 685
rect 7671 651 7679 685
rect 7743 651 7747 685
rect 7849 651 7853 685
rect 7917 651 7925 685
rect 7985 651 7997 685
rect 8053 651 8069 685
rect 8121 651 8141 685
rect 8189 651 8213 685
rect 8257 651 8285 685
rect 8325 651 8357 685
rect 8393 651 8427 685
rect 8463 651 8495 685
rect 8535 651 8563 685
rect 8607 651 8631 685
rect 8679 651 8699 685
rect 8751 651 8767 685
rect 8823 651 8835 685
rect 8895 651 8903 685
rect 8967 651 8971 685
rect 9073 651 9077 685
rect 9141 651 9149 685
rect 9209 651 9221 685
rect 9277 651 9293 685
rect 9345 651 9365 685
rect 9413 651 9437 685
rect 9481 651 9509 685
rect 9549 651 9581 685
rect 9617 651 9651 685
rect 9687 651 9719 685
rect 9759 651 9787 685
rect 9831 651 9855 685
rect 9903 651 9923 685
rect 9975 651 9991 685
rect 10047 651 10059 685
rect 10119 651 10127 685
rect 10191 651 10195 685
rect 10297 651 10301 685
rect 10365 651 10373 685
rect 10433 651 10445 685
rect 10501 651 10517 685
rect 10569 651 10589 685
rect 10637 651 10661 685
rect 10705 651 10733 685
rect 10773 651 10805 685
rect 10841 651 10877 685
rect 10911 651 11022 685
rect -322 618 11022 651
rect -322 349 11022 382
rect -322 315 -211 349
rect -177 315 -141 349
rect -105 315 -73 349
rect -33 315 -5 349
rect 39 315 63 349
rect 111 315 131 349
rect 183 315 199 349
rect 255 315 267 349
rect 327 315 335 349
rect 399 315 403 349
rect 505 315 509 349
rect 573 315 581 349
rect 641 315 653 349
rect 709 315 725 349
rect 777 315 797 349
rect 845 315 869 349
rect 913 315 941 349
rect 981 315 1013 349
rect 1049 315 1083 349
rect 1119 315 1151 349
rect 1191 315 1219 349
rect 1263 315 1287 349
rect 1335 315 1355 349
rect 1407 315 1423 349
rect 1479 315 1491 349
rect 1551 315 1559 349
rect 1623 315 1627 349
rect 1729 315 1733 349
rect 1797 315 1805 349
rect 1865 315 1877 349
rect 1933 315 1949 349
rect 2001 315 2021 349
rect 2069 315 2093 349
rect 2137 315 2165 349
rect 2205 315 2237 349
rect 2273 315 2307 349
rect 2343 315 2375 349
rect 2415 315 2443 349
rect 2487 315 2511 349
rect 2559 315 2579 349
rect 2631 315 2647 349
rect 2703 315 2715 349
rect 2775 315 2783 349
rect 2847 315 2851 349
rect 2953 315 2957 349
rect 3021 315 3029 349
rect 3089 315 3101 349
rect 3157 315 3173 349
rect 3225 315 3245 349
rect 3293 315 3317 349
rect 3361 315 3389 349
rect 3429 315 3461 349
rect 3497 315 3531 349
rect 3567 315 3599 349
rect 3639 315 3667 349
rect 3711 315 3735 349
rect 3783 315 3803 349
rect 3855 315 3871 349
rect 3927 315 3939 349
rect 3999 315 4007 349
rect 4071 315 4075 349
rect 4177 315 4181 349
rect 4245 315 4253 349
rect 4313 315 4325 349
rect 4381 315 4397 349
rect 4449 315 4469 349
rect 4517 315 4541 349
rect 4585 315 4613 349
rect 4653 315 4685 349
rect 4721 315 4755 349
rect 4791 315 4823 349
rect 4863 315 4891 349
rect 4935 315 4959 349
rect 5007 315 5027 349
rect 5079 315 5095 349
rect 5151 315 5163 349
rect 5223 315 5231 349
rect 5295 315 5299 349
rect 5401 315 5405 349
rect 5469 315 5477 349
rect 5537 315 5549 349
rect 5605 315 5621 349
rect 5673 315 5693 349
rect 5741 315 5765 349
rect 5809 315 5837 349
rect 5877 315 5909 349
rect 5945 315 5979 349
rect 6015 315 6047 349
rect 6087 315 6115 349
rect 6159 315 6183 349
rect 6231 315 6251 349
rect 6303 315 6319 349
rect 6375 315 6387 349
rect 6447 315 6455 349
rect 6519 315 6523 349
rect 6625 315 6629 349
rect 6693 315 6701 349
rect 6761 315 6773 349
rect 6829 315 6845 349
rect 6897 315 6917 349
rect 6965 315 6989 349
rect 7033 315 7061 349
rect 7101 315 7133 349
rect 7169 315 7203 349
rect 7239 315 7271 349
rect 7311 315 7339 349
rect 7383 315 7407 349
rect 7455 315 7475 349
rect 7527 315 7543 349
rect 7599 315 7611 349
rect 7671 315 7679 349
rect 7743 315 7747 349
rect 7849 315 7853 349
rect 7917 315 7925 349
rect 7985 315 7997 349
rect 8053 315 8069 349
rect 8121 315 8141 349
rect 8189 315 8213 349
rect 8257 315 8285 349
rect 8325 315 8357 349
rect 8393 315 8427 349
rect 8463 315 8495 349
rect 8535 315 8563 349
rect 8607 315 8631 349
rect 8679 315 8699 349
rect 8751 315 8767 349
rect 8823 315 8835 349
rect 8895 315 8903 349
rect 8967 315 8971 349
rect 9073 315 9077 349
rect 9141 315 9149 349
rect 9209 315 9221 349
rect 9277 315 9293 349
rect 9345 315 9365 349
rect 9413 315 9437 349
rect 9481 315 9509 349
rect 9549 315 9581 349
rect 9617 315 9651 349
rect 9687 315 9719 349
rect 9759 315 9787 349
rect 9831 315 9855 349
rect 9903 315 9923 349
rect 9975 315 9991 349
rect 10047 315 10059 349
rect 10119 315 10127 349
rect 10191 315 10195 349
rect 10297 315 10301 349
rect 10365 315 10373 349
rect 10433 315 10445 349
rect 10501 315 10517 349
rect 10569 315 10589 349
rect 10637 315 10661 349
rect 10705 315 10733 349
rect 10773 315 10805 349
rect 10841 315 10877 349
rect 10911 315 11022 349
rect -322 282 11022 315
rect -322 193 -222 282
rect -322 159 -289 193
rect -255 159 -222 193
rect -322 125 -222 159
rect -322 67 -289 125
rect -255 67 -222 125
rect -322 57 -222 67
rect -322 -5 -289 57
rect -255 -5 -222 57
rect -322 -11 -222 -5
rect -322 -77 -289 -11
rect -255 -77 -222 -11
rect -322 -79 -222 -77
rect -322 -113 -289 -79
rect -255 -113 -222 -79
rect -322 -115 -222 -113
rect -322 -181 -289 -115
rect -255 -181 -222 -115
rect -322 -187 -222 -181
rect -322 -249 -289 -187
rect -255 -249 -222 -187
rect -322 -259 -222 -249
rect -322 -317 -289 -259
rect -255 -317 -222 -259
rect -322 -331 -222 -317
rect -322 -385 -289 -331
rect -255 -385 -222 -331
rect -322 -403 -222 -385
rect -322 -453 -289 -403
rect -255 -453 -222 -403
rect -322 -475 -222 -453
rect -322 -521 -289 -475
rect -255 -521 -222 -475
rect -322 -547 -222 -521
rect -322 -589 -289 -547
rect -255 -589 -222 -547
rect -322 -619 -222 -589
rect -322 -657 -289 -619
rect -255 -657 -222 -619
rect -322 -691 -222 -657
rect -322 -725 -289 -691
rect -255 -725 -222 -691
rect -322 -759 -222 -725
rect -322 -797 -289 -759
rect -255 -797 -222 -759
rect -322 -827 -222 -797
rect -322 -869 -289 -827
rect -255 -869 -222 -827
rect -322 -895 -222 -869
rect -322 -941 -289 -895
rect -255 -941 -222 -895
rect -322 -963 -222 -941
rect -322 -1013 -289 -963
rect -255 -1013 -222 -963
rect -322 -1031 -222 -1013
rect -322 -1085 -289 -1031
rect -255 -1085 -222 -1031
rect -322 -1099 -222 -1085
rect -322 -1157 -289 -1099
rect -255 -1157 -222 -1099
rect -322 -1167 -222 -1157
rect -322 -1229 -289 -1167
rect -255 -1229 -222 -1167
rect -322 -1235 -222 -1229
rect -322 -1301 -289 -1235
rect -255 -1301 -222 -1235
rect -322 -1303 -222 -1301
rect -322 -1337 -289 -1303
rect -255 -1337 -222 -1303
rect -322 -1339 -222 -1337
rect -322 -1405 -289 -1339
rect -255 -1405 -222 -1339
rect -322 -1411 -222 -1405
rect -322 -1473 -289 -1411
rect -255 -1473 -222 -1411
rect -322 -1483 -222 -1473
rect -322 -1541 -289 -1483
rect -255 -1541 -222 -1483
rect -322 -1555 -222 -1541
rect -322 -1609 -289 -1555
rect -255 -1609 -222 -1555
rect -322 -1627 -222 -1609
rect -322 -1677 -289 -1627
rect -255 -1677 -222 -1627
rect -322 -1699 -222 -1677
rect -322 -1745 -289 -1699
rect -255 -1745 -222 -1699
rect -322 -1771 -222 -1745
rect -322 -1813 -289 -1771
rect -255 -1813 -222 -1771
rect -322 -1843 -222 -1813
rect -322 -1881 -289 -1843
rect -255 -1881 -222 -1843
rect -322 -1915 -222 -1881
rect -322 -1949 -289 -1915
rect -255 -1949 -222 -1915
rect -322 -1983 -222 -1949
rect -322 -2021 -289 -1983
rect -255 -2021 -222 -1983
rect -322 -2051 -222 -2021
rect -322 -2093 -289 -2051
rect -255 -2093 -222 -2051
rect -322 -2119 -222 -2093
rect -322 -2165 -289 -2119
rect -255 -2165 -222 -2119
rect -322 -2187 -222 -2165
rect -322 -2237 -289 -2187
rect -255 -2237 -222 -2187
rect -322 -2255 -222 -2237
rect -322 -2309 -289 -2255
rect -255 -2309 -222 -2255
rect -322 -2323 -222 -2309
rect -322 -2381 -289 -2323
rect -255 -2381 -222 -2323
rect -322 -2391 -222 -2381
rect -322 -2453 -289 -2391
rect -255 -2453 -222 -2391
rect -322 -2459 -222 -2453
rect -322 -2525 -289 -2459
rect -255 -2525 -222 -2459
rect -322 -2527 -222 -2525
rect -322 -2561 -289 -2527
rect -255 -2561 -222 -2527
rect -322 -2563 -222 -2561
rect -322 -2629 -289 -2563
rect -255 -2629 -222 -2563
rect -322 -2635 -222 -2629
rect -322 -2697 -289 -2635
rect -255 -2697 -222 -2635
rect -322 -2707 -222 -2697
rect -322 -2765 -289 -2707
rect -255 -2765 -222 -2707
rect -322 -2799 -222 -2765
rect -322 -2833 -289 -2799
rect -255 -2833 -222 -2799
rect -322 -2922 -222 -2833
rect 10922 193 11022 282
rect 10922 159 10955 193
rect 10989 159 11022 193
rect 10922 125 11022 159
rect 10922 67 10955 125
rect 10989 67 11022 125
rect 10922 57 11022 67
rect 10922 -5 10955 57
rect 10989 -5 11022 57
rect 10922 -11 11022 -5
rect 10922 -77 10955 -11
rect 10989 -77 11022 -11
rect 10922 -79 11022 -77
rect 10922 -113 10955 -79
rect 10989 -113 11022 -79
rect 10922 -115 11022 -113
rect 10922 -181 10955 -115
rect 10989 -181 11022 -115
rect 10922 -187 11022 -181
rect 10922 -249 10955 -187
rect 10989 -249 11022 -187
rect 10922 -259 11022 -249
rect 10922 -317 10955 -259
rect 10989 -317 11022 -259
rect 10922 -331 11022 -317
rect 10922 -385 10955 -331
rect 10989 -385 11022 -331
rect 10922 -403 11022 -385
rect 10922 -453 10955 -403
rect 10989 -453 11022 -403
rect 10922 -475 11022 -453
rect 10922 -521 10955 -475
rect 10989 -521 11022 -475
rect 10922 -547 11022 -521
rect 10922 -589 10955 -547
rect 10989 -589 11022 -547
rect 10922 -619 11022 -589
rect 10922 -657 10955 -619
rect 10989 -657 11022 -619
rect 10922 -691 11022 -657
rect 10922 -725 10955 -691
rect 10989 -725 11022 -691
rect 10922 -759 11022 -725
rect 10922 -797 10955 -759
rect 10989 -797 11022 -759
rect 10922 -827 11022 -797
rect 10922 -869 10955 -827
rect 10989 -869 11022 -827
rect 10922 -895 11022 -869
rect 10922 -941 10955 -895
rect 10989 -941 11022 -895
rect 10922 -963 11022 -941
rect 10922 -1013 10955 -963
rect 10989 -1013 11022 -963
rect 10922 -1031 11022 -1013
rect 10922 -1085 10955 -1031
rect 10989 -1085 11022 -1031
rect 10922 -1099 11022 -1085
rect 10922 -1157 10955 -1099
rect 10989 -1157 11022 -1099
rect 10922 -1167 11022 -1157
rect 10922 -1229 10955 -1167
rect 10989 -1229 11022 -1167
rect 10922 -1235 11022 -1229
rect 10922 -1301 10955 -1235
rect 10989 -1301 11022 -1235
rect 10922 -1303 11022 -1301
rect 10922 -1337 10955 -1303
rect 10989 -1337 11022 -1303
rect 10922 -1339 11022 -1337
rect 10922 -1405 10955 -1339
rect 10989 -1405 11022 -1339
rect 10922 -1411 11022 -1405
rect 10922 -1473 10955 -1411
rect 10989 -1473 11022 -1411
rect 10922 -1483 11022 -1473
rect 10922 -1541 10955 -1483
rect 10989 -1541 11022 -1483
rect 10922 -1555 11022 -1541
rect 10922 -1609 10955 -1555
rect 10989 -1609 11022 -1555
rect 10922 -1627 11022 -1609
rect 10922 -1677 10955 -1627
rect 10989 -1677 11022 -1627
rect 10922 -1699 11022 -1677
rect 10922 -1745 10955 -1699
rect 10989 -1745 11022 -1699
rect 10922 -1771 11022 -1745
rect 10922 -1813 10955 -1771
rect 10989 -1813 11022 -1771
rect 10922 -1843 11022 -1813
rect 10922 -1881 10955 -1843
rect 10989 -1881 11022 -1843
rect 10922 -1915 11022 -1881
rect 10922 -1949 10955 -1915
rect 10989 -1949 11022 -1915
rect 10922 -1983 11022 -1949
rect 10922 -2021 10955 -1983
rect 10989 -2021 11022 -1983
rect 10922 -2051 11022 -2021
rect 10922 -2093 10955 -2051
rect 10989 -2093 11022 -2051
rect 10922 -2119 11022 -2093
rect 10922 -2165 10955 -2119
rect 10989 -2165 11022 -2119
rect 10922 -2187 11022 -2165
rect 10922 -2237 10955 -2187
rect 10989 -2237 11022 -2187
rect 10922 -2255 11022 -2237
rect 10922 -2309 10955 -2255
rect 10989 -2309 11022 -2255
rect 10922 -2323 11022 -2309
rect 10922 -2381 10955 -2323
rect 10989 -2381 11022 -2323
rect 10922 -2391 11022 -2381
rect 10922 -2453 10955 -2391
rect 10989 -2453 11022 -2391
rect 10922 -2459 11022 -2453
rect 10922 -2525 10955 -2459
rect 10989 -2525 11022 -2459
rect 10922 -2527 11022 -2525
rect 10922 -2561 10955 -2527
rect 10989 -2561 11022 -2527
rect 10922 -2563 11022 -2561
rect 10922 -2629 10955 -2563
rect 10989 -2629 11022 -2563
rect 10922 -2635 11022 -2629
rect 10922 -2697 10955 -2635
rect 10989 -2697 11022 -2635
rect 10922 -2707 11022 -2697
rect 10922 -2765 10955 -2707
rect 10989 -2765 11022 -2707
rect 10922 -2799 11022 -2765
rect 10922 -2833 10955 -2799
rect 10989 -2833 11022 -2799
rect 10922 -2922 11022 -2833
rect -322 -2955 11022 -2922
rect -322 -2989 -211 -2955
rect -177 -2989 -141 -2955
rect -105 -2989 -73 -2955
rect -33 -2989 -5 -2955
rect 39 -2989 63 -2955
rect 111 -2989 131 -2955
rect 183 -2989 199 -2955
rect 255 -2989 267 -2955
rect 327 -2989 335 -2955
rect 399 -2989 403 -2955
rect 505 -2989 509 -2955
rect 573 -2989 581 -2955
rect 641 -2989 653 -2955
rect 709 -2989 725 -2955
rect 777 -2989 797 -2955
rect 845 -2989 869 -2955
rect 913 -2989 941 -2955
rect 981 -2989 1013 -2955
rect 1049 -2989 1083 -2955
rect 1119 -2989 1151 -2955
rect 1191 -2989 1219 -2955
rect 1263 -2989 1287 -2955
rect 1335 -2989 1355 -2955
rect 1407 -2989 1423 -2955
rect 1479 -2989 1491 -2955
rect 1551 -2989 1559 -2955
rect 1623 -2989 1627 -2955
rect 1729 -2989 1733 -2955
rect 1797 -2989 1805 -2955
rect 1865 -2989 1877 -2955
rect 1933 -2989 1949 -2955
rect 2001 -2989 2021 -2955
rect 2069 -2989 2093 -2955
rect 2137 -2989 2165 -2955
rect 2205 -2989 2237 -2955
rect 2273 -2989 2307 -2955
rect 2343 -2989 2375 -2955
rect 2415 -2989 2443 -2955
rect 2487 -2989 2511 -2955
rect 2559 -2989 2579 -2955
rect 2631 -2989 2647 -2955
rect 2703 -2989 2715 -2955
rect 2775 -2989 2783 -2955
rect 2847 -2989 2851 -2955
rect 2953 -2989 2957 -2955
rect 3021 -2989 3029 -2955
rect 3089 -2989 3101 -2955
rect 3157 -2989 3173 -2955
rect 3225 -2989 3245 -2955
rect 3293 -2989 3317 -2955
rect 3361 -2989 3389 -2955
rect 3429 -2989 3461 -2955
rect 3497 -2989 3531 -2955
rect 3567 -2989 3599 -2955
rect 3639 -2989 3667 -2955
rect 3711 -2989 3735 -2955
rect 3783 -2989 3803 -2955
rect 3855 -2989 3871 -2955
rect 3927 -2989 3939 -2955
rect 3999 -2989 4007 -2955
rect 4071 -2989 4075 -2955
rect 4177 -2989 4181 -2955
rect 4245 -2989 4253 -2955
rect 4313 -2989 4325 -2955
rect 4381 -2989 4397 -2955
rect 4449 -2989 4469 -2955
rect 4517 -2989 4541 -2955
rect 4585 -2989 4613 -2955
rect 4653 -2989 4685 -2955
rect 4721 -2989 4755 -2955
rect 4791 -2989 4823 -2955
rect 4863 -2989 4891 -2955
rect 4935 -2989 4959 -2955
rect 5007 -2989 5027 -2955
rect 5079 -2989 5095 -2955
rect 5151 -2989 5163 -2955
rect 5223 -2989 5231 -2955
rect 5295 -2989 5299 -2955
rect 5401 -2989 5405 -2955
rect 5469 -2989 5477 -2955
rect 5537 -2989 5549 -2955
rect 5605 -2989 5621 -2955
rect 5673 -2989 5693 -2955
rect 5741 -2989 5765 -2955
rect 5809 -2989 5837 -2955
rect 5877 -2989 5909 -2955
rect 5945 -2989 5979 -2955
rect 6015 -2989 6047 -2955
rect 6087 -2989 6115 -2955
rect 6159 -2989 6183 -2955
rect 6231 -2989 6251 -2955
rect 6303 -2989 6319 -2955
rect 6375 -2989 6387 -2955
rect 6447 -2989 6455 -2955
rect 6519 -2989 6523 -2955
rect 6625 -2989 6629 -2955
rect 6693 -2989 6701 -2955
rect 6761 -2989 6773 -2955
rect 6829 -2989 6845 -2955
rect 6897 -2989 6917 -2955
rect 6965 -2989 6989 -2955
rect 7033 -2989 7061 -2955
rect 7101 -2989 7133 -2955
rect 7169 -2989 7203 -2955
rect 7239 -2989 7271 -2955
rect 7311 -2989 7339 -2955
rect 7383 -2989 7407 -2955
rect 7455 -2989 7475 -2955
rect 7527 -2989 7543 -2955
rect 7599 -2989 7611 -2955
rect 7671 -2989 7679 -2955
rect 7743 -2989 7747 -2955
rect 7849 -2989 7853 -2955
rect 7917 -2989 7925 -2955
rect 7985 -2989 7997 -2955
rect 8053 -2989 8069 -2955
rect 8121 -2989 8141 -2955
rect 8189 -2989 8213 -2955
rect 8257 -2989 8285 -2955
rect 8325 -2989 8357 -2955
rect 8393 -2989 8427 -2955
rect 8463 -2989 8495 -2955
rect 8535 -2989 8563 -2955
rect 8607 -2989 8631 -2955
rect 8679 -2989 8699 -2955
rect 8751 -2989 8767 -2955
rect 8823 -2989 8835 -2955
rect 8895 -2989 8903 -2955
rect 8967 -2989 8971 -2955
rect 9073 -2989 9077 -2955
rect 9141 -2989 9149 -2955
rect 9209 -2989 9221 -2955
rect 9277 -2989 9293 -2955
rect 9345 -2989 9365 -2955
rect 9413 -2989 9437 -2955
rect 9481 -2989 9509 -2955
rect 9549 -2989 9581 -2955
rect 9617 -2989 9651 -2955
rect 9687 -2989 9719 -2955
rect 9759 -2989 9787 -2955
rect 9831 -2989 9855 -2955
rect 9903 -2989 9923 -2955
rect 9975 -2989 9991 -2955
rect 10047 -2989 10059 -2955
rect 10119 -2989 10127 -2955
rect 10191 -2989 10195 -2955
rect 10297 -2989 10301 -2955
rect 10365 -2989 10373 -2955
rect 10433 -2989 10445 -2955
rect 10501 -2989 10517 -2955
rect 10569 -2989 10589 -2955
rect 10637 -2989 10661 -2955
rect 10705 -2989 10733 -2955
rect 10773 -2989 10805 -2955
rect 10841 -2989 10877 -2955
rect 10911 -2989 11022 -2955
rect -322 -3022 11022 -2989
<< viali >>
rect -211 2335 -177 2369
rect -139 2335 -107 2369
rect -107 2335 -105 2369
rect -67 2335 -39 2369
rect -39 2335 -33 2369
rect 5 2335 29 2369
rect 29 2335 39 2369
rect 77 2335 97 2369
rect 97 2335 111 2369
rect 149 2335 165 2369
rect 165 2335 183 2369
rect 221 2335 233 2369
rect 233 2335 255 2369
rect 293 2335 301 2369
rect 301 2335 327 2369
rect 365 2335 369 2369
rect 369 2335 399 2369
rect 437 2335 471 2369
rect 509 2335 539 2369
rect 539 2335 543 2369
rect 581 2335 607 2369
rect 607 2335 615 2369
rect 653 2335 675 2369
rect 675 2335 687 2369
rect 725 2335 743 2369
rect 743 2335 759 2369
rect 797 2335 811 2369
rect 811 2335 831 2369
rect 869 2335 879 2369
rect 879 2335 903 2369
rect 941 2335 947 2369
rect 947 2335 975 2369
rect 1013 2335 1015 2369
rect 1015 2335 1047 2369
rect 1085 2335 1117 2369
rect 1117 2335 1119 2369
rect 1157 2335 1185 2369
rect 1185 2335 1191 2369
rect 1229 2335 1253 2369
rect 1253 2335 1263 2369
rect 1301 2335 1321 2369
rect 1321 2335 1335 2369
rect 1373 2335 1389 2369
rect 1389 2335 1407 2369
rect 1445 2335 1457 2369
rect 1457 2335 1479 2369
rect 1517 2335 1525 2369
rect 1525 2335 1551 2369
rect 1589 2335 1593 2369
rect 1593 2335 1623 2369
rect 1661 2335 1695 2369
rect 1733 2335 1763 2369
rect 1763 2335 1767 2369
rect 1805 2335 1831 2369
rect 1831 2335 1839 2369
rect 1877 2335 1899 2369
rect 1899 2335 1911 2369
rect 1949 2335 1967 2369
rect 1967 2335 1983 2369
rect 2021 2335 2035 2369
rect 2035 2335 2055 2369
rect 2093 2335 2103 2369
rect 2103 2335 2127 2369
rect 2165 2335 2171 2369
rect 2171 2335 2199 2369
rect 2237 2335 2239 2369
rect 2239 2335 2271 2369
rect 2309 2335 2341 2369
rect 2341 2335 2343 2369
rect 2381 2335 2409 2369
rect 2409 2335 2415 2369
rect 2453 2335 2477 2369
rect 2477 2335 2487 2369
rect 2525 2335 2545 2369
rect 2545 2335 2559 2369
rect 2597 2335 2613 2369
rect 2613 2335 2631 2369
rect 2669 2335 2681 2369
rect 2681 2335 2703 2369
rect 2741 2335 2749 2369
rect 2749 2335 2775 2369
rect 2813 2335 2817 2369
rect 2817 2335 2847 2369
rect 2885 2335 2919 2369
rect 2957 2335 2987 2369
rect 2987 2335 2991 2369
rect 3029 2335 3055 2369
rect 3055 2335 3063 2369
rect 3101 2335 3123 2369
rect 3123 2335 3135 2369
rect 3173 2335 3191 2369
rect 3191 2335 3207 2369
rect 3245 2335 3259 2369
rect 3259 2335 3279 2369
rect 3317 2335 3327 2369
rect 3327 2335 3351 2369
rect 3389 2335 3395 2369
rect 3395 2335 3423 2369
rect 3461 2335 3463 2369
rect 3463 2335 3495 2369
rect 3533 2335 3565 2369
rect 3565 2335 3567 2369
rect 3605 2335 3633 2369
rect 3633 2335 3639 2369
rect 3677 2335 3701 2369
rect 3701 2335 3711 2369
rect 3749 2335 3769 2369
rect 3769 2335 3783 2369
rect 3821 2335 3837 2369
rect 3837 2335 3855 2369
rect 3893 2335 3905 2369
rect 3905 2335 3927 2369
rect 3965 2335 3973 2369
rect 3973 2335 3999 2369
rect 4037 2335 4041 2369
rect 4041 2335 4071 2369
rect 4109 2335 4143 2369
rect 4181 2335 4211 2369
rect 4211 2335 4215 2369
rect 4253 2335 4279 2369
rect 4279 2335 4287 2369
rect 4325 2335 4347 2369
rect 4347 2335 4359 2369
rect 4397 2335 4415 2369
rect 4415 2335 4431 2369
rect 4469 2335 4483 2369
rect 4483 2335 4503 2369
rect 4541 2335 4551 2369
rect 4551 2335 4575 2369
rect 4613 2335 4619 2369
rect 4619 2335 4647 2369
rect 4685 2335 4687 2369
rect 4687 2335 4719 2369
rect 4757 2335 4789 2369
rect 4789 2335 4791 2369
rect 4829 2335 4857 2369
rect 4857 2335 4863 2369
rect 4901 2335 4925 2369
rect 4925 2335 4935 2369
rect 4973 2335 4993 2369
rect 4993 2335 5007 2369
rect 5045 2335 5061 2369
rect 5061 2335 5079 2369
rect 5117 2335 5129 2369
rect 5129 2335 5151 2369
rect 5189 2335 5197 2369
rect 5197 2335 5223 2369
rect 5261 2335 5265 2369
rect 5265 2335 5295 2369
rect 5333 2335 5367 2369
rect 5405 2335 5435 2369
rect 5435 2335 5439 2369
rect 5477 2335 5503 2369
rect 5503 2335 5511 2369
rect 5549 2335 5571 2369
rect 5571 2335 5583 2369
rect 5621 2335 5639 2369
rect 5639 2335 5655 2369
rect 5693 2335 5707 2369
rect 5707 2335 5727 2369
rect 5765 2335 5775 2369
rect 5775 2335 5799 2369
rect 5837 2335 5843 2369
rect 5843 2335 5871 2369
rect 5909 2335 5911 2369
rect 5911 2335 5943 2369
rect 5981 2335 6013 2369
rect 6013 2335 6015 2369
rect 6053 2335 6081 2369
rect 6081 2335 6087 2369
rect 6125 2335 6149 2369
rect 6149 2335 6159 2369
rect 6197 2335 6217 2369
rect 6217 2335 6231 2369
rect 6269 2335 6285 2369
rect 6285 2335 6303 2369
rect 6341 2335 6353 2369
rect 6353 2335 6375 2369
rect 6413 2335 6421 2369
rect 6421 2335 6447 2369
rect 6485 2335 6489 2369
rect 6489 2335 6519 2369
rect 6557 2335 6591 2369
rect 6629 2335 6659 2369
rect 6659 2335 6663 2369
rect 6701 2335 6727 2369
rect 6727 2335 6735 2369
rect 6773 2335 6795 2369
rect 6795 2335 6807 2369
rect 6845 2335 6863 2369
rect 6863 2335 6879 2369
rect 6917 2335 6931 2369
rect 6931 2335 6951 2369
rect 6989 2335 6999 2369
rect 6999 2335 7023 2369
rect 7061 2335 7067 2369
rect 7067 2335 7095 2369
rect 7133 2335 7135 2369
rect 7135 2335 7167 2369
rect 7205 2335 7237 2369
rect 7237 2335 7239 2369
rect 7277 2335 7305 2369
rect 7305 2335 7311 2369
rect 7349 2335 7373 2369
rect 7373 2335 7383 2369
rect 7421 2335 7441 2369
rect 7441 2335 7455 2369
rect 7493 2335 7509 2369
rect 7509 2335 7527 2369
rect 7565 2335 7577 2369
rect 7577 2335 7599 2369
rect 7637 2335 7645 2369
rect 7645 2335 7671 2369
rect 7709 2335 7713 2369
rect 7713 2335 7743 2369
rect 7781 2335 7815 2369
rect 7853 2335 7883 2369
rect 7883 2335 7887 2369
rect 7925 2335 7951 2369
rect 7951 2335 7959 2369
rect 7997 2335 8019 2369
rect 8019 2335 8031 2369
rect 8069 2335 8087 2369
rect 8087 2335 8103 2369
rect 8141 2335 8155 2369
rect 8155 2335 8175 2369
rect 8213 2335 8223 2369
rect 8223 2335 8247 2369
rect 8285 2335 8291 2369
rect 8291 2335 8319 2369
rect 8357 2335 8359 2369
rect 8359 2335 8391 2369
rect 8429 2335 8461 2369
rect 8461 2335 8463 2369
rect 8501 2335 8529 2369
rect 8529 2335 8535 2369
rect 8573 2335 8597 2369
rect 8597 2335 8607 2369
rect 8645 2335 8665 2369
rect 8665 2335 8679 2369
rect 8717 2335 8733 2369
rect 8733 2335 8751 2369
rect 8789 2335 8801 2369
rect 8801 2335 8823 2369
rect 8861 2335 8869 2369
rect 8869 2335 8895 2369
rect 8933 2335 8937 2369
rect 8937 2335 8967 2369
rect 9005 2335 9039 2369
rect 9077 2335 9107 2369
rect 9107 2335 9111 2369
rect 9149 2335 9175 2369
rect 9175 2335 9183 2369
rect 9221 2335 9243 2369
rect 9243 2335 9255 2369
rect 9293 2335 9311 2369
rect 9311 2335 9327 2369
rect 9365 2335 9379 2369
rect 9379 2335 9399 2369
rect 9437 2335 9447 2369
rect 9447 2335 9471 2369
rect 9509 2335 9515 2369
rect 9515 2335 9543 2369
rect 9581 2335 9583 2369
rect 9583 2335 9615 2369
rect 9653 2335 9685 2369
rect 9685 2335 9687 2369
rect 9725 2335 9753 2369
rect 9753 2335 9759 2369
rect 9797 2335 9821 2369
rect 9821 2335 9831 2369
rect 9869 2335 9889 2369
rect 9889 2335 9903 2369
rect 9941 2335 9957 2369
rect 9957 2335 9975 2369
rect 10013 2335 10025 2369
rect 10025 2335 10047 2369
rect 10085 2335 10093 2369
rect 10093 2335 10119 2369
rect 10157 2335 10161 2369
rect 10161 2335 10191 2369
rect 10229 2335 10263 2369
rect 10301 2335 10331 2369
rect 10331 2335 10335 2369
rect 10373 2335 10399 2369
rect 10399 2335 10407 2369
rect 10445 2335 10467 2369
rect 10467 2335 10479 2369
rect 10517 2335 10535 2369
rect 10535 2335 10551 2369
rect 10589 2335 10603 2369
rect 10603 2335 10623 2369
rect 10661 2335 10671 2369
rect 10671 2335 10695 2369
rect 10733 2335 10739 2369
rect 10739 2335 10767 2369
rect 10805 2335 10807 2369
rect 10807 2335 10839 2369
rect 10877 2335 10911 2369
rect -289 2207 -255 2211
rect -289 2177 -255 2207
rect -289 2105 -255 2139
rect -289 2037 -255 2067
rect -289 2033 -255 2037
rect -289 1969 -255 1995
rect -289 1961 -255 1969
rect -289 1901 -255 1923
rect -289 1889 -255 1901
rect -289 1833 -255 1851
rect -289 1817 -255 1833
rect -289 1765 -255 1779
rect -289 1745 -255 1765
rect -289 1697 -255 1707
rect -289 1673 -255 1697
rect -289 1629 -255 1635
rect -289 1601 -255 1629
rect -289 1561 -255 1563
rect -289 1529 -255 1561
rect -289 1459 -255 1491
rect -289 1457 -255 1459
rect -289 1391 -255 1419
rect -289 1385 -255 1391
rect -289 1323 -255 1347
rect -289 1313 -255 1323
rect -289 1255 -255 1275
rect -289 1241 -255 1255
rect -289 1187 -255 1203
rect -289 1169 -255 1187
rect -289 1119 -255 1131
rect -289 1097 -255 1119
rect -289 1051 -255 1059
rect -289 1025 -255 1051
rect -289 983 -255 987
rect -289 953 -255 983
rect -289 881 -255 915
rect -289 813 -255 843
rect -289 809 -255 813
rect 10955 2207 10989 2211
rect 10955 2177 10989 2207
rect 10955 2105 10989 2139
rect 10955 2037 10989 2067
rect 10955 2033 10989 2037
rect 10955 1969 10989 1995
rect 10955 1961 10989 1969
rect 10955 1901 10989 1923
rect 10955 1889 10989 1901
rect 10955 1833 10989 1851
rect 10955 1817 10989 1833
rect 10955 1765 10989 1779
rect 10955 1745 10989 1765
rect 10955 1697 10989 1707
rect 10955 1673 10989 1697
rect 10955 1629 10989 1635
rect 10955 1601 10989 1629
rect 10955 1561 10989 1563
rect 10955 1529 10989 1561
rect 10955 1459 10989 1491
rect 10955 1457 10989 1459
rect 10955 1391 10989 1419
rect 10955 1385 10989 1391
rect 10955 1323 10989 1347
rect 10955 1313 10989 1323
rect 10955 1255 10989 1275
rect 10955 1241 10989 1255
rect 10955 1187 10989 1203
rect 10955 1169 10989 1187
rect 10955 1119 10989 1131
rect 10955 1097 10989 1119
rect 10955 1051 10989 1059
rect 10955 1025 10989 1051
rect 10955 983 10989 987
rect 10955 953 10989 983
rect 10955 881 10989 915
rect 10955 813 10989 843
rect 10955 809 10989 813
rect -211 651 -177 685
rect -139 651 -107 685
rect -107 651 -105 685
rect -67 651 -39 685
rect -39 651 -33 685
rect 5 651 29 685
rect 29 651 39 685
rect 77 651 97 685
rect 97 651 111 685
rect 149 651 165 685
rect 165 651 183 685
rect 221 651 233 685
rect 233 651 255 685
rect 293 651 301 685
rect 301 651 327 685
rect 365 651 369 685
rect 369 651 399 685
rect 437 651 471 685
rect 509 651 539 685
rect 539 651 543 685
rect 581 651 607 685
rect 607 651 615 685
rect 653 651 675 685
rect 675 651 687 685
rect 725 651 743 685
rect 743 651 759 685
rect 797 651 811 685
rect 811 651 831 685
rect 869 651 879 685
rect 879 651 903 685
rect 941 651 947 685
rect 947 651 975 685
rect 1013 651 1015 685
rect 1015 651 1047 685
rect 1085 651 1117 685
rect 1117 651 1119 685
rect 1157 651 1185 685
rect 1185 651 1191 685
rect 1229 651 1253 685
rect 1253 651 1263 685
rect 1301 651 1321 685
rect 1321 651 1335 685
rect 1373 651 1389 685
rect 1389 651 1407 685
rect 1445 651 1457 685
rect 1457 651 1479 685
rect 1517 651 1525 685
rect 1525 651 1551 685
rect 1589 651 1593 685
rect 1593 651 1623 685
rect 1661 651 1695 685
rect 1733 651 1763 685
rect 1763 651 1767 685
rect 1805 651 1831 685
rect 1831 651 1839 685
rect 1877 651 1899 685
rect 1899 651 1911 685
rect 1949 651 1967 685
rect 1967 651 1983 685
rect 2021 651 2035 685
rect 2035 651 2055 685
rect 2093 651 2103 685
rect 2103 651 2127 685
rect 2165 651 2171 685
rect 2171 651 2199 685
rect 2237 651 2239 685
rect 2239 651 2271 685
rect 2309 651 2341 685
rect 2341 651 2343 685
rect 2381 651 2409 685
rect 2409 651 2415 685
rect 2453 651 2477 685
rect 2477 651 2487 685
rect 2525 651 2545 685
rect 2545 651 2559 685
rect 2597 651 2613 685
rect 2613 651 2631 685
rect 2669 651 2681 685
rect 2681 651 2703 685
rect 2741 651 2749 685
rect 2749 651 2775 685
rect 2813 651 2817 685
rect 2817 651 2847 685
rect 2885 651 2919 685
rect 2957 651 2987 685
rect 2987 651 2991 685
rect 3029 651 3055 685
rect 3055 651 3063 685
rect 3101 651 3123 685
rect 3123 651 3135 685
rect 3173 651 3191 685
rect 3191 651 3207 685
rect 3245 651 3259 685
rect 3259 651 3279 685
rect 3317 651 3327 685
rect 3327 651 3351 685
rect 3389 651 3395 685
rect 3395 651 3423 685
rect 3461 651 3463 685
rect 3463 651 3495 685
rect 3533 651 3565 685
rect 3565 651 3567 685
rect 3605 651 3633 685
rect 3633 651 3639 685
rect 3677 651 3701 685
rect 3701 651 3711 685
rect 3749 651 3769 685
rect 3769 651 3783 685
rect 3821 651 3837 685
rect 3837 651 3855 685
rect 3893 651 3905 685
rect 3905 651 3927 685
rect 3965 651 3973 685
rect 3973 651 3999 685
rect 4037 651 4041 685
rect 4041 651 4071 685
rect 4109 651 4143 685
rect 4181 651 4211 685
rect 4211 651 4215 685
rect 4253 651 4279 685
rect 4279 651 4287 685
rect 4325 651 4347 685
rect 4347 651 4359 685
rect 4397 651 4415 685
rect 4415 651 4431 685
rect 4469 651 4483 685
rect 4483 651 4503 685
rect 4541 651 4551 685
rect 4551 651 4575 685
rect 4613 651 4619 685
rect 4619 651 4647 685
rect 4685 651 4687 685
rect 4687 651 4719 685
rect 4757 651 4789 685
rect 4789 651 4791 685
rect 4829 651 4857 685
rect 4857 651 4863 685
rect 4901 651 4925 685
rect 4925 651 4935 685
rect 4973 651 4993 685
rect 4993 651 5007 685
rect 5045 651 5061 685
rect 5061 651 5079 685
rect 5117 651 5129 685
rect 5129 651 5151 685
rect 5189 651 5197 685
rect 5197 651 5223 685
rect 5261 651 5265 685
rect 5265 651 5295 685
rect 5333 651 5367 685
rect 5405 651 5435 685
rect 5435 651 5439 685
rect 5477 651 5503 685
rect 5503 651 5511 685
rect 5549 651 5571 685
rect 5571 651 5583 685
rect 5621 651 5639 685
rect 5639 651 5655 685
rect 5693 651 5707 685
rect 5707 651 5727 685
rect 5765 651 5775 685
rect 5775 651 5799 685
rect 5837 651 5843 685
rect 5843 651 5871 685
rect 5909 651 5911 685
rect 5911 651 5943 685
rect 5981 651 6013 685
rect 6013 651 6015 685
rect 6053 651 6081 685
rect 6081 651 6087 685
rect 6125 651 6149 685
rect 6149 651 6159 685
rect 6197 651 6217 685
rect 6217 651 6231 685
rect 6269 651 6285 685
rect 6285 651 6303 685
rect 6341 651 6353 685
rect 6353 651 6375 685
rect 6413 651 6421 685
rect 6421 651 6447 685
rect 6485 651 6489 685
rect 6489 651 6519 685
rect 6557 651 6591 685
rect 6629 651 6659 685
rect 6659 651 6663 685
rect 6701 651 6727 685
rect 6727 651 6735 685
rect 6773 651 6795 685
rect 6795 651 6807 685
rect 6845 651 6863 685
rect 6863 651 6879 685
rect 6917 651 6931 685
rect 6931 651 6951 685
rect 6989 651 6999 685
rect 6999 651 7023 685
rect 7061 651 7067 685
rect 7067 651 7095 685
rect 7133 651 7135 685
rect 7135 651 7167 685
rect 7205 651 7237 685
rect 7237 651 7239 685
rect 7277 651 7305 685
rect 7305 651 7311 685
rect 7349 651 7373 685
rect 7373 651 7383 685
rect 7421 651 7441 685
rect 7441 651 7455 685
rect 7493 651 7509 685
rect 7509 651 7527 685
rect 7565 651 7577 685
rect 7577 651 7599 685
rect 7637 651 7645 685
rect 7645 651 7671 685
rect 7709 651 7713 685
rect 7713 651 7743 685
rect 7781 651 7815 685
rect 7853 651 7883 685
rect 7883 651 7887 685
rect 7925 651 7951 685
rect 7951 651 7959 685
rect 7997 651 8019 685
rect 8019 651 8031 685
rect 8069 651 8087 685
rect 8087 651 8103 685
rect 8141 651 8155 685
rect 8155 651 8175 685
rect 8213 651 8223 685
rect 8223 651 8247 685
rect 8285 651 8291 685
rect 8291 651 8319 685
rect 8357 651 8359 685
rect 8359 651 8391 685
rect 8429 651 8461 685
rect 8461 651 8463 685
rect 8501 651 8529 685
rect 8529 651 8535 685
rect 8573 651 8597 685
rect 8597 651 8607 685
rect 8645 651 8665 685
rect 8665 651 8679 685
rect 8717 651 8733 685
rect 8733 651 8751 685
rect 8789 651 8801 685
rect 8801 651 8823 685
rect 8861 651 8869 685
rect 8869 651 8895 685
rect 8933 651 8937 685
rect 8937 651 8967 685
rect 9005 651 9039 685
rect 9077 651 9107 685
rect 9107 651 9111 685
rect 9149 651 9175 685
rect 9175 651 9183 685
rect 9221 651 9243 685
rect 9243 651 9255 685
rect 9293 651 9311 685
rect 9311 651 9327 685
rect 9365 651 9379 685
rect 9379 651 9399 685
rect 9437 651 9447 685
rect 9447 651 9471 685
rect 9509 651 9515 685
rect 9515 651 9543 685
rect 9581 651 9583 685
rect 9583 651 9615 685
rect 9653 651 9685 685
rect 9685 651 9687 685
rect 9725 651 9753 685
rect 9753 651 9759 685
rect 9797 651 9821 685
rect 9821 651 9831 685
rect 9869 651 9889 685
rect 9889 651 9903 685
rect 9941 651 9957 685
rect 9957 651 9975 685
rect 10013 651 10025 685
rect 10025 651 10047 685
rect 10085 651 10093 685
rect 10093 651 10119 685
rect 10157 651 10161 685
rect 10161 651 10191 685
rect 10229 651 10263 685
rect 10301 651 10331 685
rect 10331 651 10335 685
rect 10373 651 10399 685
rect 10399 651 10407 685
rect 10445 651 10467 685
rect 10467 651 10479 685
rect 10517 651 10535 685
rect 10535 651 10551 685
rect 10589 651 10603 685
rect 10603 651 10623 685
rect 10661 651 10671 685
rect 10671 651 10695 685
rect 10733 651 10739 685
rect 10739 651 10767 685
rect 10805 651 10807 685
rect 10807 651 10839 685
rect 10877 651 10911 685
rect -211 315 -177 349
rect -139 315 -107 349
rect -107 315 -105 349
rect -67 315 -39 349
rect -39 315 -33 349
rect 5 315 29 349
rect 29 315 39 349
rect 77 315 97 349
rect 97 315 111 349
rect 149 315 165 349
rect 165 315 183 349
rect 221 315 233 349
rect 233 315 255 349
rect 293 315 301 349
rect 301 315 327 349
rect 365 315 369 349
rect 369 315 399 349
rect 437 315 471 349
rect 509 315 539 349
rect 539 315 543 349
rect 581 315 607 349
rect 607 315 615 349
rect 653 315 675 349
rect 675 315 687 349
rect 725 315 743 349
rect 743 315 759 349
rect 797 315 811 349
rect 811 315 831 349
rect 869 315 879 349
rect 879 315 903 349
rect 941 315 947 349
rect 947 315 975 349
rect 1013 315 1015 349
rect 1015 315 1047 349
rect 1085 315 1117 349
rect 1117 315 1119 349
rect 1157 315 1185 349
rect 1185 315 1191 349
rect 1229 315 1253 349
rect 1253 315 1263 349
rect 1301 315 1321 349
rect 1321 315 1335 349
rect 1373 315 1389 349
rect 1389 315 1407 349
rect 1445 315 1457 349
rect 1457 315 1479 349
rect 1517 315 1525 349
rect 1525 315 1551 349
rect 1589 315 1593 349
rect 1593 315 1623 349
rect 1661 315 1695 349
rect 1733 315 1763 349
rect 1763 315 1767 349
rect 1805 315 1831 349
rect 1831 315 1839 349
rect 1877 315 1899 349
rect 1899 315 1911 349
rect 1949 315 1967 349
rect 1967 315 1983 349
rect 2021 315 2035 349
rect 2035 315 2055 349
rect 2093 315 2103 349
rect 2103 315 2127 349
rect 2165 315 2171 349
rect 2171 315 2199 349
rect 2237 315 2239 349
rect 2239 315 2271 349
rect 2309 315 2341 349
rect 2341 315 2343 349
rect 2381 315 2409 349
rect 2409 315 2415 349
rect 2453 315 2477 349
rect 2477 315 2487 349
rect 2525 315 2545 349
rect 2545 315 2559 349
rect 2597 315 2613 349
rect 2613 315 2631 349
rect 2669 315 2681 349
rect 2681 315 2703 349
rect 2741 315 2749 349
rect 2749 315 2775 349
rect 2813 315 2817 349
rect 2817 315 2847 349
rect 2885 315 2919 349
rect 2957 315 2987 349
rect 2987 315 2991 349
rect 3029 315 3055 349
rect 3055 315 3063 349
rect 3101 315 3123 349
rect 3123 315 3135 349
rect 3173 315 3191 349
rect 3191 315 3207 349
rect 3245 315 3259 349
rect 3259 315 3279 349
rect 3317 315 3327 349
rect 3327 315 3351 349
rect 3389 315 3395 349
rect 3395 315 3423 349
rect 3461 315 3463 349
rect 3463 315 3495 349
rect 3533 315 3565 349
rect 3565 315 3567 349
rect 3605 315 3633 349
rect 3633 315 3639 349
rect 3677 315 3701 349
rect 3701 315 3711 349
rect 3749 315 3769 349
rect 3769 315 3783 349
rect 3821 315 3837 349
rect 3837 315 3855 349
rect 3893 315 3905 349
rect 3905 315 3927 349
rect 3965 315 3973 349
rect 3973 315 3999 349
rect 4037 315 4041 349
rect 4041 315 4071 349
rect 4109 315 4143 349
rect 4181 315 4211 349
rect 4211 315 4215 349
rect 4253 315 4279 349
rect 4279 315 4287 349
rect 4325 315 4347 349
rect 4347 315 4359 349
rect 4397 315 4415 349
rect 4415 315 4431 349
rect 4469 315 4483 349
rect 4483 315 4503 349
rect 4541 315 4551 349
rect 4551 315 4575 349
rect 4613 315 4619 349
rect 4619 315 4647 349
rect 4685 315 4687 349
rect 4687 315 4719 349
rect 4757 315 4789 349
rect 4789 315 4791 349
rect 4829 315 4857 349
rect 4857 315 4863 349
rect 4901 315 4925 349
rect 4925 315 4935 349
rect 4973 315 4993 349
rect 4993 315 5007 349
rect 5045 315 5061 349
rect 5061 315 5079 349
rect 5117 315 5129 349
rect 5129 315 5151 349
rect 5189 315 5197 349
rect 5197 315 5223 349
rect 5261 315 5265 349
rect 5265 315 5295 349
rect 5333 315 5367 349
rect 5405 315 5435 349
rect 5435 315 5439 349
rect 5477 315 5503 349
rect 5503 315 5511 349
rect 5549 315 5571 349
rect 5571 315 5583 349
rect 5621 315 5639 349
rect 5639 315 5655 349
rect 5693 315 5707 349
rect 5707 315 5727 349
rect 5765 315 5775 349
rect 5775 315 5799 349
rect 5837 315 5843 349
rect 5843 315 5871 349
rect 5909 315 5911 349
rect 5911 315 5943 349
rect 5981 315 6013 349
rect 6013 315 6015 349
rect 6053 315 6081 349
rect 6081 315 6087 349
rect 6125 315 6149 349
rect 6149 315 6159 349
rect 6197 315 6217 349
rect 6217 315 6231 349
rect 6269 315 6285 349
rect 6285 315 6303 349
rect 6341 315 6353 349
rect 6353 315 6375 349
rect 6413 315 6421 349
rect 6421 315 6447 349
rect 6485 315 6489 349
rect 6489 315 6519 349
rect 6557 315 6591 349
rect 6629 315 6659 349
rect 6659 315 6663 349
rect 6701 315 6727 349
rect 6727 315 6735 349
rect 6773 315 6795 349
rect 6795 315 6807 349
rect 6845 315 6863 349
rect 6863 315 6879 349
rect 6917 315 6931 349
rect 6931 315 6951 349
rect 6989 315 6999 349
rect 6999 315 7023 349
rect 7061 315 7067 349
rect 7067 315 7095 349
rect 7133 315 7135 349
rect 7135 315 7167 349
rect 7205 315 7237 349
rect 7237 315 7239 349
rect 7277 315 7305 349
rect 7305 315 7311 349
rect 7349 315 7373 349
rect 7373 315 7383 349
rect 7421 315 7441 349
rect 7441 315 7455 349
rect 7493 315 7509 349
rect 7509 315 7527 349
rect 7565 315 7577 349
rect 7577 315 7599 349
rect 7637 315 7645 349
rect 7645 315 7671 349
rect 7709 315 7713 349
rect 7713 315 7743 349
rect 7781 315 7815 349
rect 7853 315 7883 349
rect 7883 315 7887 349
rect 7925 315 7951 349
rect 7951 315 7959 349
rect 7997 315 8019 349
rect 8019 315 8031 349
rect 8069 315 8087 349
rect 8087 315 8103 349
rect 8141 315 8155 349
rect 8155 315 8175 349
rect 8213 315 8223 349
rect 8223 315 8247 349
rect 8285 315 8291 349
rect 8291 315 8319 349
rect 8357 315 8359 349
rect 8359 315 8391 349
rect 8429 315 8461 349
rect 8461 315 8463 349
rect 8501 315 8529 349
rect 8529 315 8535 349
rect 8573 315 8597 349
rect 8597 315 8607 349
rect 8645 315 8665 349
rect 8665 315 8679 349
rect 8717 315 8733 349
rect 8733 315 8751 349
rect 8789 315 8801 349
rect 8801 315 8823 349
rect 8861 315 8869 349
rect 8869 315 8895 349
rect 8933 315 8937 349
rect 8937 315 8967 349
rect 9005 315 9039 349
rect 9077 315 9107 349
rect 9107 315 9111 349
rect 9149 315 9175 349
rect 9175 315 9183 349
rect 9221 315 9243 349
rect 9243 315 9255 349
rect 9293 315 9311 349
rect 9311 315 9327 349
rect 9365 315 9379 349
rect 9379 315 9399 349
rect 9437 315 9447 349
rect 9447 315 9471 349
rect 9509 315 9515 349
rect 9515 315 9543 349
rect 9581 315 9583 349
rect 9583 315 9615 349
rect 9653 315 9685 349
rect 9685 315 9687 349
rect 9725 315 9753 349
rect 9753 315 9759 349
rect 9797 315 9821 349
rect 9821 315 9831 349
rect 9869 315 9889 349
rect 9889 315 9903 349
rect 9941 315 9957 349
rect 9957 315 9975 349
rect 10013 315 10025 349
rect 10025 315 10047 349
rect 10085 315 10093 349
rect 10093 315 10119 349
rect 10157 315 10161 349
rect 10161 315 10191 349
rect 10229 315 10263 349
rect 10301 315 10331 349
rect 10331 315 10335 349
rect 10373 315 10399 349
rect 10399 315 10407 349
rect 10445 315 10467 349
rect 10467 315 10479 349
rect 10517 315 10535 349
rect 10535 315 10551 349
rect 10589 315 10603 349
rect 10603 315 10623 349
rect 10661 315 10671 349
rect 10671 315 10695 349
rect 10733 315 10739 349
rect 10739 315 10767 349
rect 10805 315 10807 349
rect 10807 315 10839 349
rect 10877 315 10911 349
rect -289 91 -255 101
rect -289 67 -255 91
rect -289 23 -255 29
rect -289 -5 -255 23
rect -289 -45 -255 -43
rect -289 -77 -255 -45
rect -289 -147 -255 -115
rect -289 -149 -255 -147
rect -289 -215 -255 -187
rect -289 -221 -255 -215
rect -289 -283 -255 -259
rect -289 -293 -255 -283
rect -289 -351 -255 -331
rect -289 -365 -255 -351
rect -289 -419 -255 -403
rect -289 -437 -255 -419
rect -289 -487 -255 -475
rect -289 -509 -255 -487
rect -289 -555 -255 -547
rect -289 -581 -255 -555
rect -289 -623 -255 -619
rect -289 -653 -255 -623
rect -289 -725 -255 -691
rect -289 -793 -255 -763
rect -289 -797 -255 -793
rect -289 -861 -255 -835
rect -289 -869 -255 -861
rect -289 -929 -255 -907
rect -289 -941 -255 -929
rect -289 -997 -255 -979
rect -289 -1013 -255 -997
rect -289 -1065 -255 -1051
rect -289 -1085 -255 -1065
rect -289 -1133 -255 -1123
rect -289 -1157 -255 -1133
rect -289 -1201 -255 -1195
rect -289 -1229 -255 -1201
rect -289 -1269 -255 -1267
rect -289 -1301 -255 -1269
rect -289 -1371 -255 -1339
rect -289 -1373 -255 -1371
rect -289 -1439 -255 -1411
rect -289 -1445 -255 -1439
rect -289 -1507 -255 -1483
rect -289 -1517 -255 -1507
rect -289 -1575 -255 -1555
rect -289 -1589 -255 -1575
rect -289 -1643 -255 -1627
rect -289 -1661 -255 -1643
rect -289 -1711 -255 -1699
rect -289 -1733 -255 -1711
rect -289 -1779 -255 -1771
rect -289 -1805 -255 -1779
rect -289 -1847 -255 -1843
rect -289 -1877 -255 -1847
rect -289 -1949 -255 -1915
rect -289 -2017 -255 -1987
rect -289 -2021 -255 -2017
rect -289 -2085 -255 -2059
rect -289 -2093 -255 -2085
rect -289 -2153 -255 -2131
rect -289 -2165 -255 -2153
rect -289 -2221 -255 -2203
rect -289 -2237 -255 -2221
rect -289 -2289 -255 -2275
rect -289 -2309 -255 -2289
rect -289 -2357 -255 -2347
rect -289 -2381 -255 -2357
rect -289 -2425 -255 -2419
rect -289 -2453 -255 -2425
rect -289 -2493 -255 -2491
rect -289 -2525 -255 -2493
rect -289 -2595 -255 -2563
rect -289 -2597 -255 -2595
rect -289 -2663 -255 -2635
rect -289 -2669 -255 -2663
rect -289 -2731 -255 -2707
rect -289 -2741 -255 -2731
rect 10955 91 10989 101
rect 10955 67 10989 91
rect 10955 23 10989 29
rect 10955 -5 10989 23
rect 10955 -45 10989 -43
rect 10955 -77 10989 -45
rect 10955 -147 10989 -115
rect 10955 -149 10989 -147
rect 10955 -215 10989 -187
rect 10955 -221 10989 -215
rect 10955 -283 10989 -259
rect 10955 -293 10989 -283
rect 10955 -351 10989 -331
rect 10955 -365 10989 -351
rect 10955 -419 10989 -403
rect 10955 -437 10989 -419
rect 10955 -487 10989 -475
rect 10955 -509 10989 -487
rect 10955 -555 10989 -547
rect 10955 -581 10989 -555
rect 10955 -623 10989 -619
rect 10955 -653 10989 -623
rect 10955 -725 10989 -691
rect 10955 -793 10989 -763
rect 10955 -797 10989 -793
rect 10955 -861 10989 -835
rect 10955 -869 10989 -861
rect 10955 -929 10989 -907
rect 10955 -941 10989 -929
rect 10955 -997 10989 -979
rect 10955 -1013 10989 -997
rect 10955 -1065 10989 -1051
rect 10955 -1085 10989 -1065
rect 10955 -1133 10989 -1123
rect 10955 -1157 10989 -1133
rect 10955 -1201 10989 -1195
rect 10955 -1229 10989 -1201
rect 10955 -1269 10989 -1267
rect 10955 -1301 10989 -1269
rect 10955 -1371 10989 -1339
rect 10955 -1373 10989 -1371
rect 10955 -1439 10989 -1411
rect 10955 -1445 10989 -1439
rect 10955 -1507 10989 -1483
rect 10955 -1517 10989 -1507
rect 10955 -1575 10989 -1555
rect 10955 -1589 10989 -1575
rect 10955 -1643 10989 -1627
rect 10955 -1661 10989 -1643
rect 10955 -1711 10989 -1699
rect 10955 -1733 10989 -1711
rect 10955 -1779 10989 -1771
rect 10955 -1805 10989 -1779
rect 10955 -1847 10989 -1843
rect 10955 -1877 10989 -1847
rect 10955 -1949 10989 -1915
rect 10955 -2017 10989 -1987
rect 10955 -2021 10989 -2017
rect 10955 -2085 10989 -2059
rect 10955 -2093 10989 -2085
rect 10955 -2153 10989 -2131
rect 10955 -2165 10989 -2153
rect 10955 -2221 10989 -2203
rect 10955 -2237 10989 -2221
rect 10955 -2289 10989 -2275
rect 10955 -2309 10989 -2289
rect 10955 -2357 10989 -2347
rect 10955 -2381 10989 -2357
rect 10955 -2425 10989 -2419
rect 10955 -2453 10989 -2425
rect 10955 -2493 10989 -2491
rect 10955 -2525 10989 -2493
rect 10955 -2595 10989 -2563
rect 10955 -2597 10989 -2595
rect 10955 -2663 10989 -2635
rect 10955 -2669 10989 -2663
rect 10955 -2731 10989 -2707
rect 10955 -2741 10989 -2731
rect -211 -2989 -177 -2955
rect -139 -2989 -107 -2955
rect -107 -2989 -105 -2955
rect -67 -2989 -39 -2955
rect -39 -2989 -33 -2955
rect 5 -2989 29 -2955
rect 29 -2989 39 -2955
rect 77 -2989 97 -2955
rect 97 -2989 111 -2955
rect 149 -2989 165 -2955
rect 165 -2989 183 -2955
rect 221 -2989 233 -2955
rect 233 -2989 255 -2955
rect 293 -2989 301 -2955
rect 301 -2989 327 -2955
rect 365 -2989 369 -2955
rect 369 -2989 399 -2955
rect 437 -2989 471 -2955
rect 509 -2989 539 -2955
rect 539 -2989 543 -2955
rect 581 -2989 607 -2955
rect 607 -2989 615 -2955
rect 653 -2989 675 -2955
rect 675 -2989 687 -2955
rect 725 -2989 743 -2955
rect 743 -2989 759 -2955
rect 797 -2989 811 -2955
rect 811 -2989 831 -2955
rect 869 -2989 879 -2955
rect 879 -2989 903 -2955
rect 941 -2989 947 -2955
rect 947 -2989 975 -2955
rect 1013 -2989 1015 -2955
rect 1015 -2989 1047 -2955
rect 1085 -2989 1117 -2955
rect 1117 -2989 1119 -2955
rect 1157 -2989 1185 -2955
rect 1185 -2989 1191 -2955
rect 1229 -2989 1253 -2955
rect 1253 -2989 1263 -2955
rect 1301 -2989 1321 -2955
rect 1321 -2989 1335 -2955
rect 1373 -2989 1389 -2955
rect 1389 -2989 1407 -2955
rect 1445 -2989 1457 -2955
rect 1457 -2989 1479 -2955
rect 1517 -2989 1525 -2955
rect 1525 -2989 1551 -2955
rect 1589 -2989 1593 -2955
rect 1593 -2989 1623 -2955
rect 1661 -2989 1695 -2955
rect 1733 -2989 1763 -2955
rect 1763 -2989 1767 -2955
rect 1805 -2989 1831 -2955
rect 1831 -2989 1839 -2955
rect 1877 -2989 1899 -2955
rect 1899 -2989 1911 -2955
rect 1949 -2989 1967 -2955
rect 1967 -2989 1983 -2955
rect 2021 -2989 2035 -2955
rect 2035 -2989 2055 -2955
rect 2093 -2989 2103 -2955
rect 2103 -2989 2127 -2955
rect 2165 -2989 2171 -2955
rect 2171 -2989 2199 -2955
rect 2237 -2989 2239 -2955
rect 2239 -2989 2271 -2955
rect 2309 -2989 2341 -2955
rect 2341 -2989 2343 -2955
rect 2381 -2989 2409 -2955
rect 2409 -2989 2415 -2955
rect 2453 -2989 2477 -2955
rect 2477 -2989 2487 -2955
rect 2525 -2989 2545 -2955
rect 2545 -2989 2559 -2955
rect 2597 -2989 2613 -2955
rect 2613 -2989 2631 -2955
rect 2669 -2989 2681 -2955
rect 2681 -2989 2703 -2955
rect 2741 -2989 2749 -2955
rect 2749 -2989 2775 -2955
rect 2813 -2989 2817 -2955
rect 2817 -2989 2847 -2955
rect 2885 -2989 2919 -2955
rect 2957 -2989 2987 -2955
rect 2987 -2989 2991 -2955
rect 3029 -2989 3055 -2955
rect 3055 -2989 3063 -2955
rect 3101 -2989 3123 -2955
rect 3123 -2989 3135 -2955
rect 3173 -2989 3191 -2955
rect 3191 -2989 3207 -2955
rect 3245 -2989 3259 -2955
rect 3259 -2989 3279 -2955
rect 3317 -2989 3327 -2955
rect 3327 -2989 3351 -2955
rect 3389 -2989 3395 -2955
rect 3395 -2989 3423 -2955
rect 3461 -2989 3463 -2955
rect 3463 -2989 3495 -2955
rect 3533 -2989 3565 -2955
rect 3565 -2989 3567 -2955
rect 3605 -2989 3633 -2955
rect 3633 -2989 3639 -2955
rect 3677 -2989 3701 -2955
rect 3701 -2989 3711 -2955
rect 3749 -2989 3769 -2955
rect 3769 -2989 3783 -2955
rect 3821 -2989 3837 -2955
rect 3837 -2989 3855 -2955
rect 3893 -2989 3905 -2955
rect 3905 -2989 3927 -2955
rect 3965 -2989 3973 -2955
rect 3973 -2989 3999 -2955
rect 4037 -2989 4041 -2955
rect 4041 -2989 4071 -2955
rect 4109 -2989 4143 -2955
rect 4181 -2989 4211 -2955
rect 4211 -2989 4215 -2955
rect 4253 -2989 4279 -2955
rect 4279 -2989 4287 -2955
rect 4325 -2989 4347 -2955
rect 4347 -2989 4359 -2955
rect 4397 -2989 4415 -2955
rect 4415 -2989 4431 -2955
rect 4469 -2989 4483 -2955
rect 4483 -2989 4503 -2955
rect 4541 -2989 4551 -2955
rect 4551 -2989 4575 -2955
rect 4613 -2989 4619 -2955
rect 4619 -2989 4647 -2955
rect 4685 -2989 4687 -2955
rect 4687 -2989 4719 -2955
rect 4757 -2989 4789 -2955
rect 4789 -2989 4791 -2955
rect 4829 -2989 4857 -2955
rect 4857 -2989 4863 -2955
rect 4901 -2989 4925 -2955
rect 4925 -2989 4935 -2955
rect 4973 -2989 4993 -2955
rect 4993 -2989 5007 -2955
rect 5045 -2989 5061 -2955
rect 5061 -2989 5079 -2955
rect 5117 -2989 5129 -2955
rect 5129 -2989 5151 -2955
rect 5189 -2989 5197 -2955
rect 5197 -2989 5223 -2955
rect 5261 -2989 5265 -2955
rect 5265 -2989 5295 -2955
rect 5333 -2989 5367 -2955
rect 5405 -2989 5435 -2955
rect 5435 -2989 5439 -2955
rect 5477 -2989 5503 -2955
rect 5503 -2989 5511 -2955
rect 5549 -2989 5571 -2955
rect 5571 -2989 5583 -2955
rect 5621 -2989 5639 -2955
rect 5639 -2989 5655 -2955
rect 5693 -2989 5707 -2955
rect 5707 -2989 5727 -2955
rect 5765 -2989 5775 -2955
rect 5775 -2989 5799 -2955
rect 5837 -2989 5843 -2955
rect 5843 -2989 5871 -2955
rect 5909 -2989 5911 -2955
rect 5911 -2989 5943 -2955
rect 5981 -2989 6013 -2955
rect 6013 -2989 6015 -2955
rect 6053 -2989 6081 -2955
rect 6081 -2989 6087 -2955
rect 6125 -2989 6149 -2955
rect 6149 -2989 6159 -2955
rect 6197 -2989 6217 -2955
rect 6217 -2989 6231 -2955
rect 6269 -2989 6285 -2955
rect 6285 -2989 6303 -2955
rect 6341 -2989 6353 -2955
rect 6353 -2989 6375 -2955
rect 6413 -2989 6421 -2955
rect 6421 -2989 6447 -2955
rect 6485 -2989 6489 -2955
rect 6489 -2989 6519 -2955
rect 6557 -2989 6591 -2955
rect 6629 -2989 6659 -2955
rect 6659 -2989 6663 -2955
rect 6701 -2989 6727 -2955
rect 6727 -2989 6735 -2955
rect 6773 -2989 6795 -2955
rect 6795 -2989 6807 -2955
rect 6845 -2989 6863 -2955
rect 6863 -2989 6879 -2955
rect 6917 -2989 6931 -2955
rect 6931 -2989 6951 -2955
rect 6989 -2989 6999 -2955
rect 6999 -2989 7023 -2955
rect 7061 -2989 7067 -2955
rect 7067 -2989 7095 -2955
rect 7133 -2989 7135 -2955
rect 7135 -2989 7167 -2955
rect 7205 -2989 7237 -2955
rect 7237 -2989 7239 -2955
rect 7277 -2989 7305 -2955
rect 7305 -2989 7311 -2955
rect 7349 -2989 7373 -2955
rect 7373 -2989 7383 -2955
rect 7421 -2989 7441 -2955
rect 7441 -2989 7455 -2955
rect 7493 -2989 7509 -2955
rect 7509 -2989 7527 -2955
rect 7565 -2989 7577 -2955
rect 7577 -2989 7599 -2955
rect 7637 -2989 7645 -2955
rect 7645 -2989 7671 -2955
rect 7709 -2989 7713 -2955
rect 7713 -2989 7743 -2955
rect 7781 -2989 7815 -2955
rect 7853 -2989 7883 -2955
rect 7883 -2989 7887 -2955
rect 7925 -2989 7951 -2955
rect 7951 -2989 7959 -2955
rect 7997 -2989 8019 -2955
rect 8019 -2989 8031 -2955
rect 8069 -2989 8087 -2955
rect 8087 -2989 8103 -2955
rect 8141 -2989 8155 -2955
rect 8155 -2989 8175 -2955
rect 8213 -2989 8223 -2955
rect 8223 -2989 8247 -2955
rect 8285 -2989 8291 -2955
rect 8291 -2989 8319 -2955
rect 8357 -2989 8359 -2955
rect 8359 -2989 8391 -2955
rect 8429 -2989 8461 -2955
rect 8461 -2989 8463 -2955
rect 8501 -2989 8529 -2955
rect 8529 -2989 8535 -2955
rect 8573 -2989 8597 -2955
rect 8597 -2989 8607 -2955
rect 8645 -2989 8665 -2955
rect 8665 -2989 8679 -2955
rect 8717 -2989 8733 -2955
rect 8733 -2989 8751 -2955
rect 8789 -2989 8801 -2955
rect 8801 -2989 8823 -2955
rect 8861 -2989 8869 -2955
rect 8869 -2989 8895 -2955
rect 8933 -2989 8937 -2955
rect 8937 -2989 8967 -2955
rect 9005 -2989 9039 -2955
rect 9077 -2989 9107 -2955
rect 9107 -2989 9111 -2955
rect 9149 -2989 9175 -2955
rect 9175 -2989 9183 -2955
rect 9221 -2989 9243 -2955
rect 9243 -2989 9255 -2955
rect 9293 -2989 9311 -2955
rect 9311 -2989 9327 -2955
rect 9365 -2989 9379 -2955
rect 9379 -2989 9399 -2955
rect 9437 -2989 9447 -2955
rect 9447 -2989 9471 -2955
rect 9509 -2989 9515 -2955
rect 9515 -2989 9543 -2955
rect 9581 -2989 9583 -2955
rect 9583 -2989 9615 -2955
rect 9653 -2989 9685 -2955
rect 9685 -2989 9687 -2955
rect 9725 -2989 9753 -2955
rect 9753 -2989 9759 -2955
rect 9797 -2989 9821 -2955
rect 9821 -2989 9831 -2955
rect 9869 -2989 9889 -2955
rect 9889 -2989 9903 -2955
rect 9941 -2989 9957 -2955
rect 9957 -2989 9975 -2955
rect 10013 -2989 10025 -2955
rect 10025 -2989 10047 -2955
rect 10085 -2989 10093 -2955
rect 10093 -2989 10119 -2955
rect 10157 -2989 10161 -2955
rect 10161 -2989 10191 -2955
rect 10229 -2989 10263 -2955
rect 10301 -2989 10331 -2955
rect 10331 -2989 10335 -2955
rect 10373 -2989 10399 -2955
rect 10399 -2989 10407 -2955
rect 10445 -2989 10467 -2955
rect 10467 -2989 10479 -2955
rect 10517 -2989 10535 -2955
rect 10535 -2989 10551 -2955
rect 10589 -2989 10603 -2955
rect 10603 -2989 10623 -2955
rect 10661 -2989 10671 -2955
rect 10671 -2989 10695 -2955
rect 10733 -2989 10739 -2955
rect 10739 -2989 10767 -2955
rect 10805 -2989 10807 -2955
rect 10807 -2989 10839 -2955
rect 10877 -2989 10911 -2955
<< metal1 >>
rect -328 2369 11028 2408
rect -328 2335 -211 2369
rect -177 2335 -139 2369
rect -105 2335 -67 2369
rect -33 2335 5 2369
rect 39 2335 77 2369
rect 111 2335 149 2369
rect 183 2335 221 2369
rect 255 2335 293 2369
rect 327 2335 365 2369
rect 399 2335 437 2369
rect 471 2335 509 2369
rect 543 2335 581 2369
rect 615 2335 653 2369
rect 687 2335 725 2369
rect 759 2335 797 2369
rect 831 2335 869 2369
rect 903 2335 941 2369
rect 975 2335 1013 2369
rect 1047 2335 1085 2369
rect 1119 2335 1157 2369
rect 1191 2335 1229 2369
rect 1263 2335 1301 2369
rect 1335 2335 1373 2369
rect 1407 2335 1445 2369
rect 1479 2335 1517 2369
rect 1551 2335 1589 2369
rect 1623 2335 1661 2369
rect 1695 2335 1733 2369
rect 1767 2335 1805 2369
rect 1839 2335 1877 2369
rect 1911 2335 1949 2369
rect 1983 2335 2021 2369
rect 2055 2335 2093 2369
rect 2127 2335 2165 2369
rect 2199 2335 2237 2369
rect 2271 2335 2309 2369
rect 2343 2335 2381 2369
rect 2415 2335 2453 2369
rect 2487 2335 2525 2369
rect 2559 2335 2597 2369
rect 2631 2335 2669 2369
rect 2703 2335 2741 2369
rect 2775 2335 2813 2369
rect 2847 2335 2885 2369
rect 2919 2335 2957 2369
rect 2991 2335 3029 2369
rect 3063 2335 3101 2369
rect 3135 2335 3173 2369
rect 3207 2335 3245 2369
rect 3279 2335 3317 2369
rect 3351 2335 3389 2369
rect 3423 2335 3461 2369
rect 3495 2335 3533 2369
rect 3567 2335 3605 2369
rect 3639 2335 3677 2369
rect 3711 2335 3749 2369
rect 3783 2335 3821 2369
rect 3855 2335 3893 2369
rect 3927 2335 3965 2369
rect 3999 2335 4037 2369
rect 4071 2335 4109 2369
rect 4143 2335 4181 2369
rect 4215 2335 4253 2369
rect 4287 2335 4325 2369
rect 4359 2335 4397 2369
rect 4431 2335 4469 2369
rect 4503 2335 4541 2369
rect 4575 2335 4613 2369
rect 4647 2335 4685 2369
rect 4719 2335 4757 2369
rect 4791 2335 4829 2369
rect 4863 2335 4901 2369
rect 4935 2335 4973 2369
rect 5007 2335 5045 2369
rect 5079 2335 5117 2369
rect 5151 2335 5189 2369
rect 5223 2335 5261 2369
rect 5295 2335 5333 2369
rect 5367 2335 5405 2369
rect 5439 2335 5477 2369
rect 5511 2335 5549 2369
rect 5583 2335 5621 2369
rect 5655 2335 5693 2369
rect 5727 2335 5765 2369
rect 5799 2335 5837 2369
rect 5871 2335 5909 2369
rect 5943 2335 5981 2369
rect 6015 2335 6053 2369
rect 6087 2335 6125 2369
rect 6159 2335 6197 2369
rect 6231 2335 6269 2369
rect 6303 2335 6341 2369
rect 6375 2335 6413 2369
rect 6447 2335 6485 2369
rect 6519 2335 6557 2369
rect 6591 2335 6629 2369
rect 6663 2335 6701 2369
rect 6735 2335 6773 2369
rect 6807 2335 6845 2369
rect 6879 2335 6917 2369
rect 6951 2335 6989 2369
rect 7023 2335 7061 2369
rect 7095 2335 7133 2369
rect 7167 2335 7205 2369
rect 7239 2335 7277 2369
rect 7311 2335 7349 2369
rect 7383 2335 7421 2369
rect 7455 2335 7493 2369
rect 7527 2335 7565 2369
rect 7599 2335 7637 2369
rect 7671 2335 7709 2369
rect 7743 2335 7781 2369
rect 7815 2335 7853 2369
rect 7887 2335 7925 2369
rect 7959 2335 7997 2369
rect 8031 2335 8069 2369
rect 8103 2335 8141 2369
rect 8175 2335 8213 2369
rect 8247 2335 8285 2369
rect 8319 2335 8357 2369
rect 8391 2335 8429 2369
rect 8463 2335 8501 2369
rect 8535 2335 8573 2369
rect 8607 2335 8645 2369
rect 8679 2335 8717 2369
rect 8751 2335 8789 2369
rect 8823 2335 8861 2369
rect 8895 2335 8933 2369
rect 8967 2335 9005 2369
rect 9039 2335 9077 2369
rect 9111 2335 9149 2369
rect 9183 2335 9221 2369
rect 9255 2335 9293 2369
rect 9327 2335 9365 2369
rect 9399 2335 9437 2369
rect 9471 2335 9509 2369
rect 9543 2335 9581 2369
rect 9615 2335 9653 2369
rect 9687 2335 9725 2369
rect 9759 2335 9797 2369
rect 9831 2335 9869 2369
rect 9903 2335 9941 2369
rect 9975 2335 10013 2369
rect 10047 2335 10085 2369
rect 10119 2335 10157 2369
rect 10191 2335 10229 2369
rect 10263 2335 10301 2369
rect 10335 2335 10373 2369
rect 10407 2335 10445 2369
rect 10479 2335 10517 2369
rect 10551 2335 10589 2369
rect 10623 2335 10661 2369
rect 10695 2335 10733 2369
rect 10767 2335 10805 2369
rect 10839 2335 10877 2369
rect 10911 2335 11028 2369
rect -328 2296 11028 2335
rect -328 2268 394 2296
rect -328 2211 -198 2268
rect -328 2177 -289 2211
rect -255 2177 -198 2211
rect -328 2139 -198 2177
rect -328 2105 -289 2139
rect -255 2105 -198 2139
rect -328 2067 -198 2105
rect -328 2033 -289 2067
rect -255 2033 -198 2067
rect -328 2024 -198 2033
rect 366 2024 394 2268
rect -328 1996 394 2024
rect 10306 2268 11028 2296
rect 10306 2024 10334 2268
rect 10898 2211 11028 2268
rect 10898 2177 10955 2211
rect 10989 2177 11028 2211
rect 10898 2139 11028 2177
rect 10898 2105 10955 2139
rect 10989 2105 11028 2139
rect 10898 2067 11028 2105
rect 10898 2033 10955 2067
rect 10989 2033 11028 2067
rect 10898 2024 11028 2033
rect 10306 1996 11028 2024
rect -328 1995 -216 1996
rect -328 1961 -289 1995
rect -255 1961 -216 1995
rect -328 1923 -216 1961
rect 10916 1995 11028 1996
rect 10916 1961 10955 1995
rect 10989 1961 11028 1995
rect -328 1889 -289 1923
rect -255 1889 -216 1923
rect -328 1851 -216 1889
rect -328 1817 -289 1851
rect -255 1817 -216 1851
rect -328 1779 -216 1817
rect -328 1745 -289 1779
rect -255 1745 -216 1779
rect -328 1707 -216 1745
rect 3466 1892 7322 1950
rect 3466 1776 3514 1892
rect 7278 1776 7322 1892
rect 3466 1720 7322 1776
rect 10916 1923 11028 1961
rect 10916 1889 10955 1923
rect 10989 1889 11028 1923
rect 10916 1851 11028 1889
rect 10916 1817 10955 1851
rect 10989 1817 11028 1851
rect 10916 1779 11028 1817
rect 10916 1745 10955 1779
rect 10989 1745 11028 1779
rect -328 1673 -289 1707
rect -255 1673 -216 1707
rect -328 1635 -216 1673
rect -328 1601 -289 1635
rect -255 1601 -216 1635
rect -328 1563 -216 1601
rect -328 1529 -289 1563
rect -255 1529 -216 1563
rect -328 1491 -216 1529
rect -328 1457 -289 1491
rect -255 1457 -216 1491
rect -328 1419 -216 1457
rect -328 1385 -289 1419
rect -255 1385 -216 1419
rect -328 1347 -216 1385
rect -328 1313 -289 1347
rect -255 1313 -216 1347
rect -328 1275 -216 1313
rect -328 1241 -289 1275
rect -255 1241 -216 1275
rect -328 1203 -216 1241
rect -328 1169 -289 1203
rect -255 1169 -216 1203
rect -328 1131 -216 1169
rect -328 1097 -289 1131
rect -255 1097 -216 1131
rect -328 1059 -216 1097
rect -328 1025 -289 1059
rect -255 1025 -216 1059
rect -328 987 -216 1025
rect -328 953 -289 987
rect -255 953 -216 987
rect -328 915 -216 953
rect -328 881 -289 915
rect -255 881 -216 915
rect -328 843 -216 881
rect -328 809 -289 843
rect -255 809 -216 843
rect -328 724 -216 809
rect 3504 1503 3564 1720
rect 3640 1503 3700 1720
rect 3504 1443 3700 1503
rect 3504 956 3564 1443
rect 3640 1336 3700 1443
rect 4022 1248 4082 1720
rect 4412 1498 4472 1720
rect 4538 1498 4598 1720
rect 4412 1438 4598 1498
rect 4412 1334 4472 1438
rect 3636 956 3696 1042
rect 3504 896 3696 956
rect 3504 724 3564 896
rect 3636 724 3696 896
rect 3764 952 3824 1142
rect 3896 952 3956 1042
rect 4152 952 4212 1042
rect 3764 948 4218 952
rect 3764 896 4156 948
rect 4208 896 4218 948
rect 3764 892 4218 896
rect 4280 838 4340 1125
rect 4280 786 4284 838
rect 4336 786 4340 838
rect 4280 776 4340 786
rect 4538 724 4598 1438
rect 4926 1503 4986 1720
rect 5054 1503 5114 1720
rect 5178 1503 5238 1720
rect 5302 1612 5374 1616
rect 5302 1560 5312 1612
rect 5364 1560 5374 1612
rect 5302 1556 5374 1560
rect 4926 1443 5238 1503
rect 4926 1336 4986 1443
rect 4668 952 4728 1042
rect 4662 948 4734 952
rect 4662 896 4672 948
rect 4724 896 4734 948
rect 4662 892 4734 896
rect 4794 836 4854 1157
rect 4794 784 4798 836
rect 4850 784 4854 836
rect 4794 774 4854 784
rect 4926 956 4986 1042
rect 5054 956 5114 1443
rect 5178 1332 5238 1443
rect 5308 1238 5368 1556
rect 5568 1248 5628 1720
rect 5958 1497 6018 1720
rect 6086 1497 6146 1720
rect 6218 1497 6278 1720
rect 5958 1437 6278 1497
rect 5958 1334 6018 1437
rect 5182 956 5242 1042
rect 4926 896 5242 956
rect 4926 724 4986 896
rect 5054 724 5114 896
rect 5182 724 5242 896
rect 5440 950 5500 1046
rect 5700 950 5760 1040
rect 5826 950 5886 1140
rect 5440 890 5886 950
rect 5956 950 6016 1044
rect 6086 950 6146 1437
rect 6218 1336 6278 1437
rect 6340 1490 6412 1494
rect 6340 1438 6350 1490
rect 6402 1438 6412 1490
rect 6340 1434 6412 1438
rect 6210 950 6270 1042
rect 5956 890 6270 950
rect 5700 834 5760 890
rect 5700 782 5704 834
rect 5756 782 5760 834
rect 5700 772 5760 782
rect 5956 724 6016 890
rect 6086 724 6146 890
rect 6210 724 6270 890
rect 6346 948 6406 1434
rect 6472 948 6532 1049
rect 6346 888 6532 948
rect 6602 724 6662 1720
rect 6988 1496 7048 1720
rect 7118 1496 7178 1720
rect 6988 1436 7178 1496
rect 6988 1336 7048 1436
rect 6736 948 6796 1045
rect 6864 948 6924 1148
rect 6736 888 6924 948
rect 6864 836 6924 888
rect 6988 952 7048 1044
rect 7118 952 7178 1436
rect 6988 892 7178 952
rect 6858 832 6930 836
rect 6858 780 6868 832
rect 6920 780 6930 832
rect 6858 776 6930 780
rect 6988 724 7048 892
rect 7118 724 7178 892
rect 10916 1707 11028 1745
rect 10916 1673 10955 1707
rect 10989 1673 11028 1707
rect 10916 1635 11028 1673
rect 10916 1601 10955 1635
rect 10989 1601 11028 1635
rect 10916 1563 11028 1601
rect 10916 1529 10955 1563
rect 10989 1529 11028 1563
rect 10916 1491 11028 1529
rect 10916 1457 10955 1491
rect 10989 1457 11028 1491
rect 10916 1419 11028 1457
rect 10916 1385 10955 1419
rect 10989 1385 11028 1419
rect 10916 1347 11028 1385
rect 10916 1313 10955 1347
rect 10989 1313 11028 1347
rect 10916 1275 11028 1313
rect 10916 1241 10955 1275
rect 10989 1241 11028 1275
rect 10916 1203 11028 1241
rect 10916 1169 10955 1203
rect 10989 1169 11028 1203
rect 10916 1131 11028 1169
rect 10916 1097 10955 1131
rect 10989 1097 11028 1131
rect 10916 1059 11028 1097
rect 10916 1025 10955 1059
rect 10989 1025 11028 1059
rect 10916 987 11028 1025
rect 10916 953 10955 987
rect 10989 953 11028 987
rect 10916 915 11028 953
rect 10916 881 10955 915
rect 10989 881 11028 915
rect 10916 843 11028 881
rect 10916 809 10955 843
rect 10989 809 11028 843
rect 10916 724 11028 809
rect -328 685 11028 724
rect -328 651 -211 685
rect -177 651 -139 685
rect -105 651 -67 685
rect -33 651 5 685
rect 39 651 77 685
rect 111 651 149 685
rect 183 651 221 685
rect 255 651 293 685
rect 327 651 365 685
rect 399 651 437 685
rect 471 651 509 685
rect 543 651 581 685
rect 615 651 653 685
rect 687 651 725 685
rect 759 651 797 685
rect 831 651 869 685
rect 903 651 941 685
rect 975 651 1013 685
rect 1047 651 1085 685
rect 1119 651 1157 685
rect 1191 651 1229 685
rect 1263 651 1301 685
rect 1335 651 1373 685
rect 1407 651 1445 685
rect 1479 651 1517 685
rect 1551 651 1589 685
rect 1623 651 1661 685
rect 1695 651 1733 685
rect 1767 651 1805 685
rect 1839 651 1877 685
rect 1911 651 1949 685
rect 1983 651 2021 685
rect 2055 651 2093 685
rect 2127 651 2165 685
rect 2199 651 2237 685
rect 2271 651 2309 685
rect 2343 651 2381 685
rect 2415 651 2453 685
rect 2487 651 2525 685
rect 2559 651 2597 685
rect 2631 651 2669 685
rect 2703 651 2741 685
rect 2775 651 2813 685
rect 2847 651 2885 685
rect 2919 651 2957 685
rect 2991 651 3029 685
rect 3063 651 3101 685
rect 3135 651 3173 685
rect 3207 651 3245 685
rect 3279 651 3317 685
rect 3351 651 3389 685
rect 3423 651 3461 685
rect 3495 651 3533 685
rect 3567 651 3605 685
rect 3639 651 3677 685
rect 3711 651 3749 685
rect 3783 651 3821 685
rect 3855 651 3893 685
rect 3927 651 3965 685
rect 3999 651 4037 685
rect 4071 651 4109 685
rect 4143 651 4181 685
rect 4215 651 4253 685
rect 4287 651 4325 685
rect 4359 651 4397 685
rect 4431 651 4469 685
rect 4503 651 4541 685
rect 4575 651 4613 685
rect 4647 651 4685 685
rect 4719 651 4757 685
rect 4791 651 4829 685
rect 4863 651 4901 685
rect 4935 651 4973 685
rect 5007 651 5045 685
rect 5079 651 5117 685
rect 5151 651 5189 685
rect 5223 651 5261 685
rect 5295 651 5333 685
rect 5367 651 5405 685
rect 5439 651 5477 685
rect 5511 651 5549 685
rect 5583 651 5621 685
rect 5655 651 5693 685
rect 5727 651 5765 685
rect 5799 651 5837 685
rect 5871 651 5909 685
rect 5943 651 5981 685
rect 6015 651 6053 685
rect 6087 651 6125 685
rect 6159 651 6197 685
rect 6231 651 6269 685
rect 6303 651 6341 685
rect 6375 651 6413 685
rect 6447 651 6485 685
rect 6519 651 6557 685
rect 6591 651 6629 685
rect 6663 651 6701 685
rect 6735 651 6773 685
rect 6807 651 6845 685
rect 6879 651 6917 685
rect 6951 651 6989 685
rect 7023 651 7061 685
rect 7095 651 7133 685
rect 7167 651 7205 685
rect 7239 651 7277 685
rect 7311 651 7349 685
rect 7383 651 7421 685
rect 7455 651 7493 685
rect 7527 651 7565 685
rect 7599 651 7637 685
rect 7671 651 7709 685
rect 7743 651 7781 685
rect 7815 651 7853 685
rect 7887 651 7925 685
rect 7959 651 7997 685
rect 8031 651 8069 685
rect 8103 651 8141 685
rect 8175 651 8213 685
rect 8247 651 8285 685
rect 8319 651 8357 685
rect 8391 651 8429 685
rect 8463 651 8501 685
rect 8535 651 8573 685
rect 8607 651 8645 685
rect 8679 651 8717 685
rect 8751 651 8789 685
rect 8823 651 8861 685
rect 8895 651 8933 685
rect 8967 651 9005 685
rect 9039 651 9077 685
rect 9111 651 9149 685
rect 9183 651 9221 685
rect 9255 651 9293 685
rect 9327 651 9365 685
rect 9399 651 9437 685
rect 9471 651 9509 685
rect 9543 651 9581 685
rect 9615 651 9653 685
rect 9687 651 9725 685
rect 9759 651 9797 685
rect 9831 651 9869 685
rect 9903 651 9941 685
rect 9975 651 10013 685
rect 10047 651 10085 685
rect 10119 651 10157 685
rect 10191 651 10229 685
rect 10263 651 10301 685
rect 10335 651 10373 685
rect 10407 651 10445 685
rect 10479 651 10517 685
rect 10551 651 10589 685
rect 10623 651 10661 685
rect 10695 651 10733 685
rect 10767 651 10805 685
rect 10839 651 10877 685
rect 10911 651 11028 685
rect -328 612 11028 651
rect 3052 524 3112 530
rect 5700 524 5760 530
rect 8088 524 8148 530
rect 3052 520 8148 524
rect 3052 468 3056 520
rect 3108 468 5704 520
rect 5756 468 8092 520
rect 8144 468 8148 520
rect 3052 464 8148 468
rect 3052 458 3112 464
rect 5700 458 5760 464
rect 8088 458 8148 464
rect -328 349 11028 388
rect -328 315 -211 349
rect -177 315 -139 349
rect -105 315 -67 349
rect -33 315 5 349
rect 39 315 77 349
rect 111 315 149 349
rect 183 315 221 349
rect 255 315 293 349
rect 327 315 365 349
rect 399 315 437 349
rect 471 315 509 349
rect 543 315 581 349
rect 615 315 653 349
rect 687 315 725 349
rect 759 315 797 349
rect 831 315 869 349
rect 903 315 941 349
rect 975 315 1013 349
rect 1047 315 1085 349
rect 1119 315 1157 349
rect 1191 315 1229 349
rect 1263 315 1301 349
rect 1335 315 1373 349
rect 1407 315 1445 349
rect 1479 315 1517 349
rect 1551 315 1589 349
rect 1623 315 1661 349
rect 1695 315 1733 349
rect 1767 315 1805 349
rect 1839 315 1877 349
rect 1911 315 1949 349
rect 1983 315 2021 349
rect 2055 315 2093 349
rect 2127 315 2165 349
rect 2199 315 2237 349
rect 2271 315 2309 349
rect 2343 315 2381 349
rect 2415 315 2453 349
rect 2487 315 2525 349
rect 2559 315 2597 349
rect 2631 315 2669 349
rect 2703 315 2741 349
rect 2775 315 2813 349
rect 2847 315 2885 349
rect 2919 315 2957 349
rect 2991 315 3029 349
rect 3063 315 3101 349
rect 3135 315 3173 349
rect 3207 315 3245 349
rect 3279 315 3317 349
rect 3351 315 3389 349
rect 3423 315 3461 349
rect 3495 315 3533 349
rect 3567 315 3605 349
rect 3639 315 3677 349
rect 3711 315 3749 349
rect 3783 315 3821 349
rect 3855 315 3893 349
rect 3927 315 3965 349
rect 3999 315 4037 349
rect 4071 315 4109 349
rect 4143 315 4181 349
rect 4215 315 4253 349
rect 4287 315 4325 349
rect 4359 315 4397 349
rect 4431 315 4469 349
rect 4503 315 4541 349
rect 4575 315 4613 349
rect 4647 315 4685 349
rect 4719 315 4757 349
rect 4791 315 4829 349
rect 4863 315 4901 349
rect 4935 315 4973 349
rect 5007 315 5045 349
rect 5079 315 5117 349
rect 5151 315 5189 349
rect 5223 315 5261 349
rect 5295 315 5333 349
rect 5367 315 5405 349
rect 5439 315 5477 349
rect 5511 315 5549 349
rect 5583 315 5621 349
rect 5655 315 5693 349
rect 5727 315 5765 349
rect 5799 315 5837 349
rect 5871 315 5909 349
rect 5943 315 5981 349
rect 6015 315 6053 349
rect 6087 315 6125 349
rect 6159 315 6197 349
rect 6231 315 6269 349
rect 6303 315 6341 349
rect 6375 315 6413 349
rect 6447 315 6485 349
rect 6519 315 6557 349
rect 6591 315 6629 349
rect 6663 315 6701 349
rect 6735 315 6773 349
rect 6807 315 6845 349
rect 6879 315 6917 349
rect 6951 315 6989 349
rect 7023 315 7061 349
rect 7095 315 7133 349
rect 7167 315 7205 349
rect 7239 315 7277 349
rect 7311 315 7349 349
rect 7383 315 7421 349
rect 7455 315 7493 349
rect 7527 315 7565 349
rect 7599 315 7637 349
rect 7671 315 7709 349
rect 7743 315 7781 349
rect 7815 315 7853 349
rect 7887 315 7925 349
rect 7959 315 7997 349
rect 8031 315 8069 349
rect 8103 315 8141 349
rect 8175 315 8213 349
rect 8247 315 8285 349
rect 8319 315 8357 349
rect 8391 315 8429 349
rect 8463 315 8501 349
rect 8535 315 8573 349
rect 8607 315 8645 349
rect 8679 315 8717 349
rect 8751 315 8789 349
rect 8823 315 8861 349
rect 8895 315 8933 349
rect 8967 315 9005 349
rect 9039 315 9077 349
rect 9111 315 9149 349
rect 9183 315 9221 349
rect 9255 315 9293 349
rect 9327 315 9365 349
rect 9399 315 9437 349
rect 9471 315 9509 349
rect 9543 315 9581 349
rect 9615 315 9653 349
rect 9687 315 9725 349
rect 9759 315 9797 349
rect 9831 315 9869 349
rect 9903 315 9941 349
rect 9975 315 10013 349
rect 10047 315 10085 349
rect 10119 315 10157 349
rect 10191 315 10229 349
rect 10263 315 10301 349
rect 10335 315 10373 349
rect 10407 315 10445 349
rect 10479 315 10517 349
rect 10551 315 10589 349
rect 10623 315 10661 349
rect 10695 315 10733 349
rect 10767 315 10805 349
rect 10839 315 10877 349
rect 10911 315 11028 349
rect -328 276 11028 315
rect -328 101 -216 276
rect -328 67 -289 101
rect -255 67 -216 101
rect -328 29 -216 67
rect -328 -5 -289 29
rect -255 4 -216 29
rect 726 4 786 276
rect 852 4 912 276
rect 1488 226 1560 230
rect 1488 174 1498 226
rect 1550 174 1560 226
rect 1488 170 1560 174
rect 2524 226 2596 230
rect 2524 174 2534 226
rect 2586 174 2596 226
rect 2524 170 2596 174
rect 974 110 1046 114
rect 974 58 984 110
rect 1036 58 1046 110
rect 974 54 1046 58
rect -255 -5 912 4
rect -328 -43 912 -5
rect -328 -77 -289 -43
rect -255 -56 912 -43
rect -255 -77 -216 -56
rect -328 -115 -216 -77
rect -328 -149 -289 -115
rect -255 -149 -216 -115
rect -328 -187 -216 -149
rect -328 -221 -289 -187
rect -255 -221 -216 -187
rect -328 -259 -216 -221
rect -328 -293 -289 -259
rect -255 -293 -216 -259
rect -328 -331 -216 -293
rect -328 -365 -289 -331
rect -255 -365 -216 -331
rect -328 -403 -216 -365
rect -328 -437 -289 -403
rect -255 -437 -216 -403
rect -328 -475 -216 -437
rect -328 -509 -289 -475
rect -255 -509 -216 -475
rect -328 -547 -216 -509
rect -328 -581 -289 -547
rect -255 -581 -216 -547
rect -328 -619 -216 -581
rect -328 -653 -289 -619
rect -255 -653 -216 -619
rect -328 -691 -216 -653
rect -328 -725 -289 -691
rect -255 -725 -216 -691
rect -328 -728 -216 -725
rect 726 -728 786 -56
rect 852 -140 912 -56
rect 980 -240 1040 54
rect 1364 0 1436 4
rect 1364 -52 1374 0
rect 1426 -52 1436 0
rect 1364 -56 1436 -52
rect 1370 -146 1430 -56
rect 1494 -236 1554 170
rect 2006 110 2078 114
rect 2006 58 2016 110
rect 2068 58 2078 110
rect 2006 54 2078 58
rect 1618 0 1690 4
rect 1618 -52 1628 0
rect 1680 -52 1690 0
rect 1618 -56 1690 -52
rect 1624 -142 1684 -56
rect 2012 -250 2072 54
rect 2390 0 2462 4
rect 2390 -52 2400 0
rect 2452 -52 2462 0
rect 2390 -56 2462 -52
rect 2396 -150 2456 -56
rect 2530 -240 2590 170
rect 3042 110 3114 114
rect 3042 58 3052 110
rect 3104 58 3114 110
rect 3042 54 3114 58
rect 2652 0 2724 4
rect 2652 -52 2662 0
rect 2714 -52 2724 0
rect 2652 -56 2724 -52
rect 2658 -142 2718 -56
rect 3048 -246 3108 54
rect 3172 4 3232 276
rect 3306 4 3366 276
rect 4022 4 4082 276
rect 4146 4 4206 276
rect 4784 232 4856 236
rect 4784 180 4794 232
rect 4846 180 4856 232
rect 4784 176 4856 180
rect 5820 232 5892 236
rect 5820 180 5830 232
rect 5882 180 5892 232
rect 5820 176 5892 180
rect 4270 116 4342 120
rect 4270 64 4280 116
rect 4332 64 4342 116
rect 4270 60 4342 64
rect 3172 -56 4206 4
rect 3172 -138 3232 -56
rect 852 -728 912 -622
rect 1110 -726 1170 -618
rect -328 -763 912 -728
rect -328 -797 -289 -763
rect -255 -788 912 -763
rect 1104 -730 1176 -726
rect 1104 -782 1114 -730
rect 1166 -782 1176 -730
rect 1104 -786 1176 -782
rect -255 -797 -216 -788
rect -328 -835 -216 -797
rect -328 -869 -289 -835
rect -255 -869 -216 -835
rect -328 -907 -216 -869
rect 26 -840 98 -836
rect 26 -892 36 -840
rect 88 -892 98 -840
rect 26 -896 98 -892
rect -328 -941 -289 -907
rect -255 -941 -216 -907
rect -328 -979 -216 -941
rect -328 -1013 -289 -979
rect -255 -1013 -216 -979
rect -328 -1051 -216 -1013
rect -328 -1085 -289 -1051
rect -255 -1085 -216 -1051
rect -328 -1123 -216 -1085
rect -328 -1157 -289 -1123
rect -255 -1157 -216 -1123
rect -328 -1195 -216 -1157
rect -328 -1229 -289 -1195
rect -255 -1229 -216 -1195
rect -328 -1267 -216 -1229
rect -328 -1301 -289 -1267
rect -255 -1301 -216 -1267
rect -328 -1339 -216 -1301
rect -328 -1373 -289 -1339
rect -255 -1373 -216 -1339
rect -328 -1411 -216 -1373
rect -328 -1445 -289 -1411
rect -255 -1445 -216 -1411
rect -328 -1483 -216 -1445
rect -328 -1517 -289 -1483
rect -255 -1517 -216 -1483
rect -328 -1555 -216 -1517
rect -328 -1589 -289 -1555
rect -255 -1589 -216 -1555
rect -328 -1627 -216 -1589
rect -328 -1661 -289 -1627
rect -255 -1661 -216 -1627
rect -328 -1699 -216 -1661
rect -328 -1733 -289 -1699
rect -255 -1733 -216 -1699
rect -328 -1771 -216 -1733
rect -328 -1805 -289 -1771
rect -255 -1805 -216 -1771
rect -328 -1843 -216 -1805
rect -328 -1877 -289 -1843
rect -255 -1877 -216 -1843
rect -328 -1915 -216 -1877
rect -328 -1949 -289 -1915
rect -255 -1949 -216 -1915
rect -328 -1987 -216 -1949
rect -328 -2021 -289 -1987
rect -255 -2021 -216 -1987
rect -328 -2059 -216 -2021
rect -328 -2093 -289 -2059
rect -255 -2093 -216 -2059
rect -328 -2131 -216 -2093
rect -328 -2165 -289 -2131
rect -255 -2165 -216 -2131
rect -328 -2203 -216 -2165
rect 32 -2170 92 -896
rect 172 -1082 232 -788
rect 1240 -840 1300 -546
rect 1752 -836 1812 -546
rect 1886 -726 1946 -622
rect 2140 -726 2200 -620
rect 1880 -730 1952 -726
rect 1880 -782 1890 -730
rect 1942 -782 1952 -730
rect 1880 -786 1952 -782
rect 2134 -730 2206 -726
rect 2134 -782 2144 -730
rect 2196 -782 2206 -730
rect 2134 -786 2206 -782
rect 2272 -836 2332 -542
rect 2788 -836 2848 -542
rect 2918 -726 2978 -622
rect 2912 -730 2984 -726
rect 2912 -782 2922 -730
rect 2974 -782 2984 -730
rect 2912 -786 2984 -782
rect 3172 -728 3232 -616
rect 3306 -728 3366 -56
rect 4022 -728 4082 -56
rect 4146 -144 4206 -56
rect 4276 -234 4336 60
rect 4660 6 4732 10
rect 4660 -46 4670 6
rect 4722 -46 4732 6
rect 4660 -50 4732 -46
rect 4666 -140 4726 -50
rect 4790 -230 4850 176
rect 5302 116 5374 120
rect 5302 64 5312 116
rect 5364 64 5374 116
rect 5302 60 5374 64
rect 4914 6 4986 10
rect 4914 -46 4924 6
rect 4976 -46 4986 6
rect 4914 -50 4986 -46
rect 4920 -136 4980 -50
rect 5308 -244 5368 60
rect 5686 6 5758 10
rect 5686 -46 5696 6
rect 5748 -46 5758 6
rect 5686 -50 5758 -46
rect 5692 -144 5752 -50
rect 5826 -234 5886 176
rect 6338 116 6410 120
rect 6338 64 6348 116
rect 6400 64 6410 116
rect 6338 60 6410 64
rect 5948 6 6020 10
rect 5948 -46 5958 6
rect 6010 -46 6020 6
rect 5948 -50 6020 -46
rect 5954 -136 6014 -50
rect 6344 -240 6404 60
rect 6470 10 6530 276
rect 6602 10 6662 276
rect 7318 10 7378 276
rect 7442 10 7502 276
rect 8080 226 8152 230
rect 8080 174 8090 226
rect 8142 174 8152 226
rect 8080 170 8152 174
rect 9116 226 9188 230
rect 9116 174 9126 226
rect 9178 174 9188 226
rect 9116 170 9188 174
rect 7566 110 7638 114
rect 7566 58 7576 110
rect 7628 58 7638 110
rect 7566 54 7638 58
rect 6470 -50 7502 10
rect 6470 -144 6530 -50
rect 4148 -728 4208 -616
rect 4406 -720 4466 -612
rect 1240 -892 1244 -840
rect 1296 -892 1300 -840
rect 1240 -902 1300 -892
rect 1746 -840 1818 -836
rect 1746 -892 1756 -840
rect 1808 -892 1818 -840
rect 1746 -896 1818 -892
rect 2266 -840 2338 -836
rect 2266 -892 2276 -840
rect 2328 -892 2338 -840
rect 2266 -896 2338 -892
rect 2782 -840 2854 -836
rect 2782 -892 2792 -840
rect 2844 -892 2854 -840
rect 2782 -896 2854 -892
rect 2918 -958 2978 -786
rect 3172 -788 4208 -728
rect 4400 -724 4472 -720
rect 4400 -776 4410 -724
rect 4462 -776 4472 -724
rect 4400 -780 4472 -776
rect 2912 -962 2984 -958
rect 2912 -1014 2922 -962
rect 2974 -1014 2984 -962
rect 2912 -1018 2984 -1014
rect 172 -1142 654 -1082
rect 1024 -1086 1096 -1082
rect 1024 -1138 1034 -1086
rect 1086 -1138 1096 -1086
rect 1024 -1142 1096 -1138
rect 172 -1632 232 -1142
rect 594 -1246 654 -1142
rect 1030 -1336 1090 -1142
rect 596 -1632 656 -1524
rect 1456 -1626 1516 -1524
rect 172 -1692 656 -1632
rect 1026 -1630 1516 -1626
rect 1026 -1682 1036 -1630
rect 1088 -1682 1516 -1630
rect 1026 -1686 1516 -1682
rect 172 -2162 232 -1692
rect 596 -1792 656 -1692
rect 1032 -1890 1092 -1686
rect 1456 -1786 1516 -1686
rect 592 -2162 652 -2070
rect -328 -2237 -289 -2203
rect -255 -2237 -216 -2203
rect 26 -2174 98 -2170
rect 26 -2226 36 -2174
rect 88 -2226 98 -2174
rect 26 -2230 98 -2226
rect 172 -2222 652 -2162
rect -328 -2275 -216 -2237
rect -328 -2309 -289 -2275
rect -255 -2309 -216 -2275
rect -328 -2347 -216 -2309
rect 172 -2336 232 -2222
rect 592 -2336 652 -2222
rect 1890 -2336 1950 -1394
rect 2314 -1626 2374 -1520
rect 2748 -1626 2808 -1424
rect 2308 -1628 2380 -1626
rect 2308 -1680 2318 -1628
rect 2370 -1680 2380 -1628
rect 2308 -1686 2380 -1680
rect 2742 -1630 2814 -1626
rect 2742 -1682 2752 -1630
rect 2804 -1682 2814 -1630
rect 2742 -1686 2814 -1682
rect 3178 -1628 3238 -1520
rect 3178 -1680 3182 -1628
rect 3234 -1680 3238 -1628
rect 2314 -1788 2374 -1686
rect 2748 -1866 2808 -1686
rect 3178 -1788 3238 -1680
rect 3606 -2336 3666 -788
rect 4536 -834 4596 -540
rect 4536 -886 4540 -834
rect 4592 -886 4596 -834
rect 4536 -1082 4596 -886
rect 4798 -958 4858 -478
rect 5048 -830 5108 -540
rect 5182 -720 5242 -616
rect 5436 -720 5496 -614
rect 5176 -724 5248 -720
rect 5176 -776 5186 -724
rect 5238 -776 5248 -724
rect 5176 -780 5248 -776
rect 5430 -724 5502 -720
rect 5430 -776 5440 -724
rect 5492 -776 5502 -724
rect 5430 -780 5502 -776
rect 5568 -830 5628 -536
rect 6084 -830 6144 -536
rect 6214 -720 6274 -616
rect 6208 -724 6280 -720
rect 6208 -776 6218 -724
rect 6270 -776 6280 -724
rect 6208 -780 6280 -776
rect 6468 -722 6528 -610
rect 6602 -722 6662 -50
rect 7318 -722 7378 -50
rect 7442 -140 7502 -50
rect 7572 -240 7632 54
rect 7956 0 8028 4
rect 7956 -52 7966 0
rect 8018 -52 8028 0
rect 7956 -56 8028 -52
rect 7962 -146 8022 -56
rect 8086 -236 8146 170
rect 8598 110 8670 114
rect 8598 58 8608 110
rect 8660 58 8670 110
rect 8598 54 8670 58
rect 8210 0 8282 4
rect 8210 -52 8220 0
rect 8272 -52 8282 0
rect 8210 -56 8282 -52
rect 8216 -142 8276 -56
rect 8604 -250 8664 54
rect 8982 0 9054 4
rect 8982 -52 8992 0
rect 9044 -52 9054 0
rect 8982 -56 9054 -52
rect 8988 -150 9048 -56
rect 9122 -240 9182 170
rect 9634 110 9706 114
rect 9634 58 9644 110
rect 9696 58 9706 110
rect 9634 54 9706 58
rect 9244 0 9316 4
rect 9244 -52 9254 0
rect 9306 -52 9316 0
rect 9244 -56 9316 -52
rect 9250 -142 9310 -56
rect 9640 -246 9700 54
rect 9766 2 9826 276
rect 9898 2 9958 276
rect 10916 101 11028 276
rect 10916 67 10955 101
rect 10989 67 11028 101
rect 10916 29 11028 67
rect 10916 2 10955 29
rect 9766 -5 10955 2
rect 10989 -5 11028 29
rect 9766 -43 11028 -5
rect 9766 -58 10955 -43
rect 9766 -140 9826 -58
rect 7444 -722 7504 -618
rect 6468 -782 7504 -722
rect 7702 -726 7762 -618
rect 7696 -730 7768 -726
rect 7696 -782 7706 -730
rect 7758 -782 7768 -730
rect 5042 -834 5114 -830
rect 5042 -886 5052 -834
rect 5104 -886 5114 -834
rect 5042 -890 5114 -886
rect 5562 -834 5634 -830
rect 5562 -886 5572 -834
rect 5624 -886 5634 -834
rect 5562 -890 5634 -886
rect 6078 -834 6150 -830
rect 6078 -886 6088 -834
rect 6140 -886 6150 -834
rect 6078 -890 6150 -886
rect 4792 -962 4864 -958
rect 4792 -1014 4802 -962
rect 4854 -1014 4864 -962
rect 4792 -1018 4864 -1014
rect 4458 -1086 4596 -1082
rect 4458 -1138 4468 -1086
rect 4520 -1138 4596 -1086
rect 4458 -1142 4596 -1138
rect 4894 -1140 5818 -1080
rect 4464 -1340 4524 -1142
rect 4894 -1248 4954 -1140
rect 4038 -1628 4098 -1520
rect 4896 -1624 4956 -1520
rect 5320 -1624 5380 -1140
rect 5758 -1248 5818 -1140
rect 5756 -1624 5816 -1520
rect 4038 -1680 4042 -1628
rect 4094 -1680 4098 -1628
rect 4038 -1788 4098 -1680
rect 4462 -1630 4534 -1626
rect 4462 -1682 4472 -1630
rect 4524 -1682 4534 -1630
rect 4462 -1686 4534 -1682
rect 4896 -1684 5816 -1624
rect 6184 -1626 6244 -1426
rect 6610 -1626 6670 -1520
rect 4468 -1890 4528 -1686
rect 4896 -1788 4956 -1684
rect 4894 -2168 4954 -2064
rect 5320 -2168 5380 -1684
rect 5756 -1788 5816 -1684
rect 6178 -1630 6250 -1626
rect 6178 -1682 6188 -1630
rect 6240 -1682 6250 -1630
rect 6178 -1686 6250 -1682
rect 6604 -1628 6676 -1626
rect 6604 -1680 6614 -1628
rect 6666 -1680 6676 -1628
rect 6604 -1686 6676 -1680
rect 6610 -1788 6670 -1686
rect 5756 -2168 5816 -2062
rect 4894 -2228 5816 -2168
rect 6180 -2170 6240 -1984
rect 4894 -2336 4954 -2228
rect 5320 -2336 5380 -2228
rect 5756 -2336 5816 -2228
rect 6174 -2174 6246 -2170
rect 6174 -2226 6184 -2174
rect 6236 -2226 6246 -2174
rect 6174 -2230 6246 -2226
rect 7038 -2336 7098 -782
rect 7696 -786 7768 -782
rect 7832 -836 7892 -546
rect 8344 -836 8404 -546
rect 8478 -726 8538 -622
rect 8732 -726 8792 -620
rect 8472 -730 8544 -726
rect 8472 -782 8482 -730
rect 8534 -782 8544 -730
rect 8472 -786 8544 -782
rect 8726 -730 8798 -726
rect 8726 -782 8736 -730
rect 8788 -782 8798 -730
rect 8726 -786 8798 -782
rect 8864 -836 8924 -542
rect 9380 -836 9440 -542
rect 9510 -726 9570 -622
rect 9504 -730 9576 -726
rect 9504 -782 9514 -730
rect 9566 -782 9576 -730
rect 9504 -786 9576 -782
rect 9764 -728 9824 -616
rect 9898 -728 9958 -58
rect 10916 -77 10955 -58
rect 10989 -77 11028 -43
rect 10916 -115 11028 -77
rect 10916 -149 10955 -115
rect 10989 -149 11028 -115
rect 10916 -187 11028 -149
rect 10916 -221 10955 -187
rect 10989 -221 11028 -187
rect 10916 -259 11028 -221
rect 10916 -293 10955 -259
rect 10989 -293 11028 -259
rect 10916 -331 11028 -293
rect 10916 -365 10955 -331
rect 10989 -365 11028 -331
rect 10916 -403 11028 -365
rect 10916 -437 10955 -403
rect 10989 -437 11028 -403
rect 10916 -475 11028 -437
rect 10916 -509 10955 -475
rect 10989 -509 11028 -475
rect 10916 -547 11028 -509
rect 10916 -581 10955 -547
rect 10989 -581 11028 -547
rect 10916 -619 11028 -581
rect 10916 -653 10955 -619
rect 10989 -653 11028 -619
rect 10916 -691 11028 -653
rect 10916 -725 10955 -691
rect 10989 -725 11028 -691
rect 10916 -728 11028 -725
rect 9764 -763 11028 -728
rect 9764 -788 10955 -763
rect 7826 -840 7898 -836
rect 7826 -892 7836 -840
rect 7888 -892 7898 -840
rect 7826 -896 7898 -892
rect 8338 -840 8410 -836
rect 8338 -892 8348 -840
rect 8400 -892 8410 -840
rect 8338 -896 8410 -892
rect 8858 -840 8930 -836
rect 8858 -892 8868 -840
rect 8920 -892 8930 -840
rect 8858 -896 8930 -892
rect 9374 -840 9446 -836
rect 9374 -892 9384 -840
rect 9436 -892 9446 -840
rect 9374 -896 9446 -892
rect 9608 -970 9680 -966
rect 9608 -1022 9618 -970
rect 9670 -1022 9680 -970
rect 9608 -1026 9680 -1022
rect 9614 -1332 9674 -1026
rect 10044 -1096 10104 -788
rect 10468 -1096 10528 -788
rect 10916 -797 10955 -788
rect 10989 -797 11028 -763
rect 10916 -835 11028 -797
rect 10594 -840 10666 -836
rect 10594 -892 10604 -840
rect 10656 -892 10666 -840
rect 10594 -896 10666 -892
rect 10916 -869 10955 -835
rect 10989 -869 11028 -835
rect 10044 -1156 10528 -1096
rect 10044 -1246 10104 -1156
rect 7468 -1628 7528 -1520
rect 7896 -1626 7956 -1410
rect 7468 -1680 7472 -1628
rect 7524 -1680 7528 -1628
rect 7468 -1788 7528 -1680
rect 7890 -1630 7962 -1626
rect 7890 -1682 7900 -1630
rect 7952 -1682 7962 -1630
rect 7890 -1686 7962 -1682
rect 8322 -1628 8382 -1520
rect 8322 -1680 8326 -1628
rect 8378 -1680 8382 -1628
rect 7896 -1880 7956 -1686
rect 8322 -1788 8382 -1680
rect 8756 -2336 8816 -1418
rect 9186 -1620 9246 -1520
rect 9186 -1630 9248 -1620
rect 9186 -1682 9192 -1630
rect 9244 -1682 9248 -1630
rect 9186 -1692 9248 -1682
rect 10042 -1630 10102 -1520
rect 10468 -1630 10528 -1156
rect 10042 -1690 10528 -1630
rect 9186 -1788 9246 -1692
rect 10042 -1788 10102 -1690
rect 9612 -2164 9672 -1982
rect 10044 -2164 10104 -2066
rect 10468 -2164 10528 -1690
rect 10600 -2164 10660 -896
rect 10916 -907 11028 -869
rect 10916 -941 10955 -907
rect 10989 -941 11028 -907
rect 10916 -979 11028 -941
rect 10916 -1013 10955 -979
rect 10989 -1013 11028 -979
rect 10916 -1051 11028 -1013
rect 10916 -1085 10955 -1051
rect 10989 -1085 11028 -1051
rect 10916 -1123 11028 -1085
rect 10916 -1157 10955 -1123
rect 10989 -1157 11028 -1123
rect 10916 -1195 11028 -1157
rect 10916 -1229 10955 -1195
rect 10989 -1229 11028 -1195
rect 10916 -1267 11028 -1229
rect 10916 -1301 10955 -1267
rect 10989 -1301 11028 -1267
rect 10916 -1339 11028 -1301
rect 10916 -1373 10955 -1339
rect 10989 -1373 11028 -1339
rect 10916 -1411 11028 -1373
rect 10916 -1445 10955 -1411
rect 10989 -1445 11028 -1411
rect 10916 -1483 11028 -1445
rect 10916 -1517 10955 -1483
rect 10989 -1517 11028 -1483
rect 10916 -1555 11028 -1517
rect 10916 -1589 10955 -1555
rect 10989 -1589 11028 -1555
rect 10916 -1627 11028 -1589
rect 10916 -1661 10955 -1627
rect 10989 -1661 11028 -1627
rect 10916 -1699 11028 -1661
rect 10916 -1733 10955 -1699
rect 10989 -1733 11028 -1699
rect 10916 -1771 11028 -1733
rect 10916 -1805 10955 -1771
rect 10989 -1805 11028 -1771
rect 10916 -1843 11028 -1805
rect 10916 -1877 10955 -1843
rect 10989 -1877 11028 -1843
rect 10916 -1915 11028 -1877
rect 10916 -1949 10955 -1915
rect 10989 -1949 11028 -1915
rect 10916 -1987 11028 -1949
rect 10916 -2021 10955 -1987
rect 10989 -2021 11028 -1987
rect 10916 -2059 11028 -2021
rect 10916 -2093 10955 -2059
rect 10989 -2093 11028 -2059
rect 10916 -2131 11028 -2093
rect 9606 -2168 9678 -2164
rect 9606 -2220 9616 -2168
rect 9668 -2220 9678 -2168
rect 9606 -2224 9678 -2220
rect 10044 -2224 10528 -2164
rect 10594 -2168 10666 -2164
rect 10594 -2220 10604 -2168
rect 10656 -2220 10666 -2168
rect 10594 -2224 10666 -2220
rect 10916 -2165 10955 -2131
rect 10989 -2165 11028 -2131
rect 10916 -2203 11028 -2165
rect 10044 -2336 10104 -2224
rect 10468 -2336 10528 -2224
rect 10916 -2237 10955 -2203
rect 10989 -2237 11028 -2203
rect 10916 -2275 11028 -2237
rect 10916 -2309 10955 -2275
rect 10989 -2309 11028 -2275
rect -328 -2381 -289 -2347
rect -255 -2381 -216 -2347
rect -328 -2419 -216 -2381
rect -328 -2453 -289 -2419
rect -255 -2453 -216 -2419
rect -328 -2491 -216 -2453
rect -328 -2525 -289 -2491
rect -255 -2525 -216 -2491
rect -328 -2563 -216 -2525
rect -66 -2413 10708 -2336
rect -66 -2465 18 -2413
rect 70 -2465 82 -2413
rect 134 -2465 146 -2413
rect 198 -2465 210 -2413
rect 262 -2465 274 -2413
rect 326 -2465 338 -2413
rect 390 -2465 402 -2413
rect 454 -2465 466 -2413
rect 518 -2465 530 -2413
rect 582 -2465 594 -2413
rect 646 -2465 658 -2413
rect 710 -2465 722 -2413
rect 774 -2465 786 -2413
rect 838 -2465 850 -2413
rect 902 -2465 914 -2413
rect 966 -2465 978 -2413
rect 1030 -2465 1042 -2413
rect 1094 -2465 1106 -2413
rect 1158 -2465 1170 -2413
rect 1222 -2465 1234 -2413
rect 1286 -2465 1298 -2413
rect 1350 -2465 1362 -2413
rect 1414 -2465 1426 -2413
rect 1478 -2465 1490 -2413
rect 1542 -2465 1554 -2413
rect 1606 -2465 1618 -2413
rect 1670 -2465 1682 -2413
rect 1734 -2465 1746 -2413
rect 1798 -2465 1810 -2413
rect 1862 -2465 1874 -2413
rect 1926 -2465 1938 -2413
rect 1990 -2465 2002 -2413
rect 2054 -2465 2066 -2413
rect 2118 -2465 2130 -2413
rect 2182 -2465 2194 -2413
rect 2246 -2465 2258 -2413
rect 2310 -2465 2322 -2413
rect 2374 -2465 2386 -2413
rect 2438 -2465 2450 -2413
rect 2502 -2465 2514 -2413
rect 2566 -2465 2578 -2413
rect 2630 -2465 2642 -2413
rect 2694 -2465 2706 -2413
rect 2758 -2465 2770 -2413
rect 2822 -2465 2834 -2413
rect 2886 -2465 2898 -2413
rect 2950 -2465 2962 -2413
rect 3014 -2465 3026 -2413
rect 3078 -2465 3090 -2413
rect 3142 -2465 3154 -2413
rect 3206 -2465 3218 -2413
rect 3270 -2465 3282 -2413
rect 3334 -2465 3346 -2413
rect 3398 -2465 3410 -2413
rect 3462 -2465 3474 -2413
rect 3526 -2465 3538 -2413
rect 3590 -2465 3602 -2413
rect 3654 -2465 3666 -2413
rect 3718 -2465 3730 -2413
rect 3782 -2465 3794 -2413
rect 3846 -2465 3858 -2413
rect 3910 -2465 3922 -2413
rect 3974 -2465 3986 -2413
rect 4038 -2465 4050 -2413
rect 4102 -2465 4114 -2413
rect 4166 -2465 4178 -2413
rect 4230 -2465 4242 -2413
rect 4294 -2465 4306 -2413
rect 4358 -2465 4370 -2413
rect 4422 -2465 4434 -2413
rect 4486 -2465 4498 -2413
rect 4550 -2465 4562 -2413
rect 4614 -2465 4626 -2413
rect 4678 -2465 4690 -2413
rect 4742 -2465 4754 -2413
rect 4806 -2465 4818 -2413
rect 4870 -2465 4882 -2413
rect 4934 -2465 4946 -2413
rect 4998 -2465 5010 -2413
rect 5062 -2465 5074 -2413
rect 5126 -2465 5138 -2413
rect 5190 -2465 5202 -2413
rect 5254 -2465 5266 -2413
rect 5318 -2465 5330 -2413
rect 5382 -2465 5394 -2413
rect 5446 -2465 5458 -2413
rect 5510 -2465 5522 -2413
rect 5574 -2465 5586 -2413
rect 5638 -2465 5650 -2413
rect 5702 -2465 5714 -2413
rect 5766 -2465 5778 -2413
rect 5830 -2465 5842 -2413
rect 5894 -2465 5906 -2413
rect 5958 -2465 5970 -2413
rect 6022 -2465 6034 -2413
rect 6086 -2465 6098 -2413
rect 6150 -2465 6162 -2413
rect 6214 -2465 6226 -2413
rect 6278 -2465 6290 -2413
rect 6342 -2465 6354 -2413
rect 6406 -2465 6418 -2413
rect 6470 -2465 6482 -2413
rect 6534 -2465 6546 -2413
rect 6598 -2465 6610 -2413
rect 6662 -2465 6674 -2413
rect 6726 -2465 6738 -2413
rect 6790 -2465 6802 -2413
rect 6854 -2465 6866 -2413
rect 6918 -2465 6930 -2413
rect 6982 -2465 6994 -2413
rect 7046 -2465 7058 -2413
rect 7110 -2465 7122 -2413
rect 7174 -2465 7186 -2413
rect 7238 -2465 7250 -2413
rect 7302 -2465 7314 -2413
rect 7366 -2465 7378 -2413
rect 7430 -2465 7442 -2413
rect 7494 -2465 7506 -2413
rect 7558 -2465 7570 -2413
rect 7622 -2465 7634 -2413
rect 7686 -2465 7698 -2413
rect 7750 -2465 7762 -2413
rect 7814 -2465 7826 -2413
rect 7878 -2465 7890 -2413
rect 7942 -2465 7954 -2413
rect 8006 -2465 8018 -2413
rect 8070 -2465 8082 -2413
rect 8134 -2465 8146 -2413
rect 8198 -2465 8210 -2413
rect 8262 -2465 8274 -2413
rect 8326 -2465 8338 -2413
rect 8390 -2465 8402 -2413
rect 8454 -2465 8466 -2413
rect 8518 -2465 8530 -2413
rect 8582 -2465 8594 -2413
rect 8646 -2465 8658 -2413
rect 8710 -2465 8722 -2413
rect 8774 -2465 8786 -2413
rect 8838 -2465 8850 -2413
rect 8902 -2465 8914 -2413
rect 8966 -2465 8978 -2413
rect 9030 -2465 9042 -2413
rect 9094 -2465 9106 -2413
rect 9158 -2465 9170 -2413
rect 9222 -2465 9234 -2413
rect 9286 -2465 9298 -2413
rect 9350 -2465 9362 -2413
rect 9414 -2465 9426 -2413
rect 9478 -2465 9490 -2413
rect 9542 -2465 9554 -2413
rect 9606 -2465 9618 -2413
rect 9670 -2465 9682 -2413
rect 9734 -2465 9746 -2413
rect 9798 -2465 9810 -2413
rect 9862 -2465 9874 -2413
rect 9926 -2465 9938 -2413
rect 9990 -2465 10002 -2413
rect 10054 -2465 10066 -2413
rect 10118 -2465 10130 -2413
rect 10182 -2465 10194 -2413
rect 10246 -2465 10258 -2413
rect 10310 -2465 10322 -2413
rect 10374 -2465 10386 -2413
rect 10438 -2465 10450 -2413
rect 10502 -2465 10514 -2413
rect 10566 -2465 10578 -2413
rect 10630 -2465 10708 -2413
rect -66 -2550 10708 -2465
rect 10916 -2347 11028 -2309
rect 10916 -2381 10955 -2347
rect 10989 -2381 11028 -2347
rect 10916 -2419 11028 -2381
rect 10916 -2453 10955 -2419
rect 10989 -2453 11028 -2419
rect 10916 -2491 11028 -2453
rect 10916 -2525 10955 -2491
rect 10989 -2525 11028 -2491
rect -328 -2597 -289 -2563
rect -255 -2597 -216 -2563
rect -328 -2616 -216 -2597
rect 10916 -2563 11028 -2525
rect 10916 -2597 10955 -2563
rect 10989 -2597 11028 -2563
rect 10916 -2616 11028 -2597
rect -328 -2635 394 -2616
rect -328 -2669 -289 -2635
rect -255 -2644 394 -2635
rect -255 -2669 -198 -2644
rect -328 -2707 -198 -2669
rect -328 -2741 -289 -2707
rect -255 -2741 -198 -2707
rect -328 -2888 -198 -2741
rect 366 -2888 394 -2644
rect -328 -2916 394 -2888
rect 10306 -2635 11028 -2616
rect 10306 -2644 10955 -2635
rect 10306 -2888 10334 -2644
rect 10898 -2669 10955 -2644
rect 10989 -2669 11028 -2635
rect 10898 -2707 11028 -2669
rect 10898 -2741 10955 -2707
rect 10989 -2741 11028 -2707
rect 10898 -2888 11028 -2741
rect 10306 -2916 11028 -2888
rect -328 -2955 11028 -2916
rect -328 -2989 -211 -2955
rect -177 -2989 -139 -2955
rect -105 -2989 -67 -2955
rect -33 -2989 5 -2955
rect 39 -2989 77 -2955
rect 111 -2989 149 -2955
rect 183 -2989 221 -2955
rect 255 -2989 293 -2955
rect 327 -2989 365 -2955
rect 399 -2989 437 -2955
rect 471 -2989 509 -2955
rect 543 -2989 581 -2955
rect 615 -2989 653 -2955
rect 687 -2989 725 -2955
rect 759 -2989 797 -2955
rect 831 -2989 869 -2955
rect 903 -2989 941 -2955
rect 975 -2989 1013 -2955
rect 1047 -2989 1085 -2955
rect 1119 -2989 1157 -2955
rect 1191 -2989 1229 -2955
rect 1263 -2989 1301 -2955
rect 1335 -2989 1373 -2955
rect 1407 -2989 1445 -2955
rect 1479 -2989 1517 -2955
rect 1551 -2989 1589 -2955
rect 1623 -2989 1661 -2955
rect 1695 -2989 1733 -2955
rect 1767 -2989 1805 -2955
rect 1839 -2989 1877 -2955
rect 1911 -2989 1949 -2955
rect 1983 -2989 2021 -2955
rect 2055 -2989 2093 -2955
rect 2127 -2989 2165 -2955
rect 2199 -2989 2237 -2955
rect 2271 -2989 2309 -2955
rect 2343 -2989 2381 -2955
rect 2415 -2989 2453 -2955
rect 2487 -2989 2525 -2955
rect 2559 -2989 2597 -2955
rect 2631 -2989 2669 -2955
rect 2703 -2989 2741 -2955
rect 2775 -2989 2813 -2955
rect 2847 -2989 2885 -2955
rect 2919 -2989 2957 -2955
rect 2991 -2989 3029 -2955
rect 3063 -2989 3101 -2955
rect 3135 -2989 3173 -2955
rect 3207 -2989 3245 -2955
rect 3279 -2989 3317 -2955
rect 3351 -2989 3389 -2955
rect 3423 -2989 3461 -2955
rect 3495 -2989 3533 -2955
rect 3567 -2989 3605 -2955
rect 3639 -2989 3677 -2955
rect 3711 -2989 3749 -2955
rect 3783 -2989 3821 -2955
rect 3855 -2989 3893 -2955
rect 3927 -2989 3965 -2955
rect 3999 -2989 4037 -2955
rect 4071 -2989 4109 -2955
rect 4143 -2989 4181 -2955
rect 4215 -2989 4253 -2955
rect 4287 -2989 4325 -2955
rect 4359 -2989 4397 -2955
rect 4431 -2989 4469 -2955
rect 4503 -2989 4541 -2955
rect 4575 -2989 4613 -2955
rect 4647 -2989 4685 -2955
rect 4719 -2989 4757 -2955
rect 4791 -2989 4829 -2955
rect 4863 -2989 4901 -2955
rect 4935 -2989 4973 -2955
rect 5007 -2989 5045 -2955
rect 5079 -2989 5117 -2955
rect 5151 -2989 5189 -2955
rect 5223 -2989 5261 -2955
rect 5295 -2989 5333 -2955
rect 5367 -2989 5405 -2955
rect 5439 -2989 5477 -2955
rect 5511 -2989 5549 -2955
rect 5583 -2989 5621 -2955
rect 5655 -2989 5693 -2955
rect 5727 -2989 5765 -2955
rect 5799 -2989 5837 -2955
rect 5871 -2989 5909 -2955
rect 5943 -2989 5981 -2955
rect 6015 -2989 6053 -2955
rect 6087 -2989 6125 -2955
rect 6159 -2989 6197 -2955
rect 6231 -2989 6269 -2955
rect 6303 -2989 6341 -2955
rect 6375 -2989 6413 -2955
rect 6447 -2989 6485 -2955
rect 6519 -2989 6557 -2955
rect 6591 -2989 6629 -2955
rect 6663 -2989 6701 -2955
rect 6735 -2989 6773 -2955
rect 6807 -2989 6845 -2955
rect 6879 -2989 6917 -2955
rect 6951 -2989 6989 -2955
rect 7023 -2989 7061 -2955
rect 7095 -2989 7133 -2955
rect 7167 -2989 7205 -2955
rect 7239 -2989 7277 -2955
rect 7311 -2989 7349 -2955
rect 7383 -2989 7421 -2955
rect 7455 -2989 7493 -2955
rect 7527 -2989 7565 -2955
rect 7599 -2989 7637 -2955
rect 7671 -2989 7709 -2955
rect 7743 -2989 7781 -2955
rect 7815 -2989 7853 -2955
rect 7887 -2989 7925 -2955
rect 7959 -2989 7997 -2955
rect 8031 -2989 8069 -2955
rect 8103 -2989 8141 -2955
rect 8175 -2989 8213 -2955
rect 8247 -2989 8285 -2955
rect 8319 -2989 8357 -2955
rect 8391 -2989 8429 -2955
rect 8463 -2989 8501 -2955
rect 8535 -2989 8573 -2955
rect 8607 -2989 8645 -2955
rect 8679 -2989 8717 -2955
rect 8751 -2989 8789 -2955
rect 8823 -2989 8861 -2955
rect 8895 -2989 8933 -2955
rect 8967 -2989 9005 -2955
rect 9039 -2989 9077 -2955
rect 9111 -2989 9149 -2955
rect 9183 -2989 9221 -2955
rect 9255 -2989 9293 -2955
rect 9327 -2989 9365 -2955
rect 9399 -2989 9437 -2955
rect 9471 -2989 9509 -2955
rect 9543 -2989 9581 -2955
rect 9615 -2989 9653 -2955
rect 9687 -2989 9725 -2955
rect 9759 -2989 9797 -2955
rect 9831 -2989 9869 -2955
rect 9903 -2989 9941 -2955
rect 9975 -2989 10013 -2955
rect 10047 -2989 10085 -2955
rect 10119 -2989 10157 -2955
rect 10191 -2989 10229 -2955
rect 10263 -2989 10301 -2955
rect 10335 -2989 10373 -2955
rect 10407 -2989 10445 -2955
rect 10479 -2989 10517 -2955
rect 10551 -2989 10589 -2955
rect 10623 -2989 10661 -2955
rect 10695 -2989 10733 -2955
rect 10767 -2989 10805 -2955
rect 10839 -2989 10877 -2955
rect 10911 -2989 11028 -2955
rect -328 -3028 11028 -2989
<< via1 >>
rect -198 2024 366 2268
rect 10334 2024 10898 2268
rect 3514 1776 7278 1892
rect 4156 896 4208 948
rect 4284 786 4336 838
rect 5312 1560 5364 1612
rect 4672 896 4724 948
rect 4798 784 4850 836
rect 6350 1438 6402 1490
rect 5704 782 5756 834
rect 6868 780 6920 832
rect 3056 468 3108 520
rect 5704 468 5756 520
rect 8092 468 8144 520
rect 1498 174 1550 226
rect 2534 174 2586 226
rect 984 58 1036 110
rect 1374 -52 1426 0
rect 2016 58 2068 110
rect 1628 -52 1680 0
rect 2400 -52 2452 0
rect 3052 58 3104 110
rect 2662 -52 2714 0
rect 4794 180 4846 232
rect 5830 180 5882 232
rect 4280 64 4332 116
rect 1114 -782 1166 -730
rect 36 -892 88 -840
rect 1890 -782 1942 -730
rect 2144 -782 2196 -730
rect 2922 -782 2974 -730
rect 4670 -46 4722 6
rect 5312 64 5364 116
rect 4924 -46 4976 6
rect 5696 -46 5748 6
rect 6348 64 6400 116
rect 5958 -46 6010 6
rect 8090 174 8142 226
rect 9126 174 9178 226
rect 7576 58 7628 110
rect 1244 -892 1296 -840
rect 1756 -892 1808 -840
rect 2276 -892 2328 -840
rect 2792 -892 2844 -840
rect 4410 -776 4462 -724
rect 2922 -1014 2974 -962
rect 1034 -1138 1086 -1086
rect 1036 -1682 1088 -1630
rect 36 -2226 88 -2174
rect 2318 -1680 2370 -1628
rect 2752 -1682 2804 -1630
rect 3182 -1680 3234 -1628
rect 4540 -886 4592 -834
rect 5186 -776 5238 -724
rect 5440 -776 5492 -724
rect 6218 -776 6270 -724
rect 7966 -52 8018 0
rect 8608 58 8660 110
rect 8220 -52 8272 0
rect 8992 -52 9044 0
rect 9644 58 9696 110
rect 9254 -52 9306 0
rect 7706 -782 7758 -730
rect 5052 -886 5104 -834
rect 5572 -886 5624 -834
rect 6088 -886 6140 -834
rect 4802 -1014 4854 -962
rect 4468 -1138 4520 -1086
rect 4042 -1680 4094 -1628
rect 4472 -1682 4524 -1630
rect 6188 -1682 6240 -1630
rect 6614 -1680 6666 -1628
rect 6184 -2226 6236 -2174
rect 8482 -782 8534 -730
rect 8736 -782 8788 -730
rect 9514 -782 9566 -730
rect 7836 -892 7888 -840
rect 8348 -892 8400 -840
rect 8868 -892 8920 -840
rect 9384 -892 9436 -840
rect 9618 -1022 9670 -970
rect 10604 -892 10656 -840
rect 7472 -1680 7524 -1628
rect 7900 -1682 7952 -1630
rect 8326 -1680 8378 -1628
rect 9192 -1682 9244 -1630
rect 9616 -2220 9668 -2168
rect 10604 -2220 10656 -2168
rect 18 -2465 70 -2413
rect 82 -2465 134 -2413
rect 146 -2465 198 -2413
rect 210 -2465 262 -2413
rect 274 -2465 326 -2413
rect 338 -2465 390 -2413
rect 402 -2465 454 -2413
rect 466 -2465 518 -2413
rect 530 -2465 582 -2413
rect 594 -2465 646 -2413
rect 658 -2465 710 -2413
rect 722 -2465 774 -2413
rect 786 -2465 838 -2413
rect 850 -2465 902 -2413
rect 914 -2465 966 -2413
rect 978 -2465 1030 -2413
rect 1042 -2465 1094 -2413
rect 1106 -2465 1158 -2413
rect 1170 -2465 1222 -2413
rect 1234 -2465 1286 -2413
rect 1298 -2465 1350 -2413
rect 1362 -2465 1414 -2413
rect 1426 -2465 1478 -2413
rect 1490 -2465 1542 -2413
rect 1554 -2465 1606 -2413
rect 1618 -2465 1670 -2413
rect 1682 -2465 1734 -2413
rect 1746 -2465 1798 -2413
rect 1810 -2465 1862 -2413
rect 1874 -2465 1926 -2413
rect 1938 -2465 1990 -2413
rect 2002 -2465 2054 -2413
rect 2066 -2465 2118 -2413
rect 2130 -2465 2182 -2413
rect 2194 -2465 2246 -2413
rect 2258 -2465 2310 -2413
rect 2322 -2465 2374 -2413
rect 2386 -2465 2438 -2413
rect 2450 -2465 2502 -2413
rect 2514 -2465 2566 -2413
rect 2578 -2465 2630 -2413
rect 2642 -2465 2694 -2413
rect 2706 -2465 2758 -2413
rect 2770 -2465 2822 -2413
rect 2834 -2465 2886 -2413
rect 2898 -2465 2950 -2413
rect 2962 -2465 3014 -2413
rect 3026 -2465 3078 -2413
rect 3090 -2465 3142 -2413
rect 3154 -2465 3206 -2413
rect 3218 -2465 3270 -2413
rect 3282 -2465 3334 -2413
rect 3346 -2465 3398 -2413
rect 3410 -2465 3462 -2413
rect 3474 -2465 3526 -2413
rect 3538 -2465 3590 -2413
rect 3602 -2465 3654 -2413
rect 3666 -2465 3718 -2413
rect 3730 -2465 3782 -2413
rect 3794 -2465 3846 -2413
rect 3858 -2465 3910 -2413
rect 3922 -2465 3974 -2413
rect 3986 -2465 4038 -2413
rect 4050 -2465 4102 -2413
rect 4114 -2465 4166 -2413
rect 4178 -2465 4230 -2413
rect 4242 -2465 4294 -2413
rect 4306 -2465 4358 -2413
rect 4370 -2465 4422 -2413
rect 4434 -2465 4486 -2413
rect 4498 -2465 4550 -2413
rect 4562 -2465 4614 -2413
rect 4626 -2465 4678 -2413
rect 4690 -2465 4742 -2413
rect 4754 -2465 4806 -2413
rect 4818 -2465 4870 -2413
rect 4882 -2465 4934 -2413
rect 4946 -2465 4998 -2413
rect 5010 -2465 5062 -2413
rect 5074 -2465 5126 -2413
rect 5138 -2465 5190 -2413
rect 5202 -2465 5254 -2413
rect 5266 -2465 5318 -2413
rect 5330 -2465 5382 -2413
rect 5394 -2465 5446 -2413
rect 5458 -2465 5510 -2413
rect 5522 -2465 5574 -2413
rect 5586 -2465 5638 -2413
rect 5650 -2465 5702 -2413
rect 5714 -2465 5766 -2413
rect 5778 -2465 5830 -2413
rect 5842 -2465 5894 -2413
rect 5906 -2465 5958 -2413
rect 5970 -2465 6022 -2413
rect 6034 -2465 6086 -2413
rect 6098 -2465 6150 -2413
rect 6162 -2465 6214 -2413
rect 6226 -2465 6278 -2413
rect 6290 -2465 6342 -2413
rect 6354 -2465 6406 -2413
rect 6418 -2465 6470 -2413
rect 6482 -2465 6534 -2413
rect 6546 -2465 6598 -2413
rect 6610 -2465 6662 -2413
rect 6674 -2465 6726 -2413
rect 6738 -2465 6790 -2413
rect 6802 -2465 6854 -2413
rect 6866 -2465 6918 -2413
rect 6930 -2465 6982 -2413
rect 6994 -2465 7046 -2413
rect 7058 -2465 7110 -2413
rect 7122 -2465 7174 -2413
rect 7186 -2465 7238 -2413
rect 7250 -2465 7302 -2413
rect 7314 -2465 7366 -2413
rect 7378 -2465 7430 -2413
rect 7442 -2465 7494 -2413
rect 7506 -2465 7558 -2413
rect 7570 -2465 7622 -2413
rect 7634 -2465 7686 -2413
rect 7698 -2465 7750 -2413
rect 7762 -2465 7814 -2413
rect 7826 -2465 7878 -2413
rect 7890 -2465 7942 -2413
rect 7954 -2465 8006 -2413
rect 8018 -2465 8070 -2413
rect 8082 -2465 8134 -2413
rect 8146 -2465 8198 -2413
rect 8210 -2465 8262 -2413
rect 8274 -2465 8326 -2413
rect 8338 -2465 8390 -2413
rect 8402 -2465 8454 -2413
rect 8466 -2465 8518 -2413
rect 8530 -2465 8582 -2413
rect 8594 -2465 8646 -2413
rect 8658 -2465 8710 -2413
rect 8722 -2465 8774 -2413
rect 8786 -2465 8838 -2413
rect 8850 -2465 8902 -2413
rect 8914 -2465 8966 -2413
rect 8978 -2465 9030 -2413
rect 9042 -2465 9094 -2413
rect 9106 -2465 9158 -2413
rect 9170 -2465 9222 -2413
rect 9234 -2465 9286 -2413
rect 9298 -2465 9350 -2413
rect 9362 -2465 9414 -2413
rect 9426 -2465 9478 -2413
rect 9490 -2465 9542 -2413
rect 9554 -2465 9606 -2413
rect 9618 -2465 9670 -2413
rect 9682 -2465 9734 -2413
rect 9746 -2465 9798 -2413
rect 9810 -2465 9862 -2413
rect 9874 -2465 9926 -2413
rect 9938 -2465 9990 -2413
rect 10002 -2465 10054 -2413
rect 10066 -2465 10118 -2413
rect 10130 -2465 10182 -2413
rect 10194 -2465 10246 -2413
rect 10258 -2465 10310 -2413
rect 10322 -2465 10374 -2413
rect 10386 -2465 10438 -2413
rect 10450 -2465 10502 -2413
rect 10514 -2465 10566 -2413
rect 10578 -2465 10630 -2413
rect -198 -2888 366 -2644
rect 10334 -2888 10898 -2644
<< metal2 >>
rect -216 2294 384 2306
rect -216 2268 -184 2294
rect 352 2268 384 2294
rect -216 2024 -198 2268
rect 366 2024 384 2268
rect -216 1998 -184 2024
rect 352 1998 384 2024
rect -216 1986 384 1998
rect 10316 2294 10916 2306
rect 10316 2268 10348 2294
rect 10884 2268 10916 2294
rect 10316 2024 10334 2268
rect 10898 2024 10916 2268
rect 10316 1998 10348 2024
rect 10884 1998 10916 2024
rect 10316 1986 10916 1998
rect 3466 1902 7322 1950
rect 3466 1892 3528 1902
rect 7264 1892 7322 1902
rect 3466 1776 3514 1892
rect 7278 1776 7322 1892
rect 3466 1766 3528 1776
rect 7264 1766 7322 1776
rect 3466 1720 7322 1766
rect 5308 1616 5368 1622
rect 602 1612 5368 1616
rect 602 1560 5312 1612
rect 5364 1560 5368 1612
rect 602 1556 5368 1560
rect 602 168 662 1556
rect 5308 1550 5368 1556
rect 6346 1494 6406 1500
rect 2532 1490 6406 1494
rect 2532 1438 6350 1490
rect 6402 1438 6406 1490
rect 2532 1434 6406 1438
rect 2532 236 2592 1434
rect 6346 1428 6406 1434
rect 4152 952 4212 958
rect 4668 952 4728 958
rect 4152 948 10792 952
rect 4152 896 4156 948
rect 4208 896 4672 948
rect 4724 896 10792 948
rect 4152 892 10792 896
rect 4152 886 4212 892
rect 4668 886 4728 892
rect 4274 838 4346 842
rect 4274 786 4284 838
rect 4336 786 4346 838
rect 4274 782 4346 786
rect 4788 836 4860 840
rect 4788 784 4798 836
rect 4850 784 4860 836
rect 3046 520 3118 524
rect 3046 468 3056 520
rect 3108 468 3118 520
rect 3046 464 3118 468
rect -84 108 662 168
rect 1494 230 1554 236
rect 2530 230 2592 236
rect 1494 226 2592 230
rect 1494 174 1498 226
rect 1550 174 2534 226
rect 2586 174 2592 226
rect 1494 170 2592 174
rect 1494 164 1554 170
rect 2530 164 2590 170
rect 3052 120 3112 464
rect 4280 126 4340 782
rect 4788 780 4860 784
rect 5694 834 5766 838
rect 5694 782 5704 834
rect 5756 782 5766 834
rect 4794 242 4854 780
rect 5694 778 5766 782
rect 6864 836 6924 842
rect 6864 832 7632 836
rect 6864 780 6868 832
rect 6920 780 7632 832
rect 5700 524 5760 778
rect 6864 776 7632 780
rect 6864 770 6924 776
rect 5694 520 5766 524
rect 5694 468 5704 520
rect 5756 468 5766 520
rect 5694 464 5766 468
rect 4790 236 4854 242
rect 5826 236 5886 242
rect 4790 232 5886 236
rect 4790 180 4794 232
rect 4846 180 5830 232
rect 5882 180 5886 232
rect 4790 176 5886 180
rect 4790 170 4850 176
rect 5826 170 5886 176
rect 980 114 1040 120
rect 2012 114 2072 120
rect 3048 114 3112 120
rect 980 110 3112 114
rect -84 -1626 -24 108
rect 980 58 984 110
rect 1036 58 2016 110
rect 2068 58 3052 110
rect 3104 58 3112 110
rect 980 54 3112 58
rect 4276 120 4340 126
rect 5308 120 5368 126
rect 6344 120 6404 126
rect 4276 116 7262 120
rect 4276 64 4280 116
rect 4332 64 5312 116
rect 5364 64 6348 116
rect 6400 64 7262 116
rect 4276 60 7262 64
rect 4276 54 4336 60
rect 5308 54 5368 60
rect 6344 54 6404 60
rect 980 48 1040 54
rect 2012 48 2072 54
rect 3048 48 3108 54
rect 4666 10 4726 16
rect 4920 10 4980 16
rect 5692 10 5752 16
rect 5954 10 6014 16
rect 1370 4 1430 10
rect 1624 4 1684 10
rect 2396 4 2456 10
rect 2658 4 2718 10
rect 4666 6 6014 10
rect 1370 0 3716 4
rect 1370 -52 1374 0
rect 1426 -52 1628 0
rect 1680 -52 2400 0
rect 2452 -52 2662 0
rect 2714 -52 3716 0
rect 1370 -56 3716 -52
rect 4666 -46 4670 6
rect 4722 -46 4924 6
rect 4976 -46 5696 6
rect 5748 -46 5958 6
rect 6010 -46 6014 6
rect 4666 -50 6014 -46
rect 4666 -56 4726 -50
rect 4920 -56 4980 -50
rect 5692 -56 5752 -50
rect 5954 -56 6014 -50
rect 7202 4 7262 60
rect 7572 114 7632 776
rect 8082 520 8154 524
rect 8082 468 8092 520
rect 8144 468 8154 520
rect 8082 464 8154 468
rect 8088 236 8148 464
rect 8086 230 8148 236
rect 9122 230 9182 236
rect 8086 226 9182 230
rect 8086 174 8090 226
rect 8142 174 9126 226
rect 9178 174 9182 226
rect 8086 170 9182 174
rect 8086 164 8146 170
rect 9122 164 9182 170
rect 8604 114 8664 120
rect 9640 114 9700 120
rect 7572 110 9700 114
rect 7572 58 7576 110
rect 7628 58 8608 110
rect 8660 58 9644 110
rect 9696 58 9700 110
rect 7572 54 9700 58
rect 7572 48 7632 54
rect 8604 48 8664 54
rect 9640 48 9700 54
rect 7962 4 8022 10
rect 8216 4 8276 10
rect 8988 4 9048 10
rect 9250 4 9310 10
rect 7202 0 9310 4
rect 7202 -52 7966 0
rect 8018 -52 8220 0
rect 8272 -52 8992 0
rect 9044 -52 9254 0
rect 9306 -52 9310 0
rect 7202 -56 9310 -52
rect 1370 -62 1430 -56
rect 1624 -62 1684 -56
rect 2396 -62 2456 -56
rect 2658 -62 2718 -56
rect 1110 -726 1170 -720
rect 1886 -726 1946 -720
rect 2140 -726 2200 -720
rect 2918 -726 2978 -720
rect 1110 -730 2978 -726
rect 1110 -782 1114 -730
rect 1166 -782 1890 -730
rect 1942 -782 2144 -730
rect 2196 -782 2922 -730
rect 2974 -782 2978 -730
rect 1110 -786 2978 -782
rect 1110 -792 1170 -786
rect 1886 -792 1946 -786
rect 2140 -792 2200 -786
rect 2918 -792 2978 -786
rect 32 -836 92 -830
rect 1752 -836 1812 -830
rect 2272 -836 2332 -830
rect 2788 -836 2848 -830
rect 32 -840 2848 -836
rect 3656 -838 3716 -56
rect 7962 -62 8022 -56
rect 8216 -62 8276 -56
rect 8988 -62 9048 -56
rect 9250 -62 9310 -56
rect 4406 -720 4466 -714
rect 5182 -720 5242 -714
rect 5436 -720 5496 -714
rect 6214 -720 6274 -714
rect 4406 -724 6274 -720
rect 4406 -776 4410 -724
rect 4462 -776 5186 -724
rect 5238 -776 5440 -724
rect 5492 -776 6218 -724
rect 6270 -776 6274 -724
rect 4406 -780 6274 -776
rect 4406 -786 4466 -780
rect 5182 -786 5242 -780
rect 5436 -786 5496 -780
rect 6214 -786 6274 -780
rect 7702 -726 7762 -720
rect 8478 -726 8538 -720
rect 8732 -726 8792 -720
rect 9510 -726 9570 -720
rect 7702 -730 9570 -726
rect 7702 -782 7706 -730
rect 7758 -782 8482 -730
rect 8534 -782 8736 -730
rect 8788 -782 9514 -730
rect 9566 -782 9570 -730
rect 7702 -786 9570 -782
rect 7702 -792 7764 -786
rect 8478 -792 8538 -786
rect 8732 -792 8792 -786
rect 9510 -792 9570 -786
rect 5048 -830 5108 -824
rect 5568 -830 5628 -824
rect 6084 -830 6144 -824
rect 4530 -834 6144 -830
rect 32 -892 36 -840
rect 88 -892 1244 -840
rect 1296 -892 1756 -840
rect 1808 -892 2276 -840
rect 2328 -892 2792 -840
rect 2844 -892 2848 -840
rect 32 -896 2848 -892
rect 32 -902 92 -896
rect 1752 -902 1812 -896
rect 2272 -902 2332 -896
rect 2788 -902 2848 -896
rect 3647 -840 3725 -838
rect 3647 -896 3658 -840
rect 3714 -896 3725 -840
rect 4530 -886 4540 -834
rect 4592 -886 5052 -834
rect 5104 -886 5572 -834
rect 5624 -886 6088 -834
rect 6140 -886 6144 -834
rect 7704 -840 7764 -792
rect 7832 -836 7892 -830
rect 8344 -836 8404 -830
rect 8864 -836 8924 -830
rect 9380 -836 9440 -830
rect 10600 -836 10660 -830
rect 7832 -840 10660 -836
rect 4530 -890 6144 -886
rect 5048 -896 5108 -890
rect 5568 -896 5628 -890
rect 6084 -896 6144 -890
rect 7697 -896 7706 -840
rect 7762 -896 7771 -840
rect 7832 -892 7836 -840
rect 7888 -892 8348 -840
rect 8400 -892 8868 -840
rect 8920 -892 9384 -840
rect 9436 -892 10604 -840
rect 10656 -892 10660 -840
rect 7832 -896 10660 -892
rect 3647 -898 3725 -896
rect 7704 -898 7764 -896
rect 7832 -902 7892 -896
rect 8344 -902 8404 -896
rect 8864 -902 8924 -896
rect 9380 -902 9440 -896
rect 10600 -902 10660 -896
rect 2918 -958 2978 -952
rect 4798 -958 4858 -952
rect 2918 -962 4858 -958
rect 2918 -1014 2922 -962
rect 2974 -1014 4802 -962
rect 4854 -1014 4858 -962
rect 2918 -1018 4858 -1014
rect 2918 -1024 2978 -1018
rect 4798 -1024 4858 -1018
rect 9614 -966 9674 -960
rect 10732 -966 10792 892
rect 9614 -970 10792 -966
rect 9614 -1022 9618 -970
rect 9670 -1022 10792 -970
rect 9614 -1026 10792 -1022
rect 9614 -1032 9674 -1026
rect 1030 -1082 1090 -1076
rect 4464 -1082 4524 -1076
rect 1030 -1086 4524 -1082
rect 1030 -1138 1034 -1086
rect 1086 -1138 4468 -1086
rect 4520 -1138 4524 -1086
rect 1030 -1142 4524 -1138
rect 1030 -1148 1090 -1142
rect 4464 -1148 4524 -1142
rect 1032 -1626 1092 -1620
rect -84 -1630 1092 -1626
rect -84 -1682 1036 -1630
rect 1088 -1682 1092 -1630
rect -84 -1686 1092 -1682
rect 1032 -1692 1092 -1686
rect 2314 -1626 2374 -1620
rect 2748 -1626 2808 -1620
rect 4468 -1626 4528 -1620
rect 6184 -1626 6244 -1620
rect 6610 -1626 6670 -1620
rect 7896 -1626 7956 -1620
rect 2314 -1628 9254 -1626
rect 2314 -1680 2318 -1628
rect 2370 -1630 3182 -1628
rect 2370 -1680 2752 -1630
rect 2314 -1682 2752 -1680
rect 2804 -1680 3182 -1630
rect 3234 -1680 4042 -1628
rect 4094 -1630 6614 -1628
rect 4094 -1680 4472 -1630
rect 2804 -1682 4472 -1680
rect 4524 -1682 6188 -1630
rect 6240 -1680 6614 -1630
rect 6666 -1680 7472 -1628
rect 7524 -1630 8326 -1628
rect 7524 -1680 7900 -1630
rect 6240 -1682 7900 -1680
rect 7952 -1680 8326 -1630
rect 8378 -1630 9254 -1628
rect 8378 -1680 9192 -1630
rect 7952 -1682 9192 -1680
rect 9244 -1682 9254 -1630
rect 2314 -1686 9254 -1682
rect 2314 -1692 2374 -1686
rect 2748 -1692 2808 -1686
rect 4468 -1692 4528 -1686
rect 6184 -1692 6244 -1686
rect 6610 -1692 6670 -1686
rect 7896 -1692 7956 -1686
rect 9612 -2164 9672 -2158
rect 10600 -2164 10660 -2158
rect 32 -2170 92 -2164
rect 6180 -2170 6240 -2164
rect 32 -2174 6240 -2170
rect 32 -2226 36 -2174
rect 88 -2226 6184 -2174
rect 6236 -2226 6240 -2174
rect 32 -2230 6240 -2226
rect 9612 -2168 10660 -2164
rect 9612 -2220 9616 -2168
rect 9668 -2220 10604 -2168
rect 10656 -2220 10660 -2168
rect 9612 -2224 10660 -2220
rect 9612 -2230 9672 -2224
rect 10600 -2230 10660 -2224
rect 32 -2236 92 -2230
rect 6180 -2236 6240 -2230
rect -66 -2411 10708 -2336
rect -66 -2467 16 -2411
rect 72 -2413 96 -2411
rect 152 -2413 176 -2411
rect 232 -2413 256 -2411
rect 312 -2413 336 -2411
rect 392 -2413 416 -2411
rect 472 -2413 496 -2411
rect 552 -2413 576 -2411
rect 632 -2413 656 -2411
rect 712 -2413 736 -2411
rect 792 -2413 816 -2411
rect 872 -2413 896 -2411
rect 952 -2413 976 -2411
rect 1032 -2413 1056 -2411
rect 1112 -2413 1136 -2411
rect 1192 -2413 1216 -2411
rect 1272 -2413 1296 -2411
rect 1352 -2413 1376 -2411
rect 1432 -2413 1456 -2411
rect 1512 -2413 1536 -2411
rect 1592 -2413 1616 -2411
rect 1672 -2413 1696 -2411
rect 1752 -2413 1776 -2411
rect 1832 -2413 1856 -2411
rect 1912 -2413 1936 -2411
rect 1992 -2413 2016 -2411
rect 2072 -2413 2096 -2411
rect 2152 -2413 2176 -2411
rect 2232 -2413 2256 -2411
rect 2312 -2413 2336 -2411
rect 2392 -2413 2416 -2411
rect 2472 -2413 2496 -2411
rect 2552 -2413 2576 -2411
rect 2632 -2413 2656 -2411
rect 2712 -2413 2736 -2411
rect 2792 -2413 2816 -2411
rect 2872 -2413 2896 -2411
rect 2952 -2413 2976 -2411
rect 3032 -2413 3056 -2411
rect 3112 -2413 3136 -2411
rect 3192 -2413 3216 -2411
rect 3272 -2413 3296 -2411
rect 3352 -2413 3376 -2411
rect 3432 -2413 3456 -2411
rect 3512 -2413 3536 -2411
rect 3592 -2413 3616 -2411
rect 3672 -2413 3696 -2411
rect 3752 -2413 3776 -2411
rect 3832 -2413 3856 -2411
rect 3912 -2413 3936 -2411
rect 3992 -2413 4016 -2411
rect 4072 -2413 4096 -2411
rect 4152 -2413 4176 -2411
rect 4232 -2413 4256 -2411
rect 4312 -2413 4336 -2411
rect 4392 -2413 4416 -2411
rect 4472 -2413 4496 -2411
rect 4552 -2413 4576 -2411
rect 4632 -2413 4656 -2411
rect 4712 -2413 4736 -2411
rect 4792 -2413 4816 -2411
rect 4872 -2413 4896 -2411
rect 4952 -2413 4976 -2411
rect 5032 -2413 5056 -2411
rect 5112 -2413 5136 -2411
rect 5192 -2413 5216 -2411
rect 5272 -2413 5296 -2411
rect 5352 -2413 5376 -2411
rect 5432 -2413 5456 -2411
rect 5512 -2413 5536 -2411
rect 5592 -2413 5616 -2411
rect 5672 -2413 5696 -2411
rect 5752 -2413 5776 -2411
rect 5832 -2413 5856 -2411
rect 5912 -2413 5936 -2411
rect 5992 -2413 6016 -2411
rect 6072 -2413 6096 -2411
rect 6152 -2413 6176 -2411
rect 6232 -2413 6256 -2411
rect 6312 -2413 6336 -2411
rect 6392 -2413 6416 -2411
rect 6472 -2413 6496 -2411
rect 6552 -2413 6576 -2411
rect 6632 -2413 6656 -2411
rect 6712 -2413 6736 -2411
rect 6792 -2413 6816 -2411
rect 6872 -2413 6896 -2411
rect 6952 -2413 6976 -2411
rect 7032 -2413 7056 -2411
rect 7112 -2413 7136 -2411
rect 7192 -2413 7216 -2411
rect 7272 -2413 7296 -2411
rect 7352 -2413 7376 -2411
rect 7432 -2413 7456 -2411
rect 7512 -2413 7536 -2411
rect 7592 -2413 7616 -2411
rect 7672 -2413 7696 -2411
rect 7752 -2413 7776 -2411
rect 7832 -2413 7856 -2411
rect 7912 -2413 7936 -2411
rect 7992 -2413 8016 -2411
rect 8072 -2413 8096 -2411
rect 8152 -2413 8176 -2411
rect 8232 -2413 8256 -2411
rect 8312 -2413 8336 -2411
rect 8392 -2413 8416 -2411
rect 8472 -2413 8496 -2411
rect 8552 -2413 8576 -2411
rect 8632 -2413 8656 -2411
rect 8712 -2413 8736 -2411
rect 8792 -2413 8816 -2411
rect 8872 -2413 8896 -2411
rect 8952 -2413 8976 -2411
rect 9032 -2413 9056 -2411
rect 9112 -2413 9136 -2411
rect 9192 -2413 9216 -2411
rect 9272 -2413 9296 -2411
rect 9352 -2413 9376 -2411
rect 9432 -2413 9456 -2411
rect 9512 -2413 9536 -2411
rect 9592 -2413 9616 -2411
rect 9672 -2413 9696 -2411
rect 9752 -2413 9776 -2411
rect 9832 -2413 9856 -2411
rect 9912 -2413 9936 -2411
rect 9992 -2413 10016 -2411
rect 10072 -2413 10096 -2411
rect 10152 -2413 10176 -2411
rect 10232 -2413 10256 -2411
rect 10312 -2413 10336 -2411
rect 10392 -2413 10416 -2411
rect 10472 -2413 10496 -2411
rect 10552 -2413 10576 -2411
rect 72 -2465 82 -2413
rect 326 -2465 336 -2413
rect 392 -2465 402 -2413
rect 646 -2465 656 -2413
rect 712 -2465 722 -2413
rect 966 -2465 976 -2413
rect 1032 -2465 1042 -2413
rect 1286 -2465 1296 -2413
rect 1352 -2465 1362 -2413
rect 1606 -2465 1616 -2413
rect 1672 -2465 1682 -2413
rect 1926 -2465 1936 -2413
rect 1992 -2465 2002 -2413
rect 2246 -2465 2256 -2413
rect 2312 -2465 2322 -2413
rect 2566 -2465 2576 -2413
rect 2632 -2465 2642 -2413
rect 2886 -2465 2896 -2413
rect 2952 -2465 2962 -2413
rect 3206 -2465 3216 -2413
rect 3272 -2465 3282 -2413
rect 3526 -2465 3536 -2413
rect 3592 -2465 3602 -2413
rect 3846 -2465 3856 -2413
rect 3912 -2465 3922 -2413
rect 4166 -2465 4176 -2413
rect 4232 -2465 4242 -2413
rect 4486 -2465 4496 -2413
rect 4552 -2465 4562 -2413
rect 4806 -2465 4816 -2413
rect 4872 -2465 4882 -2413
rect 5126 -2465 5136 -2413
rect 5192 -2465 5202 -2413
rect 5446 -2465 5456 -2413
rect 5512 -2465 5522 -2413
rect 5766 -2465 5776 -2413
rect 5832 -2465 5842 -2413
rect 6086 -2465 6096 -2413
rect 6152 -2465 6162 -2413
rect 6406 -2465 6416 -2413
rect 6472 -2465 6482 -2413
rect 6726 -2465 6736 -2413
rect 6792 -2465 6802 -2413
rect 7046 -2465 7056 -2413
rect 7112 -2465 7122 -2413
rect 7366 -2465 7376 -2413
rect 7432 -2465 7442 -2413
rect 7686 -2465 7696 -2413
rect 7752 -2465 7762 -2413
rect 8006 -2465 8016 -2413
rect 8072 -2465 8082 -2413
rect 8326 -2465 8336 -2413
rect 8392 -2465 8402 -2413
rect 8646 -2465 8656 -2413
rect 8712 -2465 8722 -2413
rect 8966 -2465 8976 -2413
rect 9032 -2465 9042 -2413
rect 9286 -2465 9296 -2413
rect 9352 -2465 9362 -2413
rect 9606 -2465 9616 -2413
rect 9672 -2465 9682 -2413
rect 9926 -2465 9936 -2413
rect 9992 -2465 10002 -2413
rect 10246 -2465 10256 -2413
rect 10312 -2465 10322 -2413
rect 10566 -2465 10576 -2413
rect 72 -2467 96 -2465
rect 152 -2467 176 -2465
rect 232 -2467 256 -2465
rect 312 -2467 336 -2465
rect 392 -2467 416 -2465
rect 472 -2467 496 -2465
rect 552 -2467 576 -2465
rect 632 -2467 656 -2465
rect 712 -2467 736 -2465
rect 792 -2467 816 -2465
rect 872 -2467 896 -2465
rect 952 -2467 976 -2465
rect 1032 -2467 1056 -2465
rect 1112 -2467 1136 -2465
rect 1192 -2467 1216 -2465
rect 1272 -2467 1296 -2465
rect 1352 -2467 1376 -2465
rect 1432 -2467 1456 -2465
rect 1512 -2467 1536 -2465
rect 1592 -2467 1616 -2465
rect 1672 -2467 1696 -2465
rect 1752 -2467 1776 -2465
rect 1832 -2467 1856 -2465
rect 1912 -2467 1936 -2465
rect 1992 -2467 2016 -2465
rect 2072 -2467 2096 -2465
rect 2152 -2467 2176 -2465
rect 2232 -2467 2256 -2465
rect 2312 -2467 2336 -2465
rect 2392 -2467 2416 -2465
rect 2472 -2467 2496 -2465
rect 2552 -2467 2576 -2465
rect 2632 -2467 2656 -2465
rect 2712 -2467 2736 -2465
rect 2792 -2467 2816 -2465
rect 2872 -2467 2896 -2465
rect 2952 -2467 2976 -2465
rect 3032 -2467 3056 -2465
rect 3112 -2467 3136 -2465
rect 3192 -2467 3216 -2465
rect 3272 -2467 3296 -2465
rect 3352 -2467 3376 -2465
rect 3432 -2467 3456 -2465
rect 3512 -2467 3536 -2465
rect 3592 -2467 3616 -2465
rect 3672 -2467 3696 -2465
rect 3752 -2467 3776 -2465
rect 3832 -2467 3856 -2465
rect 3912 -2467 3936 -2465
rect 3992 -2467 4016 -2465
rect 4072 -2467 4096 -2465
rect 4152 -2467 4176 -2465
rect 4232 -2467 4256 -2465
rect 4312 -2467 4336 -2465
rect 4392 -2467 4416 -2465
rect 4472 -2467 4496 -2465
rect 4552 -2467 4576 -2465
rect 4632 -2467 4656 -2465
rect 4712 -2467 4736 -2465
rect 4792 -2467 4816 -2465
rect 4872 -2467 4896 -2465
rect 4952 -2467 4976 -2465
rect 5032 -2467 5056 -2465
rect 5112 -2467 5136 -2465
rect 5192 -2467 5216 -2465
rect 5272 -2467 5296 -2465
rect 5352 -2467 5376 -2465
rect 5432 -2467 5456 -2465
rect 5512 -2467 5536 -2465
rect 5592 -2467 5616 -2465
rect 5672 -2467 5696 -2465
rect 5752 -2467 5776 -2465
rect 5832 -2467 5856 -2465
rect 5912 -2467 5936 -2465
rect 5992 -2467 6016 -2465
rect 6072 -2467 6096 -2465
rect 6152 -2467 6176 -2465
rect 6232 -2467 6256 -2465
rect 6312 -2467 6336 -2465
rect 6392 -2467 6416 -2465
rect 6472 -2467 6496 -2465
rect 6552 -2467 6576 -2465
rect 6632 -2467 6656 -2465
rect 6712 -2467 6736 -2465
rect 6792 -2467 6816 -2465
rect 6872 -2467 6896 -2465
rect 6952 -2467 6976 -2465
rect 7032 -2467 7056 -2465
rect 7112 -2467 7136 -2465
rect 7192 -2467 7216 -2465
rect 7272 -2467 7296 -2465
rect 7352 -2467 7376 -2465
rect 7432 -2467 7456 -2465
rect 7512 -2467 7536 -2465
rect 7592 -2467 7616 -2465
rect 7672 -2467 7696 -2465
rect 7752 -2467 7776 -2465
rect 7832 -2467 7856 -2465
rect 7912 -2467 7936 -2465
rect 7992 -2467 8016 -2465
rect 8072 -2467 8096 -2465
rect 8152 -2467 8176 -2465
rect 8232 -2467 8256 -2465
rect 8312 -2467 8336 -2465
rect 8392 -2467 8416 -2465
rect 8472 -2467 8496 -2465
rect 8552 -2467 8576 -2465
rect 8632 -2467 8656 -2465
rect 8712 -2467 8736 -2465
rect 8792 -2467 8816 -2465
rect 8872 -2467 8896 -2465
rect 8952 -2467 8976 -2465
rect 9032 -2467 9056 -2465
rect 9112 -2467 9136 -2465
rect 9192 -2467 9216 -2465
rect 9272 -2467 9296 -2465
rect 9352 -2467 9376 -2465
rect 9432 -2467 9456 -2465
rect 9512 -2467 9536 -2465
rect 9592 -2467 9616 -2465
rect 9672 -2467 9696 -2465
rect 9752 -2467 9776 -2465
rect 9832 -2467 9856 -2465
rect 9912 -2467 9936 -2465
rect 9992 -2467 10016 -2465
rect 10072 -2467 10096 -2465
rect 10152 -2467 10176 -2465
rect 10232 -2467 10256 -2465
rect 10312 -2467 10336 -2465
rect 10392 -2467 10416 -2465
rect 10472 -2467 10496 -2465
rect 10552 -2467 10576 -2465
rect 10632 -2467 10708 -2411
rect -66 -2550 10708 -2467
rect -216 -2618 384 -2606
rect -216 -2644 -184 -2618
rect 352 -2644 384 -2618
rect -216 -2888 -198 -2644
rect 366 -2888 384 -2644
rect -216 -2914 -184 -2888
rect 352 -2914 384 -2888
rect -216 -2926 384 -2914
rect 10316 -2618 10916 -2606
rect 10316 -2644 10348 -2618
rect 10884 -2644 10916 -2618
rect 10316 -2888 10334 -2644
rect 10898 -2888 10916 -2644
rect 10316 -2914 10348 -2888
rect 10884 -2914 10916 -2888
rect 10316 -2926 10916 -2914
<< via2 >>
rect -184 2268 352 2294
rect -184 2024 352 2268
rect -184 1998 352 2024
rect 10348 2268 10884 2294
rect 10348 2024 10884 2268
rect 10348 1998 10884 2024
rect 3528 1892 7264 1902
rect 3528 1776 7264 1892
rect 3528 1766 7264 1776
rect 3658 -896 3714 -840
rect 7706 -896 7762 -840
rect 16 -2413 72 -2411
rect 96 -2413 152 -2411
rect 176 -2413 232 -2411
rect 256 -2413 312 -2411
rect 336 -2413 392 -2411
rect 416 -2413 472 -2411
rect 496 -2413 552 -2411
rect 576 -2413 632 -2411
rect 656 -2413 712 -2411
rect 736 -2413 792 -2411
rect 816 -2413 872 -2411
rect 896 -2413 952 -2411
rect 976 -2413 1032 -2411
rect 1056 -2413 1112 -2411
rect 1136 -2413 1192 -2411
rect 1216 -2413 1272 -2411
rect 1296 -2413 1352 -2411
rect 1376 -2413 1432 -2411
rect 1456 -2413 1512 -2411
rect 1536 -2413 1592 -2411
rect 1616 -2413 1672 -2411
rect 1696 -2413 1752 -2411
rect 1776 -2413 1832 -2411
rect 1856 -2413 1912 -2411
rect 1936 -2413 1992 -2411
rect 2016 -2413 2072 -2411
rect 2096 -2413 2152 -2411
rect 2176 -2413 2232 -2411
rect 2256 -2413 2312 -2411
rect 2336 -2413 2392 -2411
rect 2416 -2413 2472 -2411
rect 2496 -2413 2552 -2411
rect 2576 -2413 2632 -2411
rect 2656 -2413 2712 -2411
rect 2736 -2413 2792 -2411
rect 2816 -2413 2872 -2411
rect 2896 -2413 2952 -2411
rect 2976 -2413 3032 -2411
rect 3056 -2413 3112 -2411
rect 3136 -2413 3192 -2411
rect 3216 -2413 3272 -2411
rect 3296 -2413 3352 -2411
rect 3376 -2413 3432 -2411
rect 3456 -2413 3512 -2411
rect 3536 -2413 3592 -2411
rect 3616 -2413 3672 -2411
rect 3696 -2413 3752 -2411
rect 3776 -2413 3832 -2411
rect 3856 -2413 3912 -2411
rect 3936 -2413 3992 -2411
rect 4016 -2413 4072 -2411
rect 4096 -2413 4152 -2411
rect 4176 -2413 4232 -2411
rect 4256 -2413 4312 -2411
rect 4336 -2413 4392 -2411
rect 4416 -2413 4472 -2411
rect 4496 -2413 4552 -2411
rect 4576 -2413 4632 -2411
rect 4656 -2413 4712 -2411
rect 4736 -2413 4792 -2411
rect 4816 -2413 4872 -2411
rect 4896 -2413 4952 -2411
rect 4976 -2413 5032 -2411
rect 5056 -2413 5112 -2411
rect 5136 -2413 5192 -2411
rect 5216 -2413 5272 -2411
rect 5296 -2413 5352 -2411
rect 5376 -2413 5432 -2411
rect 5456 -2413 5512 -2411
rect 5536 -2413 5592 -2411
rect 5616 -2413 5672 -2411
rect 5696 -2413 5752 -2411
rect 5776 -2413 5832 -2411
rect 5856 -2413 5912 -2411
rect 5936 -2413 5992 -2411
rect 6016 -2413 6072 -2411
rect 6096 -2413 6152 -2411
rect 6176 -2413 6232 -2411
rect 6256 -2413 6312 -2411
rect 6336 -2413 6392 -2411
rect 6416 -2413 6472 -2411
rect 6496 -2413 6552 -2411
rect 6576 -2413 6632 -2411
rect 6656 -2413 6712 -2411
rect 6736 -2413 6792 -2411
rect 6816 -2413 6872 -2411
rect 6896 -2413 6952 -2411
rect 6976 -2413 7032 -2411
rect 7056 -2413 7112 -2411
rect 7136 -2413 7192 -2411
rect 7216 -2413 7272 -2411
rect 7296 -2413 7352 -2411
rect 7376 -2413 7432 -2411
rect 7456 -2413 7512 -2411
rect 7536 -2413 7592 -2411
rect 7616 -2413 7672 -2411
rect 7696 -2413 7752 -2411
rect 7776 -2413 7832 -2411
rect 7856 -2413 7912 -2411
rect 7936 -2413 7992 -2411
rect 8016 -2413 8072 -2411
rect 8096 -2413 8152 -2411
rect 8176 -2413 8232 -2411
rect 8256 -2413 8312 -2411
rect 8336 -2413 8392 -2411
rect 8416 -2413 8472 -2411
rect 8496 -2413 8552 -2411
rect 8576 -2413 8632 -2411
rect 8656 -2413 8712 -2411
rect 8736 -2413 8792 -2411
rect 8816 -2413 8872 -2411
rect 8896 -2413 8952 -2411
rect 8976 -2413 9032 -2411
rect 9056 -2413 9112 -2411
rect 9136 -2413 9192 -2411
rect 9216 -2413 9272 -2411
rect 9296 -2413 9352 -2411
rect 9376 -2413 9432 -2411
rect 9456 -2413 9512 -2411
rect 9536 -2413 9592 -2411
rect 9616 -2413 9672 -2411
rect 9696 -2413 9752 -2411
rect 9776 -2413 9832 -2411
rect 9856 -2413 9912 -2411
rect 9936 -2413 9992 -2411
rect 10016 -2413 10072 -2411
rect 10096 -2413 10152 -2411
rect 10176 -2413 10232 -2411
rect 10256 -2413 10312 -2411
rect 10336 -2413 10392 -2411
rect 10416 -2413 10472 -2411
rect 10496 -2413 10552 -2411
rect 10576 -2413 10632 -2411
rect 16 -2465 18 -2413
rect 18 -2465 70 -2413
rect 70 -2465 72 -2413
rect 96 -2465 134 -2413
rect 134 -2465 146 -2413
rect 146 -2465 152 -2413
rect 176 -2465 198 -2413
rect 198 -2465 210 -2413
rect 210 -2465 232 -2413
rect 256 -2465 262 -2413
rect 262 -2465 274 -2413
rect 274 -2465 312 -2413
rect 336 -2465 338 -2413
rect 338 -2465 390 -2413
rect 390 -2465 392 -2413
rect 416 -2465 454 -2413
rect 454 -2465 466 -2413
rect 466 -2465 472 -2413
rect 496 -2465 518 -2413
rect 518 -2465 530 -2413
rect 530 -2465 552 -2413
rect 576 -2465 582 -2413
rect 582 -2465 594 -2413
rect 594 -2465 632 -2413
rect 656 -2465 658 -2413
rect 658 -2465 710 -2413
rect 710 -2465 712 -2413
rect 736 -2465 774 -2413
rect 774 -2465 786 -2413
rect 786 -2465 792 -2413
rect 816 -2465 838 -2413
rect 838 -2465 850 -2413
rect 850 -2465 872 -2413
rect 896 -2465 902 -2413
rect 902 -2465 914 -2413
rect 914 -2465 952 -2413
rect 976 -2465 978 -2413
rect 978 -2465 1030 -2413
rect 1030 -2465 1032 -2413
rect 1056 -2465 1094 -2413
rect 1094 -2465 1106 -2413
rect 1106 -2465 1112 -2413
rect 1136 -2465 1158 -2413
rect 1158 -2465 1170 -2413
rect 1170 -2465 1192 -2413
rect 1216 -2465 1222 -2413
rect 1222 -2465 1234 -2413
rect 1234 -2465 1272 -2413
rect 1296 -2465 1298 -2413
rect 1298 -2465 1350 -2413
rect 1350 -2465 1352 -2413
rect 1376 -2465 1414 -2413
rect 1414 -2465 1426 -2413
rect 1426 -2465 1432 -2413
rect 1456 -2465 1478 -2413
rect 1478 -2465 1490 -2413
rect 1490 -2465 1512 -2413
rect 1536 -2465 1542 -2413
rect 1542 -2465 1554 -2413
rect 1554 -2465 1592 -2413
rect 1616 -2465 1618 -2413
rect 1618 -2465 1670 -2413
rect 1670 -2465 1672 -2413
rect 1696 -2465 1734 -2413
rect 1734 -2465 1746 -2413
rect 1746 -2465 1752 -2413
rect 1776 -2465 1798 -2413
rect 1798 -2465 1810 -2413
rect 1810 -2465 1832 -2413
rect 1856 -2465 1862 -2413
rect 1862 -2465 1874 -2413
rect 1874 -2465 1912 -2413
rect 1936 -2465 1938 -2413
rect 1938 -2465 1990 -2413
rect 1990 -2465 1992 -2413
rect 2016 -2465 2054 -2413
rect 2054 -2465 2066 -2413
rect 2066 -2465 2072 -2413
rect 2096 -2465 2118 -2413
rect 2118 -2465 2130 -2413
rect 2130 -2465 2152 -2413
rect 2176 -2465 2182 -2413
rect 2182 -2465 2194 -2413
rect 2194 -2465 2232 -2413
rect 2256 -2465 2258 -2413
rect 2258 -2465 2310 -2413
rect 2310 -2465 2312 -2413
rect 2336 -2465 2374 -2413
rect 2374 -2465 2386 -2413
rect 2386 -2465 2392 -2413
rect 2416 -2465 2438 -2413
rect 2438 -2465 2450 -2413
rect 2450 -2465 2472 -2413
rect 2496 -2465 2502 -2413
rect 2502 -2465 2514 -2413
rect 2514 -2465 2552 -2413
rect 2576 -2465 2578 -2413
rect 2578 -2465 2630 -2413
rect 2630 -2465 2632 -2413
rect 2656 -2465 2694 -2413
rect 2694 -2465 2706 -2413
rect 2706 -2465 2712 -2413
rect 2736 -2465 2758 -2413
rect 2758 -2465 2770 -2413
rect 2770 -2465 2792 -2413
rect 2816 -2465 2822 -2413
rect 2822 -2465 2834 -2413
rect 2834 -2465 2872 -2413
rect 2896 -2465 2898 -2413
rect 2898 -2465 2950 -2413
rect 2950 -2465 2952 -2413
rect 2976 -2465 3014 -2413
rect 3014 -2465 3026 -2413
rect 3026 -2465 3032 -2413
rect 3056 -2465 3078 -2413
rect 3078 -2465 3090 -2413
rect 3090 -2465 3112 -2413
rect 3136 -2465 3142 -2413
rect 3142 -2465 3154 -2413
rect 3154 -2465 3192 -2413
rect 3216 -2465 3218 -2413
rect 3218 -2465 3270 -2413
rect 3270 -2465 3272 -2413
rect 3296 -2465 3334 -2413
rect 3334 -2465 3346 -2413
rect 3346 -2465 3352 -2413
rect 3376 -2465 3398 -2413
rect 3398 -2465 3410 -2413
rect 3410 -2465 3432 -2413
rect 3456 -2465 3462 -2413
rect 3462 -2465 3474 -2413
rect 3474 -2465 3512 -2413
rect 3536 -2465 3538 -2413
rect 3538 -2465 3590 -2413
rect 3590 -2465 3592 -2413
rect 3616 -2465 3654 -2413
rect 3654 -2465 3666 -2413
rect 3666 -2465 3672 -2413
rect 3696 -2465 3718 -2413
rect 3718 -2465 3730 -2413
rect 3730 -2465 3752 -2413
rect 3776 -2465 3782 -2413
rect 3782 -2465 3794 -2413
rect 3794 -2465 3832 -2413
rect 3856 -2465 3858 -2413
rect 3858 -2465 3910 -2413
rect 3910 -2465 3912 -2413
rect 3936 -2465 3974 -2413
rect 3974 -2465 3986 -2413
rect 3986 -2465 3992 -2413
rect 4016 -2465 4038 -2413
rect 4038 -2465 4050 -2413
rect 4050 -2465 4072 -2413
rect 4096 -2465 4102 -2413
rect 4102 -2465 4114 -2413
rect 4114 -2465 4152 -2413
rect 4176 -2465 4178 -2413
rect 4178 -2465 4230 -2413
rect 4230 -2465 4232 -2413
rect 4256 -2465 4294 -2413
rect 4294 -2465 4306 -2413
rect 4306 -2465 4312 -2413
rect 4336 -2465 4358 -2413
rect 4358 -2465 4370 -2413
rect 4370 -2465 4392 -2413
rect 4416 -2465 4422 -2413
rect 4422 -2465 4434 -2413
rect 4434 -2465 4472 -2413
rect 4496 -2465 4498 -2413
rect 4498 -2465 4550 -2413
rect 4550 -2465 4552 -2413
rect 4576 -2465 4614 -2413
rect 4614 -2465 4626 -2413
rect 4626 -2465 4632 -2413
rect 4656 -2465 4678 -2413
rect 4678 -2465 4690 -2413
rect 4690 -2465 4712 -2413
rect 4736 -2465 4742 -2413
rect 4742 -2465 4754 -2413
rect 4754 -2465 4792 -2413
rect 4816 -2465 4818 -2413
rect 4818 -2465 4870 -2413
rect 4870 -2465 4872 -2413
rect 4896 -2465 4934 -2413
rect 4934 -2465 4946 -2413
rect 4946 -2465 4952 -2413
rect 4976 -2465 4998 -2413
rect 4998 -2465 5010 -2413
rect 5010 -2465 5032 -2413
rect 5056 -2465 5062 -2413
rect 5062 -2465 5074 -2413
rect 5074 -2465 5112 -2413
rect 5136 -2465 5138 -2413
rect 5138 -2465 5190 -2413
rect 5190 -2465 5192 -2413
rect 5216 -2465 5254 -2413
rect 5254 -2465 5266 -2413
rect 5266 -2465 5272 -2413
rect 5296 -2465 5318 -2413
rect 5318 -2465 5330 -2413
rect 5330 -2465 5352 -2413
rect 5376 -2465 5382 -2413
rect 5382 -2465 5394 -2413
rect 5394 -2465 5432 -2413
rect 5456 -2465 5458 -2413
rect 5458 -2465 5510 -2413
rect 5510 -2465 5512 -2413
rect 5536 -2465 5574 -2413
rect 5574 -2465 5586 -2413
rect 5586 -2465 5592 -2413
rect 5616 -2465 5638 -2413
rect 5638 -2465 5650 -2413
rect 5650 -2465 5672 -2413
rect 5696 -2465 5702 -2413
rect 5702 -2465 5714 -2413
rect 5714 -2465 5752 -2413
rect 5776 -2465 5778 -2413
rect 5778 -2465 5830 -2413
rect 5830 -2465 5832 -2413
rect 5856 -2465 5894 -2413
rect 5894 -2465 5906 -2413
rect 5906 -2465 5912 -2413
rect 5936 -2465 5958 -2413
rect 5958 -2465 5970 -2413
rect 5970 -2465 5992 -2413
rect 6016 -2465 6022 -2413
rect 6022 -2465 6034 -2413
rect 6034 -2465 6072 -2413
rect 6096 -2465 6098 -2413
rect 6098 -2465 6150 -2413
rect 6150 -2465 6152 -2413
rect 6176 -2465 6214 -2413
rect 6214 -2465 6226 -2413
rect 6226 -2465 6232 -2413
rect 6256 -2465 6278 -2413
rect 6278 -2465 6290 -2413
rect 6290 -2465 6312 -2413
rect 6336 -2465 6342 -2413
rect 6342 -2465 6354 -2413
rect 6354 -2465 6392 -2413
rect 6416 -2465 6418 -2413
rect 6418 -2465 6470 -2413
rect 6470 -2465 6472 -2413
rect 6496 -2465 6534 -2413
rect 6534 -2465 6546 -2413
rect 6546 -2465 6552 -2413
rect 6576 -2465 6598 -2413
rect 6598 -2465 6610 -2413
rect 6610 -2465 6632 -2413
rect 6656 -2465 6662 -2413
rect 6662 -2465 6674 -2413
rect 6674 -2465 6712 -2413
rect 6736 -2465 6738 -2413
rect 6738 -2465 6790 -2413
rect 6790 -2465 6792 -2413
rect 6816 -2465 6854 -2413
rect 6854 -2465 6866 -2413
rect 6866 -2465 6872 -2413
rect 6896 -2465 6918 -2413
rect 6918 -2465 6930 -2413
rect 6930 -2465 6952 -2413
rect 6976 -2465 6982 -2413
rect 6982 -2465 6994 -2413
rect 6994 -2465 7032 -2413
rect 7056 -2465 7058 -2413
rect 7058 -2465 7110 -2413
rect 7110 -2465 7112 -2413
rect 7136 -2465 7174 -2413
rect 7174 -2465 7186 -2413
rect 7186 -2465 7192 -2413
rect 7216 -2465 7238 -2413
rect 7238 -2465 7250 -2413
rect 7250 -2465 7272 -2413
rect 7296 -2465 7302 -2413
rect 7302 -2465 7314 -2413
rect 7314 -2465 7352 -2413
rect 7376 -2465 7378 -2413
rect 7378 -2465 7430 -2413
rect 7430 -2465 7432 -2413
rect 7456 -2465 7494 -2413
rect 7494 -2465 7506 -2413
rect 7506 -2465 7512 -2413
rect 7536 -2465 7558 -2413
rect 7558 -2465 7570 -2413
rect 7570 -2465 7592 -2413
rect 7616 -2465 7622 -2413
rect 7622 -2465 7634 -2413
rect 7634 -2465 7672 -2413
rect 7696 -2465 7698 -2413
rect 7698 -2465 7750 -2413
rect 7750 -2465 7752 -2413
rect 7776 -2465 7814 -2413
rect 7814 -2465 7826 -2413
rect 7826 -2465 7832 -2413
rect 7856 -2465 7878 -2413
rect 7878 -2465 7890 -2413
rect 7890 -2465 7912 -2413
rect 7936 -2465 7942 -2413
rect 7942 -2465 7954 -2413
rect 7954 -2465 7992 -2413
rect 8016 -2465 8018 -2413
rect 8018 -2465 8070 -2413
rect 8070 -2465 8072 -2413
rect 8096 -2465 8134 -2413
rect 8134 -2465 8146 -2413
rect 8146 -2465 8152 -2413
rect 8176 -2465 8198 -2413
rect 8198 -2465 8210 -2413
rect 8210 -2465 8232 -2413
rect 8256 -2465 8262 -2413
rect 8262 -2465 8274 -2413
rect 8274 -2465 8312 -2413
rect 8336 -2465 8338 -2413
rect 8338 -2465 8390 -2413
rect 8390 -2465 8392 -2413
rect 8416 -2465 8454 -2413
rect 8454 -2465 8466 -2413
rect 8466 -2465 8472 -2413
rect 8496 -2465 8518 -2413
rect 8518 -2465 8530 -2413
rect 8530 -2465 8552 -2413
rect 8576 -2465 8582 -2413
rect 8582 -2465 8594 -2413
rect 8594 -2465 8632 -2413
rect 8656 -2465 8658 -2413
rect 8658 -2465 8710 -2413
rect 8710 -2465 8712 -2413
rect 8736 -2465 8774 -2413
rect 8774 -2465 8786 -2413
rect 8786 -2465 8792 -2413
rect 8816 -2465 8838 -2413
rect 8838 -2465 8850 -2413
rect 8850 -2465 8872 -2413
rect 8896 -2465 8902 -2413
rect 8902 -2465 8914 -2413
rect 8914 -2465 8952 -2413
rect 8976 -2465 8978 -2413
rect 8978 -2465 9030 -2413
rect 9030 -2465 9032 -2413
rect 9056 -2465 9094 -2413
rect 9094 -2465 9106 -2413
rect 9106 -2465 9112 -2413
rect 9136 -2465 9158 -2413
rect 9158 -2465 9170 -2413
rect 9170 -2465 9192 -2413
rect 9216 -2465 9222 -2413
rect 9222 -2465 9234 -2413
rect 9234 -2465 9272 -2413
rect 9296 -2465 9298 -2413
rect 9298 -2465 9350 -2413
rect 9350 -2465 9352 -2413
rect 9376 -2465 9414 -2413
rect 9414 -2465 9426 -2413
rect 9426 -2465 9432 -2413
rect 9456 -2465 9478 -2413
rect 9478 -2465 9490 -2413
rect 9490 -2465 9512 -2413
rect 9536 -2465 9542 -2413
rect 9542 -2465 9554 -2413
rect 9554 -2465 9592 -2413
rect 9616 -2465 9618 -2413
rect 9618 -2465 9670 -2413
rect 9670 -2465 9672 -2413
rect 9696 -2465 9734 -2413
rect 9734 -2465 9746 -2413
rect 9746 -2465 9752 -2413
rect 9776 -2465 9798 -2413
rect 9798 -2465 9810 -2413
rect 9810 -2465 9832 -2413
rect 9856 -2465 9862 -2413
rect 9862 -2465 9874 -2413
rect 9874 -2465 9912 -2413
rect 9936 -2465 9938 -2413
rect 9938 -2465 9990 -2413
rect 9990 -2465 9992 -2413
rect 10016 -2465 10054 -2413
rect 10054 -2465 10066 -2413
rect 10066 -2465 10072 -2413
rect 10096 -2465 10118 -2413
rect 10118 -2465 10130 -2413
rect 10130 -2465 10152 -2413
rect 10176 -2465 10182 -2413
rect 10182 -2465 10194 -2413
rect 10194 -2465 10232 -2413
rect 10256 -2465 10258 -2413
rect 10258 -2465 10310 -2413
rect 10310 -2465 10312 -2413
rect 10336 -2465 10374 -2413
rect 10374 -2465 10386 -2413
rect 10386 -2465 10392 -2413
rect 10416 -2465 10438 -2413
rect 10438 -2465 10450 -2413
rect 10450 -2465 10472 -2413
rect 10496 -2465 10502 -2413
rect 10502 -2465 10514 -2413
rect 10514 -2465 10552 -2413
rect 10576 -2465 10578 -2413
rect 10578 -2465 10630 -2413
rect 10630 -2465 10632 -2413
rect 16 -2467 72 -2465
rect 96 -2467 152 -2465
rect 176 -2467 232 -2465
rect 256 -2467 312 -2465
rect 336 -2467 392 -2465
rect 416 -2467 472 -2465
rect 496 -2467 552 -2465
rect 576 -2467 632 -2465
rect 656 -2467 712 -2465
rect 736 -2467 792 -2465
rect 816 -2467 872 -2465
rect 896 -2467 952 -2465
rect 976 -2467 1032 -2465
rect 1056 -2467 1112 -2465
rect 1136 -2467 1192 -2465
rect 1216 -2467 1272 -2465
rect 1296 -2467 1352 -2465
rect 1376 -2467 1432 -2465
rect 1456 -2467 1512 -2465
rect 1536 -2467 1592 -2465
rect 1616 -2467 1672 -2465
rect 1696 -2467 1752 -2465
rect 1776 -2467 1832 -2465
rect 1856 -2467 1912 -2465
rect 1936 -2467 1992 -2465
rect 2016 -2467 2072 -2465
rect 2096 -2467 2152 -2465
rect 2176 -2467 2232 -2465
rect 2256 -2467 2312 -2465
rect 2336 -2467 2392 -2465
rect 2416 -2467 2472 -2465
rect 2496 -2467 2552 -2465
rect 2576 -2467 2632 -2465
rect 2656 -2467 2712 -2465
rect 2736 -2467 2792 -2465
rect 2816 -2467 2872 -2465
rect 2896 -2467 2952 -2465
rect 2976 -2467 3032 -2465
rect 3056 -2467 3112 -2465
rect 3136 -2467 3192 -2465
rect 3216 -2467 3272 -2465
rect 3296 -2467 3352 -2465
rect 3376 -2467 3432 -2465
rect 3456 -2467 3512 -2465
rect 3536 -2467 3592 -2465
rect 3616 -2467 3672 -2465
rect 3696 -2467 3752 -2465
rect 3776 -2467 3832 -2465
rect 3856 -2467 3912 -2465
rect 3936 -2467 3992 -2465
rect 4016 -2467 4072 -2465
rect 4096 -2467 4152 -2465
rect 4176 -2467 4232 -2465
rect 4256 -2467 4312 -2465
rect 4336 -2467 4392 -2465
rect 4416 -2467 4472 -2465
rect 4496 -2467 4552 -2465
rect 4576 -2467 4632 -2465
rect 4656 -2467 4712 -2465
rect 4736 -2467 4792 -2465
rect 4816 -2467 4872 -2465
rect 4896 -2467 4952 -2465
rect 4976 -2467 5032 -2465
rect 5056 -2467 5112 -2465
rect 5136 -2467 5192 -2465
rect 5216 -2467 5272 -2465
rect 5296 -2467 5352 -2465
rect 5376 -2467 5432 -2465
rect 5456 -2467 5512 -2465
rect 5536 -2467 5592 -2465
rect 5616 -2467 5672 -2465
rect 5696 -2467 5752 -2465
rect 5776 -2467 5832 -2465
rect 5856 -2467 5912 -2465
rect 5936 -2467 5992 -2465
rect 6016 -2467 6072 -2465
rect 6096 -2467 6152 -2465
rect 6176 -2467 6232 -2465
rect 6256 -2467 6312 -2465
rect 6336 -2467 6392 -2465
rect 6416 -2467 6472 -2465
rect 6496 -2467 6552 -2465
rect 6576 -2467 6632 -2465
rect 6656 -2467 6712 -2465
rect 6736 -2467 6792 -2465
rect 6816 -2467 6872 -2465
rect 6896 -2467 6952 -2465
rect 6976 -2467 7032 -2465
rect 7056 -2467 7112 -2465
rect 7136 -2467 7192 -2465
rect 7216 -2467 7272 -2465
rect 7296 -2467 7352 -2465
rect 7376 -2467 7432 -2465
rect 7456 -2467 7512 -2465
rect 7536 -2467 7592 -2465
rect 7616 -2467 7672 -2465
rect 7696 -2467 7752 -2465
rect 7776 -2467 7832 -2465
rect 7856 -2467 7912 -2465
rect 7936 -2467 7992 -2465
rect 8016 -2467 8072 -2465
rect 8096 -2467 8152 -2465
rect 8176 -2467 8232 -2465
rect 8256 -2467 8312 -2465
rect 8336 -2467 8392 -2465
rect 8416 -2467 8472 -2465
rect 8496 -2467 8552 -2465
rect 8576 -2467 8632 -2465
rect 8656 -2467 8712 -2465
rect 8736 -2467 8792 -2465
rect 8816 -2467 8872 -2465
rect 8896 -2467 8952 -2465
rect 8976 -2467 9032 -2465
rect 9056 -2467 9112 -2465
rect 9136 -2467 9192 -2465
rect 9216 -2467 9272 -2465
rect 9296 -2467 9352 -2465
rect 9376 -2467 9432 -2465
rect 9456 -2467 9512 -2465
rect 9536 -2467 9592 -2465
rect 9616 -2467 9672 -2465
rect 9696 -2467 9752 -2465
rect 9776 -2467 9832 -2465
rect 9856 -2467 9912 -2465
rect 9936 -2467 9992 -2465
rect 10016 -2467 10072 -2465
rect 10096 -2467 10152 -2465
rect 10176 -2467 10232 -2465
rect 10256 -2467 10312 -2465
rect 10336 -2467 10392 -2465
rect 10416 -2467 10472 -2465
rect 10496 -2467 10552 -2465
rect 10576 -2467 10632 -2465
rect -184 -2644 352 -2618
rect -184 -2888 352 -2644
rect -184 -2914 352 -2888
rect 10348 -2644 10884 -2618
rect 10348 -2888 10884 -2644
rect 10348 -2914 10884 -2888
<< metal3 >>
rect -226 2294 394 2301
rect -226 2258 -184 2294
rect 352 2258 394 2294
rect -226 2034 -188 2258
rect 356 2034 394 2258
rect -226 1998 -184 2034
rect 352 1998 394 2034
rect -226 1991 394 1998
rect 10306 2294 10926 2301
rect 10306 2258 10348 2294
rect 10884 2258 10926 2294
rect 10306 2034 10344 2258
rect 10888 2034 10926 2258
rect 10306 1998 10348 2034
rect 10884 1998 10926 2034
rect 10306 1991 10926 1998
rect 3466 1906 7322 1950
rect 3466 1762 3524 1906
rect 7268 1762 7322 1906
rect 3466 1720 7322 1762
rect 3628 -840 7786 -820
rect 3628 -896 3658 -840
rect 3714 -896 7706 -840
rect 7762 -896 7786 -840
rect 3628 -920 7786 -896
rect -66 -2407 10708 -2336
rect -66 -2471 12 -2407
rect 76 -2471 92 -2407
rect 156 -2471 172 -2407
rect 236 -2471 252 -2407
rect 316 -2471 332 -2407
rect 396 -2471 412 -2407
rect 476 -2471 492 -2407
rect 556 -2471 572 -2407
rect 636 -2471 652 -2407
rect 716 -2471 732 -2407
rect 796 -2471 812 -2407
rect 876 -2471 892 -2407
rect 956 -2471 972 -2407
rect 1036 -2471 1052 -2407
rect 1116 -2471 1132 -2407
rect 1196 -2471 1212 -2407
rect 1276 -2471 1292 -2407
rect 1356 -2471 1372 -2407
rect 1436 -2471 1452 -2407
rect 1516 -2471 1532 -2407
rect 1596 -2471 1612 -2407
rect 1676 -2471 1692 -2407
rect 1756 -2471 1772 -2407
rect 1836 -2471 1852 -2407
rect 1916 -2471 1932 -2407
rect 1996 -2471 2012 -2407
rect 2076 -2471 2092 -2407
rect 2156 -2471 2172 -2407
rect 2236 -2471 2252 -2407
rect 2316 -2471 2332 -2407
rect 2396 -2471 2412 -2407
rect 2476 -2471 2492 -2407
rect 2556 -2471 2572 -2407
rect 2636 -2471 2652 -2407
rect 2716 -2471 2732 -2407
rect 2796 -2471 2812 -2407
rect 2876 -2471 2892 -2407
rect 2956 -2471 2972 -2407
rect 3036 -2471 3052 -2407
rect 3116 -2471 3132 -2407
rect 3196 -2471 3212 -2407
rect 3276 -2471 3292 -2407
rect 3356 -2471 3372 -2407
rect 3436 -2471 3452 -2407
rect 3516 -2471 3532 -2407
rect 3596 -2471 3612 -2407
rect 3676 -2471 3692 -2407
rect 3756 -2471 3772 -2407
rect 3836 -2471 3852 -2407
rect 3916 -2471 3932 -2407
rect 3996 -2471 4012 -2407
rect 4076 -2471 4092 -2407
rect 4156 -2471 4172 -2407
rect 4236 -2471 4252 -2407
rect 4316 -2471 4332 -2407
rect 4396 -2471 4412 -2407
rect 4476 -2471 4492 -2407
rect 4556 -2471 4572 -2407
rect 4636 -2471 4652 -2407
rect 4716 -2471 4732 -2407
rect 4796 -2471 4812 -2407
rect 4876 -2471 4892 -2407
rect 4956 -2471 4972 -2407
rect 5036 -2471 5052 -2407
rect 5116 -2471 5132 -2407
rect 5196 -2471 5212 -2407
rect 5276 -2471 5292 -2407
rect 5356 -2471 5372 -2407
rect 5436 -2471 5452 -2407
rect 5516 -2471 5532 -2407
rect 5596 -2471 5612 -2407
rect 5676 -2471 5692 -2407
rect 5756 -2471 5772 -2407
rect 5836 -2471 5852 -2407
rect 5916 -2471 5932 -2407
rect 5996 -2471 6012 -2407
rect 6076 -2471 6092 -2407
rect 6156 -2471 6172 -2407
rect 6236 -2471 6252 -2407
rect 6316 -2471 6332 -2407
rect 6396 -2471 6412 -2407
rect 6476 -2471 6492 -2407
rect 6556 -2471 6572 -2407
rect 6636 -2471 6652 -2407
rect 6716 -2471 6732 -2407
rect 6796 -2471 6812 -2407
rect 6876 -2471 6892 -2407
rect 6956 -2471 6972 -2407
rect 7036 -2471 7052 -2407
rect 7116 -2471 7132 -2407
rect 7196 -2471 7212 -2407
rect 7276 -2471 7292 -2407
rect 7356 -2471 7372 -2407
rect 7436 -2471 7452 -2407
rect 7516 -2471 7532 -2407
rect 7596 -2471 7612 -2407
rect 7676 -2471 7692 -2407
rect 7756 -2471 7772 -2407
rect 7836 -2471 7852 -2407
rect 7916 -2471 7932 -2407
rect 7996 -2471 8012 -2407
rect 8076 -2471 8092 -2407
rect 8156 -2471 8172 -2407
rect 8236 -2471 8252 -2407
rect 8316 -2471 8332 -2407
rect 8396 -2471 8412 -2407
rect 8476 -2471 8492 -2407
rect 8556 -2471 8572 -2407
rect 8636 -2471 8652 -2407
rect 8716 -2471 8732 -2407
rect 8796 -2471 8812 -2407
rect 8876 -2471 8892 -2407
rect 8956 -2471 8972 -2407
rect 9036 -2471 9052 -2407
rect 9116 -2471 9132 -2407
rect 9196 -2471 9212 -2407
rect 9276 -2471 9292 -2407
rect 9356 -2471 9372 -2407
rect 9436 -2471 9452 -2407
rect 9516 -2471 9532 -2407
rect 9596 -2471 9612 -2407
rect 9676 -2471 9692 -2407
rect 9756 -2471 9772 -2407
rect 9836 -2471 9852 -2407
rect 9916 -2471 9932 -2407
rect 9996 -2471 10012 -2407
rect 10076 -2471 10092 -2407
rect 10156 -2471 10172 -2407
rect 10236 -2471 10252 -2407
rect 10316 -2471 10332 -2407
rect 10396 -2471 10412 -2407
rect 10476 -2471 10492 -2407
rect 10556 -2471 10572 -2407
rect 10636 -2471 10708 -2407
rect -66 -2550 10708 -2471
rect -226 -2618 394 -2611
rect -226 -2654 -184 -2618
rect 352 -2654 394 -2618
rect -226 -2878 -188 -2654
rect 356 -2878 394 -2654
rect -226 -2914 -184 -2878
rect 352 -2914 394 -2878
rect -226 -2921 394 -2914
rect 10306 -2618 10926 -2611
rect 10306 -2654 10348 -2618
rect 10884 -2654 10926 -2618
rect 10306 -2878 10344 -2654
rect 10888 -2878 10926 -2654
rect 10306 -2914 10348 -2878
rect 10884 -2914 10926 -2878
rect 10306 -2921 10926 -2914
<< via3 >>
rect -188 2034 -184 2258
rect -184 2034 352 2258
rect 352 2034 356 2258
rect 10344 2034 10348 2258
rect 10348 2034 10884 2258
rect 10884 2034 10888 2258
rect 3524 1902 7268 1906
rect 3524 1766 3528 1902
rect 3528 1766 7264 1902
rect 7264 1766 7268 1902
rect 3524 1762 7268 1766
rect 12 -2411 76 -2407
rect 12 -2467 16 -2411
rect 16 -2467 72 -2411
rect 72 -2467 76 -2411
rect 12 -2471 76 -2467
rect 92 -2411 156 -2407
rect 92 -2467 96 -2411
rect 96 -2467 152 -2411
rect 152 -2467 156 -2411
rect 92 -2471 156 -2467
rect 172 -2411 236 -2407
rect 172 -2467 176 -2411
rect 176 -2467 232 -2411
rect 232 -2467 236 -2411
rect 172 -2471 236 -2467
rect 252 -2411 316 -2407
rect 252 -2467 256 -2411
rect 256 -2467 312 -2411
rect 312 -2467 316 -2411
rect 252 -2471 316 -2467
rect 332 -2411 396 -2407
rect 332 -2467 336 -2411
rect 336 -2467 392 -2411
rect 392 -2467 396 -2411
rect 332 -2471 396 -2467
rect 412 -2411 476 -2407
rect 412 -2467 416 -2411
rect 416 -2467 472 -2411
rect 472 -2467 476 -2411
rect 412 -2471 476 -2467
rect 492 -2411 556 -2407
rect 492 -2467 496 -2411
rect 496 -2467 552 -2411
rect 552 -2467 556 -2411
rect 492 -2471 556 -2467
rect 572 -2411 636 -2407
rect 572 -2467 576 -2411
rect 576 -2467 632 -2411
rect 632 -2467 636 -2411
rect 572 -2471 636 -2467
rect 652 -2411 716 -2407
rect 652 -2467 656 -2411
rect 656 -2467 712 -2411
rect 712 -2467 716 -2411
rect 652 -2471 716 -2467
rect 732 -2411 796 -2407
rect 732 -2467 736 -2411
rect 736 -2467 792 -2411
rect 792 -2467 796 -2411
rect 732 -2471 796 -2467
rect 812 -2411 876 -2407
rect 812 -2467 816 -2411
rect 816 -2467 872 -2411
rect 872 -2467 876 -2411
rect 812 -2471 876 -2467
rect 892 -2411 956 -2407
rect 892 -2467 896 -2411
rect 896 -2467 952 -2411
rect 952 -2467 956 -2411
rect 892 -2471 956 -2467
rect 972 -2411 1036 -2407
rect 972 -2467 976 -2411
rect 976 -2467 1032 -2411
rect 1032 -2467 1036 -2411
rect 972 -2471 1036 -2467
rect 1052 -2411 1116 -2407
rect 1052 -2467 1056 -2411
rect 1056 -2467 1112 -2411
rect 1112 -2467 1116 -2411
rect 1052 -2471 1116 -2467
rect 1132 -2411 1196 -2407
rect 1132 -2467 1136 -2411
rect 1136 -2467 1192 -2411
rect 1192 -2467 1196 -2411
rect 1132 -2471 1196 -2467
rect 1212 -2411 1276 -2407
rect 1212 -2467 1216 -2411
rect 1216 -2467 1272 -2411
rect 1272 -2467 1276 -2411
rect 1212 -2471 1276 -2467
rect 1292 -2411 1356 -2407
rect 1292 -2467 1296 -2411
rect 1296 -2467 1352 -2411
rect 1352 -2467 1356 -2411
rect 1292 -2471 1356 -2467
rect 1372 -2411 1436 -2407
rect 1372 -2467 1376 -2411
rect 1376 -2467 1432 -2411
rect 1432 -2467 1436 -2411
rect 1372 -2471 1436 -2467
rect 1452 -2411 1516 -2407
rect 1452 -2467 1456 -2411
rect 1456 -2467 1512 -2411
rect 1512 -2467 1516 -2411
rect 1452 -2471 1516 -2467
rect 1532 -2411 1596 -2407
rect 1532 -2467 1536 -2411
rect 1536 -2467 1592 -2411
rect 1592 -2467 1596 -2411
rect 1532 -2471 1596 -2467
rect 1612 -2411 1676 -2407
rect 1612 -2467 1616 -2411
rect 1616 -2467 1672 -2411
rect 1672 -2467 1676 -2411
rect 1612 -2471 1676 -2467
rect 1692 -2411 1756 -2407
rect 1692 -2467 1696 -2411
rect 1696 -2467 1752 -2411
rect 1752 -2467 1756 -2411
rect 1692 -2471 1756 -2467
rect 1772 -2411 1836 -2407
rect 1772 -2467 1776 -2411
rect 1776 -2467 1832 -2411
rect 1832 -2467 1836 -2411
rect 1772 -2471 1836 -2467
rect 1852 -2411 1916 -2407
rect 1852 -2467 1856 -2411
rect 1856 -2467 1912 -2411
rect 1912 -2467 1916 -2411
rect 1852 -2471 1916 -2467
rect 1932 -2411 1996 -2407
rect 1932 -2467 1936 -2411
rect 1936 -2467 1992 -2411
rect 1992 -2467 1996 -2411
rect 1932 -2471 1996 -2467
rect 2012 -2411 2076 -2407
rect 2012 -2467 2016 -2411
rect 2016 -2467 2072 -2411
rect 2072 -2467 2076 -2411
rect 2012 -2471 2076 -2467
rect 2092 -2411 2156 -2407
rect 2092 -2467 2096 -2411
rect 2096 -2467 2152 -2411
rect 2152 -2467 2156 -2411
rect 2092 -2471 2156 -2467
rect 2172 -2411 2236 -2407
rect 2172 -2467 2176 -2411
rect 2176 -2467 2232 -2411
rect 2232 -2467 2236 -2411
rect 2172 -2471 2236 -2467
rect 2252 -2411 2316 -2407
rect 2252 -2467 2256 -2411
rect 2256 -2467 2312 -2411
rect 2312 -2467 2316 -2411
rect 2252 -2471 2316 -2467
rect 2332 -2411 2396 -2407
rect 2332 -2467 2336 -2411
rect 2336 -2467 2392 -2411
rect 2392 -2467 2396 -2411
rect 2332 -2471 2396 -2467
rect 2412 -2411 2476 -2407
rect 2412 -2467 2416 -2411
rect 2416 -2467 2472 -2411
rect 2472 -2467 2476 -2411
rect 2412 -2471 2476 -2467
rect 2492 -2411 2556 -2407
rect 2492 -2467 2496 -2411
rect 2496 -2467 2552 -2411
rect 2552 -2467 2556 -2411
rect 2492 -2471 2556 -2467
rect 2572 -2411 2636 -2407
rect 2572 -2467 2576 -2411
rect 2576 -2467 2632 -2411
rect 2632 -2467 2636 -2411
rect 2572 -2471 2636 -2467
rect 2652 -2411 2716 -2407
rect 2652 -2467 2656 -2411
rect 2656 -2467 2712 -2411
rect 2712 -2467 2716 -2411
rect 2652 -2471 2716 -2467
rect 2732 -2411 2796 -2407
rect 2732 -2467 2736 -2411
rect 2736 -2467 2792 -2411
rect 2792 -2467 2796 -2411
rect 2732 -2471 2796 -2467
rect 2812 -2411 2876 -2407
rect 2812 -2467 2816 -2411
rect 2816 -2467 2872 -2411
rect 2872 -2467 2876 -2411
rect 2812 -2471 2876 -2467
rect 2892 -2411 2956 -2407
rect 2892 -2467 2896 -2411
rect 2896 -2467 2952 -2411
rect 2952 -2467 2956 -2411
rect 2892 -2471 2956 -2467
rect 2972 -2411 3036 -2407
rect 2972 -2467 2976 -2411
rect 2976 -2467 3032 -2411
rect 3032 -2467 3036 -2411
rect 2972 -2471 3036 -2467
rect 3052 -2411 3116 -2407
rect 3052 -2467 3056 -2411
rect 3056 -2467 3112 -2411
rect 3112 -2467 3116 -2411
rect 3052 -2471 3116 -2467
rect 3132 -2411 3196 -2407
rect 3132 -2467 3136 -2411
rect 3136 -2467 3192 -2411
rect 3192 -2467 3196 -2411
rect 3132 -2471 3196 -2467
rect 3212 -2411 3276 -2407
rect 3212 -2467 3216 -2411
rect 3216 -2467 3272 -2411
rect 3272 -2467 3276 -2411
rect 3212 -2471 3276 -2467
rect 3292 -2411 3356 -2407
rect 3292 -2467 3296 -2411
rect 3296 -2467 3352 -2411
rect 3352 -2467 3356 -2411
rect 3292 -2471 3356 -2467
rect 3372 -2411 3436 -2407
rect 3372 -2467 3376 -2411
rect 3376 -2467 3432 -2411
rect 3432 -2467 3436 -2411
rect 3372 -2471 3436 -2467
rect 3452 -2411 3516 -2407
rect 3452 -2467 3456 -2411
rect 3456 -2467 3512 -2411
rect 3512 -2467 3516 -2411
rect 3452 -2471 3516 -2467
rect 3532 -2411 3596 -2407
rect 3532 -2467 3536 -2411
rect 3536 -2467 3592 -2411
rect 3592 -2467 3596 -2411
rect 3532 -2471 3596 -2467
rect 3612 -2411 3676 -2407
rect 3612 -2467 3616 -2411
rect 3616 -2467 3672 -2411
rect 3672 -2467 3676 -2411
rect 3612 -2471 3676 -2467
rect 3692 -2411 3756 -2407
rect 3692 -2467 3696 -2411
rect 3696 -2467 3752 -2411
rect 3752 -2467 3756 -2411
rect 3692 -2471 3756 -2467
rect 3772 -2411 3836 -2407
rect 3772 -2467 3776 -2411
rect 3776 -2467 3832 -2411
rect 3832 -2467 3836 -2411
rect 3772 -2471 3836 -2467
rect 3852 -2411 3916 -2407
rect 3852 -2467 3856 -2411
rect 3856 -2467 3912 -2411
rect 3912 -2467 3916 -2411
rect 3852 -2471 3916 -2467
rect 3932 -2411 3996 -2407
rect 3932 -2467 3936 -2411
rect 3936 -2467 3992 -2411
rect 3992 -2467 3996 -2411
rect 3932 -2471 3996 -2467
rect 4012 -2411 4076 -2407
rect 4012 -2467 4016 -2411
rect 4016 -2467 4072 -2411
rect 4072 -2467 4076 -2411
rect 4012 -2471 4076 -2467
rect 4092 -2411 4156 -2407
rect 4092 -2467 4096 -2411
rect 4096 -2467 4152 -2411
rect 4152 -2467 4156 -2411
rect 4092 -2471 4156 -2467
rect 4172 -2411 4236 -2407
rect 4172 -2467 4176 -2411
rect 4176 -2467 4232 -2411
rect 4232 -2467 4236 -2411
rect 4172 -2471 4236 -2467
rect 4252 -2411 4316 -2407
rect 4252 -2467 4256 -2411
rect 4256 -2467 4312 -2411
rect 4312 -2467 4316 -2411
rect 4252 -2471 4316 -2467
rect 4332 -2411 4396 -2407
rect 4332 -2467 4336 -2411
rect 4336 -2467 4392 -2411
rect 4392 -2467 4396 -2411
rect 4332 -2471 4396 -2467
rect 4412 -2411 4476 -2407
rect 4412 -2467 4416 -2411
rect 4416 -2467 4472 -2411
rect 4472 -2467 4476 -2411
rect 4412 -2471 4476 -2467
rect 4492 -2411 4556 -2407
rect 4492 -2467 4496 -2411
rect 4496 -2467 4552 -2411
rect 4552 -2467 4556 -2411
rect 4492 -2471 4556 -2467
rect 4572 -2411 4636 -2407
rect 4572 -2467 4576 -2411
rect 4576 -2467 4632 -2411
rect 4632 -2467 4636 -2411
rect 4572 -2471 4636 -2467
rect 4652 -2411 4716 -2407
rect 4652 -2467 4656 -2411
rect 4656 -2467 4712 -2411
rect 4712 -2467 4716 -2411
rect 4652 -2471 4716 -2467
rect 4732 -2411 4796 -2407
rect 4732 -2467 4736 -2411
rect 4736 -2467 4792 -2411
rect 4792 -2467 4796 -2411
rect 4732 -2471 4796 -2467
rect 4812 -2411 4876 -2407
rect 4812 -2467 4816 -2411
rect 4816 -2467 4872 -2411
rect 4872 -2467 4876 -2411
rect 4812 -2471 4876 -2467
rect 4892 -2411 4956 -2407
rect 4892 -2467 4896 -2411
rect 4896 -2467 4952 -2411
rect 4952 -2467 4956 -2411
rect 4892 -2471 4956 -2467
rect 4972 -2411 5036 -2407
rect 4972 -2467 4976 -2411
rect 4976 -2467 5032 -2411
rect 5032 -2467 5036 -2411
rect 4972 -2471 5036 -2467
rect 5052 -2411 5116 -2407
rect 5052 -2467 5056 -2411
rect 5056 -2467 5112 -2411
rect 5112 -2467 5116 -2411
rect 5052 -2471 5116 -2467
rect 5132 -2411 5196 -2407
rect 5132 -2467 5136 -2411
rect 5136 -2467 5192 -2411
rect 5192 -2467 5196 -2411
rect 5132 -2471 5196 -2467
rect 5212 -2411 5276 -2407
rect 5212 -2467 5216 -2411
rect 5216 -2467 5272 -2411
rect 5272 -2467 5276 -2411
rect 5212 -2471 5276 -2467
rect 5292 -2411 5356 -2407
rect 5292 -2467 5296 -2411
rect 5296 -2467 5352 -2411
rect 5352 -2467 5356 -2411
rect 5292 -2471 5356 -2467
rect 5372 -2411 5436 -2407
rect 5372 -2467 5376 -2411
rect 5376 -2467 5432 -2411
rect 5432 -2467 5436 -2411
rect 5372 -2471 5436 -2467
rect 5452 -2411 5516 -2407
rect 5452 -2467 5456 -2411
rect 5456 -2467 5512 -2411
rect 5512 -2467 5516 -2411
rect 5452 -2471 5516 -2467
rect 5532 -2411 5596 -2407
rect 5532 -2467 5536 -2411
rect 5536 -2467 5592 -2411
rect 5592 -2467 5596 -2411
rect 5532 -2471 5596 -2467
rect 5612 -2411 5676 -2407
rect 5612 -2467 5616 -2411
rect 5616 -2467 5672 -2411
rect 5672 -2467 5676 -2411
rect 5612 -2471 5676 -2467
rect 5692 -2411 5756 -2407
rect 5692 -2467 5696 -2411
rect 5696 -2467 5752 -2411
rect 5752 -2467 5756 -2411
rect 5692 -2471 5756 -2467
rect 5772 -2411 5836 -2407
rect 5772 -2467 5776 -2411
rect 5776 -2467 5832 -2411
rect 5832 -2467 5836 -2411
rect 5772 -2471 5836 -2467
rect 5852 -2411 5916 -2407
rect 5852 -2467 5856 -2411
rect 5856 -2467 5912 -2411
rect 5912 -2467 5916 -2411
rect 5852 -2471 5916 -2467
rect 5932 -2411 5996 -2407
rect 5932 -2467 5936 -2411
rect 5936 -2467 5992 -2411
rect 5992 -2467 5996 -2411
rect 5932 -2471 5996 -2467
rect 6012 -2411 6076 -2407
rect 6012 -2467 6016 -2411
rect 6016 -2467 6072 -2411
rect 6072 -2467 6076 -2411
rect 6012 -2471 6076 -2467
rect 6092 -2411 6156 -2407
rect 6092 -2467 6096 -2411
rect 6096 -2467 6152 -2411
rect 6152 -2467 6156 -2411
rect 6092 -2471 6156 -2467
rect 6172 -2411 6236 -2407
rect 6172 -2467 6176 -2411
rect 6176 -2467 6232 -2411
rect 6232 -2467 6236 -2411
rect 6172 -2471 6236 -2467
rect 6252 -2411 6316 -2407
rect 6252 -2467 6256 -2411
rect 6256 -2467 6312 -2411
rect 6312 -2467 6316 -2411
rect 6252 -2471 6316 -2467
rect 6332 -2411 6396 -2407
rect 6332 -2467 6336 -2411
rect 6336 -2467 6392 -2411
rect 6392 -2467 6396 -2411
rect 6332 -2471 6396 -2467
rect 6412 -2411 6476 -2407
rect 6412 -2467 6416 -2411
rect 6416 -2467 6472 -2411
rect 6472 -2467 6476 -2411
rect 6412 -2471 6476 -2467
rect 6492 -2411 6556 -2407
rect 6492 -2467 6496 -2411
rect 6496 -2467 6552 -2411
rect 6552 -2467 6556 -2411
rect 6492 -2471 6556 -2467
rect 6572 -2411 6636 -2407
rect 6572 -2467 6576 -2411
rect 6576 -2467 6632 -2411
rect 6632 -2467 6636 -2411
rect 6572 -2471 6636 -2467
rect 6652 -2411 6716 -2407
rect 6652 -2467 6656 -2411
rect 6656 -2467 6712 -2411
rect 6712 -2467 6716 -2411
rect 6652 -2471 6716 -2467
rect 6732 -2411 6796 -2407
rect 6732 -2467 6736 -2411
rect 6736 -2467 6792 -2411
rect 6792 -2467 6796 -2411
rect 6732 -2471 6796 -2467
rect 6812 -2411 6876 -2407
rect 6812 -2467 6816 -2411
rect 6816 -2467 6872 -2411
rect 6872 -2467 6876 -2411
rect 6812 -2471 6876 -2467
rect 6892 -2411 6956 -2407
rect 6892 -2467 6896 -2411
rect 6896 -2467 6952 -2411
rect 6952 -2467 6956 -2411
rect 6892 -2471 6956 -2467
rect 6972 -2411 7036 -2407
rect 6972 -2467 6976 -2411
rect 6976 -2467 7032 -2411
rect 7032 -2467 7036 -2411
rect 6972 -2471 7036 -2467
rect 7052 -2411 7116 -2407
rect 7052 -2467 7056 -2411
rect 7056 -2467 7112 -2411
rect 7112 -2467 7116 -2411
rect 7052 -2471 7116 -2467
rect 7132 -2411 7196 -2407
rect 7132 -2467 7136 -2411
rect 7136 -2467 7192 -2411
rect 7192 -2467 7196 -2411
rect 7132 -2471 7196 -2467
rect 7212 -2411 7276 -2407
rect 7212 -2467 7216 -2411
rect 7216 -2467 7272 -2411
rect 7272 -2467 7276 -2411
rect 7212 -2471 7276 -2467
rect 7292 -2411 7356 -2407
rect 7292 -2467 7296 -2411
rect 7296 -2467 7352 -2411
rect 7352 -2467 7356 -2411
rect 7292 -2471 7356 -2467
rect 7372 -2411 7436 -2407
rect 7372 -2467 7376 -2411
rect 7376 -2467 7432 -2411
rect 7432 -2467 7436 -2411
rect 7372 -2471 7436 -2467
rect 7452 -2411 7516 -2407
rect 7452 -2467 7456 -2411
rect 7456 -2467 7512 -2411
rect 7512 -2467 7516 -2411
rect 7452 -2471 7516 -2467
rect 7532 -2411 7596 -2407
rect 7532 -2467 7536 -2411
rect 7536 -2467 7592 -2411
rect 7592 -2467 7596 -2411
rect 7532 -2471 7596 -2467
rect 7612 -2411 7676 -2407
rect 7612 -2467 7616 -2411
rect 7616 -2467 7672 -2411
rect 7672 -2467 7676 -2411
rect 7612 -2471 7676 -2467
rect 7692 -2411 7756 -2407
rect 7692 -2467 7696 -2411
rect 7696 -2467 7752 -2411
rect 7752 -2467 7756 -2411
rect 7692 -2471 7756 -2467
rect 7772 -2411 7836 -2407
rect 7772 -2467 7776 -2411
rect 7776 -2467 7832 -2411
rect 7832 -2467 7836 -2411
rect 7772 -2471 7836 -2467
rect 7852 -2411 7916 -2407
rect 7852 -2467 7856 -2411
rect 7856 -2467 7912 -2411
rect 7912 -2467 7916 -2411
rect 7852 -2471 7916 -2467
rect 7932 -2411 7996 -2407
rect 7932 -2467 7936 -2411
rect 7936 -2467 7992 -2411
rect 7992 -2467 7996 -2411
rect 7932 -2471 7996 -2467
rect 8012 -2411 8076 -2407
rect 8012 -2467 8016 -2411
rect 8016 -2467 8072 -2411
rect 8072 -2467 8076 -2411
rect 8012 -2471 8076 -2467
rect 8092 -2411 8156 -2407
rect 8092 -2467 8096 -2411
rect 8096 -2467 8152 -2411
rect 8152 -2467 8156 -2411
rect 8092 -2471 8156 -2467
rect 8172 -2411 8236 -2407
rect 8172 -2467 8176 -2411
rect 8176 -2467 8232 -2411
rect 8232 -2467 8236 -2411
rect 8172 -2471 8236 -2467
rect 8252 -2411 8316 -2407
rect 8252 -2467 8256 -2411
rect 8256 -2467 8312 -2411
rect 8312 -2467 8316 -2411
rect 8252 -2471 8316 -2467
rect 8332 -2411 8396 -2407
rect 8332 -2467 8336 -2411
rect 8336 -2467 8392 -2411
rect 8392 -2467 8396 -2411
rect 8332 -2471 8396 -2467
rect 8412 -2411 8476 -2407
rect 8412 -2467 8416 -2411
rect 8416 -2467 8472 -2411
rect 8472 -2467 8476 -2411
rect 8412 -2471 8476 -2467
rect 8492 -2411 8556 -2407
rect 8492 -2467 8496 -2411
rect 8496 -2467 8552 -2411
rect 8552 -2467 8556 -2411
rect 8492 -2471 8556 -2467
rect 8572 -2411 8636 -2407
rect 8572 -2467 8576 -2411
rect 8576 -2467 8632 -2411
rect 8632 -2467 8636 -2411
rect 8572 -2471 8636 -2467
rect 8652 -2411 8716 -2407
rect 8652 -2467 8656 -2411
rect 8656 -2467 8712 -2411
rect 8712 -2467 8716 -2411
rect 8652 -2471 8716 -2467
rect 8732 -2411 8796 -2407
rect 8732 -2467 8736 -2411
rect 8736 -2467 8792 -2411
rect 8792 -2467 8796 -2411
rect 8732 -2471 8796 -2467
rect 8812 -2411 8876 -2407
rect 8812 -2467 8816 -2411
rect 8816 -2467 8872 -2411
rect 8872 -2467 8876 -2411
rect 8812 -2471 8876 -2467
rect 8892 -2411 8956 -2407
rect 8892 -2467 8896 -2411
rect 8896 -2467 8952 -2411
rect 8952 -2467 8956 -2411
rect 8892 -2471 8956 -2467
rect 8972 -2411 9036 -2407
rect 8972 -2467 8976 -2411
rect 8976 -2467 9032 -2411
rect 9032 -2467 9036 -2411
rect 8972 -2471 9036 -2467
rect 9052 -2411 9116 -2407
rect 9052 -2467 9056 -2411
rect 9056 -2467 9112 -2411
rect 9112 -2467 9116 -2411
rect 9052 -2471 9116 -2467
rect 9132 -2411 9196 -2407
rect 9132 -2467 9136 -2411
rect 9136 -2467 9192 -2411
rect 9192 -2467 9196 -2411
rect 9132 -2471 9196 -2467
rect 9212 -2411 9276 -2407
rect 9212 -2467 9216 -2411
rect 9216 -2467 9272 -2411
rect 9272 -2467 9276 -2411
rect 9212 -2471 9276 -2467
rect 9292 -2411 9356 -2407
rect 9292 -2467 9296 -2411
rect 9296 -2467 9352 -2411
rect 9352 -2467 9356 -2411
rect 9292 -2471 9356 -2467
rect 9372 -2411 9436 -2407
rect 9372 -2467 9376 -2411
rect 9376 -2467 9432 -2411
rect 9432 -2467 9436 -2411
rect 9372 -2471 9436 -2467
rect 9452 -2411 9516 -2407
rect 9452 -2467 9456 -2411
rect 9456 -2467 9512 -2411
rect 9512 -2467 9516 -2411
rect 9452 -2471 9516 -2467
rect 9532 -2411 9596 -2407
rect 9532 -2467 9536 -2411
rect 9536 -2467 9592 -2411
rect 9592 -2467 9596 -2411
rect 9532 -2471 9596 -2467
rect 9612 -2411 9676 -2407
rect 9612 -2467 9616 -2411
rect 9616 -2467 9672 -2411
rect 9672 -2467 9676 -2411
rect 9612 -2471 9676 -2467
rect 9692 -2411 9756 -2407
rect 9692 -2467 9696 -2411
rect 9696 -2467 9752 -2411
rect 9752 -2467 9756 -2411
rect 9692 -2471 9756 -2467
rect 9772 -2411 9836 -2407
rect 9772 -2467 9776 -2411
rect 9776 -2467 9832 -2411
rect 9832 -2467 9836 -2411
rect 9772 -2471 9836 -2467
rect 9852 -2411 9916 -2407
rect 9852 -2467 9856 -2411
rect 9856 -2467 9912 -2411
rect 9912 -2467 9916 -2411
rect 9852 -2471 9916 -2467
rect 9932 -2411 9996 -2407
rect 9932 -2467 9936 -2411
rect 9936 -2467 9992 -2411
rect 9992 -2467 9996 -2411
rect 9932 -2471 9996 -2467
rect 10012 -2411 10076 -2407
rect 10012 -2467 10016 -2411
rect 10016 -2467 10072 -2411
rect 10072 -2467 10076 -2411
rect 10012 -2471 10076 -2467
rect 10092 -2411 10156 -2407
rect 10092 -2467 10096 -2411
rect 10096 -2467 10152 -2411
rect 10152 -2467 10156 -2411
rect 10092 -2471 10156 -2467
rect 10172 -2411 10236 -2407
rect 10172 -2467 10176 -2411
rect 10176 -2467 10232 -2411
rect 10232 -2467 10236 -2411
rect 10172 -2471 10236 -2467
rect 10252 -2411 10316 -2407
rect 10252 -2467 10256 -2411
rect 10256 -2467 10312 -2411
rect 10312 -2467 10316 -2411
rect 10252 -2471 10316 -2467
rect 10332 -2411 10396 -2407
rect 10332 -2467 10336 -2411
rect 10336 -2467 10392 -2411
rect 10392 -2467 10396 -2411
rect 10332 -2471 10396 -2467
rect 10412 -2411 10476 -2407
rect 10412 -2467 10416 -2411
rect 10416 -2467 10472 -2411
rect 10472 -2467 10476 -2411
rect 10412 -2471 10476 -2467
rect 10492 -2411 10556 -2407
rect 10492 -2467 10496 -2411
rect 10496 -2467 10552 -2411
rect 10552 -2467 10556 -2411
rect 10492 -2471 10556 -2467
rect 10572 -2411 10636 -2407
rect 10572 -2467 10576 -2411
rect 10576 -2467 10632 -2411
rect 10632 -2467 10636 -2411
rect 10572 -2471 10636 -2467
rect -188 -2878 -184 -2654
rect -184 -2878 352 -2654
rect 352 -2878 356 -2654
rect 10344 -2878 10348 -2654
rect 10348 -2878 10884 -2654
rect 10884 -2878 10888 -2654
<< metal4 >>
rect -400 2258 11100 2480
rect -400 2034 -188 2258
rect 356 2034 10344 2258
rect 10888 2034 11100 2258
rect -400 1906 11100 2034
rect -400 1762 3524 1906
rect 7268 1762 11100 1906
rect -400 1680 11100 1762
rect -400 -2407 11100 -2300
rect -400 -2471 12 -2407
rect 76 -2471 92 -2407
rect 156 -2471 172 -2407
rect 236 -2471 252 -2407
rect 316 -2471 332 -2407
rect 396 -2471 412 -2407
rect 476 -2471 492 -2407
rect 556 -2471 572 -2407
rect 636 -2471 652 -2407
rect 716 -2471 732 -2407
rect 796 -2471 812 -2407
rect 876 -2471 892 -2407
rect 956 -2471 972 -2407
rect 1036 -2471 1052 -2407
rect 1116 -2471 1132 -2407
rect 1196 -2471 1212 -2407
rect 1276 -2471 1292 -2407
rect 1356 -2471 1372 -2407
rect 1436 -2471 1452 -2407
rect 1516 -2471 1532 -2407
rect 1596 -2471 1612 -2407
rect 1676 -2471 1692 -2407
rect 1756 -2471 1772 -2407
rect 1836 -2471 1852 -2407
rect 1916 -2471 1932 -2407
rect 1996 -2471 2012 -2407
rect 2076 -2471 2092 -2407
rect 2156 -2471 2172 -2407
rect 2236 -2471 2252 -2407
rect 2316 -2471 2332 -2407
rect 2396 -2471 2412 -2407
rect 2476 -2471 2492 -2407
rect 2556 -2471 2572 -2407
rect 2636 -2471 2652 -2407
rect 2716 -2471 2732 -2407
rect 2796 -2471 2812 -2407
rect 2876 -2471 2892 -2407
rect 2956 -2471 2972 -2407
rect 3036 -2471 3052 -2407
rect 3116 -2471 3132 -2407
rect 3196 -2471 3212 -2407
rect 3276 -2471 3292 -2407
rect 3356 -2471 3372 -2407
rect 3436 -2471 3452 -2407
rect 3516 -2471 3532 -2407
rect 3596 -2471 3612 -2407
rect 3676 -2471 3692 -2407
rect 3756 -2471 3772 -2407
rect 3836 -2471 3852 -2407
rect 3916 -2471 3932 -2407
rect 3996 -2471 4012 -2407
rect 4076 -2471 4092 -2407
rect 4156 -2471 4172 -2407
rect 4236 -2471 4252 -2407
rect 4316 -2471 4332 -2407
rect 4396 -2471 4412 -2407
rect 4476 -2471 4492 -2407
rect 4556 -2471 4572 -2407
rect 4636 -2471 4652 -2407
rect 4716 -2471 4732 -2407
rect 4796 -2471 4812 -2407
rect 4876 -2471 4892 -2407
rect 4956 -2471 4972 -2407
rect 5036 -2471 5052 -2407
rect 5116 -2471 5132 -2407
rect 5196 -2471 5212 -2407
rect 5276 -2471 5292 -2407
rect 5356 -2471 5372 -2407
rect 5436 -2471 5452 -2407
rect 5516 -2471 5532 -2407
rect 5596 -2471 5612 -2407
rect 5676 -2471 5692 -2407
rect 5756 -2471 5772 -2407
rect 5836 -2471 5852 -2407
rect 5916 -2471 5932 -2407
rect 5996 -2471 6012 -2407
rect 6076 -2471 6092 -2407
rect 6156 -2471 6172 -2407
rect 6236 -2471 6252 -2407
rect 6316 -2471 6332 -2407
rect 6396 -2471 6412 -2407
rect 6476 -2471 6492 -2407
rect 6556 -2471 6572 -2407
rect 6636 -2471 6652 -2407
rect 6716 -2471 6732 -2407
rect 6796 -2471 6812 -2407
rect 6876 -2471 6892 -2407
rect 6956 -2471 6972 -2407
rect 7036 -2471 7052 -2407
rect 7116 -2471 7132 -2407
rect 7196 -2471 7212 -2407
rect 7276 -2471 7292 -2407
rect 7356 -2471 7372 -2407
rect 7436 -2471 7452 -2407
rect 7516 -2471 7532 -2407
rect 7596 -2471 7612 -2407
rect 7676 -2471 7692 -2407
rect 7756 -2471 7772 -2407
rect 7836 -2471 7852 -2407
rect 7916 -2471 7932 -2407
rect 7996 -2471 8012 -2407
rect 8076 -2471 8092 -2407
rect 8156 -2471 8172 -2407
rect 8236 -2471 8252 -2407
rect 8316 -2471 8332 -2407
rect 8396 -2471 8412 -2407
rect 8476 -2471 8492 -2407
rect 8556 -2471 8572 -2407
rect 8636 -2471 8652 -2407
rect 8716 -2471 8732 -2407
rect 8796 -2471 8812 -2407
rect 8876 -2471 8892 -2407
rect 8956 -2471 8972 -2407
rect 9036 -2471 9052 -2407
rect 9116 -2471 9132 -2407
rect 9196 -2471 9212 -2407
rect 9276 -2471 9292 -2407
rect 9356 -2471 9372 -2407
rect 9436 -2471 9452 -2407
rect 9516 -2471 9532 -2407
rect 9596 -2471 9612 -2407
rect 9676 -2471 9692 -2407
rect 9756 -2471 9772 -2407
rect 9836 -2471 9852 -2407
rect 9916 -2471 9932 -2407
rect 9996 -2471 10012 -2407
rect 10076 -2471 10092 -2407
rect 10156 -2471 10172 -2407
rect 10236 -2471 10252 -2407
rect 10316 -2471 10332 -2407
rect 10396 -2471 10412 -2407
rect 10476 -2471 10492 -2407
rect 10556 -2471 10572 -2407
rect 10636 -2471 11100 -2407
rect -400 -2654 11100 -2471
rect -400 -2878 -188 -2654
rect 356 -2878 10344 -2654
rect 10888 -2878 11100 -2654
rect -400 -3100 11100 -2878
use sky130_fd_pr__nfet_01v8_lvt_YXNJ6N  sky130_fd_pr__nfet_01v8_lvt_YXNJ6N_0
timestamp 1626486988
transform 1 0 5339 0 1 -378
box -1345 -288 1345 288
use sky130_fd_pr__pfet_01v8_HVERXA  sky130_fd_pr__pfet_01v8_HVERXA_0
timestamp 1626486988
transform 1 0 5343 0 1 1190
box -1871 -200 1871 200
use sky130_fd_pr__nfet_01v8_3YN2WN  sky130_fd_pr__nfet_01v8_3YN2WN_1
timestamp 1626486988
transform 1 0 5353 0 1 -1386
box -5203 -188 5203 188
use sky130_fd_pr__nfet_01v8_3YN2WN  sky130_fd_pr__nfet_01v8_3YN2WN_0
timestamp 1626486988
transform 1 0 5353 0 1 -1926
box -5203 -188 5203 188
use sky130_fd_pr__nfet_01v8_YXNJ6N  sky130_fd_pr__nfet_01v8_YXNJ6N_1
timestamp 1626486988
transform 1 0 8635 0 1 -378
box -1345 -288 1345 288
use sky130_fd_pr__nfet_01v8_YXNJ6N  sky130_fd_pr__nfet_01v8_YXNJ6N_0
timestamp 1626486988
transform 1 0 2043 0 1 -378
box -1345 -288 1345 288
<< labels >>
flabel metal1 s 1044 -1164 1062 -1152 1 FreeSans 600 0 0 0 vtail_diff
flabel metal1 s 9634 -1132 9650 -1116 1 FreeSans 600 0 0 0 vbiasp
flabel metal1 s 9628 -2132 9644 -2122 1 FreeSans 600 0 0 0 vcmn_tail2
flabel metal1 s 6202 -2146 6214 -2134 1 FreeSans 600 0 0 0 vcmn_tail1
flabel metal1 s 1262 -1662 1270 -1654 1 FreeSans 600 0 0 0 vcmc
flabel metal2 s 6878 -1662 6892 -1652 1 FreeSans 600 0 0 0 ibiasn
flabel metal2 s 8640 -872 8650 -858 1 FreeSans 600 0 0 0 vcmn_tail2
flabel metal2 s 8428 -30 8440 -14 1 FreeSans 600 0 0 0 vom
flabel metal2 s 8082 -768 8104 -750 1 FreeSans 600 0 0 0 vocm
flabel metal2 s 7816 84 7828 94 1 FreeSans 600 0 0 0 vcmcn2
flabel metal2 s 8638 196 8648 208 1 FreeSans 600 0 0 0 vcmcn
flabel metal2 s 4368 918 4374 930 1 FreeSans 600 0 0 0 vbiasp
flabel metal2 s 5334 -876 5352 -860 1 FreeSans 600 0 0 0 vtail_diff
flabel metal2 s 5154 -28 5172 -12 1 FreeSans 600 0 0 0 vim
flabel metal2 s 4486 84 4506 96 1 FreeSans 600 0 0 0 vom
flabel metal2 s 5310 198 5330 214 1 FreeSans 600 0 0 0 vop
flabel metal2 s 2032 190 2050 210 1 FreeSans 600 0 0 0 vcmcn1
flabel metal2 s 1136 72 1156 86 1 FreeSans 600 0 0 0 vcmcn
flabel metal2 s 1856 -42 1878 -30 1 FreeSans 600 0 0 0 vocm
flabel metal2 s 1492 -760 1510 -748 1 FreeSans 600 0 0 0 vop
flabel metal2 s 2030 -874 2050 -858 1 FreeSans 600 0 0 0 vcmn_tail1
flabel metal2 s 4684 -754 4692 -748 1 FreeSans 600 0 0 0 vip
flabel metal1 s 5328 1322 5346 1338 1 FreeSans 600 0 0 0 vcmc
flabel metal2 s 4306 554 4312 558 1 FreeSans 600 0 0 0 vom
flabel metal2 s 4818 552 4824 558 1 FreeSans 600 0 0 0 vop
flabel metal4 s -66 2456 -54 2470 1 FreeSans 600 0 0 0 VDD
flabel metal4 s 172 -3088 186 -3074 1 FreeSans 600 0 0 0 VSS
<< properties >>
string FIXED_BBOX -272 -2972 10972 332
<< end >>
