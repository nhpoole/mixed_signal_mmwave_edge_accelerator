magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< pwell >>
rect -26 -26 176 1426
<< scnmos >>
rect 60 0 90 1400
<< ndiff >>
rect 0 0 60 1400
rect 90 0 150 1400
<< poly >>
rect 60 1400 90 1426
rect 60 -26 90 0
<< locali >>
rect 8 667 42 733
rect 108 667 142 733
use contact_11  contact_11_0
timestamp 1624494425
transform 1 0 100 0 1 667
box -26 -22 76 88
use contact_11  contact_11_1
timestamp 1624494425
transform 1 0 0 0 1 667
box -26 -22 76 88
<< labels >>
rlabel poly s 75 700 75 700 4 G
rlabel locali s 25 700 25 700 4 S
rlabel locali s 125 700 125 700 4 D
<< properties >>
string FIXED_BBOX -25 -26 175 1426
<< end >>
