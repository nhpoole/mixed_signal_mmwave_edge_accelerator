magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< nwell >>
rect -54 -54 1716 454
<< scpmos >>
rect 60 0 90 400
rect 168 0 198 400
rect 276 0 306 400
rect 384 0 414 400
rect 492 0 522 400
rect 600 0 630 400
rect 708 0 738 400
rect 816 0 846 400
rect 924 0 954 400
rect 1032 0 1062 400
rect 1140 0 1170 400
rect 1248 0 1278 400
rect 1356 0 1386 400
rect 1464 0 1494 400
rect 1572 0 1602 400
<< pdiff >>
rect 0 0 60 400
rect 90 0 168 400
rect 198 0 276 400
rect 306 0 384 400
rect 414 0 492 400
rect 522 0 600 400
rect 630 0 708 400
rect 738 0 816 400
rect 846 0 924 400
rect 954 0 1032 400
rect 1062 0 1140 400
rect 1170 0 1248 400
rect 1278 0 1356 400
rect 1386 0 1464 400
rect 1494 0 1572 400
rect 1602 0 1662 400
<< poly >>
rect 60 400 90 426
rect 168 400 198 426
rect 276 400 306 426
rect 384 400 414 426
rect 492 400 522 426
rect 600 400 630 426
rect 708 400 738 426
rect 816 400 846 426
rect 924 400 954 426
rect 1032 400 1062 426
rect 1140 400 1170 426
rect 1248 400 1278 426
rect 1356 400 1386 426
rect 1464 400 1494 426
rect 1572 400 1602 426
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
rect 816 -26 846 0
rect 924 -26 954 0
rect 1032 -26 1062 0
rect 1140 -26 1170 0
rect 1248 -26 1278 0
rect 1356 -26 1386 0
rect 1464 -26 1494 0
rect 1572 -26 1602 0
rect 60 -56 1602 -26
<< locali >>
rect 8 167 42 233
rect 112 133 146 200
rect 220 167 254 233
rect 328 133 362 200
rect 436 167 470 233
rect 544 133 578 200
rect 652 167 686 233
rect 760 133 794 200
rect 868 167 902 233
rect 976 133 1010 200
rect 1084 167 1118 233
rect 1192 133 1226 200
rect 1300 167 1334 233
rect 1408 133 1442 200
rect 1516 167 1550 233
rect 1620 133 1654 200
rect 112 99 1654 133
use contact_12  contact_12_14
timestamp 1624494425
transform 1 0 104 0 1 167
box -59 -51 109 117
use contact_12  contact_12_15
timestamp 1624494425
transform 1 0 0 0 1 167
box -59 -51 109 117
use contact_12  contact_12_12
timestamp 1624494425
transform 1 0 320 0 1 167
box -59 -51 109 117
use contact_12  contact_12_13
timestamp 1624494425
transform 1 0 212 0 1 167
box -59 -51 109 117
use contact_12  contact_12_11
timestamp 1624494425
transform 1 0 428 0 1 167
box -59 -51 109 117
use contact_12  contact_12_9
timestamp 1624494425
transform 1 0 644 0 1 167
box -59 -51 109 117
use contact_12  contact_12_10
timestamp 1624494425
transform 1 0 536 0 1 167
box -59 -51 109 117
use contact_12  contact_12_8
timestamp 1624494425
transform 1 0 752 0 1 167
box -59 -51 109 117
use contact_12  contact_12_6
timestamp 1624494425
transform 1 0 968 0 1 167
box -59 -51 109 117
use contact_12  contact_12_7
timestamp 1624494425
transform 1 0 860 0 1 167
box -59 -51 109 117
use contact_12  contact_12_5
timestamp 1624494425
transform 1 0 1076 0 1 167
box -59 -51 109 117
use contact_12  contact_12_3
timestamp 1624494425
transform 1 0 1292 0 1 167
box -59 -51 109 117
use contact_12  contact_12_4
timestamp 1624494425
transform 1 0 1184 0 1 167
box -59 -51 109 117
use contact_12  contact_12_1
timestamp 1624494425
transform 1 0 1508 0 1 167
box -59 -51 109 117
use contact_12  contact_12_2
timestamp 1624494425
transform 1 0 1400 0 1 167
box -59 -51 109 117
use contact_12  contact_12_0
timestamp 1624494425
transform 1 0 1612 0 1 167
box -59 -51 109 117
<< labels >>
rlabel poly s 831 -41 831 -41 4 G
rlabel locali s 669 200 669 200 4 S
rlabel locali s 1533 200 1533 200 4 S
rlabel locali s 237 200 237 200 4 S
rlabel locali s 885 200 885 200 4 S
rlabel locali s 25 200 25 200 4 S
rlabel locali s 453 200 453 200 4 S
rlabel locali s 1101 200 1101 200 4 S
rlabel locali s 1317 200 1317 200 4 S
rlabel locali s 883 116 883 116 4 D
<< properties >>
string FIXED_BBOX -54 -56 1716 454
<< end >>
