magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -3048 -2960 3047 2960
<< metal3 >>
rect -1788 1550 -1089 1700
rect -1788 1486 -1173 1550
rect -1109 1486 -1089 1550
rect -1788 1470 -1089 1486
rect -1788 1406 -1173 1470
rect -1109 1406 -1089 1470
rect -1788 1390 -1089 1406
rect -1788 1326 -1173 1390
rect -1109 1326 -1089 1390
rect -1788 1310 -1089 1326
rect -1788 1246 -1173 1310
rect -1109 1246 -1089 1310
rect -1788 1100 -1089 1246
rect -1069 1549 -370 1700
rect -1069 1485 -454 1549
rect -390 1485 -370 1549
rect -1069 1469 -370 1485
rect -1069 1405 -454 1469
rect -390 1405 -370 1469
rect -1069 1389 -370 1405
rect -1069 1325 -454 1389
rect -390 1325 -370 1389
rect -1069 1309 -370 1325
rect -1069 1245 -454 1309
rect -390 1245 -370 1309
rect -1069 1100 -370 1245
rect -350 1549 349 1700
rect -350 1485 265 1549
rect 329 1485 349 1549
rect -350 1469 349 1485
rect -350 1405 265 1469
rect 329 1405 349 1469
rect -350 1389 349 1405
rect -350 1325 265 1389
rect 329 1325 349 1389
rect -350 1309 349 1325
rect -350 1245 265 1309
rect 329 1245 349 1309
rect -350 1100 349 1245
rect 369 1549 1068 1700
rect 369 1485 984 1549
rect 1048 1485 1068 1549
rect 369 1469 1068 1485
rect 369 1405 984 1469
rect 1048 1405 1068 1469
rect 369 1389 1068 1405
rect 369 1325 984 1389
rect 1048 1325 1068 1389
rect 369 1309 1068 1325
rect 369 1245 984 1309
rect 1048 1245 1068 1309
rect 369 1100 1068 1245
rect 1088 1549 1787 1700
rect 1088 1485 1703 1549
rect 1767 1485 1787 1549
rect 1088 1469 1787 1485
rect 1088 1405 1703 1469
rect 1767 1405 1787 1469
rect 1088 1389 1787 1405
rect 1088 1325 1703 1389
rect 1767 1325 1787 1389
rect 1088 1309 1787 1325
rect 1088 1245 1703 1309
rect 1767 1245 1787 1309
rect 1088 1100 1787 1245
rect -1788 850 -1089 1000
rect -1788 786 -1173 850
rect -1109 786 -1089 850
rect -1788 770 -1089 786
rect -1788 706 -1173 770
rect -1109 706 -1089 770
rect -1788 690 -1089 706
rect -1788 626 -1173 690
rect -1109 626 -1089 690
rect -1788 610 -1089 626
rect -1788 546 -1173 610
rect -1109 546 -1089 610
rect -1788 400 -1089 546
rect -1069 850 -370 1000
rect -1069 786 -454 850
rect -390 786 -370 850
rect -1069 770 -370 786
rect -1069 706 -454 770
rect -390 706 -370 770
rect -1069 690 -370 706
rect -1069 626 -454 690
rect -390 626 -370 690
rect -1069 610 -370 626
rect -1069 546 -454 610
rect -390 546 -370 610
rect -1069 400 -370 546
rect -350 850 349 1000
rect -350 786 265 850
rect 329 786 349 850
rect -350 770 349 786
rect -350 706 265 770
rect 329 706 349 770
rect -350 690 349 706
rect -350 626 265 690
rect 329 626 349 690
rect -350 610 349 626
rect -350 546 265 610
rect 329 546 349 610
rect -350 400 349 546
rect 369 850 1068 1000
rect 369 786 984 850
rect 1048 786 1068 850
rect 369 770 1068 786
rect 369 706 984 770
rect 1048 706 1068 770
rect 369 690 1068 706
rect 369 626 984 690
rect 1048 626 1068 690
rect 369 610 1068 626
rect 369 546 984 610
rect 1048 546 1068 610
rect 369 400 1068 546
rect 1088 850 1787 1000
rect 1088 786 1703 850
rect 1767 786 1787 850
rect 1088 770 1787 786
rect 1088 706 1703 770
rect 1767 706 1787 770
rect 1088 690 1787 706
rect 1088 626 1703 690
rect 1767 626 1787 690
rect 1088 610 1787 626
rect 1088 546 1703 610
rect 1767 546 1787 610
rect 1088 400 1787 546
rect -1788 150 -1089 300
rect -1788 86 -1173 150
rect -1109 86 -1089 150
rect -1788 70 -1089 86
rect -1788 6 -1173 70
rect -1109 6 -1089 70
rect -1788 -10 -1089 6
rect -1788 -74 -1173 -10
rect -1109 -74 -1089 -10
rect -1788 -90 -1089 -74
rect -1788 -154 -1173 -90
rect -1109 -154 -1089 -90
rect -1788 -300 -1089 -154
rect -1069 150 -370 300
rect -1069 86 -454 150
rect -390 86 -370 150
rect -1069 70 -370 86
rect -1069 6 -454 70
rect -390 6 -370 70
rect -1069 -10 -370 6
rect -1069 -74 -454 -10
rect -390 -74 -370 -10
rect -1069 -90 -370 -74
rect -1069 -154 -454 -90
rect -390 -154 -370 -90
rect -1069 -300 -370 -154
rect -350 150 349 300
rect -350 86 265 150
rect 329 86 349 150
rect -350 70 349 86
rect -350 6 265 70
rect 329 6 349 70
rect -350 -10 349 6
rect -350 -74 265 -10
rect 329 -74 349 -10
rect -350 -90 349 -74
rect -350 -154 265 -90
rect 329 -154 349 -90
rect -350 -300 349 -154
rect 369 150 1068 300
rect 369 86 984 150
rect 1048 86 1068 150
rect 369 70 1068 86
rect 369 6 984 70
rect 1048 6 1068 70
rect 369 -10 1068 6
rect 369 -74 984 -10
rect 1048 -74 1068 -10
rect 369 -90 1068 -74
rect 369 -154 984 -90
rect 1048 -154 1068 -90
rect 369 -300 1068 -154
rect 1088 150 1787 300
rect 1088 86 1703 150
rect 1767 86 1787 150
rect 1088 70 1787 86
rect 1088 6 1703 70
rect 1767 6 1787 70
rect 1088 -10 1787 6
rect 1088 -74 1703 -10
rect 1767 -74 1787 -10
rect 1088 -90 1787 -74
rect 1088 -154 1703 -90
rect 1767 -154 1787 -90
rect 1088 -300 1787 -154
rect -1788 -550 -1089 -400
rect -1788 -614 -1173 -550
rect -1109 -614 -1089 -550
rect -1788 -630 -1089 -614
rect -1788 -694 -1173 -630
rect -1109 -694 -1089 -630
rect -1788 -710 -1089 -694
rect -1788 -774 -1173 -710
rect -1109 -774 -1089 -710
rect -1788 -790 -1089 -774
rect -1788 -854 -1173 -790
rect -1109 -854 -1089 -790
rect -1788 -1000 -1089 -854
rect -1069 -550 -370 -400
rect -1069 -614 -454 -550
rect -390 -614 -370 -550
rect -1069 -630 -370 -614
rect -1069 -694 -454 -630
rect -390 -694 -370 -630
rect -1069 -710 -370 -694
rect -1069 -774 -454 -710
rect -390 -774 -370 -710
rect -1069 -790 -370 -774
rect -1069 -854 -454 -790
rect -390 -854 -370 -790
rect -1069 -1000 -370 -854
rect -350 -550 349 -400
rect -350 -614 265 -550
rect 329 -614 349 -550
rect -350 -630 349 -614
rect -350 -694 265 -630
rect 329 -694 349 -630
rect -350 -710 349 -694
rect -350 -774 265 -710
rect 329 -774 349 -710
rect -350 -790 349 -774
rect -350 -854 265 -790
rect 329 -854 349 -790
rect -350 -1000 349 -854
rect 369 -550 1068 -400
rect 369 -614 984 -550
rect 1048 -614 1068 -550
rect 369 -630 1068 -614
rect 369 -694 984 -630
rect 1048 -694 1068 -630
rect 369 -710 1068 -694
rect 369 -774 984 -710
rect 1048 -774 1068 -710
rect 369 -790 1068 -774
rect 369 -854 984 -790
rect 1048 -854 1068 -790
rect 369 -1000 1068 -854
rect 1088 -550 1787 -400
rect 1088 -614 1703 -550
rect 1767 -614 1787 -550
rect 1088 -630 1787 -614
rect 1088 -694 1703 -630
rect 1767 -694 1787 -630
rect 1088 -710 1787 -694
rect 1088 -774 1703 -710
rect 1767 -774 1787 -710
rect 1088 -790 1787 -774
rect 1088 -854 1703 -790
rect 1767 -854 1787 -790
rect 1088 -1000 1787 -854
rect -1788 -1250 -1089 -1100
rect -1788 -1314 -1173 -1250
rect -1109 -1314 -1089 -1250
rect -1788 -1330 -1089 -1314
rect -1788 -1394 -1173 -1330
rect -1109 -1394 -1089 -1330
rect -1788 -1410 -1089 -1394
rect -1788 -1474 -1173 -1410
rect -1109 -1474 -1089 -1410
rect -1788 -1490 -1089 -1474
rect -1788 -1554 -1173 -1490
rect -1109 -1554 -1089 -1490
rect -1788 -1700 -1089 -1554
rect -1069 -1250 -370 -1100
rect -1069 -1314 -454 -1250
rect -390 -1314 -370 -1250
rect -1069 -1330 -370 -1314
rect -1069 -1394 -454 -1330
rect -390 -1394 -370 -1330
rect -1069 -1410 -370 -1394
rect -1069 -1474 -454 -1410
rect -390 -1474 -370 -1410
rect -1069 -1490 -370 -1474
rect -1069 -1554 -454 -1490
rect -390 -1554 -370 -1490
rect -1069 -1700 -370 -1554
rect -350 -1250 349 -1100
rect -350 -1314 265 -1250
rect 329 -1314 349 -1250
rect -350 -1330 349 -1314
rect -350 -1394 265 -1330
rect 329 -1394 349 -1330
rect -350 -1410 349 -1394
rect -350 -1474 265 -1410
rect 329 -1474 349 -1410
rect -350 -1490 349 -1474
rect -350 -1554 265 -1490
rect 329 -1554 349 -1490
rect -350 -1700 349 -1554
rect 369 -1250 1068 -1100
rect 369 -1314 984 -1250
rect 1048 -1314 1068 -1250
rect 369 -1330 1068 -1314
rect 369 -1394 984 -1330
rect 1048 -1394 1068 -1330
rect 369 -1410 1068 -1394
rect 369 -1474 984 -1410
rect 1048 -1474 1068 -1410
rect 369 -1490 1068 -1474
rect 369 -1554 984 -1490
rect 1048 -1554 1068 -1490
rect 369 -1700 1068 -1554
rect 1088 -1250 1787 -1100
rect 1088 -1314 1703 -1250
rect 1767 -1314 1787 -1250
rect 1088 -1330 1787 -1314
rect 1088 -1394 1703 -1330
rect 1767 -1394 1787 -1330
rect 1088 -1410 1787 -1394
rect 1088 -1474 1703 -1410
rect 1767 -1474 1787 -1410
rect 1088 -1490 1787 -1474
rect 1088 -1554 1703 -1490
rect 1767 -1554 1787 -1490
rect 1088 -1700 1787 -1554
<< via3 >>
rect -1173 1486 -1109 1550
rect -1173 1406 -1109 1470
rect -1173 1326 -1109 1390
rect -1173 1246 -1109 1310
rect -454 1485 -390 1549
rect -454 1405 -390 1469
rect -454 1325 -390 1389
rect -454 1245 -390 1309
rect 265 1485 329 1549
rect 265 1405 329 1469
rect 265 1325 329 1389
rect 265 1245 329 1309
rect 984 1485 1048 1549
rect 984 1405 1048 1469
rect 984 1325 1048 1389
rect 984 1245 1048 1309
rect 1703 1485 1767 1549
rect 1703 1405 1767 1469
rect 1703 1325 1767 1389
rect 1703 1245 1767 1309
rect -1173 786 -1109 850
rect -1173 706 -1109 770
rect -1173 626 -1109 690
rect -1173 546 -1109 610
rect -454 786 -390 850
rect -454 706 -390 770
rect -454 626 -390 690
rect -454 546 -390 610
rect 265 786 329 850
rect 265 706 329 770
rect 265 626 329 690
rect 265 546 329 610
rect 984 786 1048 850
rect 984 706 1048 770
rect 984 626 1048 690
rect 984 546 1048 610
rect 1703 786 1767 850
rect 1703 706 1767 770
rect 1703 626 1767 690
rect 1703 546 1767 610
rect -1173 86 -1109 150
rect -1173 6 -1109 70
rect -1173 -74 -1109 -10
rect -1173 -154 -1109 -90
rect -454 86 -390 150
rect -454 6 -390 70
rect -454 -74 -390 -10
rect -454 -154 -390 -90
rect 265 86 329 150
rect 265 6 329 70
rect 265 -74 329 -10
rect 265 -154 329 -90
rect 984 86 1048 150
rect 984 6 1048 70
rect 984 -74 1048 -10
rect 984 -154 1048 -90
rect 1703 86 1767 150
rect 1703 6 1767 70
rect 1703 -74 1767 -10
rect 1703 -154 1767 -90
rect -1173 -614 -1109 -550
rect -1173 -694 -1109 -630
rect -1173 -774 -1109 -710
rect -1173 -854 -1109 -790
rect -454 -614 -390 -550
rect -454 -694 -390 -630
rect -454 -774 -390 -710
rect -454 -854 -390 -790
rect 265 -614 329 -550
rect 265 -694 329 -630
rect 265 -774 329 -710
rect 265 -854 329 -790
rect 984 -614 1048 -550
rect 984 -694 1048 -630
rect 984 -774 1048 -710
rect 984 -854 1048 -790
rect 1703 -614 1767 -550
rect 1703 -694 1767 -630
rect 1703 -774 1767 -710
rect 1703 -854 1767 -790
rect -1173 -1314 -1109 -1250
rect -1173 -1394 -1109 -1330
rect -1173 -1474 -1109 -1410
rect -1173 -1554 -1109 -1490
rect -454 -1314 -390 -1250
rect -454 -1394 -390 -1330
rect -454 -1474 -390 -1410
rect -454 -1554 -390 -1490
rect 265 -1314 329 -1250
rect 265 -1394 329 -1330
rect 265 -1474 329 -1410
rect 265 -1554 329 -1490
rect 984 -1314 1048 -1250
rect 984 -1394 1048 -1330
rect 984 -1474 1048 -1410
rect 984 -1554 1048 -1490
rect 1703 -1314 1767 -1250
rect 1703 -1394 1767 -1330
rect 1703 -1474 1767 -1410
rect 1703 -1554 1767 -1490
<< mimcap >>
rect -1688 1552 -1288 1600
rect -1688 1248 -1640 1552
rect -1336 1248 -1288 1552
rect -1688 1200 -1288 1248
rect -969 1552 -569 1600
rect -969 1248 -921 1552
rect -617 1248 -569 1552
rect -969 1200 -569 1248
rect -250 1552 150 1600
rect -250 1248 -202 1552
rect 102 1248 150 1552
rect -250 1200 150 1248
rect 469 1552 869 1600
rect 469 1248 517 1552
rect 821 1248 869 1552
rect 469 1200 869 1248
rect 1188 1552 1588 1600
rect 1188 1248 1236 1552
rect 1540 1248 1588 1552
rect 1188 1200 1588 1248
rect -1688 852 -1288 900
rect -1688 548 -1640 852
rect -1336 548 -1288 852
rect -1688 500 -1288 548
rect -969 852 -569 900
rect -969 548 -921 852
rect -617 548 -569 852
rect -969 500 -569 548
rect -250 852 150 900
rect -250 548 -202 852
rect 102 548 150 852
rect -250 500 150 548
rect 469 852 869 900
rect 469 548 517 852
rect 821 548 869 852
rect 469 500 869 548
rect 1188 852 1588 900
rect 1188 548 1236 852
rect 1540 548 1588 852
rect 1188 500 1588 548
rect -1688 152 -1288 200
rect -1688 -152 -1640 152
rect -1336 -152 -1288 152
rect -1688 -200 -1288 -152
rect -969 152 -569 200
rect -969 -152 -921 152
rect -617 -152 -569 152
rect -969 -200 -569 -152
rect -250 152 150 200
rect -250 -152 -202 152
rect 102 -152 150 152
rect -250 -200 150 -152
rect 469 152 869 200
rect 469 -152 517 152
rect 821 -152 869 152
rect 469 -200 869 -152
rect 1188 152 1588 200
rect 1188 -152 1236 152
rect 1540 -152 1588 152
rect 1188 -200 1588 -152
rect -1688 -548 -1288 -500
rect -1688 -852 -1640 -548
rect -1336 -852 -1288 -548
rect -1688 -900 -1288 -852
rect -969 -548 -569 -500
rect -969 -852 -921 -548
rect -617 -852 -569 -548
rect -969 -900 -569 -852
rect -250 -548 150 -500
rect -250 -852 -202 -548
rect 102 -852 150 -548
rect -250 -900 150 -852
rect 469 -548 869 -500
rect 469 -852 517 -548
rect 821 -852 869 -548
rect 469 -900 869 -852
rect 1188 -548 1588 -500
rect 1188 -852 1236 -548
rect 1540 -852 1588 -548
rect 1188 -900 1588 -852
rect -1688 -1248 -1288 -1200
rect -1688 -1552 -1640 -1248
rect -1336 -1552 -1288 -1248
rect -1688 -1600 -1288 -1552
rect -969 -1248 -569 -1200
rect -969 -1552 -921 -1248
rect -617 -1552 -569 -1248
rect -969 -1600 -569 -1552
rect -250 -1248 150 -1200
rect -250 -1552 -202 -1248
rect 102 -1552 150 -1248
rect -250 -1600 150 -1552
rect 469 -1248 869 -1200
rect 469 -1552 517 -1248
rect 821 -1552 869 -1248
rect 469 -1600 869 -1552
rect 1188 -1248 1588 -1200
rect 1188 -1552 1236 -1248
rect 1540 -1552 1588 -1248
rect 1188 -1600 1588 -1552
<< mimcapcontact >>
rect -1640 1248 -1336 1552
rect -921 1248 -617 1552
rect -202 1248 102 1552
rect 517 1248 821 1552
rect 1236 1248 1540 1552
rect -1640 548 -1336 852
rect -921 548 -617 852
rect -202 548 102 852
rect 517 548 821 852
rect 1236 548 1540 852
rect -1640 -152 -1336 152
rect -921 -152 -617 152
rect -202 -152 102 152
rect 517 -152 821 152
rect 1236 -152 1540 152
rect -1640 -852 -1336 -548
rect -921 -852 -617 -548
rect -202 -852 102 -548
rect 517 -852 821 -548
rect 1236 -852 1540 -548
rect -1640 -1552 -1336 -1248
rect -921 -1552 -617 -1248
rect -202 -1552 102 -1248
rect 517 -1552 821 -1248
rect 1236 -1552 1540 -1248
<< metal4 >>
rect -1649 1552 -1327 1561
rect -1649 1248 -1640 1552
rect -1336 1248 -1327 1552
rect -1649 1239 -1327 1248
rect -1189 1550 -1093 1600
rect -1189 1486 -1173 1550
rect -1109 1486 -1093 1550
rect -1189 1470 -1093 1486
rect -1189 1406 -1173 1470
rect -1109 1406 -1093 1470
rect -1189 1390 -1093 1406
rect -1189 1326 -1173 1390
rect -1109 1326 -1093 1390
rect -1189 1310 -1093 1326
rect -1189 1246 -1173 1310
rect -1109 1246 -1093 1310
rect -1189 1196 -1093 1246
rect -930 1552 -608 1561
rect -930 1248 -921 1552
rect -617 1248 -608 1552
rect -930 1239 -608 1248
rect -470 1549 -374 1598
rect -470 1485 -454 1549
rect -390 1485 -374 1549
rect -470 1469 -374 1485
rect -470 1405 -454 1469
rect -390 1405 -374 1469
rect -470 1389 -374 1405
rect -470 1325 -454 1389
rect -390 1325 -374 1389
rect -470 1309 -374 1325
rect -470 1245 -454 1309
rect -390 1245 -374 1309
rect -470 1196 -374 1245
rect -211 1552 111 1561
rect -211 1248 -202 1552
rect 102 1248 111 1552
rect -211 1239 111 1248
rect 249 1549 345 1598
rect 249 1485 265 1549
rect 329 1485 345 1549
rect 249 1469 345 1485
rect 249 1405 265 1469
rect 329 1405 345 1469
rect 249 1389 345 1405
rect 249 1325 265 1389
rect 329 1325 345 1389
rect 249 1309 345 1325
rect 249 1245 265 1309
rect 329 1245 345 1309
rect 249 1196 345 1245
rect 508 1552 830 1561
rect 508 1248 517 1552
rect 821 1248 830 1552
rect 508 1239 830 1248
rect 968 1549 1064 1598
rect 968 1485 984 1549
rect 1048 1485 1064 1549
rect 968 1469 1064 1485
rect 968 1405 984 1469
rect 1048 1405 1064 1469
rect 968 1389 1064 1405
rect 968 1325 984 1389
rect 1048 1325 1064 1389
rect 968 1309 1064 1325
rect 968 1245 984 1309
rect 1048 1245 1064 1309
rect 968 1196 1064 1245
rect 1227 1552 1549 1561
rect 1227 1248 1236 1552
rect 1540 1248 1549 1552
rect 1227 1239 1549 1248
rect 1687 1549 1783 1598
rect 1687 1485 1703 1549
rect 1767 1485 1783 1549
rect 1687 1469 1783 1485
rect 1687 1405 1703 1469
rect 1767 1405 1783 1469
rect 1687 1389 1783 1405
rect 1687 1325 1703 1389
rect 1767 1325 1783 1389
rect 1687 1309 1783 1325
rect 1687 1245 1703 1309
rect 1767 1245 1783 1309
rect 1687 1196 1783 1245
rect -1649 852 -1327 861
rect -1649 548 -1640 852
rect -1336 548 -1327 852
rect -1649 539 -1327 548
rect -1189 850 -1093 898
rect -1189 786 -1173 850
rect -1109 786 -1093 850
rect -1189 770 -1093 786
rect -1189 706 -1173 770
rect -1109 706 -1093 770
rect -1189 690 -1093 706
rect -1189 626 -1173 690
rect -1109 626 -1093 690
rect -1189 610 -1093 626
rect -1189 546 -1173 610
rect -1109 546 -1093 610
rect -1189 494 -1093 546
rect -930 852 -608 861
rect -930 548 -921 852
rect -617 548 -608 852
rect -930 539 -608 548
rect -470 850 -374 898
rect -470 786 -454 850
rect -390 786 -374 850
rect -470 770 -374 786
rect -470 706 -454 770
rect -390 706 -374 770
rect -470 690 -374 706
rect -470 626 -454 690
rect -390 626 -374 690
rect -470 610 -374 626
rect -470 546 -454 610
rect -390 546 -374 610
rect -470 494 -374 546
rect -211 852 111 861
rect -211 548 -202 852
rect 102 548 111 852
rect -211 539 111 548
rect 249 850 345 898
rect 249 786 265 850
rect 329 786 345 850
rect 249 770 345 786
rect 249 706 265 770
rect 329 706 345 770
rect 249 690 345 706
rect 249 626 265 690
rect 329 626 345 690
rect 249 610 345 626
rect 249 546 265 610
rect 329 546 345 610
rect 249 494 345 546
rect 508 852 830 861
rect 508 548 517 852
rect 821 548 830 852
rect 508 539 830 548
rect 968 850 1064 898
rect 968 786 984 850
rect 1048 786 1064 850
rect 968 770 1064 786
rect 968 706 984 770
rect 1048 706 1064 770
rect 968 690 1064 706
rect 968 626 984 690
rect 1048 626 1064 690
rect 968 610 1064 626
rect 968 546 984 610
rect 1048 546 1064 610
rect 968 494 1064 546
rect 1227 852 1549 861
rect 1227 548 1236 852
rect 1540 548 1549 852
rect 1227 539 1549 548
rect 1687 850 1783 898
rect 1687 786 1703 850
rect 1767 786 1783 850
rect 1687 770 1783 786
rect 1687 706 1703 770
rect 1767 706 1783 770
rect 1687 690 1783 706
rect 1687 626 1703 690
rect 1767 626 1783 690
rect 1687 610 1783 626
rect 1687 546 1703 610
rect 1767 546 1783 610
rect 1687 494 1783 546
rect -1649 152 -1327 161
rect -1649 -152 -1640 152
rect -1336 -152 -1327 152
rect -1649 -161 -1327 -152
rect -1189 150 -1093 198
rect -1189 86 -1173 150
rect -1109 86 -1093 150
rect -1189 70 -1093 86
rect -1189 6 -1173 70
rect -1109 6 -1093 70
rect -1189 -10 -1093 6
rect -1189 -74 -1173 -10
rect -1109 -74 -1093 -10
rect -1189 -90 -1093 -74
rect -1189 -154 -1173 -90
rect -1109 -154 -1093 -90
rect -1189 -204 -1093 -154
rect -930 152 -608 161
rect -930 -152 -921 152
rect -617 -152 -608 152
rect -930 -161 -608 -152
rect -470 150 -374 198
rect -470 86 -454 150
rect -390 86 -374 150
rect -470 70 -374 86
rect -470 6 -454 70
rect -390 6 -374 70
rect -470 -10 -374 6
rect -470 -74 -454 -10
rect -390 -74 -374 -10
rect -470 -90 -374 -74
rect -470 -154 -454 -90
rect -390 -154 -374 -90
rect -470 -204 -374 -154
rect -211 152 111 161
rect -211 -152 -202 152
rect 102 -152 111 152
rect -211 -161 111 -152
rect 249 150 345 198
rect 249 86 265 150
rect 329 86 345 150
rect 249 70 345 86
rect 249 6 265 70
rect 329 6 345 70
rect 249 -10 345 6
rect 249 -74 265 -10
rect 329 -74 345 -10
rect 249 -90 345 -74
rect 249 -154 265 -90
rect 329 -154 345 -90
rect 249 -204 345 -154
rect 508 152 830 161
rect 508 -152 517 152
rect 821 -152 830 152
rect 508 -161 830 -152
rect 968 150 1064 198
rect 968 86 984 150
rect 1048 86 1064 150
rect 968 70 1064 86
rect 968 6 984 70
rect 1048 6 1064 70
rect 968 -10 1064 6
rect 968 -74 984 -10
rect 1048 -74 1064 -10
rect 968 -90 1064 -74
rect 968 -154 984 -90
rect 1048 -154 1064 -90
rect 968 -204 1064 -154
rect 1227 152 1549 161
rect 1227 -152 1236 152
rect 1540 -152 1549 152
rect 1227 -161 1549 -152
rect 1687 150 1783 198
rect 1687 86 1703 150
rect 1767 86 1783 150
rect 1687 70 1783 86
rect 1687 6 1703 70
rect 1767 6 1783 70
rect 1687 -10 1783 6
rect 1687 -74 1703 -10
rect 1767 -74 1783 -10
rect 1687 -90 1783 -74
rect 1687 -154 1703 -90
rect 1767 -154 1783 -90
rect 1687 -204 1783 -154
rect -1649 -548 -1327 -539
rect -1649 -852 -1640 -548
rect -1336 -852 -1327 -548
rect -1649 -861 -1327 -852
rect -1189 -550 -1093 -502
rect -1189 -614 -1173 -550
rect -1109 -614 -1093 -550
rect -1189 -630 -1093 -614
rect -1189 -694 -1173 -630
rect -1109 -694 -1093 -630
rect -1189 -710 -1093 -694
rect -1189 -774 -1173 -710
rect -1109 -774 -1093 -710
rect -1189 -790 -1093 -774
rect -1189 -854 -1173 -790
rect -1109 -854 -1093 -790
rect -1189 -904 -1093 -854
rect -930 -548 -608 -539
rect -930 -852 -921 -548
rect -617 -852 -608 -548
rect -930 -861 -608 -852
rect -470 -550 -374 -502
rect -470 -614 -454 -550
rect -390 -614 -374 -550
rect -470 -630 -374 -614
rect -470 -694 -454 -630
rect -390 -694 -374 -630
rect -470 -710 -374 -694
rect -470 -774 -454 -710
rect -390 -774 -374 -710
rect -470 -790 -374 -774
rect -470 -854 -454 -790
rect -390 -854 -374 -790
rect -470 -904 -374 -854
rect -211 -548 111 -539
rect -211 -852 -202 -548
rect 102 -852 111 -548
rect -211 -861 111 -852
rect 249 -550 345 -502
rect 249 -614 265 -550
rect 329 -614 345 -550
rect 249 -630 345 -614
rect 249 -694 265 -630
rect 329 -694 345 -630
rect 249 -710 345 -694
rect 249 -774 265 -710
rect 329 -774 345 -710
rect 249 -790 345 -774
rect 249 -854 265 -790
rect 329 -854 345 -790
rect 249 -904 345 -854
rect 508 -548 830 -539
rect 508 -852 517 -548
rect 821 -852 830 -548
rect 508 -861 830 -852
rect 968 -550 1064 -502
rect 968 -614 984 -550
rect 1048 -614 1064 -550
rect 968 -630 1064 -614
rect 968 -694 984 -630
rect 1048 -694 1064 -630
rect 968 -710 1064 -694
rect 968 -774 984 -710
rect 1048 -774 1064 -710
rect 968 -790 1064 -774
rect 968 -854 984 -790
rect 1048 -854 1064 -790
rect 968 -904 1064 -854
rect 1227 -548 1549 -539
rect 1227 -852 1236 -548
rect 1540 -852 1549 -548
rect 1227 -861 1549 -852
rect 1687 -550 1783 -502
rect 1687 -614 1703 -550
rect 1767 -614 1783 -550
rect 1687 -630 1783 -614
rect 1687 -694 1703 -630
rect 1767 -694 1783 -630
rect 1687 -710 1783 -694
rect 1687 -774 1703 -710
rect 1767 -774 1783 -710
rect 1687 -790 1783 -774
rect 1687 -854 1703 -790
rect 1767 -854 1783 -790
rect 1687 -904 1783 -854
rect -1649 -1248 -1327 -1239
rect -1649 -1552 -1640 -1248
rect -1336 -1552 -1327 -1248
rect -1649 -1561 -1327 -1552
rect -1189 -1250 -1093 -1202
rect -1189 -1314 -1173 -1250
rect -1109 -1314 -1093 -1250
rect -1189 -1330 -1093 -1314
rect -1189 -1394 -1173 -1330
rect -1109 -1394 -1093 -1330
rect -1189 -1410 -1093 -1394
rect -1189 -1474 -1173 -1410
rect -1109 -1474 -1093 -1410
rect -1189 -1490 -1093 -1474
rect -1189 -1554 -1173 -1490
rect -1109 -1554 -1093 -1490
rect -1189 -1604 -1093 -1554
rect -930 -1248 -608 -1239
rect -930 -1552 -921 -1248
rect -617 -1552 -608 -1248
rect -930 -1561 -608 -1552
rect -470 -1250 -374 -1202
rect -470 -1314 -454 -1250
rect -390 -1314 -374 -1250
rect -470 -1330 -374 -1314
rect -470 -1394 -454 -1330
rect -390 -1394 -374 -1330
rect -470 -1410 -374 -1394
rect -470 -1474 -454 -1410
rect -390 -1474 -374 -1410
rect -470 -1490 -374 -1474
rect -470 -1554 -454 -1490
rect -390 -1554 -374 -1490
rect -470 -1604 -374 -1554
rect -211 -1248 111 -1239
rect -211 -1552 -202 -1248
rect 102 -1552 111 -1248
rect -211 -1561 111 -1552
rect 249 -1250 345 -1202
rect 249 -1314 265 -1250
rect 329 -1314 345 -1250
rect 249 -1330 345 -1314
rect 249 -1394 265 -1330
rect 329 -1394 345 -1330
rect 249 -1410 345 -1394
rect 249 -1474 265 -1410
rect 329 -1474 345 -1410
rect 249 -1490 345 -1474
rect 249 -1554 265 -1490
rect 329 -1554 345 -1490
rect 249 -1604 345 -1554
rect 508 -1248 830 -1239
rect 508 -1552 517 -1248
rect 821 -1552 830 -1248
rect 508 -1561 830 -1552
rect 968 -1250 1064 -1202
rect 968 -1314 984 -1250
rect 1048 -1314 1064 -1250
rect 968 -1330 1064 -1314
rect 968 -1394 984 -1330
rect 1048 -1394 1064 -1330
rect 968 -1410 1064 -1394
rect 968 -1474 984 -1410
rect 1048 -1474 1064 -1410
rect 968 -1490 1064 -1474
rect 968 -1554 984 -1490
rect 1048 -1554 1064 -1490
rect 968 -1604 1064 -1554
rect 1227 -1248 1549 -1239
rect 1227 -1552 1236 -1248
rect 1540 -1552 1549 -1248
rect 1227 -1561 1549 -1552
rect 1687 -1250 1783 -1202
rect 1687 -1314 1703 -1250
rect 1767 -1314 1783 -1250
rect 1687 -1330 1783 -1314
rect 1687 -1394 1703 -1330
rect 1767 -1394 1783 -1330
rect 1687 -1410 1783 -1394
rect 1687 -1474 1703 -1410
rect 1767 -1474 1783 -1410
rect 1687 -1490 1783 -1474
rect 1687 -1554 1703 -1490
rect 1767 -1554 1783 -1490
rect 1687 -1604 1783 -1554
<< properties >>
string FIXED_BBOX 1088 1100 1688 1700
<< end >>
