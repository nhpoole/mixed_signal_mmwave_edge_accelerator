magic
tech sky130A
timestamp 1626065694
<< checkpaint >>
rect -798 -720 798 720
<< metal4 >>
rect -168 59 168 90
rect -168 -59 -139 59
rect -21 -59 21 59
rect 139 -59 168 59
rect -168 -90 168 -59
<< via4 >>
rect -139 -59 -21 59
rect 21 -59 139 59
<< metal5 >>
rect -168 59 168 90
rect -168 -59 -139 59
rect -21 -59 21 59
rect 139 -59 168 59
rect -168 -90 168 -59
<< end >>
