magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -1461 -1559 1461 1545
<< pwell >>
rect -201 -299 201 285
<< nmos >>
rect -15 -65 15 65
<< ndiff >>
rect -73 51 -15 65
rect -73 17 -61 51
rect -27 17 -15 51
rect -73 -17 -15 17
rect -73 -51 -61 -17
rect -27 -51 -15 -17
rect -73 -65 -15 -51
rect 15 51 73 65
rect 15 17 27 51
rect 61 17 73 51
rect 15 -17 73 17
rect 15 -51 27 -17
rect 61 -51 73 -17
rect 15 -65 73 -51
<< ndiffc >>
rect -61 17 -27 51
rect -61 -51 -27 -17
rect 27 17 61 51
rect 27 -51 61 -17
<< psubdiff >>
rect -175 225 -51 259
rect -17 225 17 259
rect 51 225 175 259
rect -175 85 -141 225
rect 141 85 175 225
rect -175 17 -141 51
rect -175 -51 -141 -17
rect 141 17 175 51
rect 141 -51 175 -17
rect -175 -239 -141 -85
rect 141 -239 175 -85
rect -175 -273 -51 -239
rect -17 -273 17 -239
rect 51 -273 175 -239
<< psubdiffcont >>
rect -51 225 -17 259
rect 17 225 51 259
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect -51 -273 -17 -239
rect 17 -273 51 -239
<< poly >>
rect -33 137 33 153
rect -33 103 -17 137
rect 17 103 33 137
rect -33 87 33 103
rect -15 65 15 87
rect -15 -87 15 -65
rect -33 -103 33 -87
rect -33 -137 -17 -103
rect 17 -137 33 -103
rect -33 -153 33 -137
<< polycont >>
rect -17 103 17 137
rect -17 -137 17 -103
<< locali >>
rect -175 225 -51 259
rect -17 225 17 259
rect 51 225 175 259
rect -175 85 -141 225
rect -33 103 -17 137
rect 17 103 33 137
rect 141 85 175 225
rect -175 17 -141 51
rect -175 -51 -141 -17
rect -61 53 -27 69
rect -61 -17 -27 17
rect -61 -69 -27 -53
rect 27 53 61 69
rect 27 -17 61 17
rect 27 -69 61 -53
rect 141 17 175 51
rect 141 -51 175 -17
rect -175 -239 -141 -85
rect -33 -137 -17 -103
rect 17 -137 33 -103
rect 141 -239 175 -85
rect -175 -273 -51 -239
rect -17 -273 17 -239
rect 51 -273 175 -239
<< viali >>
rect -17 103 17 137
rect -61 51 -27 53
rect -61 19 -27 51
rect -61 -51 -27 -19
rect -61 -53 -27 -51
rect 27 51 61 53
rect 27 19 61 51
rect 27 -51 61 -19
rect 27 -53 61 -51
rect -17 -137 17 -103
<< metal1 >>
rect -29 137 29 143
rect -29 103 -17 137
rect 17 103 29 137
rect -29 97 29 103
rect -67 53 -21 65
rect -67 19 -61 53
rect -27 19 -21 53
rect -67 -19 -21 19
rect -67 -53 -61 -19
rect -27 -53 -21 -19
rect -67 -65 -21 -53
rect 21 53 67 65
rect 21 19 27 53
rect 61 19 67 53
rect 21 -19 67 19
rect 21 -53 27 -19
rect 61 -53 67 -19
rect 21 -65 67 -53
rect -29 -103 29 -97
rect -29 -137 -17 -103
rect 17 -137 29 -103
rect -29 -143 29 -137
<< properties >>
string FIXED_BBOX -158 -222 158 222
<< end >>
