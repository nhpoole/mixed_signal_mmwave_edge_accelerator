magic
tech sky130A
magscale 1 2
timestamp 1622096065
<< nwell >>
rect -452 -300 452 300
<< pmos >>
rect -358 -200 -158 200
rect -100 -200 100 200
rect 158 -200 358 200
<< pdiff >>
rect -416 188 -358 200
rect -416 -188 -404 188
rect -370 -188 -358 188
rect -416 -200 -358 -188
rect -158 188 -100 200
rect -158 -188 -146 188
rect -112 -188 -100 188
rect -158 -200 -100 -188
rect 100 188 158 200
rect 100 -188 112 188
rect 146 -188 158 188
rect 100 -200 158 -188
rect 358 188 416 200
rect 358 -188 370 188
rect 404 -188 416 188
rect 358 -200 416 -188
<< pdiffc >>
rect -404 -188 -370 188
rect -146 -188 -112 188
rect 112 -188 146 188
rect 370 -188 404 188
<< poly >>
rect -324 281 -192 297
rect -324 264 -308 281
rect -358 247 -308 264
rect -208 264 -192 281
rect -66 281 66 297
rect -66 264 -50 281
rect -208 247 -158 264
rect -358 200 -158 247
rect -100 247 -50 264
rect 50 264 66 281
rect 192 281 324 297
rect 192 264 208 281
rect 50 247 100 264
rect -100 200 100 247
rect 158 247 208 264
rect 308 264 324 281
rect 308 247 358 264
rect 158 200 358 247
rect -358 -247 -158 -200
rect -358 -264 -308 -247
rect -324 -281 -308 -264
rect -208 -264 -158 -247
rect -100 -247 100 -200
rect -100 -264 -50 -247
rect -208 -281 -192 -264
rect -324 -297 -192 -281
rect -66 -281 -50 -264
rect 50 -264 100 -247
rect 158 -247 358 -200
rect 158 -264 208 -247
rect 50 -281 66 -264
rect -66 -297 66 -281
rect 192 -281 208 -264
rect 308 -264 358 -247
rect 308 -281 324 -264
rect 192 -297 324 -281
<< polycont >>
rect -308 247 -208 281
rect -50 247 50 281
rect 208 247 308 281
rect -308 -281 -208 -247
rect -50 -281 50 -247
rect 208 -281 308 -247
<< locali >>
rect -324 247 -308 281
rect -208 247 -192 281
rect -66 247 -50 281
rect 50 247 66 281
rect 192 247 208 281
rect 308 247 324 281
rect -404 188 -370 204
rect -404 -204 -370 -188
rect -146 188 -112 204
rect -146 -204 -112 -188
rect 112 188 146 204
rect 112 -204 146 -188
rect 370 188 404 204
rect 370 -204 404 -188
rect -324 -281 -308 -247
rect -208 -281 -192 -247
rect -66 -281 -50 -247
rect 50 -281 66 -247
rect 192 -281 208 -247
rect 308 -281 324 -247
<< viali >>
rect -300 247 -216 281
rect -42 247 42 281
rect 216 247 300 281
rect -404 -188 -370 188
rect -146 -188 -112 188
rect 112 -188 146 188
rect 370 -188 404 188
rect -300 -281 -216 -247
rect -42 -281 42 -247
rect 216 -281 300 -247
<< metal1 >>
rect -312 281 -204 287
rect -312 247 -300 281
rect -216 247 -204 281
rect -312 241 -204 247
rect -54 281 54 287
rect -54 247 -42 281
rect 42 247 54 281
rect -54 241 54 247
rect 204 281 312 287
rect 204 247 216 281
rect 300 247 312 281
rect 204 241 312 247
rect -410 188 -364 200
rect -410 -188 -404 188
rect -370 -188 -364 188
rect -410 -200 -364 -188
rect -152 188 -106 200
rect -152 -188 -146 188
rect -112 -188 -106 188
rect -152 -200 -106 -188
rect 106 188 152 200
rect 106 -188 112 188
rect 146 -188 152 188
rect 106 -200 152 -188
rect 364 188 410 200
rect 364 -188 370 188
rect 404 -188 410 188
rect 364 -200 410 -188
rect -312 -247 -204 -241
rect -312 -281 -300 -247
rect -216 -281 -204 -247
rect -312 -287 -204 -281
rect -54 -247 54 -241
rect -54 -281 -42 -247
rect 42 -281 54 -247
rect -54 -287 54 -281
rect 204 -247 312 -241
rect 204 -281 216 -247
rect 300 -281 312 -247
rect 204 -287 312 -281
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 2 l 1 m 1 nf 3 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
