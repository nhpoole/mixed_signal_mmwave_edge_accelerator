magic
tech sky130A
magscale 1 2
timestamp 1623661481
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 30 -17 64 17
<< locali >>
rect 22 261 66 393
rect 103 349 169 417
rect 271 349 337 417
rect 395 349 505 417
rect 607 349 673 417
rect 103 315 673 349
rect 22 215 350 261
rect 395 198 473 315
rect 517 199 711 265
rect 755 215 1093 257
rect 1219 215 1539 260
rect 1659 215 1997 256
rect 439 161 473 198
rect 439 127 1113 161
rect 1961 151 1997 215
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 19 451 741 485
rect 707 349 741 451
rect 779 383 845 527
rect 879 349 913 493
rect 954 383 1088 527
rect 1128 349 1162 493
rect 1243 383 1309 527
rect 1343 349 1377 493
rect 1411 383 1477 527
rect 1511 349 1545 493
rect 1683 383 1749 527
rect 1783 349 1817 493
rect 1851 383 1917 527
rect 1951 349 1985 493
rect 707 315 1985 349
rect 35 127 405 161
rect 1243 127 1901 161
rect 35 51 69 127
rect 103 17 169 93
rect 203 51 237 127
rect 371 93 405 127
rect 271 17 337 93
rect 371 59 757 93
rect 795 59 1561 93
rect 1599 17 1665 93
rect 1699 51 1733 127
rect 1767 17 1833 93
rect 1867 51 1901 127
rect 1937 17 2005 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< labels >>
rlabel locali s 755 215 1093 257 6 A1
port 1 nsew signal input
rlabel locali s 1219 215 1539 260 6 A2
port 2 nsew signal input
rlabel locali s 1961 151 1997 215 6 A3
port 3 nsew signal input
rlabel locali s 1659 215 1997 256 6 A3
port 3 nsew signal input
rlabel locali s 517 199 711 265 6 B1
port 4 nsew signal input
rlabel locali s 22 261 66 393 6 B2
port 5 nsew signal input
rlabel locali s 22 215 350 261 6 B2
port 5 nsew signal input
rlabel locali s 607 349 673 417 6 Y
port 6 nsew signal output
rlabel locali s 439 161 473 198 6 Y
port 6 nsew signal output
rlabel locali s 439 127 1113 161 6 Y
port 6 nsew signal output
rlabel locali s 395 349 505 417 6 Y
port 6 nsew signal output
rlabel locali s 395 198 473 315 6 Y
port 6 nsew signal output
rlabel locali s 271 349 337 417 6 Y
port 6 nsew signal output
rlabel locali s 103 349 169 417 6 Y
port 6 nsew signal output
rlabel locali s 103 315 673 349 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -48 2024 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 17 8 VNB
port 8 nsew ground bidirectional
rlabel nwell s -38 261 2062 582 6 VPB
port 9 nsew power bidirectional
rlabel metal1 s 0 496 2024 592 6 VPWR
port 10 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2024 544
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
