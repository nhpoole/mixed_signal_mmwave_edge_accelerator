magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< pwell >>
rect -26 -26 284 278
<< scnmos >>
rect 60 0 90 252
rect 168 0 198 252
<< ndiff >>
rect 0 0 60 252
rect 90 0 168 252
rect 198 0 258 252
<< poly >>
rect 60 278 198 308
rect 60 252 90 278
rect 168 252 198 278
rect 60 -26 90 0
rect 168 -26 198 0
<< locali >>
rect 8 93 42 159
rect 112 93 146 159
rect 216 93 250 159
use contact_11  contact_11_2
timestamp 1624494425
transform 1 0 0 0 1 93
box -26 -22 76 88
use contact_11  contact_11_1
timestamp 1624494425
transform 1 0 104 0 1 93
box -26 -22 76 88
use contact_11  contact_11_0
timestamp 1624494425
transform 1 0 208 0 1 93
box -26 -22 76 88
<< labels >>
rlabel poly s 129 293 129 293 4 G
rlabel locali s 25 126 25 126 4 S
rlabel locali s 233 126 233 126 4 S
rlabel locali s 129 126 129 126 4 D
<< properties >>
string FIXED_BBOX -25 -26 283 308
<< end >>
