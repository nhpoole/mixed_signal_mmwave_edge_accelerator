magic
tech sky130A
magscale 1 2
timestamp 1621829047
<< nwell >>
rect -1796 -819 1796 819
<< pmoshvt >>
rect -1600 -600 1600 600
<< pdiff >>
rect -1658 588 -1600 600
rect -1658 -588 -1646 588
rect -1612 -588 -1600 588
rect -1658 -600 -1600 -588
rect 1600 588 1658 600
rect 1600 -588 1612 588
rect 1646 -588 1658 588
rect 1600 -600 1658 -588
<< pdiffc >>
rect -1646 -588 -1612 588
rect 1612 -588 1646 588
<< nsubdiff >>
rect -1760 749 -1664 783
rect 1664 749 1760 783
rect -1760 687 -1726 749
rect 1726 687 1760 749
rect -1760 -749 -1726 -687
rect 1726 -749 1760 -687
rect -1760 -783 -1664 -749
rect 1664 -783 1760 -749
<< nsubdiffcont >>
rect -1664 749 1664 783
rect -1760 -687 -1726 687
rect 1726 -687 1760 687
rect -1664 -783 1664 -749
<< poly >>
rect -966 681 966 697
rect -966 664 -950 681
rect -1600 647 -950 664
rect 950 664 966 681
rect 950 647 1600 664
rect -1600 600 1600 647
rect -1600 -647 1600 -600
rect -1600 -664 -950 -647
rect -966 -681 -950 -664
rect 950 -664 1600 -647
rect 950 -681 966 -664
rect -966 -697 966 -681
<< polycont >>
rect -950 647 950 681
rect -950 -681 950 -647
<< locali >>
rect -1760 749 -1664 783
rect 1664 749 1760 783
rect -1760 687 -1726 749
rect 1726 687 1760 749
rect -966 647 -950 681
rect 950 647 966 681
rect -1646 588 -1612 604
rect -1646 -604 -1612 -588
rect 1612 588 1646 604
rect 1612 -604 1646 -588
rect -966 -681 -950 -647
rect 950 -681 966 -647
rect -1760 -749 -1726 -687
rect 1726 -749 1760 -687
rect -1760 -783 -1664 -749
rect 1664 -783 1760 -749
<< viali >>
rect -792 647 792 681
rect -1646 -588 -1612 588
rect 1612 -588 1646 588
rect -792 -681 792 -647
<< metal1 >>
rect -804 681 804 687
rect -804 647 -792 681
rect 792 647 804 681
rect -804 641 804 647
rect -1652 588 -1606 600
rect -1652 -588 -1646 588
rect -1612 -588 -1606 588
rect -1652 -600 -1606 -588
rect 1606 588 1652 600
rect 1606 -588 1612 588
rect 1646 -588 1652 588
rect 1606 -600 1652 -588
rect -804 -647 804 -641
rect -804 -681 -792 -647
rect 792 -681 804 -647
rect -804 -687 804 -681
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_hvt
string FIXED_BBOX -1743 -766 1743 766
string parameters w 6 l 16 m 1 nf 1 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
