magic
tech sky130A
magscale 1 2
timestamp 1620621618
<< nmoslvt >>
rect -561 -100 -501 100
rect -443 -100 -383 100
rect -325 -100 -265 100
rect -207 -100 -147 100
rect -89 -100 -29 100
rect 29 -100 89 100
rect 147 -100 207 100
rect 265 -100 325 100
rect 383 -100 443 100
rect 501 -100 561 100
<< ndiff >>
rect -619 88 -561 100
rect -619 -88 -607 88
rect -573 -88 -561 88
rect -619 -100 -561 -88
rect -501 88 -443 100
rect -501 -88 -489 88
rect -455 -88 -443 88
rect -501 -100 -443 -88
rect -383 88 -325 100
rect -383 -88 -371 88
rect -337 -88 -325 88
rect -383 -100 -325 -88
rect -265 88 -207 100
rect -265 -88 -253 88
rect -219 -88 -207 88
rect -265 -100 -207 -88
rect -147 88 -89 100
rect -147 -88 -135 88
rect -101 -88 -89 88
rect -147 -100 -89 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 89 88 147 100
rect 89 -88 101 88
rect 135 -88 147 88
rect 89 -100 147 -88
rect 207 88 265 100
rect 207 -88 219 88
rect 253 -88 265 88
rect 207 -100 265 -88
rect 325 88 383 100
rect 325 -88 337 88
rect 371 -88 383 88
rect 325 -100 383 -88
rect 443 88 501 100
rect 443 -88 455 88
rect 489 -88 501 88
rect 443 -100 501 -88
rect 561 88 619 100
rect 561 -88 573 88
rect 607 -88 619 88
rect 561 -100 619 -88
<< ndiffc >>
rect -607 -88 -573 88
rect -489 -88 -455 88
rect -371 -88 -337 88
rect -253 -88 -219 88
rect -135 -88 -101 88
rect -17 -88 17 88
rect 101 -88 135 88
rect 219 -88 253 88
rect 337 -88 371 88
rect 455 -88 489 88
rect 573 -88 607 88
<< poly >>
rect -561 100 -501 126
rect -443 100 -383 126
rect -325 100 -265 126
rect -207 100 -147 126
rect -89 100 -29 126
rect 29 100 89 126
rect 147 100 207 126
rect 265 100 325 126
rect 383 100 443 126
rect 501 100 561 126
rect -561 -126 -501 -100
rect -443 -126 -383 -100
rect -325 -126 -265 -100
rect -207 -126 -147 -100
rect -89 -126 -29 -100
rect 29 -126 89 -100
rect 147 -126 207 -100
rect 265 -126 325 -100
rect 383 -126 443 -100
rect 501 -126 561 -100
<< locali >>
rect -607 88 -573 104
rect -607 -104 -573 -88
rect -489 88 -455 104
rect -489 -104 -455 -88
rect -371 88 -337 104
rect -371 -104 -337 -88
rect -253 88 -219 104
rect -253 -104 -219 -88
rect -135 88 -101 104
rect -135 -104 -101 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 101 88 135 104
rect 101 -104 135 -88
rect 219 88 253 104
rect 219 -104 253 -88
rect 337 88 371 104
rect 337 -104 371 -88
rect 455 88 489 104
rect 455 -104 489 -88
rect 573 88 607 104
rect 573 -104 607 -88
<< viali >>
rect -607 -88 -573 88
rect -489 -88 -455 88
rect -371 -88 -337 88
rect -253 -88 -219 88
rect -135 -88 -101 88
rect -17 -88 17 88
rect 101 -88 135 88
rect 219 -88 253 88
rect 337 -88 371 88
rect 455 -88 489 88
rect 573 -88 607 88
<< metal1 >>
rect -613 88 -567 100
rect -613 -88 -607 88
rect -573 -88 -567 88
rect -613 -100 -567 -88
rect -495 88 -449 100
rect -495 -88 -489 88
rect -455 -88 -449 88
rect -495 -100 -449 -88
rect -377 88 -331 100
rect -377 -88 -371 88
rect -337 -88 -331 88
rect -377 -100 -331 -88
rect -259 88 -213 100
rect -259 -88 -253 88
rect -219 -88 -213 88
rect -259 -100 -213 -88
rect -141 88 -95 100
rect -141 -88 -135 88
rect -101 -88 -95 88
rect -141 -100 -95 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 95 88 141 100
rect 95 -88 101 88
rect 135 -88 141 88
rect 95 -100 141 -88
rect 213 88 259 100
rect 213 -88 219 88
rect 253 -88 259 88
rect 213 -100 259 -88
rect 331 88 377 100
rect 331 -88 337 88
rect 371 -88 377 88
rect 331 -100 377 -88
rect 449 88 495 100
rect 449 -88 455 88
rect 489 -88 495 88
rect 449 -100 495 -88
rect 567 88 613 100
rect 567 -88 573 88
rect 607 -88 613 88
rect 567 -100 613 -88
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string parameters w 1 l 0.3 m 1 nf 10 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
