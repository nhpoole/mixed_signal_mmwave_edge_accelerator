magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -2099 -1460 2099 1460
<< nwell >>
rect -839 -200 839 200
<< pmos >>
rect -745 -100 -545 100
rect -487 -100 -287 100
rect -229 -100 -29 100
rect 29 -100 229 100
rect 287 -100 487 100
rect 545 -100 745 100
<< pdiff >>
rect -803 85 -745 100
rect -803 51 -791 85
rect -757 51 -745 85
rect -803 17 -745 51
rect -803 -17 -791 17
rect -757 -17 -745 17
rect -803 -51 -745 -17
rect -803 -85 -791 -51
rect -757 -85 -745 -51
rect -803 -100 -745 -85
rect -545 85 -487 100
rect -545 51 -533 85
rect -499 51 -487 85
rect -545 17 -487 51
rect -545 -17 -533 17
rect -499 -17 -487 17
rect -545 -51 -487 -17
rect -545 -85 -533 -51
rect -499 -85 -487 -51
rect -545 -100 -487 -85
rect -287 85 -229 100
rect -287 51 -275 85
rect -241 51 -229 85
rect -287 17 -229 51
rect -287 -17 -275 17
rect -241 -17 -229 17
rect -287 -51 -229 -17
rect -287 -85 -275 -51
rect -241 -85 -229 -51
rect -287 -100 -229 -85
rect -29 85 29 100
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -100 29 -85
rect 229 85 287 100
rect 229 51 241 85
rect 275 51 287 85
rect 229 17 287 51
rect 229 -17 241 17
rect 275 -17 287 17
rect 229 -51 287 -17
rect 229 -85 241 -51
rect 275 -85 287 -51
rect 229 -100 287 -85
rect 487 85 545 100
rect 487 51 499 85
rect 533 51 545 85
rect 487 17 545 51
rect 487 -17 499 17
rect 533 -17 545 17
rect 487 -51 545 -17
rect 487 -85 499 -51
rect 533 -85 545 -51
rect 487 -100 545 -85
rect 745 85 803 100
rect 745 51 757 85
rect 791 51 803 85
rect 745 17 803 51
rect 745 -17 757 17
rect 791 -17 803 17
rect 745 -51 803 -17
rect 745 -85 757 -51
rect 791 -85 803 -51
rect 745 -100 803 -85
<< pdiffc >>
rect -791 51 -757 85
rect -791 -17 -757 17
rect -791 -85 -757 -51
rect -533 51 -499 85
rect -533 -17 -499 17
rect -533 -85 -499 -51
rect -275 51 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 241 51 275 85
rect 241 -17 275 17
rect 241 -85 275 -51
rect 499 51 533 85
rect 499 -17 533 17
rect 499 -85 533 -51
rect 757 51 791 85
rect 757 -17 791 17
rect 757 -85 791 -51
<< poly >>
rect -711 181 -579 197
rect -711 164 -662 181
rect -745 147 -662 164
rect -628 164 -579 181
rect -453 181 -321 197
rect -453 164 -404 181
rect -628 147 -545 164
rect -745 100 -545 147
rect -487 147 -404 164
rect -370 164 -321 181
rect -195 181 -63 197
rect -195 164 -146 181
rect -370 147 -287 164
rect -487 100 -287 147
rect -229 147 -146 164
rect -112 164 -63 181
rect 63 181 195 197
rect 63 164 112 181
rect -112 147 -29 164
rect -229 100 -29 147
rect 29 147 112 164
rect 146 164 195 181
rect 321 181 453 197
rect 321 164 370 181
rect 146 147 229 164
rect 29 100 229 147
rect 287 147 370 164
rect 404 164 453 181
rect 579 181 711 197
rect 579 164 628 181
rect 404 147 487 164
rect 287 100 487 147
rect 545 147 628 164
rect 662 164 711 181
rect 662 147 745 164
rect 545 100 745 147
rect -745 -147 -545 -100
rect -745 -164 -662 -147
rect -711 -181 -662 -164
rect -628 -164 -545 -147
rect -487 -147 -287 -100
rect -487 -164 -404 -147
rect -628 -181 -579 -164
rect -711 -197 -579 -181
rect -453 -181 -404 -164
rect -370 -164 -287 -147
rect -229 -147 -29 -100
rect -229 -164 -146 -147
rect -370 -181 -321 -164
rect -453 -197 -321 -181
rect -195 -181 -146 -164
rect -112 -164 -29 -147
rect 29 -147 229 -100
rect 29 -164 112 -147
rect -112 -181 -63 -164
rect -195 -197 -63 -181
rect 63 -181 112 -164
rect 146 -164 229 -147
rect 287 -147 487 -100
rect 287 -164 370 -147
rect 146 -181 195 -164
rect 63 -197 195 -181
rect 321 -181 370 -164
rect 404 -164 487 -147
rect 545 -147 745 -100
rect 545 -164 628 -147
rect 404 -181 453 -164
rect 321 -197 453 -181
rect 579 -181 628 -164
rect 662 -164 745 -147
rect 662 -181 711 -164
rect 579 -197 711 -181
<< polycont >>
rect -662 147 -628 181
rect -404 147 -370 181
rect -146 147 -112 181
rect 112 147 146 181
rect 370 147 404 181
rect 628 147 662 181
rect -662 -181 -628 -147
rect -404 -181 -370 -147
rect -146 -181 -112 -147
rect 112 -181 146 -147
rect 370 -181 404 -147
rect 628 -181 662 -147
<< locali >>
rect -711 147 -662 181
rect -628 147 -579 181
rect -453 147 -404 181
rect -370 147 -321 181
rect -195 147 -146 181
rect -112 147 -63 181
rect 63 147 112 181
rect 146 147 195 181
rect 321 147 370 181
rect 404 147 453 181
rect 579 147 628 181
rect 662 147 711 181
rect -791 85 -757 104
rect -791 17 -757 19
rect -791 -19 -757 -17
rect -791 -104 -757 -85
rect -533 85 -499 104
rect -533 17 -499 19
rect -533 -19 -499 -17
rect -533 -104 -499 -85
rect -275 85 -241 104
rect -275 17 -241 19
rect -275 -19 -241 -17
rect -275 -104 -241 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 241 85 275 104
rect 241 17 275 19
rect 241 -19 275 -17
rect 241 -104 275 -85
rect 499 85 533 104
rect 499 17 533 19
rect 499 -19 533 -17
rect 499 -104 533 -85
rect 757 85 791 104
rect 757 17 791 19
rect 757 -19 791 -17
rect 757 -104 791 -85
rect -711 -181 -662 -147
rect -628 -181 -579 -147
rect -453 -181 -404 -147
rect -370 -181 -321 -147
rect -195 -181 -146 -147
rect -112 -181 -63 -147
rect 63 -181 112 -147
rect 146 -181 195 -147
rect 321 -181 370 -147
rect 404 -181 453 -147
rect 579 -181 628 -147
rect 662 -181 711 -147
<< viali >>
rect -662 147 -628 181
rect -404 147 -370 181
rect -146 147 -112 181
rect 112 147 146 181
rect 370 147 404 181
rect 628 147 662 181
rect -791 51 -757 53
rect -791 19 -757 51
rect -791 -51 -757 -19
rect -791 -53 -757 -51
rect -533 51 -499 53
rect -533 19 -499 51
rect -533 -51 -499 -19
rect -533 -53 -499 -51
rect -275 51 -241 53
rect -275 19 -241 51
rect -275 -51 -241 -19
rect -275 -53 -241 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 241 51 275 53
rect 241 19 275 51
rect 241 -51 275 -19
rect 241 -53 275 -51
rect 499 51 533 53
rect 499 19 533 51
rect 499 -51 533 -19
rect 499 -53 533 -51
rect 757 51 791 53
rect 757 19 791 51
rect 757 -51 791 -19
rect 757 -53 791 -51
rect -662 -181 -628 -147
rect -404 -181 -370 -147
rect -146 -181 -112 -147
rect 112 -181 146 -147
rect 370 -181 404 -147
rect 628 -181 662 -147
<< metal1 >>
rect -699 181 -591 187
rect -699 147 -662 181
rect -628 147 -591 181
rect -699 141 -591 147
rect -441 181 -333 187
rect -441 147 -404 181
rect -370 147 -333 181
rect -441 141 -333 147
rect -183 181 -75 187
rect -183 147 -146 181
rect -112 147 -75 181
rect -183 141 -75 147
rect 75 181 183 187
rect 75 147 112 181
rect 146 147 183 181
rect 75 141 183 147
rect 333 181 441 187
rect 333 147 370 181
rect 404 147 441 181
rect 333 141 441 147
rect 591 181 699 187
rect 591 147 628 181
rect 662 147 699 181
rect 591 141 699 147
rect -797 53 -751 100
rect -797 19 -791 53
rect -757 19 -751 53
rect -797 -19 -751 19
rect -797 -53 -791 -19
rect -757 -53 -751 -19
rect -797 -100 -751 -53
rect -539 53 -493 100
rect -539 19 -533 53
rect -499 19 -493 53
rect -539 -19 -493 19
rect -539 -53 -533 -19
rect -499 -53 -493 -19
rect -539 -100 -493 -53
rect -281 53 -235 100
rect -281 19 -275 53
rect -241 19 -235 53
rect -281 -19 -235 19
rect -281 -53 -275 -19
rect -241 -53 -235 -19
rect -281 -100 -235 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 235 53 281 100
rect 235 19 241 53
rect 275 19 281 53
rect 235 -19 281 19
rect 235 -53 241 -19
rect 275 -53 281 -19
rect 235 -100 281 -53
rect 493 53 539 100
rect 493 19 499 53
rect 533 19 539 53
rect 493 -19 539 19
rect 493 -53 499 -19
rect 533 -53 539 -19
rect 493 -100 539 -53
rect 751 53 797 100
rect 751 19 757 53
rect 791 19 797 53
rect 751 -19 797 19
rect 751 -53 757 -19
rect 791 -53 797 -19
rect 751 -100 797 -53
rect -699 -147 -591 -141
rect -699 -181 -662 -147
rect -628 -181 -591 -147
rect -699 -187 -591 -181
rect -441 -147 -333 -141
rect -441 -181 -404 -147
rect -370 -181 -333 -147
rect -441 -187 -333 -181
rect -183 -147 -75 -141
rect -183 -181 -146 -147
rect -112 -181 -75 -147
rect -183 -187 -75 -181
rect 75 -147 183 -141
rect 75 -181 112 -147
rect 146 -181 183 -147
rect 75 -187 183 -181
rect 333 -147 441 -141
rect 333 -181 370 -147
rect 404 -181 441 -147
rect 333 -187 441 -181
rect 591 -147 699 -141
rect 591 -181 628 -147
rect 662 -181 699 -147
rect 591 -187 699 -181
<< end >>
