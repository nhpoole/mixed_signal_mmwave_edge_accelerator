magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -1319 -1314 1469 1424
<< nwell >>
rect -54 -54 204 164
<< scpmos >>
rect 60 0 90 110
<< pdiff >>
rect 0 0 60 110
rect 90 0 150 110
<< poly >>
rect 60 110 90 136
rect 60 -26 90 0
<< locali >>
rect 8 22 42 88
rect 108 22 142 88
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_0
timestamp 1626486988
transform 1 0 100 0 1 22
box -59 -51 109 117
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_1
timestamp 1626486988
transform 1 0 0 0 1 22
box -59 -51 109 117
<< labels >>
rlabel locali s 25 55 25 55 4 S
rlabel locali s 125 55 125 55 4 D
rlabel poly s 75 55 75 55 4 G
<< properties >>
string FIXED_BBOX -54 -54 204 164
<< end >>
