magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -3934 -4166 4581 1714
<< nwell >>
rect -2454 122 3321 444
rect -2622 -634 3320 -398
rect -2622 -730 -2260 -634
rect -2242 -730 3320 -634
rect -2622 -966 3320 -730
rect -2622 -2054 3320 -1486
rect -2622 -2896 3320 -2574
<< locali >>
rect -2214 139 -2166 146
rect -2214 105 -2207 139
rect -2173 105 -2166 139
rect -2214 98 -2166 105
rect -552 119 -504 126
rect -1962 81 -1914 88
rect -1962 47 -1955 81
rect -1921 47 -1914 81
rect -552 85 -545 119
rect -511 85 -504 119
rect -552 78 -504 85
rect -436 119 -388 126
rect -436 85 -429 119
rect -395 85 -388 119
rect -436 78 -388 85
rect -324 119 -276 126
rect -324 85 -317 119
rect -283 85 -276 119
rect -324 78 -276 85
rect -192 119 -144 126
rect -192 85 -185 119
rect -151 85 -144 119
rect -192 78 -144 85
rect -82 119 -34 126
rect -82 85 -75 119
rect -41 85 -34 119
rect -82 78 -34 85
rect 34 119 82 126
rect 34 85 41 119
rect 75 85 82 119
rect 34 78 82 85
rect 166 117 214 124
rect 166 83 173 117
rect 207 83 214 117
rect 166 76 214 83
rect -1962 40 -1914 47
rect -858 1 -810 8
rect -858 -33 -851 1
rect -817 -33 -810 1
rect -858 -40 -810 -33
rect -2584 -155 -2555 -121
rect -2521 -155 -2492 -121
rect 3190 -155 3219 -121
rect 3253 -155 3282 -121
rect -2567 -198 -2509 -155
rect 3207 -198 3265 -155
rect 1842 -247 1890 -240
rect 1842 -281 1849 -247
rect 1883 -281 1890 -247
rect 1842 -288 1890 -281
rect -1962 -323 -1914 -316
rect -1962 -357 -1955 -323
rect -1921 -357 -1914 -323
rect 736 -323 784 -316
rect -1962 -364 -1914 -357
rect -552 -361 -504 -354
rect -2218 -371 -2170 -364
rect -2218 -405 -2211 -371
rect -2177 -405 -2170 -371
rect -552 -395 -545 -361
rect -511 -395 -504 -361
rect -552 -402 -504 -395
rect -436 -361 -388 -354
rect -436 -395 -429 -361
rect -395 -395 -388 -361
rect -436 -402 -388 -395
rect -324 -361 -276 -354
rect -324 -395 -317 -361
rect -283 -395 -276 -361
rect -324 -402 -276 -395
rect -192 -361 -144 -354
rect -192 -395 -185 -361
rect -151 -395 -144 -361
rect -192 -402 -144 -395
rect -82 -361 -34 -354
rect -82 -395 -75 -361
rect -41 -395 -34 -361
rect -82 -402 -34 -395
rect 34 -361 82 -354
rect 34 -395 41 -361
rect 75 -395 82 -361
rect 34 -402 82 -395
rect 170 -359 218 -352
rect 170 -393 177 -359
rect 211 -393 218 -359
rect 736 -357 743 -323
rect 777 -357 784 -323
rect 736 -364 784 -357
rect 2146 -361 2194 -354
rect 170 -400 218 -393
rect 2146 -395 2153 -361
rect 2187 -395 2194 -361
rect 2146 -402 2194 -395
rect 2262 -361 2310 -354
rect 2262 -395 2269 -361
rect 2303 -395 2310 -361
rect 2262 -402 2310 -395
rect 2374 -361 2422 -354
rect 2374 -395 2381 -361
rect 2415 -395 2422 -361
rect 2374 -402 2422 -395
rect 2506 -361 2554 -354
rect 2506 -395 2513 -361
rect 2547 -395 2554 -361
rect 2506 -402 2554 -395
rect 2616 -361 2664 -354
rect 2616 -395 2623 -361
rect 2657 -395 2664 -361
rect 2616 -402 2664 -395
rect 2732 -361 2780 -354
rect 2732 -395 2739 -361
rect 2773 -395 2780 -361
rect 2732 -402 2780 -395
rect 2864 -359 2912 -352
rect 2864 -393 2871 -359
rect 2905 -393 2912 -359
rect 2864 -400 2912 -393
rect -2218 -412 -2170 -405
rect 480 -413 528 -406
rect 480 -447 487 -413
rect 521 -447 528 -413
rect 480 -454 528 -447
rect -858 -545 -810 -538
rect -858 -579 -851 -545
rect -817 -579 -810 -545
rect -858 -586 -810 -579
rect -2567 -665 -2509 -622
rect 3207 -665 3265 -622
rect -2584 -699 -2555 -665
rect -2521 -699 -2492 -665
rect 3190 -699 3219 -665
rect 3253 -699 3282 -665
rect -2567 -742 -2509 -699
rect 3207 -742 3265 -699
rect 1840 -785 1888 -778
rect 1840 -819 1847 -785
rect 1881 -819 1888 -785
rect 1840 -826 1888 -819
rect -2218 -917 -2170 -910
rect -2218 -951 -2211 -917
rect -2177 -951 -2170 -917
rect -2218 -958 -2170 -951
rect 480 -957 528 -950
rect -552 -969 -504 -962
rect -1962 -1007 -1914 -1000
rect -1962 -1041 -1955 -1007
rect -1921 -1041 -1914 -1007
rect -552 -1003 -545 -969
rect -511 -1003 -504 -969
rect -552 -1010 -504 -1003
rect -436 -969 -388 -962
rect -436 -1003 -429 -969
rect -395 -1003 -388 -969
rect -436 -1010 -388 -1003
rect -324 -969 -276 -962
rect -324 -1003 -317 -969
rect -283 -1003 -276 -969
rect -324 -1010 -276 -1003
rect -192 -969 -144 -962
rect -192 -1003 -185 -969
rect -151 -1003 -144 -969
rect -192 -1010 -144 -1003
rect -82 -969 -34 -962
rect -82 -1003 -75 -969
rect -41 -1003 -34 -969
rect -82 -1010 -34 -1003
rect 34 -969 82 -962
rect 34 -1003 41 -969
rect 75 -1003 82 -969
rect 34 -1010 82 -1003
rect 166 -971 218 -964
rect 166 -1005 175 -971
rect 209 -1005 218 -971
rect 480 -991 487 -957
rect 521 -991 528 -957
rect 480 -998 528 -991
rect 2146 -969 2194 -962
rect 166 -1012 218 -1005
rect 736 -1007 784 -1000
rect -1962 -1048 -1914 -1041
rect 736 -1041 743 -1007
rect 777 -1041 784 -1007
rect 2146 -1003 2153 -969
rect 2187 -1003 2194 -969
rect 2146 -1010 2194 -1003
rect 2262 -969 2310 -962
rect 2262 -1003 2269 -969
rect 2303 -1003 2310 -969
rect 2262 -1010 2310 -1003
rect 2374 -969 2422 -962
rect 2374 -1003 2381 -969
rect 2415 -1003 2422 -969
rect 2374 -1010 2422 -1003
rect 2506 -969 2554 -962
rect 2506 -1003 2513 -969
rect 2547 -1003 2554 -969
rect 2506 -1010 2554 -1003
rect 2616 -969 2664 -962
rect 2616 -1003 2623 -969
rect 2657 -1003 2664 -969
rect 2616 -1010 2664 -1003
rect 2732 -969 2780 -962
rect 2732 -1003 2739 -969
rect 2773 -1003 2780 -969
rect 2732 -1010 2780 -1003
rect 2864 -971 2912 -964
rect 2864 -1005 2871 -971
rect 2905 -1005 2912 -971
rect 2864 -1012 2912 -1005
rect 736 -1048 784 -1041
rect -858 -1089 -810 -1082
rect -858 -1123 -851 -1089
rect -817 -1123 -810 -1089
rect -858 -1130 -810 -1123
rect -2567 -1209 -2509 -1166
rect 3207 -1209 3265 -1166
rect -2584 -1243 -2555 -1209
rect -2521 -1243 -2492 -1209
rect 3190 -1243 3219 -1209
rect 3253 -1243 3282 -1209
rect -2567 -1286 -2509 -1243
rect 3207 -1286 3265 -1243
rect 1840 -1329 1888 -1322
rect 1840 -1363 1847 -1329
rect 1881 -1363 1888 -1329
rect 1840 -1370 1888 -1363
rect -1962 -1411 -1914 -1404
rect -1962 -1445 -1955 -1411
rect -1921 -1445 -1914 -1411
rect 736 -1411 784 -1404
rect -1962 -1452 -1914 -1445
rect -552 -1449 -504 -1442
rect -2218 -1461 -2170 -1454
rect -2218 -1495 -2211 -1461
rect -2177 -1495 -2170 -1461
rect -552 -1483 -545 -1449
rect -511 -1483 -504 -1449
rect -552 -1490 -504 -1483
rect -436 -1449 -388 -1442
rect -436 -1483 -429 -1449
rect -395 -1483 -388 -1449
rect -436 -1490 -388 -1483
rect -324 -1449 -276 -1442
rect -324 -1483 -317 -1449
rect -283 -1483 -276 -1449
rect -324 -1490 -276 -1483
rect -192 -1449 -144 -1442
rect -192 -1483 -185 -1449
rect -151 -1483 -144 -1449
rect -192 -1490 -144 -1483
rect -82 -1449 -34 -1442
rect -82 -1483 -75 -1449
rect -41 -1483 -34 -1449
rect -82 -1490 -34 -1483
rect 34 -1449 82 -1442
rect 34 -1483 41 -1449
rect 75 -1483 82 -1449
rect 34 -1490 82 -1483
rect 166 -1447 214 -1440
rect 166 -1481 173 -1447
rect 207 -1481 214 -1447
rect 736 -1445 743 -1411
rect 777 -1445 784 -1411
rect 736 -1452 784 -1445
rect 2146 -1449 2194 -1442
rect 166 -1488 214 -1481
rect 2146 -1483 2153 -1449
rect 2187 -1483 2194 -1449
rect 2146 -1490 2194 -1483
rect 2262 -1449 2310 -1442
rect 2262 -1483 2269 -1449
rect 2303 -1483 2310 -1449
rect 2262 -1490 2310 -1483
rect 2374 -1449 2422 -1442
rect 2374 -1483 2381 -1449
rect 2415 -1483 2422 -1449
rect 2374 -1490 2422 -1483
rect 2506 -1449 2554 -1442
rect 2506 -1483 2513 -1449
rect 2547 -1483 2554 -1449
rect 2506 -1490 2554 -1483
rect 2616 -1449 2664 -1442
rect 2616 -1483 2623 -1449
rect 2657 -1483 2664 -1449
rect 2616 -1490 2664 -1483
rect 2732 -1449 2780 -1442
rect 2732 -1483 2739 -1449
rect 2773 -1483 2780 -1449
rect 2732 -1490 2780 -1483
rect 2864 -1447 2916 -1440
rect 2864 -1481 2873 -1447
rect 2907 -1481 2916 -1447
rect 2864 -1488 2916 -1481
rect -2218 -1502 -2170 -1495
rect 480 -1501 528 -1494
rect 480 -1535 487 -1501
rect 521 -1535 528 -1501
rect 480 -1542 528 -1535
rect -858 -1633 -810 -1626
rect -858 -1667 -851 -1633
rect -817 -1667 -810 -1633
rect -858 -1674 -810 -1667
rect -2567 -1753 -2509 -1710
rect 3207 -1753 3265 -1710
rect -2584 -1787 -2555 -1753
rect -2521 -1787 -2492 -1753
rect 3190 -1787 3219 -1753
rect 3253 -1787 3282 -1753
rect -2567 -1830 -2509 -1787
rect 3207 -1830 3265 -1787
rect 1840 -1873 1888 -1866
rect 1840 -1907 1847 -1873
rect 1881 -1907 1888 -1873
rect 1840 -1914 1888 -1907
rect -2218 -2005 -2170 -1998
rect -2218 -2039 -2211 -2005
rect -2177 -2039 -2170 -2005
rect -2218 -2046 -2170 -2039
rect 480 -2047 528 -2040
rect -552 -2057 -504 -2050
rect -1962 -2095 -1914 -2088
rect -1962 -2129 -1955 -2095
rect -1921 -2129 -1914 -2095
rect -552 -2091 -545 -2057
rect -511 -2091 -504 -2057
rect -552 -2098 -504 -2091
rect -436 -2057 -388 -2050
rect -436 -2091 -429 -2057
rect -395 -2091 -388 -2057
rect -436 -2098 -388 -2091
rect -324 -2057 -276 -2050
rect -324 -2091 -317 -2057
rect -283 -2091 -276 -2057
rect -324 -2098 -276 -2091
rect -192 -2057 -144 -2050
rect -192 -2091 -185 -2057
rect -151 -2091 -144 -2057
rect -192 -2098 -144 -2091
rect -82 -2057 -34 -2050
rect -82 -2091 -75 -2057
rect -41 -2091 -34 -2057
rect -82 -2098 -34 -2091
rect 34 -2057 82 -2050
rect 34 -2091 41 -2057
rect 75 -2091 82 -2057
rect 34 -2098 82 -2091
rect 166 -2059 214 -2052
rect 166 -2093 173 -2059
rect 207 -2093 214 -2059
rect 480 -2081 487 -2047
rect 521 -2081 528 -2047
rect 480 -2088 528 -2081
rect 2146 -2057 2194 -2050
rect 166 -2100 214 -2093
rect 736 -2095 784 -2088
rect -1962 -2136 -1914 -2129
rect 736 -2129 743 -2095
rect 777 -2129 784 -2095
rect 2146 -2091 2153 -2057
rect 2187 -2091 2194 -2057
rect 2146 -2098 2194 -2091
rect 2262 -2057 2310 -2050
rect 2262 -2091 2269 -2057
rect 2303 -2091 2310 -2057
rect 2262 -2098 2310 -2091
rect 2374 -2057 2422 -2050
rect 2374 -2091 2381 -2057
rect 2415 -2091 2422 -2057
rect 2374 -2098 2422 -2091
rect 2506 -2057 2554 -2050
rect 2506 -2091 2513 -2057
rect 2547 -2091 2554 -2057
rect 2506 -2098 2554 -2091
rect 2616 -2057 2664 -2050
rect 2616 -2091 2623 -2057
rect 2657 -2091 2664 -2057
rect 2616 -2098 2664 -2091
rect 2732 -2057 2780 -2050
rect 2732 -2091 2739 -2057
rect 2773 -2091 2780 -2057
rect 2732 -2098 2780 -2091
rect 2868 -2059 2916 -2052
rect 2868 -2093 2875 -2059
rect 2909 -2093 2916 -2059
rect 2868 -2100 2916 -2093
rect 736 -2136 784 -2129
rect -858 -2175 -810 -2168
rect -858 -2209 -851 -2175
rect -817 -2209 -810 -2175
rect -858 -2216 -810 -2209
rect -2567 -2297 -2509 -2254
rect 3207 -2297 3265 -2254
rect -2584 -2331 -2555 -2297
rect -2521 -2331 -2492 -2297
rect 3190 -2331 3219 -2297
rect 3253 -2331 3282 -2297
rect -2567 -2374 -2509 -2331
rect 3207 -2374 3265 -2331
rect 1840 -2419 1888 -2412
rect 1840 -2453 1847 -2419
rect 1881 -2453 1888 -2419
rect 1840 -2460 1888 -2453
rect -1962 -2499 -1914 -2492
rect -1962 -2533 -1955 -2499
rect -1921 -2533 -1914 -2499
rect 736 -2499 784 -2492
rect -1962 -2540 -1914 -2533
rect -552 -2537 -504 -2530
rect -2218 -2547 -2170 -2540
rect -2218 -2581 -2211 -2547
rect -2177 -2581 -2170 -2547
rect -552 -2571 -545 -2537
rect -511 -2571 -504 -2537
rect -552 -2578 -504 -2571
rect -436 -2537 -388 -2530
rect -436 -2571 -429 -2537
rect -395 -2571 -388 -2537
rect -436 -2578 -388 -2571
rect -324 -2537 -276 -2530
rect -324 -2571 -317 -2537
rect -283 -2571 -276 -2537
rect -324 -2578 -276 -2571
rect -192 -2537 -144 -2530
rect -192 -2571 -185 -2537
rect -151 -2571 -144 -2537
rect -192 -2578 -144 -2571
rect -82 -2537 -34 -2530
rect -82 -2571 -75 -2537
rect -41 -2571 -34 -2537
rect -82 -2578 -34 -2571
rect 34 -2537 82 -2530
rect 34 -2571 41 -2537
rect 75 -2571 82 -2537
rect 34 -2578 82 -2571
rect 166 -2535 218 -2528
rect 166 -2569 175 -2535
rect 209 -2569 218 -2535
rect 166 -2576 218 -2569
rect 488 -2529 536 -2522
rect 488 -2563 495 -2529
rect 529 -2563 536 -2529
rect 736 -2533 743 -2499
rect 777 -2533 784 -2499
rect 736 -2540 784 -2533
rect 2146 -2537 2194 -2530
rect 488 -2570 536 -2563
rect 2146 -2571 2153 -2537
rect 2187 -2571 2194 -2537
rect 2146 -2578 2194 -2571
rect 2262 -2537 2310 -2530
rect 2262 -2571 2269 -2537
rect 2303 -2571 2310 -2537
rect 2262 -2578 2310 -2571
rect 2374 -2537 2422 -2530
rect 2374 -2571 2381 -2537
rect 2415 -2571 2422 -2537
rect 2374 -2578 2422 -2571
rect 2506 -2537 2554 -2530
rect 2506 -2571 2513 -2537
rect 2547 -2571 2554 -2537
rect 2506 -2578 2554 -2571
rect 2616 -2537 2664 -2530
rect 2616 -2571 2623 -2537
rect 2657 -2571 2664 -2537
rect 2616 -2578 2664 -2571
rect 2732 -2537 2780 -2530
rect 2732 -2571 2739 -2537
rect 2773 -2571 2780 -2537
rect 2732 -2578 2780 -2571
rect 2864 -2535 2912 -2528
rect 2864 -2569 2871 -2535
rect 2905 -2569 2912 -2535
rect 2864 -2576 2912 -2569
rect -2218 -2588 -2170 -2581
rect -858 -2719 -810 -2712
rect -858 -2753 -851 -2719
rect -817 -2753 -810 -2719
rect -858 -2760 -810 -2753
rect -2567 -2841 -2509 -2798
rect 3207 -2841 3265 -2798
rect -2584 -2875 -2555 -2841
rect -2521 -2875 -2492 -2841
rect 3190 -2875 3219 -2841
rect 3253 -2875 3282 -2841
<< viali >>
rect -2207 105 -2173 139
rect -1955 47 -1921 81
rect -545 85 -511 119
rect -429 85 -395 119
rect -317 85 -283 119
rect -185 85 -151 119
rect -75 85 -41 119
rect 41 85 75 119
rect 173 83 207 117
rect -851 -33 -817 1
rect -2555 -155 -2521 -121
rect 3219 -155 3253 -121
rect 1849 -281 1883 -247
rect -1955 -357 -1921 -323
rect -2211 -405 -2177 -371
rect -545 -395 -511 -361
rect -429 -395 -395 -361
rect -317 -395 -283 -361
rect -185 -395 -151 -361
rect -75 -395 -41 -361
rect 41 -395 75 -361
rect 177 -393 211 -359
rect 743 -357 777 -323
rect 2153 -395 2187 -361
rect 2269 -395 2303 -361
rect 2381 -395 2415 -361
rect 2513 -395 2547 -361
rect 2623 -395 2657 -361
rect 2739 -395 2773 -361
rect 2871 -393 2905 -359
rect 487 -447 521 -413
rect -851 -579 -817 -545
rect -2555 -699 -2521 -665
rect 3219 -699 3253 -665
rect 1847 -819 1881 -785
rect -2211 -951 -2177 -917
rect -1955 -1041 -1921 -1007
rect -545 -1003 -511 -969
rect -429 -1003 -395 -969
rect -317 -1003 -283 -969
rect -185 -1003 -151 -969
rect -75 -1003 -41 -969
rect 41 -1003 75 -969
rect 175 -1005 209 -971
rect 487 -991 521 -957
rect 743 -1041 777 -1007
rect 2153 -1003 2187 -969
rect 2269 -1003 2303 -969
rect 2381 -1003 2415 -969
rect 2513 -1003 2547 -969
rect 2623 -1003 2657 -969
rect 2739 -1003 2773 -969
rect 2871 -1005 2905 -971
rect -851 -1123 -817 -1089
rect -2555 -1243 -2521 -1209
rect 3219 -1243 3253 -1209
rect 1847 -1363 1881 -1329
rect -1955 -1445 -1921 -1411
rect -2211 -1495 -2177 -1461
rect -545 -1483 -511 -1449
rect -429 -1483 -395 -1449
rect -317 -1483 -283 -1449
rect -185 -1483 -151 -1449
rect -75 -1483 -41 -1449
rect 41 -1483 75 -1449
rect 173 -1481 207 -1447
rect 743 -1445 777 -1411
rect 2153 -1483 2187 -1449
rect 2269 -1483 2303 -1449
rect 2381 -1483 2415 -1449
rect 2513 -1483 2547 -1449
rect 2623 -1483 2657 -1449
rect 2739 -1483 2773 -1449
rect 2873 -1481 2907 -1447
rect 487 -1535 521 -1501
rect -851 -1667 -817 -1633
rect -2555 -1787 -2521 -1753
rect 3219 -1787 3253 -1753
rect 1847 -1907 1881 -1873
rect -2211 -2039 -2177 -2005
rect -1955 -2129 -1921 -2095
rect -545 -2091 -511 -2057
rect -429 -2091 -395 -2057
rect -317 -2091 -283 -2057
rect -185 -2091 -151 -2057
rect -75 -2091 -41 -2057
rect 41 -2091 75 -2057
rect 173 -2093 207 -2059
rect 487 -2081 521 -2047
rect 743 -2129 777 -2095
rect 2153 -2091 2187 -2057
rect 2269 -2091 2303 -2057
rect 2381 -2091 2415 -2057
rect 2513 -2091 2547 -2057
rect 2623 -2091 2657 -2057
rect 2739 -2091 2773 -2057
rect 2875 -2093 2909 -2059
rect -851 -2209 -817 -2175
rect -2555 -2331 -2521 -2297
rect 3219 -2331 3253 -2297
rect 1847 -2453 1881 -2419
rect -1955 -2533 -1921 -2499
rect -2211 -2581 -2177 -2547
rect -545 -2571 -511 -2537
rect -429 -2571 -395 -2537
rect -317 -2571 -283 -2537
rect -185 -2571 -151 -2537
rect -75 -2571 -41 -2537
rect 41 -2571 75 -2537
rect 175 -2569 209 -2535
rect 495 -2563 529 -2529
rect 743 -2533 777 -2499
rect 2153 -2571 2187 -2537
rect 2269 -2571 2303 -2537
rect 2381 -2571 2415 -2537
rect 2513 -2571 2547 -2537
rect 2623 -2571 2657 -2537
rect 2739 -2571 2773 -2537
rect 2871 -2569 2905 -2535
rect -851 -2753 -817 -2719
rect -2555 -2875 -2521 -2841
rect 3219 -2875 3253 -2841
<< metal1 >>
rect -2492 358 -2242 454
rect 242 432 3190 454
rect 242 380 314 432
rect 366 380 3190 432
rect 242 358 3190 380
rect -2674 139 -2154 152
rect -2674 105 -2207 139
rect -2173 105 -2154 139
rect -2674 92 -2154 105
rect -564 119 -376 132
rect -1968 94 -1908 100
rect -1974 90 -1902 94
rect -1974 38 -1964 90
rect -1912 38 -1902 90
rect -564 85 -545 119
rect -511 85 -429 119
rect -395 85 -376 119
rect -564 72 -376 85
rect -336 119 94 132
rect 160 130 220 136
rect -336 85 -317 119
rect -283 85 -185 119
rect -151 85 -75 119
rect -41 85 41 119
rect 75 85 94 119
rect -336 72 94 85
rect 154 126 226 130
rect 154 74 164 126
rect 216 74 226 126
rect 154 70 226 74
rect 160 64 220 70
rect -1974 34 -1902 38
rect -1968 28 -1908 34
rect -864 14 -804 20
rect -870 10 -798 14
rect -870 -42 -860 10
rect -808 -42 -798 10
rect -870 -46 -798 -42
rect -864 -52 -804 -46
rect -2584 -112 -2242 -90
rect -2584 -121 -2366 -112
rect -2584 -155 -2555 -121
rect -2521 -155 -2366 -121
rect -2584 -164 -2366 -155
rect -2314 -164 -2242 -112
rect -2584 -186 -2242 -164
rect 242 -186 456 -90
rect 2938 -112 3282 -90
rect 2938 -164 3012 -112
rect 3064 -121 3282 -112
rect 3064 -155 3219 -121
rect 3253 -155 3282 -121
rect 3064 -164 3282 -155
rect 2938 -186 3282 -164
rect 1836 -234 1896 -228
rect 1830 -238 1902 -234
rect 1830 -290 1840 -238
rect 1892 -290 1902 -238
rect 1830 -294 1902 -290
rect 1836 -300 1896 -294
rect -1968 -310 -1908 -304
rect 730 -310 790 -304
rect -1974 -314 -1902 -310
rect -2224 -358 -2164 -352
rect -2230 -362 -2158 -358
rect -2230 -414 -2220 -362
rect -2168 -414 -2158 -362
rect -1974 -366 -1964 -314
rect -1912 -366 -1902 -314
rect 724 -314 796 -310
rect -1974 -370 -1902 -366
rect -564 -361 -376 -348
rect -1968 -376 -1908 -370
rect -564 -395 -545 -361
rect -511 -395 -429 -361
rect -395 -395 -376 -361
rect -564 -408 -376 -395
rect -336 -361 94 -348
rect -336 -395 -317 -361
rect -283 -395 -185 -361
rect -151 -395 -75 -361
rect -41 -395 41 -361
rect 75 -395 94 -361
rect -336 -408 94 -395
rect 152 -350 230 -346
rect 152 -402 162 -350
rect 214 -402 230 -350
rect 724 -366 734 -314
rect 786 -366 796 -314
rect 2858 -346 2918 -340
rect 724 -370 796 -366
rect 2134 -361 2322 -348
rect 730 -376 790 -370
rect 474 -400 534 -394
rect 2134 -395 2153 -361
rect 2187 -395 2269 -361
rect 2303 -395 2322 -361
rect 152 -406 230 -402
rect 468 -404 540 -400
rect -2230 -418 -2158 -414
rect -2224 -424 -2164 -418
rect 468 -456 478 -404
rect 530 -456 540 -404
rect 2134 -408 2322 -395
rect 2362 -361 2792 -348
rect 2362 -395 2381 -361
rect 2415 -395 2513 -361
rect 2547 -395 2623 -361
rect 2657 -395 2739 -361
rect 2773 -395 2792 -361
rect 2362 -408 2792 -395
rect 2852 -350 2924 -346
rect 2852 -402 2862 -350
rect 2914 -402 2924 -350
rect 2852 -406 2924 -402
rect 2858 -412 2918 -406
rect 468 -460 540 -456
rect 474 -466 534 -460
rect -864 -532 -804 -526
rect -870 -536 -798 -532
rect -870 -588 -860 -536
rect -808 -588 -798 -536
rect -870 -592 -798 -588
rect -864 -598 -804 -592
rect -2584 -665 -2242 -634
rect -2584 -699 -2555 -665
rect -2521 -699 -2242 -665
rect -2584 -730 -2242 -699
rect 242 -656 456 -634
rect 242 -708 314 -656
rect 366 -708 456 -656
rect 242 -730 456 -708
rect 2936 -665 3282 -634
rect 2936 -699 3219 -665
rect 3253 -699 3282 -665
rect 2936 -730 3282 -699
rect 1834 -772 1894 -766
rect 1828 -776 1900 -772
rect 1828 -828 1838 -776
rect 1890 -828 1900 -776
rect 1828 -832 1900 -828
rect 1834 -838 1894 -832
rect -2224 -904 -2164 -898
rect -2230 -908 -2158 -904
rect -2230 -960 -2220 -908
rect -2168 -960 -2158 -908
rect 474 -944 534 -938
rect 468 -948 540 -944
rect -2230 -964 -2158 -960
rect -2224 -970 -2164 -964
rect -564 -969 -376 -956
rect -1968 -994 -1908 -988
rect -1974 -998 -1902 -994
rect -1974 -1050 -1964 -998
rect -1912 -1050 -1902 -998
rect -564 -1003 -545 -969
rect -511 -1003 -429 -969
rect -395 -1003 -376 -969
rect -564 -1016 -376 -1003
rect -336 -969 94 -956
rect 160 -958 220 -952
rect -336 -1003 -317 -969
rect -283 -1003 -185 -969
rect -151 -1003 -75 -969
rect -41 -1003 41 -969
rect 75 -1003 94 -969
rect -336 -1016 94 -1003
rect 154 -962 226 -958
rect 154 -1014 164 -962
rect 216 -1014 226 -962
rect 468 -1000 478 -948
rect 530 -1000 540 -948
rect 2134 -969 2322 -956
rect 730 -994 790 -988
rect 468 -1004 540 -1000
rect 724 -998 796 -994
rect 474 -1010 534 -1004
rect 154 -1018 226 -1014
rect 160 -1024 220 -1018
rect -1974 -1054 -1902 -1050
rect 724 -1050 734 -998
rect 786 -1050 796 -998
rect 2134 -1003 2153 -969
rect 2187 -1003 2269 -969
rect 2303 -1003 2322 -969
rect 2134 -1016 2322 -1003
rect 2362 -969 2792 -956
rect 2858 -958 2918 -952
rect 2362 -1003 2381 -969
rect 2415 -1003 2513 -969
rect 2547 -1003 2623 -969
rect 2657 -1003 2739 -969
rect 2773 -1003 2792 -969
rect 2362 -1016 2792 -1003
rect 2852 -962 2924 -958
rect 2852 -1014 2862 -962
rect 2914 -1014 2924 -962
rect 2852 -1018 2924 -1014
rect 2858 -1024 2918 -1018
rect 724 -1054 796 -1050
rect -1968 -1060 -1908 -1054
rect 730 -1060 790 -1054
rect -864 -1076 -804 -1070
rect -870 -1080 -798 -1076
rect -870 -1132 -860 -1080
rect -808 -1132 -798 -1080
rect -870 -1136 -798 -1132
rect -864 -1142 -804 -1136
rect -2584 -1200 -2224 -1178
rect -2584 -1209 -2366 -1200
rect -2584 -1243 -2555 -1209
rect -2521 -1243 -2366 -1209
rect -2584 -1252 -2366 -1243
rect -2314 -1252 -2224 -1200
rect -2584 -1274 -2224 -1252
rect 242 -1274 456 -1178
rect 2938 -1200 3282 -1178
rect 2938 -1252 3012 -1200
rect 3064 -1209 3282 -1200
rect 3064 -1243 3219 -1209
rect 3253 -1243 3282 -1209
rect 3064 -1252 3282 -1243
rect 2938 -1274 3282 -1252
rect 1834 -1316 1894 -1310
rect 1828 -1320 1900 -1316
rect 1828 -1372 1838 -1320
rect 1890 -1372 1900 -1320
rect 1828 -1376 1900 -1372
rect 1834 -1382 1894 -1376
rect -1968 -1398 -1908 -1392
rect 730 -1398 790 -1392
rect -1974 -1402 -1902 -1398
rect -2224 -1448 -2164 -1442
rect -2230 -1452 -2158 -1448
rect -2230 -1504 -2220 -1452
rect -2168 -1504 -2158 -1452
rect -1974 -1454 -1964 -1402
rect -1912 -1454 -1902 -1402
rect 724 -1402 796 -1398
rect 160 -1434 220 -1428
rect -1974 -1458 -1902 -1454
rect -564 -1449 -376 -1436
rect -1968 -1464 -1908 -1458
rect -564 -1483 -545 -1449
rect -511 -1483 -429 -1449
rect -395 -1483 -376 -1449
rect -564 -1496 -376 -1483
rect -336 -1449 94 -1436
rect -336 -1483 -317 -1449
rect -283 -1483 -185 -1449
rect -151 -1483 -75 -1449
rect -41 -1483 41 -1449
rect 75 -1483 94 -1449
rect -336 -1496 94 -1483
rect 154 -1438 226 -1434
rect 154 -1490 164 -1438
rect 216 -1490 226 -1438
rect 724 -1454 734 -1402
rect 786 -1454 796 -1402
rect 2858 -1434 2918 -1428
rect 724 -1458 796 -1454
rect 2134 -1449 2322 -1436
rect 730 -1464 790 -1458
rect 474 -1488 534 -1482
rect 2134 -1483 2153 -1449
rect 2187 -1483 2269 -1449
rect 2303 -1483 2322 -1449
rect 154 -1494 226 -1490
rect 468 -1492 540 -1488
rect 160 -1500 220 -1494
rect -2230 -1508 -2158 -1504
rect -2224 -1514 -2164 -1508
rect 468 -1544 478 -1492
rect 530 -1544 540 -1492
rect 2134 -1496 2322 -1483
rect 2362 -1449 2792 -1436
rect 2362 -1483 2381 -1449
rect 2415 -1483 2513 -1449
rect 2547 -1483 2623 -1449
rect 2657 -1483 2739 -1449
rect 2773 -1483 2792 -1449
rect 2362 -1496 2792 -1483
rect 2852 -1438 2924 -1434
rect 2852 -1490 2862 -1438
rect 2914 -1490 2924 -1438
rect 2852 -1494 2924 -1490
rect 2858 -1500 2918 -1494
rect 468 -1548 540 -1544
rect 474 -1554 534 -1548
rect -864 -1620 -804 -1614
rect -870 -1624 -798 -1620
rect -870 -1676 -860 -1624
rect -808 -1676 -798 -1624
rect -870 -1680 -798 -1676
rect -864 -1686 -804 -1680
rect -2584 -1753 -2242 -1722
rect -2584 -1787 -2555 -1753
rect -2521 -1787 -2242 -1753
rect -2584 -1818 -2242 -1787
rect 242 -1744 456 -1722
rect 242 -1796 314 -1744
rect 366 -1796 456 -1744
rect 242 -1818 456 -1796
rect 2936 -1753 3282 -1722
rect 2936 -1787 3219 -1753
rect 3253 -1787 3282 -1753
rect 2936 -1818 3282 -1787
rect 1834 -1860 1894 -1854
rect 1828 -1864 1900 -1860
rect 1828 -1916 1838 -1864
rect 1890 -1916 1900 -1864
rect 1828 -1920 1900 -1916
rect 1834 -1926 1894 -1920
rect -2224 -1992 -2164 -1986
rect -2230 -1996 -2158 -1992
rect -2230 -2048 -2220 -1996
rect -2168 -2048 -2158 -1996
rect 474 -2034 534 -2028
rect 468 -2038 540 -2034
rect -2230 -2052 -2158 -2048
rect -2224 -2058 -2164 -2052
rect -564 -2057 -376 -2044
rect -1968 -2082 -1908 -2076
rect -1974 -2086 -1902 -2082
rect -1974 -2138 -1964 -2086
rect -1912 -2138 -1902 -2086
rect -564 -2091 -545 -2057
rect -511 -2091 -429 -2057
rect -395 -2091 -376 -2057
rect -564 -2104 -376 -2091
rect -336 -2057 94 -2044
rect 160 -2046 220 -2040
rect -336 -2091 -317 -2057
rect -283 -2091 -185 -2057
rect -151 -2091 -75 -2057
rect -41 -2091 41 -2057
rect 75 -2091 94 -2057
rect -336 -2104 94 -2091
rect 154 -2050 226 -2046
rect 154 -2102 164 -2050
rect 216 -2102 226 -2050
rect 468 -2090 478 -2038
rect 530 -2090 540 -2038
rect 2134 -2057 2322 -2044
rect 730 -2082 790 -2076
rect 468 -2094 540 -2090
rect 724 -2086 796 -2082
rect 474 -2100 534 -2094
rect 154 -2106 226 -2102
rect 160 -2112 220 -2106
rect -1974 -2142 -1902 -2138
rect 724 -2138 734 -2086
rect 786 -2138 796 -2086
rect 2134 -2091 2153 -2057
rect 2187 -2091 2269 -2057
rect 2303 -2091 2322 -2057
rect 2134 -2104 2322 -2091
rect 2362 -2057 2792 -2044
rect 2362 -2091 2381 -2057
rect 2415 -2091 2513 -2057
rect 2547 -2091 2623 -2057
rect 2657 -2091 2739 -2057
rect 2773 -2091 2792 -2057
rect 2362 -2104 2792 -2091
rect 2850 -2050 2928 -2046
rect 2850 -2102 2860 -2050
rect 2912 -2102 2928 -2050
rect 2850 -2106 2928 -2102
rect 724 -2142 796 -2138
rect -1968 -2148 -1908 -2142
rect 730 -2148 790 -2142
rect -864 -2162 -804 -2156
rect -870 -2166 -798 -2162
rect -870 -2218 -860 -2166
rect -808 -2218 -798 -2166
rect -870 -2222 -798 -2218
rect -864 -2228 -804 -2222
rect -2584 -2288 -2224 -2266
rect -2584 -2297 -2366 -2288
rect -2584 -2331 -2555 -2297
rect -2521 -2331 -2366 -2297
rect -2584 -2340 -2366 -2331
rect -2314 -2340 -2224 -2288
rect -2584 -2362 -2224 -2340
rect 242 -2362 456 -2266
rect 2936 -2288 3282 -2266
rect 2936 -2340 3012 -2288
rect 3064 -2297 3282 -2288
rect 3064 -2331 3219 -2297
rect 3253 -2331 3282 -2297
rect 3064 -2340 3282 -2331
rect 2936 -2362 3282 -2340
rect 1834 -2406 1894 -2400
rect 1828 -2410 1900 -2406
rect 1828 -2462 1838 -2410
rect 1890 -2462 1900 -2410
rect 1828 -2466 1900 -2462
rect 1834 -2472 1894 -2466
rect -1968 -2486 -1908 -2480
rect 730 -2486 790 -2480
rect -1974 -2490 -1902 -2486
rect -2224 -2534 -2164 -2528
rect -2230 -2538 -2158 -2534
rect -2230 -2590 -2220 -2538
rect -2168 -2590 -2158 -2538
rect -1974 -2542 -1964 -2490
rect -1912 -2542 -1902 -2490
rect 724 -2490 796 -2486
rect 482 -2516 542 -2510
rect 160 -2522 220 -2516
rect 476 -2520 548 -2516
rect -1974 -2546 -1902 -2542
rect -564 -2537 -376 -2524
rect -1968 -2552 -1908 -2546
rect -564 -2571 -545 -2537
rect -511 -2571 -429 -2537
rect -395 -2571 -376 -2537
rect -564 -2584 -376 -2571
rect -336 -2537 94 -2524
rect -336 -2571 -317 -2537
rect -283 -2571 -185 -2537
rect -151 -2571 -75 -2537
rect -41 -2571 41 -2537
rect 75 -2571 94 -2537
rect -336 -2584 94 -2571
rect 154 -2526 226 -2522
rect 154 -2578 164 -2526
rect 216 -2578 226 -2526
rect 476 -2572 486 -2520
rect 538 -2572 548 -2520
rect 724 -2542 734 -2490
rect 786 -2542 796 -2490
rect 2858 -2522 2918 -2516
rect 724 -2546 796 -2542
rect 2134 -2537 2322 -2524
rect 730 -2552 790 -2546
rect 476 -2576 548 -2572
rect 2134 -2571 2153 -2537
rect 2187 -2571 2269 -2537
rect 2303 -2571 2322 -2537
rect 154 -2582 226 -2578
rect 482 -2582 542 -2576
rect 160 -2588 220 -2582
rect 2134 -2584 2322 -2571
rect 2362 -2537 2792 -2524
rect 2362 -2571 2381 -2537
rect 2415 -2571 2513 -2537
rect 2547 -2571 2623 -2537
rect 2657 -2571 2739 -2537
rect 2773 -2571 2792 -2537
rect 2362 -2584 2792 -2571
rect 2852 -2526 2924 -2522
rect 2852 -2578 2862 -2526
rect 2914 -2578 2924 -2526
rect 2852 -2582 2924 -2578
rect 2858 -2588 2918 -2582
rect -2230 -2594 -2158 -2590
rect -2224 -2600 -2164 -2594
rect -864 -2706 -804 -2700
rect -870 -2710 -798 -2706
rect -870 -2762 -860 -2710
rect -808 -2762 -798 -2710
rect -870 -2766 -798 -2762
rect -864 -2772 -804 -2766
rect -2584 -2841 -2242 -2810
rect -2584 -2875 -2555 -2841
rect -2521 -2875 -2242 -2841
rect -2584 -2906 -2242 -2875
rect 242 -2832 456 -2810
rect 242 -2884 314 -2832
rect 366 -2884 456 -2832
rect 242 -2906 456 -2884
rect 2936 -2841 3282 -2810
rect 2936 -2875 3219 -2841
rect 3253 -2875 3282 -2841
rect 2936 -2906 3282 -2875
<< via1 >>
rect 314 380 366 432
rect -1964 81 -1912 90
rect -1964 47 -1955 81
rect -1955 47 -1921 81
rect -1921 47 -1912 81
rect -1964 38 -1912 47
rect 164 117 216 126
rect 164 83 173 117
rect 173 83 207 117
rect 207 83 216 117
rect 164 74 216 83
rect -860 1 -808 10
rect -860 -33 -851 1
rect -851 -33 -817 1
rect -817 -33 -808 1
rect -860 -42 -808 -33
rect -2366 -164 -2314 -112
rect 3012 -164 3064 -112
rect 1840 -247 1892 -238
rect 1840 -281 1849 -247
rect 1849 -281 1883 -247
rect 1883 -281 1892 -247
rect 1840 -290 1892 -281
rect -2220 -371 -2168 -362
rect -2220 -405 -2211 -371
rect -2211 -405 -2177 -371
rect -2177 -405 -2168 -371
rect -2220 -414 -2168 -405
rect -1964 -323 -1912 -314
rect -1964 -357 -1955 -323
rect -1955 -357 -1921 -323
rect -1921 -357 -1912 -323
rect -1964 -366 -1912 -357
rect 162 -359 214 -350
rect 162 -393 177 -359
rect 177 -393 211 -359
rect 211 -393 214 -359
rect 162 -402 214 -393
rect 734 -323 786 -314
rect 734 -357 743 -323
rect 743 -357 777 -323
rect 777 -357 786 -323
rect 734 -366 786 -357
rect 478 -413 530 -404
rect 478 -447 487 -413
rect 487 -447 521 -413
rect 521 -447 530 -413
rect 478 -456 530 -447
rect 2862 -359 2914 -350
rect 2862 -393 2871 -359
rect 2871 -393 2905 -359
rect 2905 -393 2914 -359
rect 2862 -402 2914 -393
rect -860 -545 -808 -536
rect -860 -579 -851 -545
rect -851 -579 -817 -545
rect -817 -579 -808 -545
rect -860 -588 -808 -579
rect 314 -708 366 -656
rect 1838 -785 1890 -776
rect 1838 -819 1847 -785
rect 1847 -819 1881 -785
rect 1881 -819 1890 -785
rect 1838 -828 1890 -819
rect -2220 -917 -2168 -908
rect -2220 -951 -2211 -917
rect -2211 -951 -2177 -917
rect -2177 -951 -2168 -917
rect -2220 -960 -2168 -951
rect -1964 -1007 -1912 -998
rect -1964 -1041 -1955 -1007
rect -1955 -1041 -1921 -1007
rect -1921 -1041 -1912 -1007
rect -1964 -1050 -1912 -1041
rect 164 -971 216 -962
rect 164 -1005 175 -971
rect 175 -1005 209 -971
rect 209 -1005 216 -971
rect 164 -1014 216 -1005
rect 478 -957 530 -948
rect 478 -991 487 -957
rect 487 -991 521 -957
rect 521 -991 530 -957
rect 478 -1000 530 -991
rect 734 -1007 786 -998
rect 734 -1041 743 -1007
rect 743 -1041 777 -1007
rect 777 -1041 786 -1007
rect 734 -1050 786 -1041
rect 2862 -971 2914 -962
rect 2862 -1005 2871 -971
rect 2871 -1005 2905 -971
rect 2905 -1005 2914 -971
rect 2862 -1014 2914 -1005
rect -860 -1089 -808 -1080
rect -860 -1123 -851 -1089
rect -851 -1123 -817 -1089
rect -817 -1123 -808 -1089
rect -860 -1132 -808 -1123
rect -2366 -1252 -2314 -1200
rect 3012 -1252 3064 -1200
rect 1838 -1329 1890 -1320
rect 1838 -1363 1847 -1329
rect 1847 -1363 1881 -1329
rect 1881 -1363 1890 -1329
rect 1838 -1372 1890 -1363
rect -2220 -1461 -2168 -1452
rect -2220 -1495 -2211 -1461
rect -2211 -1495 -2177 -1461
rect -2177 -1495 -2168 -1461
rect -2220 -1504 -2168 -1495
rect -1964 -1411 -1912 -1402
rect -1964 -1445 -1955 -1411
rect -1955 -1445 -1921 -1411
rect -1921 -1445 -1912 -1411
rect -1964 -1454 -1912 -1445
rect 164 -1447 216 -1438
rect 164 -1481 173 -1447
rect 173 -1481 207 -1447
rect 207 -1481 216 -1447
rect 164 -1490 216 -1481
rect 734 -1411 786 -1402
rect 734 -1445 743 -1411
rect 743 -1445 777 -1411
rect 777 -1445 786 -1411
rect 734 -1454 786 -1445
rect 478 -1501 530 -1492
rect 478 -1535 487 -1501
rect 487 -1535 521 -1501
rect 521 -1535 530 -1501
rect 478 -1544 530 -1535
rect 2862 -1447 2914 -1438
rect 2862 -1481 2873 -1447
rect 2873 -1481 2907 -1447
rect 2907 -1481 2914 -1447
rect 2862 -1490 2914 -1481
rect -860 -1633 -808 -1624
rect -860 -1667 -851 -1633
rect -851 -1667 -817 -1633
rect -817 -1667 -808 -1633
rect -860 -1676 -808 -1667
rect 314 -1796 366 -1744
rect 1838 -1873 1890 -1864
rect 1838 -1907 1847 -1873
rect 1847 -1907 1881 -1873
rect 1881 -1907 1890 -1873
rect 1838 -1916 1890 -1907
rect -2220 -2005 -2168 -1996
rect -2220 -2039 -2211 -2005
rect -2211 -2039 -2177 -2005
rect -2177 -2039 -2168 -2005
rect -2220 -2048 -2168 -2039
rect -1964 -2095 -1912 -2086
rect -1964 -2129 -1955 -2095
rect -1955 -2129 -1921 -2095
rect -1921 -2129 -1912 -2095
rect -1964 -2138 -1912 -2129
rect 164 -2059 216 -2050
rect 164 -2093 173 -2059
rect 173 -2093 207 -2059
rect 207 -2093 216 -2059
rect 164 -2102 216 -2093
rect 478 -2047 530 -2038
rect 478 -2081 487 -2047
rect 487 -2081 521 -2047
rect 521 -2081 530 -2047
rect 478 -2090 530 -2081
rect 734 -2095 786 -2086
rect 734 -2129 743 -2095
rect 743 -2129 777 -2095
rect 777 -2129 786 -2095
rect 734 -2138 786 -2129
rect 2860 -2059 2912 -2050
rect 2860 -2093 2875 -2059
rect 2875 -2093 2909 -2059
rect 2909 -2093 2912 -2059
rect 2860 -2102 2912 -2093
rect -860 -2175 -808 -2166
rect -860 -2209 -851 -2175
rect -851 -2209 -817 -2175
rect -817 -2209 -808 -2175
rect -860 -2218 -808 -2209
rect -2366 -2340 -2314 -2288
rect 3012 -2340 3064 -2288
rect 1838 -2419 1890 -2410
rect 1838 -2453 1847 -2419
rect 1847 -2453 1881 -2419
rect 1881 -2453 1890 -2419
rect 1838 -2462 1890 -2453
rect -2220 -2547 -2168 -2538
rect -2220 -2581 -2211 -2547
rect -2211 -2581 -2177 -2547
rect -2177 -2581 -2168 -2547
rect -2220 -2590 -2168 -2581
rect -1964 -2499 -1912 -2490
rect -1964 -2533 -1955 -2499
rect -1955 -2533 -1921 -2499
rect -1921 -2533 -1912 -2499
rect -1964 -2542 -1912 -2533
rect 164 -2535 216 -2526
rect 164 -2569 175 -2535
rect 175 -2569 209 -2535
rect 209 -2569 216 -2535
rect 164 -2578 216 -2569
rect 486 -2529 538 -2520
rect 486 -2563 495 -2529
rect 495 -2563 529 -2529
rect 529 -2563 538 -2529
rect 486 -2572 538 -2563
rect 734 -2499 786 -2490
rect 734 -2533 743 -2499
rect 743 -2533 777 -2499
rect 777 -2533 786 -2499
rect 734 -2542 786 -2533
rect 2862 -2535 2914 -2526
rect 2862 -2569 2871 -2535
rect 2871 -2569 2905 -2535
rect 2905 -2569 2914 -2535
rect 2862 -2578 2914 -2569
rect -860 -2719 -808 -2710
rect -860 -2753 -851 -2719
rect -851 -2753 -817 -2719
rect -817 -2753 -808 -2719
rect -860 -2762 -808 -2753
rect 314 -2884 366 -2832
<< metal2 >>
rect 280 434 400 454
rect 280 378 312 434
rect 368 378 400 434
rect 280 358 400 378
rect -1968 126 226 130
rect -1968 90 164 126
rect -1968 38 -1964 90
rect -1912 74 164 90
rect 216 74 226 126
rect -1912 70 226 74
rect -1912 38 -1908 70
rect -1968 28 -1908 38
rect -864 10 -804 20
rect -864 -42 -860 10
rect -808 -42 -804 10
rect -2400 -110 -2280 -90
rect -864 -106 -804 -42
rect -2400 -166 -2368 -110
rect -2312 -166 -2280 -110
rect -2400 -186 -2280 -166
rect -2224 -166 -804 -106
rect -2224 -362 -2164 -166
rect 1836 -234 1896 104
rect 2978 -110 3098 -90
rect 2978 -166 3010 -110
rect 3066 -166 3098 -110
rect 2978 -186 3098 -166
rect 1830 -238 1902 -234
rect 1830 -290 1840 -238
rect 1892 -290 1902 -238
rect 1830 -294 1902 -290
rect -2224 -414 -2220 -362
rect -2168 -414 -2164 -362
rect -1968 -314 -1908 -304
rect -1968 -366 -1964 -314
rect -1912 -346 -1908 -314
rect 730 -314 790 -304
rect 158 -346 224 -340
rect -1912 -350 224 -346
rect -1912 -366 162 -350
rect -1968 -402 162 -366
rect 214 -402 224 -350
rect 730 -366 734 -314
rect 786 -346 790 -314
rect 786 -350 2924 -346
rect 786 -366 2862 -350
rect -1968 -406 224 -402
rect 158 -412 224 -406
rect 474 -404 534 -394
rect -2224 -424 -2164 -414
rect 474 -456 478 -404
rect 530 -456 534 -404
rect 730 -402 2862 -366
rect 2914 -402 2924 -350
rect 730 -406 2924 -402
rect -864 -536 -804 -526
rect -864 -588 -860 -536
rect -808 -588 -804 -536
rect -864 -652 -804 -588
rect -2224 -712 -804 -652
rect 280 -654 400 -634
rect 280 -710 312 -654
rect 368 -710 400 -654
rect -2224 -908 -2164 -712
rect 280 -730 400 -710
rect 474 -652 534 -456
rect 474 -712 1894 -652
rect 1834 -776 1894 -712
rect 1834 -828 1838 -776
rect 1890 -828 1894 -776
rect 1834 -838 1894 -828
rect -2224 -960 -2220 -908
rect -2168 -960 -2164 -908
rect 474 -948 534 -938
rect -2224 -970 -2164 -960
rect -1968 -962 226 -958
rect -1968 -998 164 -962
rect -1968 -1050 -1964 -998
rect -1912 -1014 164 -998
rect 216 -1014 226 -962
rect -1912 -1018 226 -1014
rect 474 -1000 478 -948
rect 530 -1000 534 -948
rect -1912 -1050 -1908 -1018
rect -1968 -1060 -1908 -1050
rect -864 -1080 -804 -1070
rect -864 -1132 -860 -1080
rect -808 -1132 -804 -1080
rect -2400 -1198 -2280 -1178
rect -864 -1196 -804 -1132
rect -2400 -1254 -2368 -1198
rect -2312 -1254 -2280 -1198
rect -2400 -1274 -2280 -1254
rect -2224 -1256 -804 -1196
rect 474 -1196 534 -1000
rect 730 -962 2924 -958
rect 730 -998 2862 -962
rect 730 -1050 734 -998
rect 786 -1014 2862 -998
rect 2914 -1014 2924 -962
rect 786 -1018 2924 -1014
rect 786 -1050 790 -1018
rect 730 -1060 790 -1050
rect 474 -1256 1894 -1196
rect -2224 -1452 -2164 -1256
rect 1834 -1320 1894 -1256
rect 2978 -1198 3098 -1178
rect 2978 -1254 3010 -1198
rect 3066 -1254 3098 -1198
rect 2978 -1274 3098 -1254
rect 1834 -1372 1838 -1320
rect 1890 -1372 1894 -1320
rect 1834 -1382 1894 -1372
rect -2224 -1504 -2220 -1452
rect -2168 -1504 -2164 -1452
rect -1968 -1402 -1908 -1392
rect -1968 -1454 -1964 -1402
rect -1912 -1434 -1908 -1402
rect 730 -1402 790 -1392
rect -1912 -1438 226 -1434
rect -1912 -1454 164 -1438
rect -1968 -1490 164 -1454
rect 216 -1490 226 -1438
rect 730 -1454 734 -1402
rect 786 -1434 790 -1402
rect 786 -1438 2924 -1434
rect 786 -1454 2862 -1438
rect -1968 -1494 226 -1490
rect 474 -1492 534 -1482
rect -2224 -1514 -2164 -1504
rect 474 -1544 478 -1492
rect 530 -1544 534 -1492
rect 730 -1490 2862 -1454
rect 2914 -1490 2924 -1438
rect 730 -1494 2924 -1490
rect -864 -1624 -804 -1614
rect -864 -1676 -860 -1624
rect -808 -1676 -804 -1624
rect -864 -1740 -804 -1676
rect -2224 -1800 -804 -1740
rect 280 -1742 400 -1722
rect 280 -1798 312 -1742
rect 368 -1798 400 -1742
rect -2224 -1996 -2164 -1800
rect 280 -1818 400 -1798
rect 474 -1740 534 -1544
rect 474 -1800 1894 -1740
rect 1834 -1864 1894 -1800
rect 1834 -1916 1838 -1864
rect 1890 -1916 1894 -1864
rect 1834 -1926 1894 -1916
rect -2224 -2048 -2220 -1996
rect -2168 -2048 -2164 -1996
rect 474 -2038 534 -2028
rect -2224 -2058 -2164 -2048
rect -1968 -2050 226 -2046
rect -1968 -2086 164 -2050
rect -1968 -2138 -1964 -2086
rect -1912 -2102 164 -2086
rect 216 -2102 226 -2050
rect -1912 -2106 226 -2102
rect 474 -2090 478 -2038
rect 530 -2090 534 -2038
rect 2856 -2046 2922 -2040
rect -1912 -2138 -1908 -2106
rect -1968 -2148 -1908 -2138
rect -864 -2166 -804 -2156
rect -864 -2218 -860 -2166
rect -808 -2218 -804 -2166
rect -2400 -2286 -2280 -2266
rect -864 -2282 -804 -2218
rect -2400 -2342 -2368 -2286
rect -2312 -2342 -2280 -2286
rect -2400 -2362 -2280 -2342
rect -2224 -2342 -804 -2282
rect 474 -2286 534 -2090
rect 730 -2050 2922 -2046
rect 730 -2086 2860 -2050
rect 730 -2138 734 -2086
rect 786 -2102 2860 -2086
rect 2912 -2102 2922 -2050
rect 786 -2106 2922 -2102
rect 786 -2138 790 -2106
rect 2856 -2112 2922 -2106
rect 730 -2148 790 -2138
rect 2978 -2286 3098 -2266
rect -2224 -2538 -2164 -2342
rect 474 -2346 1894 -2286
rect 1834 -2410 1894 -2346
rect 2978 -2342 3010 -2286
rect 3066 -2342 3098 -2286
rect 2978 -2362 3098 -2342
rect 1834 -2462 1838 -2410
rect 1890 -2462 1894 -2410
rect 1834 -2472 1894 -2462
rect -2224 -2590 -2220 -2538
rect -2168 -2590 -2164 -2538
rect -1968 -2490 -1908 -2480
rect -1968 -2542 -1964 -2490
rect -1912 -2522 -1908 -2490
rect 730 -2490 790 -2480
rect 482 -2516 542 -2510
rect 376 -2520 542 -2516
rect -1912 -2526 226 -2522
rect -1912 -2542 164 -2526
rect -1968 -2578 164 -2542
rect 216 -2578 226 -2526
rect -1968 -2582 226 -2578
rect 376 -2572 486 -2520
rect 538 -2572 542 -2520
rect 376 -2576 542 -2572
rect -2224 -2600 -2164 -2590
rect -864 -2706 -804 -2700
rect 376 -2706 436 -2576
rect 482 -2582 542 -2576
rect 730 -2542 734 -2490
rect 786 -2522 790 -2490
rect 786 -2526 2924 -2522
rect 786 -2542 2862 -2526
rect 730 -2578 2862 -2542
rect 2914 -2578 2924 -2526
rect 730 -2582 2924 -2578
rect -864 -2710 436 -2706
rect -864 -2762 -860 -2710
rect -808 -2762 436 -2710
rect -864 -2766 436 -2762
rect -864 -2772 -804 -2766
rect 280 -2830 400 -2810
rect 280 -2886 312 -2830
rect 368 -2886 400 -2830
rect 280 -2906 400 -2886
<< via2 >>
rect 312 432 368 434
rect 312 380 314 432
rect 314 380 366 432
rect 366 380 368 432
rect 312 378 368 380
rect -2368 -112 -2312 -110
rect -2368 -164 -2366 -112
rect -2366 -164 -2314 -112
rect -2314 -164 -2312 -112
rect -2368 -166 -2312 -164
rect 3010 -112 3066 -110
rect 3010 -164 3012 -112
rect 3012 -164 3064 -112
rect 3064 -164 3066 -112
rect 3010 -166 3066 -164
rect 312 -656 368 -654
rect 312 -708 314 -656
rect 314 -708 366 -656
rect 366 -708 368 -656
rect 312 -710 368 -708
rect -2368 -1200 -2312 -1198
rect -2368 -1252 -2366 -1200
rect -2366 -1252 -2314 -1200
rect -2314 -1252 -2312 -1200
rect -2368 -1254 -2312 -1252
rect 3010 -1200 3066 -1198
rect 3010 -1252 3012 -1200
rect 3012 -1252 3064 -1200
rect 3064 -1252 3066 -1200
rect 3010 -1254 3066 -1252
rect 312 -1744 368 -1742
rect 312 -1796 314 -1744
rect 314 -1796 366 -1744
rect 366 -1796 368 -1744
rect 312 -1798 368 -1796
rect -2368 -2288 -2312 -2286
rect -2368 -2340 -2366 -2288
rect -2366 -2340 -2314 -2288
rect -2314 -2340 -2312 -2288
rect -2368 -2342 -2312 -2340
rect 3010 -2288 3066 -2286
rect 3010 -2340 3012 -2288
rect 3012 -2340 3064 -2288
rect 3064 -2340 3066 -2288
rect 3010 -2342 3066 -2340
rect 312 -2832 368 -2830
rect 312 -2884 314 -2832
rect 314 -2884 366 -2832
rect 366 -2884 368 -2832
rect 312 -2886 368 -2884
<< metal3 >>
rect 280 438 400 454
rect 280 374 308 438
rect 372 374 400 438
rect 280 358 400 374
rect -2400 -106 -2280 -90
rect -2400 -170 -2372 -106
rect -2308 -170 -2280 -106
rect -2400 -186 -2280 -170
rect 2978 -106 3098 -90
rect 2978 -170 3006 -106
rect 3070 -170 3098 -106
rect 2978 -186 3098 -170
rect 280 -650 400 -634
rect 280 -714 308 -650
rect 372 -714 400 -650
rect 280 -730 400 -714
rect -2400 -1194 -2280 -1178
rect -2400 -1258 -2372 -1194
rect -2308 -1258 -2280 -1194
rect -2400 -1274 -2280 -1258
rect 2978 -1194 3098 -1178
rect 2978 -1258 3006 -1194
rect 3070 -1258 3098 -1194
rect 2978 -1274 3098 -1258
rect 280 -1738 400 -1722
rect 280 -1802 308 -1738
rect 372 -1802 400 -1738
rect 280 -1818 400 -1802
rect -2400 -2282 -2280 -2266
rect -2400 -2346 -2372 -2282
rect -2308 -2346 -2280 -2282
rect -2400 -2362 -2280 -2346
rect 2978 -2282 3098 -2266
rect 2978 -2346 3006 -2282
rect 3070 -2346 3098 -2282
rect 2978 -2362 3098 -2346
rect 280 -2826 400 -2810
rect 280 -2890 308 -2826
rect 372 -2890 400 -2826
rect 280 -2906 400 -2890
<< via3 >>
rect 308 434 372 438
rect 308 378 312 434
rect 312 378 368 434
rect 368 378 372 434
rect 308 374 372 378
rect -2372 -110 -2308 -106
rect -2372 -166 -2368 -110
rect -2368 -166 -2312 -110
rect -2312 -166 -2308 -110
rect -2372 -170 -2308 -166
rect 3006 -110 3070 -106
rect 3006 -166 3010 -110
rect 3010 -166 3066 -110
rect 3066 -166 3070 -110
rect 3006 -170 3070 -166
rect 308 -654 372 -650
rect 308 -710 312 -654
rect 312 -710 368 -654
rect 368 -710 372 -654
rect 308 -714 372 -710
rect -2372 -1198 -2308 -1194
rect -2372 -1254 -2368 -1198
rect -2368 -1254 -2312 -1198
rect -2312 -1254 -2308 -1198
rect -2372 -1258 -2308 -1254
rect 3006 -1198 3070 -1194
rect 3006 -1254 3010 -1198
rect 3010 -1254 3066 -1198
rect 3066 -1254 3070 -1198
rect 3006 -1258 3070 -1254
rect 308 -1742 372 -1738
rect 308 -1798 312 -1742
rect 312 -1798 368 -1742
rect 368 -1798 372 -1742
rect 308 -1802 372 -1798
rect -2372 -2286 -2308 -2282
rect -2372 -2342 -2368 -2286
rect -2368 -2342 -2312 -2286
rect -2312 -2342 -2308 -2286
rect -2372 -2346 -2308 -2342
rect 3006 -2286 3070 -2282
rect 3006 -2342 3010 -2286
rect 3010 -2342 3066 -2286
rect 3066 -2342 3070 -2286
rect 3006 -2346 3070 -2342
rect 308 -2830 372 -2826
rect 308 -2886 312 -2830
rect 312 -2886 368 -2830
rect 368 -2886 372 -2830
rect 308 -2890 372 -2886
<< metal4 >>
rect -2400 -106 -2280 454
rect -2400 -170 -2372 -106
rect -2308 -170 -2280 -106
rect -2400 -1194 -2280 -170
rect -2400 -1258 -2372 -1194
rect -2308 -1258 -2280 -1194
rect -2400 -2282 -2280 -1258
rect -2400 -2346 -2372 -2282
rect -2308 -2346 -2280 -2282
rect -2400 -2906 -2280 -2346
rect 280 438 400 454
rect 280 374 308 438
rect 372 374 400 438
rect 280 -650 400 374
rect 280 -714 308 -650
rect 372 -714 400 -650
rect 280 -1738 400 -714
rect 280 -1802 308 -1738
rect 372 -1802 400 -1738
rect 280 -2826 400 -1802
rect 280 -2890 308 -2826
rect 372 -2890 400 -2826
rect 280 -2906 400 -2890
rect 2978 -106 3098 454
rect 2978 -170 3006 -106
rect 3070 -170 3098 -106
rect 2978 -1194 3098 -170
rect 2978 -1258 3006 -1194
rect 3070 -1258 3098 -1194
rect 2978 -2282 3098 -1258
rect 2978 -2346 3006 -2282
rect 3070 -2346 3098 -2282
rect 2978 -2906 3098 -2346
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1626486988
transform 1 0 -2584 0 -1 -2314
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1626486988
transform 1 0 -2584 0 1 -2314
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_0
timestamp 1626486988
transform 1 0 -2242 0 -1 -2314
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_1
timestamp 1626486988
transform 1 0 -2242 0 1 -2314
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_1
timestamp 1626486988
transform 1 0 -218 0 -1 -2314
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0
timestamp 1626486988
transform 1 0 -218 0 1 -2314
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1626486988
transform 1 0 -494 0 1 -2314
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0
timestamp 1626486988
transform 1 0 -494 0 -1 -2314
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_2
timestamp 1626486988
transform 1 0 456 0 -1 -2314
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_3
timestamp 1626486988
transform 1 0 456 0 1 -2314
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_3
timestamp 1626486988
transform 1 0 2480 0 -1 -2314
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_2
timestamp 1626486988
transform 1 0 2480 0 1 -2314
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1626486988
transform 1 0 2204 0 1 -2314
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1626486988
transform 1 0 2204 0 -1 -2314
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1626486988
transform -1 0 3282 0 -1 -2314
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1626486988
transform -1 0 3282 0 1 -2314
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1626486988
transform 1 0 -2584 0 -1 -1226
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_4
timestamp 1626486988
transform 1 0 -2242 0 -1 -1226
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_4
timestamp 1626486988
transform 1 0 -218 0 -1 -1226
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4
timestamp 1626486988
transform 1 0 -494 0 -1 -1226
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_5
timestamp 1626486988
transform 1 0 456 0 -1 -1226
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_5
timestamp 1626486988
transform 1 0 2480 0 -1 -1226
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_5
timestamp 1626486988
transform 1 0 2204 0 -1 -1226
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1626486988
transform -1 0 3282 0 -1 -1226
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1626486988
transform 1 0 -2584 0 1 -1226
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_6
timestamp 1626486988
transform 1 0 -2242 0 1 -1226
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_6
timestamp 1626486988
transform 1 0 -218 0 1 -1226
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_6
timestamp 1626486988
transform 1 0 -494 0 1 -1226
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_7
timestamp 1626486988
transform 1 0 456 0 1 -1226
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_7
timestamp 1626486988
transform 1 0 2480 0 1 -1226
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_7
timestamp 1626486988
transform 1 0 2204 0 1 -1226
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1626486988
transform -1 0 3282 0 1 -1226
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1626486988
transform 1 0 -2584 0 -1 -138
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_8
timestamp 1626486988
transform 1 0 -2242 0 -1 -138
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_8
timestamp 1626486988
transform 1 0 -218 0 -1 -138
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_8
timestamp 1626486988
transform 1 0 -494 0 -1 -138
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_9
timestamp 1626486988
transform 1 0 456 0 -1 -138
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_9
timestamp 1626486988
transform 1 0 2480 0 -1 -138
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_9
timestamp 1626486988
transform 1 0 2204 0 -1 -138
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1626486988
transform -1 0 3282 0 -1 -138
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1626486988
transform 1 0 -2584 0 1 -138
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_10
timestamp 1626486988
transform 1 0 -2242 0 1 -138
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_10
timestamp 1626486988
transform 1 0 -218 0 1 -138
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_10
timestamp 1626486988
transform 1 0 -494 0 1 -138
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1626486988
transform -1 0 3282 0 1 -138
box -38 -48 130 592
<< labels >>
flabel metal1 s -2660 116 -2654 122 1 FreeSans 600 0 0 0 vin
flabel metal4 s -2348 -374 -2344 -370 1 FreeSans 600 0 0 0 VSS
flabel metal4 s 332 -378 342 -370 1 FreeSans 600 0 0 0 VDD
flabel metal2 s 1856 80 1866 88 1 FreeSans 600 0 0 0 vout
flabel metal1 s 3210 -1244 3261 -1206 0 FreeSans 250 180 0 0 VGND
port 1 nsew
flabel metal1 s 3210 -1246 3261 -1208 0 FreeSans 250 180 0 0 VGND
port 1 nsew
flabel metal1 s 3210 -2332 3261 -2294 0 FreeSans 250 180 0 0 VGND
port 1 nsew
flabel metal1 s 3210 -2334 3261 -2296 0 FreeSans 250 180 0 0 VGND
port 1 nsew
flabel metal1 s -2563 -2334 -2512 -2296 0 FreeSans 250 0 0 0 VGND
port 1 nsew
flabel metal1 s -2563 -2332 -2512 -2294 0 FreeSans 250 0 0 0 VGND
port 1 nsew
flabel metal1 s -2563 -1246 -2512 -1208 0 FreeSans 250 0 0 0 VGND
port 1 nsew
flabel metal1 s -2563 -1244 -2512 -1206 0 FreeSans 250 0 0 0 VGND
port 1 nsew
flabel metal1 s -2563 -158 -2512 -120 0 FreeSans 250 0 0 0 VGND
port 1 nsew
flabel metal1 s 3210 -158 3261 -120 0 FreeSans 250 180 0 0 VGND
port 1 nsew
flabel metal1 s -2562 -691 -2509 -662 0 FreeSans 250 0 0 0 VPWR
port 2 nsew
flabel metal1 s -2562 -702 -2509 -673 0 FreeSans 250 0 0 0 VPWR
port 2 nsew
flabel metal1 s -2562 -1779 -2509 -1750 0 FreeSans 250 0 0 0 VPWR
port 2 nsew
flabel metal1 s -2562 -1790 -2509 -1761 0 FreeSans 250 0 0 0 VPWR
port 2 nsew
flabel metal1 s -2562 -2867 -2509 -2838 0 FreeSans 250 0 0 0 VPWR
port 2 nsew
flabel metal1 s 3207 -2867 3260 -2838 0 FreeSans 250 180 0 0 VPWR
port 2 nsew
flabel metal1 s 3207 -1790 3260 -1761 0 FreeSans 250 180 0 0 VPWR
port 2 nsew
flabel metal1 s 3207 -1779 3260 -1750 0 FreeSans 250 180 0 0 VPWR
port 2 nsew
flabel metal1 s 3207 -702 3260 -673 0 FreeSans 250 180 0 0 VPWR
port 2 nsew
flabel metal1 s 3207 -691 3260 -662 0 FreeSans 250 180 0 0 VPWR
port 2 nsew
<< end >>
