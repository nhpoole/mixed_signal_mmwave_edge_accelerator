magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< metal3 >>
rect -1150 272 1149 300
rect -1150 -272 1065 272
rect 1129 -272 1149 272
rect -1150 -300 1149 -272
<< via3 >>
rect 1065 -272 1129 272
<< mimcap >>
rect -1050 160 950 200
rect -1050 -160 -1010 160
rect 910 -160 950 160
rect -1050 -200 950 -160
<< mimcapcontact >>
rect -1010 -160 910 160
<< metal4 >>
rect 1049 272 1145 288
rect -1011 160 911 161
rect -1011 -160 -1010 160
rect 910 -160 911 160
rect -1011 -161 911 -160
rect 1049 -272 1065 272
rect 1129 -272 1145 272
rect 1049 -288 1145 -272
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX -1150 -300 1050 300
string parameters w 10.00 l 2.00 val 44.56 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
