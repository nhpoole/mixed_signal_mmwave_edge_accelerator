magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -2210 -2160 2098 2160
<< metal3 >>
rect -950 -900 838 900
<< mimcap >>
rect -850 752 750 800
rect -850 -752 -802 752
rect 702 -752 750 752
rect -850 -800 750 -752
<< mimcapcontact >>
rect -802 -752 702 752
<< metal4 >>
rect -811 752 711 761
rect -811 -752 -802 752
rect 702 -752 711 752
rect -811 -761 711 -752
<< properties >>
string FIXED_BBOX -950 -900 850 900
<< end >>
