.lib ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt
.param vdsn=0.9 vgsn=0.6 vdp=0.9 vgp=1.2 vdd=1.8

.control
save all
save @m.xm2.msky130_fd_pr__nfet_01v8[gm] @m.xm3.msky130_fd_pr__nfet_01v8_lvt[gm] @m.xm6.msky130_fd_pr__nfet_03v3_nvt[gm]
save @m.xm2.msky130_fd_pr__nfet_01v8[vth] @m.xm3.msky130_fd_pr__nfet_01v8_lvt[vth] @m.xm6.msky130_fd_pr__nfet_03v3_nvt[vth]
save @m.xm2.msky130_fd_pr__nfet_01v8[id] @m.xm3.msky130_fd_pr__nfet_01v8_lvt[id] @m.xm6.msky130_fd_pr__nfet_03v3_nvt[id]
save @m.xm2.msky130_fd_pr__nfet_01v8[cgg] @m.xm3.msky130_fd_pr__nfet_01v8_lvt[cgg] @m.xm6.msky130_fd_pr__nfet_03v3_nvt[cgg]
save @m.xm1.msky130_fd_pr__pfet_01v8[gm] @m.xm4.msky130_fd_pr__pfet_01v8_lvt[gm] @m.xm5.msky130_fd_pr__pfet_01v8_hvt[gm]
save @m.xm1.msky130_fd_pr__pfet_01v8[vth] @m.xm4.msky130_fd_pr__pfet_01v8_lvt[vth] @m.xm5.msky130_fd_pr__pfet_01v8_hvt[vth]
save @m.xm1.msky130_fd_pr__pfet_01v8[id] @m.xm4.msky130_fd_pr__pfet_01v8_lvt[id] @m.xm5.msky130_fd_pr__pfet_01v8_hvt[id]
save @m.xm1.msky130_fd_pr__pfet_01v8[cgg] @m.xm4.msky130_fd_pr__pfet_01v8_lvt[cgg] @m.xm5.msky130_fd_pr__pfet_01v8_hvt[cgg]
op
dc vgsn 0.2 1.8 0.05
run
write char_nmos.raw
dc vgp 0 1.6 0.05
run
write char_pmos.raw
* print all
quit
.endc