magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -1260 -1260 108530 70542
<< locali >>
rect 95030 61087 95193 61121
rect 11993 60847 12156 60881
rect 95030 60847 95193 60881
rect 11993 60297 12156 60331
rect 95030 60297 95193 60331
rect 11993 60057 12156 60091
rect 95030 60057 95193 60091
rect 11993 59507 12156 59541
rect 95030 59507 95193 59541
rect 11993 59267 12156 59301
rect 95030 59267 95193 59301
rect 11993 58717 12156 58751
rect 95030 58717 95193 58751
rect 11993 58477 12156 58511
rect 95030 58477 95193 58511
rect 11993 57927 12156 57961
rect 95030 57927 95193 57961
rect 11993 57687 12156 57721
rect 95030 57687 95193 57721
rect 11993 57137 12156 57171
rect 95030 57137 95193 57171
rect 11993 56897 12156 56931
rect 95030 56897 95193 56931
rect 11993 56347 12156 56381
rect 95030 56347 95193 56381
rect 11993 56107 12156 56141
rect 95030 56107 95193 56141
rect 11993 55557 12156 55591
rect 95030 55557 95193 55591
rect 11993 55317 12156 55351
rect 95030 55317 95193 55351
rect 11993 54767 12156 54801
rect 95030 54767 95193 54801
rect 11993 54527 12156 54561
rect 95030 54527 95193 54561
rect 11993 53977 12156 54011
rect 95030 53977 95193 54011
rect 11993 53737 12156 53771
rect 95030 53737 95193 53771
rect 11993 53187 12156 53221
rect 95030 53187 95193 53221
rect 11993 52947 12156 52981
rect 95030 52947 95193 52981
rect 11993 52397 12156 52431
rect 95030 52397 95193 52431
rect 11993 52157 12156 52191
rect 95030 52157 95193 52191
rect 11993 51607 12156 51641
rect 95030 51607 95193 51641
rect 11993 51367 12156 51401
rect 95030 51367 95193 51401
rect 11993 50817 12156 50851
rect 95030 50817 95193 50851
rect 11993 50577 12156 50611
rect 95030 50577 95193 50611
rect 11993 50027 12156 50061
rect 95030 50027 95193 50061
rect 11993 49787 12156 49821
rect 95030 49787 95193 49821
rect 11993 49237 12156 49271
rect 95030 49237 95193 49271
rect 11993 48997 12156 49031
rect 95030 48997 95193 49031
rect 11993 48447 12156 48481
rect 95030 48447 95193 48481
rect 11993 48207 12156 48241
rect 95030 48207 95193 48241
rect 11993 47657 12156 47691
rect 95030 47657 95193 47691
rect 11993 47417 12156 47451
rect 95030 47417 95193 47451
rect 11993 46867 12156 46901
rect 95030 46867 95193 46901
rect 11993 46627 12156 46661
rect 95030 46627 95193 46661
rect 11993 46077 12156 46111
rect 95030 46077 95193 46111
rect 11993 45837 12156 45871
rect 95030 45837 95193 45871
rect 11993 45287 12156 45321
rect 95030 45287 95193 45321
rect 11993 45047 12156 45081
rect 95030 45047 95193 45081
rect 11993 44497 12156 44531
rect 95030 44497 95193 44531
rect 11993 44257 12156 44291
rect 95030 44257 95193 44291
rect 11993 43707 12156 43741
rect 95030 43707 95193 43741
rect 11993 43467 12156 43501
rect 95030 43467 95193 43501
rect 11993 42917 12156 42951
rect 95030 42917 95193 42951
rect 11993 42677 12156 42711
rect 95030 42677 95193 42711
rect 11993 42127 12156 42161
rect 95030 42127 95193 42161
rect 11993 41887 12156 41921
rect 95030 41887 95193 41921
rect 11993 41337 12156 41371
rect 95030 41337 95193 41371
rect 11993 41097 12156 41131
rect 95030 41097 95193 41131
rect 11993 40547 12156 40581
rect 95030 40547 95193 40581
rect 11993 40307 12156 40341
rect 95030 40307 95193 40341
rect 11993 39757 12156 39791
rect 95030 39757 95193 39791
rect 11993 39517 12156 39551
rect 95030 39517 95193 39551
rect 11993 38967 12156 39001
rect 95030 38967 95193 39001
rect 11993 38727 12156 38761
rect 95030 38727 95193 38761
rect 11993 38177 12156 38211
rect 95030 38177 95193 38211
rect 11993 37937 12156 37971
rect 95030 37937 95193 37971
rect 11993 37387 12156 37421
rect 95030 37387 95193 37421
rect 11993 37147 12156 37181
rect 95030 37147 95193 37181
rect 11993 36597 12156 36631
rect 95030 36597 95193 36631
rect 11993 36357 12156 36391
rect 95030 36357 95193 36391
rect 11993 35807 12156 35841
rect 95030 35807 95193 35841
rect 11993 35567 12156 35601
rect 95030 35567 95193 35601
rect 11993 35017 12156 35051
rect 95030 35017 95193 35051
rect 11993 34777 12156 34811
rect 95030 34777 95193 34811
rect 11993 34227 12156 34261
rect 95030 34227 95193 34261
rect 11993 33987 12156 34021
rect 95030 33987 95193 34021
rect 11993 33437 12156 33471
rect 95030 33437 95193 33471
rect 11993 33197 12156 33231
rect 95030 33197 95193 33231
rect 11993 32647 12156 32681
rect 95030 32647 95193 32681
rect 11993 32407 12156 32441
rect 95030 32407 95193 32441
rect 11993 31857 12156 31891
rect 95030 31857 95193 31891
rect 11993 31617 12156 31651
rect 95030 31617 95193 31651
rect 11993 31067 12156 31101
rect 95030 31067 95193 31101
rect 11993 30827 12156 30861
rect 95030 30827 95193 30861
rect 11993 30277 12156 30311
rect 95030 30277 95193 30311
rect 11993 30037 12156 30071
rect 95030 30037 95193 30071
rect 11993 29487 12156 29521
rect 95030 29487 95193 29521
rect 11993 29247 12156 29281
rect 95030 29247 95193 29281
rect 11993 28697 12156 28731
rect 95030 28697 95193 28731
rect 11993 28457 12156 28491
rect 95030 28457 95193 28491
rect 11993 27907 12156 27941
rect 95030 27907 95193 27941
rect 11993 27667 12156 27701
rect 95030 27667 95193 27701
rect 11993 27117 12156 27151
rect 95030 27117 95193 27151
rect 11993 26877 12156 26911
rect 95030 26877 95193 26911
rect 11993 26327 12156 26361
rect 95030 26327 95193 26361
rect 11993 26087 12156 26121
rect 95030 26087 95193 26121
rect 11993 25537 12156 25571
rect 95030 25537 95193 25571
rect 11993 25297 12156 25331
rect 95030 25297 95193 25331
rect 11993 24747 12156 24781
rect 95030 24747 95193 24781
rect 11993 24507 12156 24541
rect 95030 24507 95193 24541
rect 11993 23957 12156 23991
rect 95030 23957 95193 23991
rect 11993 23717 12156 23751
rect 95030 23717 95193 23751
rect 11993 23167 12156 23201
rect 95030 23167 95193 23201
rect 11993 22927 12156 22961
rect 95030 22927 95193 22961
rect 11993 22377 12156 22411
rect 95030 22377 95193 22411
rect 11993 22137 12156 22171
rect 95030 22137 95193 22171
rect 11993 21587 12156 21621
rect 95030 21587 95193 21621
rect 11993 21347 12156 21381
rect 95030 21347 95193 21381
rect 11993 20797 12156 20831
rect 95030 20797 95193 20831
rect 11993 20557 12156 20591
rect 95030 20557 95193 20591
rect 11993 20007 12156 20041
rect 95030 20007 95193 20041
rect 11993 19767 12156 19801
rect 95030 19767 95193 19801
rect 11993 19217 12156 19251
rect 95030 19217 95193 19251
rect 11993 18977 12156 19011
rect 95030 18977 95193 19011
rect 11993 18427 12156 18461
rect 95030 18427 95193 18461
rect 11993 18187 12156 18221
rect 95030 18187 95193 18221
rect 11993 17637 12156 17671
rect 95030 17637 95193 17671
rect 11993 17397 12156 17431
rect 95030 17397 95193 17431
rect 11993 16847 12156 16881
rect 95030 16847 95193 16881
rect 11993 16607 12156 16641
rect 95030 16607 95193 16641
rect 11993 16057 12156 16091
rect 95030 16057 95193 16091
rect 11993 15817 12156 15851
rect 95030 15817 95193 15851
rect 11993 15267 12156 15301
rect 95030 15267 95193 15301
rect 11993 15027 12156 15061
rect 95030 15027 95193 15061
rect 11993 14477 12156 14511
rect 95030 14477 95193 14511
rect 11993 14237 12156 14271
rect 95030 14237 95193 14271
rect 11993 13687 12156 13721
rect 95030 13687 95193 13721
rect 11993 13447 12156 13481
rect 95030 13447 95193 13481
rect 11993 12897 12156 12931
rect 95030 12897 95193 12931
rect 11993 12657 12156 12691
rect 95030 12657 95193 12691
rect 11993 12107 12156 12141
rect 95030 12107 95193 12141
rect 11993 11867 12156 11901
rect 95030 11867 95193 11901
rect 11993 11317 12156 11351
rect 95030 11317 95193 11351
rect 11993 11077 12156 11111
rect 95030 11077 95193 11111
rect 11993 10527 12156 10561
rect 95030 10527 95193 10561
rect 11993 10287 12156 10321
<< metal1 >>
rect 99828 68503 99892 68555
rect 101898 68500 101944 68558
rect 13761 67470 13807 67724
rect 16257 67470 16303 67724
rect 18753 67470 18799 67724
rect 21249 67470 21295 67724
rect 23745 67470 23791 67724
rect 26241 67470 26287 67724
rect 28737 67470 28783 67724
rect 31233 67470 31279 67724
rect 33729 67470 33775 67724
rect 36225 67470 36271 67724
rect 38721 67470 38767 67724
rect 41217 67470 41263 67724
rect 43713 67470 43759 67724
rect 46209 67470 46255 67724
rect 48705 67470 48751 67724
rect 51201 67470 51247 67724
rect 53697 67470 53743 67724
rect 56193 67470 56239 67724
rect 58689 67470 58735 67724
rect 61185 67470 61231 67724
rect 63681 67470 63727 67724
rect 66177 67470 66223 67724
rect 68673 67470 68719 67724
rect 71169 67470 71215 67724
rect 73665 67470 73711 67724
rect 76161 67470 76207 67724
rect 78657 67470 78703 67724
rect 81153 67470 81199 67724
rect 83649 67470 83695 67724
rect 86145 67470 86191 67724
rect 88641 67470 88687 67724
rect 91137 67470 91183 67724
rect 99828 67013 99892 67065
rect 101774 67010 101820 67068
rect 99828 65675 99892 65727
rect 99828 64185 99892 64237
rect 93595 62780 93623 62904
rect 13723 61914 13751 62026
rect 14187 61914 14215 62026
rect 13723 61886 13983 61914
rect 13955 61774 13983 61886
rect 14027 61886 14215 61914
rect 14347 61914 14375 62026
rect 14811 61914 14839 62026
rect 14347 61886 14535 61914
rect 14027 61774 14055 61886
rect 14507 61774 14535 61886
rect 14579 61886 14839 61914
rect 14971 61914 14999 62026
rect 15435 61914 15463 62026
rect 14971 61886 15231 61914
rect 14579 61774 14607 61886
rect 15203 61774 15231 61886
rect 15275 61886 15463 61914
rect 15595 61914 15623 62026
rect 16059 61914 16087 62026
rect 15595 61886 15783 61914
rect 15275 61774 15303 61886
rect 15755 61774 15783 61886
rect 15827 61886 16087 61914
rect 16219 61914 16247 62026
rect 16683 61914 16711 62026
rect 16219 61886 16479 61914
rect 15827 61774 15855 61886
rect 16451 61774 16479 61886
rect 16523 61886 16711 61914
rect 16843 61914 16871 62026
rect 17307 61914 17335 62026
rect 16843 61886 17031 61914
rect 16523 61774 16551 61886
rect 17003 61774 17031 61886
rect 17075 61886 17335 61914
rect 17467 61914 17495 62026
rect 17931 61914 17959 62026
rect 17467 61886 17727 61914
rect 17075 61774 17103 61886
rect 17699 61774 17727 61886
rect 17771 61886 17959 61914
rect 18091 61914 18119 62026
rect 18555 61914 18583 62026
rect 18091 61886 18279 61914
rect 17771 61774 17799 61886
rect 18251 61774 18279 61886
rect 18323 61886 18583 61914
rect 18715 61914 18743 62026
rect 19179 61914 19207 62026
rect 18715 61886 18975 61914
rect 18323 61774 18351 61886
rect 18947 61774 18975 61886
rect 19019 61886 19207 61914
rect 19339 61914 19367 62026
rect 19803 61914 19831 62026
rect 19339 61886 19527 61914
rect 19019 61774 19047 61886
rect 19499 61774 19527 61886
rect 19571 61886 19831 61914
rect 19963 61914 19991 62026
rect 20427 61914 20455 62026
rect 19963 61886 20223 61914
rect 19571 61774 19599 61886
rect 20195 61774 20223 61886
rect 20267 61886 20455 61914
rect 20587 61914 20615 62026
rect 21051 61914 21079 62026
rect 20587 61886 20775 61914
rect 20267 61774 20295 61886
rect 20747 61774 20775 61886
rect 20819 61886 21079 61914
rect 21211 61914 21239 62026
rect 21675 61914 21703 62026
rect 21211 61886 21471 61914
rect 20819 61774 20847 61886
rect 21443 61774 21471 61886
rect 21515 61886 21703 61914
rect 21835 61914 21863 62026
rect 22299 61914 22327 62026
rect 21835 61886 22023 61914
rect 21515 61774 21543 61886
rect 21995 61774 22023 61886
rect 22067 61886 22327 61914
rect 22459 61914 22487 62026
rect 22923 61914 22951 62026
rect 22459 61886 22719 61914
rect 22067 61774 22095 61886
rect 22691 61774 22719 61886
rect 22763 61886 22951 61914
rect 23083 61914 23111 62026
rect 23547 61914 23575 62026
rect 23083 61886 23271 61914
rect 22763 61774 22791 61886
rect 23243 61774 23271 61886
rect 23315 61886 23575 61914
rect 23707 61914 23735 62026
rect 24171 61914 24199 62026
rect 23707 61886 23967 61914
rect 23315 61774 23343 61886
rect 23939 61774 23967 61886
rect 24011 61886 24199 61914
rect 24331 61914 24359 62026
rect 24795 61914 24823 62026
rect 24331 61886 24519 61914
rect 24011 61774 24039 61886
rect 24491 61774 24519 61886
rect 24563 61886 24823 61914
rect 24955 61914 24983 62026
rect 25419 61914 25447 62026
rect 24955 61886 25215 61914
rect 24563 61774 24591 61886
rect 25187 61774 25215 61886
rect 25259 61886 25447 61914
rect 25579 61914 25607 62026
rect 26043 61914 26071 62026
rect 25579 61886 25767 61914
rect 25259 61774 25287 61886
rect 25739 61774 25767 61886
rect 25811 61886 26071 61914
rect 26203 61914 26231 62026
rect 26667 61914 26695 62026
rect 26203 61886 26463 61914
rect 25811 61774 25839 61886
rect 26435 61774 26463 61886
rect 26507 61886 26695 61914
rect 26827 61914 26855 62026
rect 27291 61914 27319 62026
rect 26827 61886 27015 61914
rect 26507 61774 26535 61886
rect 26987 61774 27015 61886
rect 27059 61886 27319 61914
rect 27451 61914 27479 62026
rect 27915 61914 27943 62026
rect 27451 61886 27711 61914
rect 27059 61774 27087 61886
rect 27683 61774 27711 61886
rect 27755 61886 27943 61914
rect 28075 61914 28103 62026
rect 28539 61914 28567 62026
rect 28075 61886 28263 61914
rect 27755 61774 27783 61886
rect 28235 61774 28263 61886
rect 28307 61886 28567 61914
rect 28699 61914 28727 62026
rect 29163 61914 29191 62026
rect 28699 61886 28959 61914
rect 28307 61774 28335 61886
rect 28931 61774 28959 61886
rect 29003 61886 29191 61914
rect 29323 61914 29351 62026
rect 29787 61914 29815 62026
rect 29323 61886 29511 61914
rect 29003 61774 29031 61886
rect 29483 61774 29511 61886
rect 29555 61886 29815 61914
rect 29947 61914 29975 62026
rect 30411 61914 30439 62026
rect 29947 61886 30207 61914
rect 29555 61774 29583 61886
rect 30179 61774 30207 61886
rect 30251 61886 30439 61914
rect 30571 61914 30599 62026
rect 31035 61914 31063 62026
rect 30571 61886 30759 61914
rect 30251 61774 30279 61886
rect 30731 61774 30759 61886
rect 30803 61886 31063 61914
rect 31195 61914 31223 62026
rect 31659 61914 31687 62026
rect 31195 61886 31455 61914
rect 30803 61774 30831 61886
rect 31427 61774 31455 61886
rect 31499 61886 31687 61914
rect 31819 61914 31847 62026
rect 32283 61914 32311 62026
rect 31819 61886 32007 61914
rect 31499 61774 31527 61886
rect 31979 61774 32007 61886
rect 32051 61886 32311 61914
rect 32443 61914 32471 62026
rect 32907 61914 32935 62026
rect 32443 61886 32703 61914
rect 32051 61774 32079 61886
rect 32675 61774 32703 61886
rect 32747 61886 32935 61914
rect 33067 61914 33095 62026
rect 33531 61914 33559 62026
rect 33067 61886 33255 61914
rect 32747 61774 32775 61886
rect 33227 61774 33255 61886
rect 33299 61886 33559 61914
rect 33691 61914 33719 62026
rect 34155 61914 34183 62026
rect 33691 61886 33951 61914
rect 33299 61774 33327 61886
rect 33923 61774 33951 61886
rect 33995 61886 34183 61914
rect 34315 61914 34343 62026
rect 34779 61914 34807 62026
rect 34315 61886 34503 61914
rect 33995 61774 34023 61886
rect 34475 61774 34503 61886
rect 34547 61886 34807 61914
rect 34939 61914 34967 62026
rect 35403 61914 35431 62026
rect 34939 61886 35199 61914
rect 34547 61774 34575 61886
rect 35171 61774 35199 61886
rect 35243 61886 35431 61914
rect 35563 61914 35591 62026
rect 36027 61914 36055 62026
rect 35563 61886 35751 61914
rect 35243 61774 35271 61886
rect 35723 61774 35751 61886
rect 35795 61886 36055 61914
rect 36187 61914 36215 62026
rect 36651 61914 36679 62026
rect 36187 61886 36447 61914
rect 35795 61774 35823 61886
rect 36419 61774 36447 61886
rect 36491 61886 36679 61914
rect 36811 61914 36839 62026
rect 37275 61914 37303 62026
rect 36811 61886 36999 61914
rect 36491 61774 36519 61886
rect 36971 61774 36999 61886
rect 37043 61886 37303 61914
rect 37435 61914 37463 62026
rect 37899 61914 37927 62026
rect 37435 61886 37695 61914
rect 37043 61774 37071 61886
rect 37667 61774 37695 61886
rect 37739 61886 37927 61914
rect 38059 61914 38087 62026
rect 38523 61914 38551 62026
rect 38059 61886 38247 61914
rect 37739 61774 37767 61886
rect 38219 61774 38247 61886
rect 38291 61886 38551 61914
rect 38683 61914 38711 62026
rect 39147 61914 39175 62026
rect 38683 61886 38943 61914
rect 38291 61774 38319 61886
rect 38915 61774 38943 61886
rect 38987 61886 39175 61914
rect 39307 61914 39335 62026
rect 39771 61914 39799 62026
rect 39307 61886 39495 61914
rect 38987 61774 39015 61886
rect 39467 61774 39495 61886
rect 39539 61886 39799 61914
rect 39931 61914 39959 62026
rect 40395 61914 40423 62026
rect 39931 61886 40191 61914
rect 39539 61774 39567 61886
rect 40163 61774 40191 61886
rect 40235 61886 40423 61914
rect 40555 61914 40583 62026
rect 41019 61914 41047 62026
rect 40555 61886 40743 61914
rect 40235 61774 40263 61886
rect 40715 61774 40743 61886
rect 40787 61886 41047 61914
rect 41179 61914 41207 62026
rect 41643 61914 41671 62026
rect 41179 61886 41439 61914
rect 40787 61774 40815 61886
rect 41411 61774 41439 61886
rect 41483 61886 41671 61914
rect 41803 61914 41831 62026
rect 42267 61914 42295 62026
rect 41803 61886 41991 61914
rect 41483 61774 41511 61886
rect 41963 61774 41991 61886
rect 42035 61886 42295 61914
rect 42427 61914 42455 62026
rect 42891 61914 42919 62026
rect 42427 61886 42687 61914
rect 42035 61774 42063 61886
rect 42659 61774 42687 61886
rect 42731 61886 42919 61914
rect 43051 61914 43079 62026
rect 43515 61914 43543 62026
rect 43051 61886 43239 61914
rect 42731 61774 42759 61886
rect 43211 61774 43239 61886
rect 43283 61886 43543 61914
rect 43675 61914 43703 62026
rect 44139 61914 44167 62026
rect 43675 61886 43935 61914
rect 43283 61774 43311 61886
rect 43907 61774 43935 61886
rect 43979 61886 44167 61914
rect 44299 61914 44327 62026
rect 44763 61914 44791 62026
rect 44299 61886 44487 61914
rect 43979 61774 44007 61886
rect 44459 61774 44487 61886
rect 44531 61886 44791 61914
rect 44923 61914 44951 62026
rect 45387 61914 45415 62026
rect 44923 61886 45183 61914
rect 44531 61774 44559 61886
rect 45155 61774 45183 61886
rect 45227 61886 45415 61914
rect 45547 61914 45575 62026
rect 46011 61914 46039 62026
rect 45547 61886 45735 61914
rect 45227 61774 45255 61886
rect 45707 61774 45735 61886
rect 45779 61886 46039 61914
rect 46171 61914 46199 62026
rect 46635 61914 46663 62026
rect 46171 61886 46431 61914
rect 45779 61774 45807 61886
rect 46403 61774 46431 61886
rect 46475 61886 46663 61914
rect 46795 61914 46823 62026
rect 47259 61914 47287 62026
rect 46795 61886 46983 61914
rect 46475 61774 46503 61886
rect 46955 61774 46983 61886
rect 47027 61886 47287 61914
rect 47419 61914 47447 62026
rect 47883 61914 47911 62026
rect 47419 61886 47679 61914
rect 47027 61774 47055 61886
rect 47651 61774 47679 61886
rect 47723 61886 47911 61914
rect 48043 61914 48071 62026
rect 48507 61914 48535 62026
rect 48043 61886 48231 61914
rect 47723 61774 47751 61886
rect 48203 61774 48231 61886
rect 48275 61886 48535 61914
rect 48667 61914 48695 62026
rect 49131 61914 49159 62026
rect 48667 61886 48927 61914
rect 48275 61774 48303 61886
rect 48899 61774 48927 61886
rect 48971 61886 49159 61914
rect 49291 61914 49319 62026
rect 49755 61914 49783 62026
rect 49291 61886 49479 61914
rect 48971 61774 48999 61886
rect 49451 61774 49479 61886
rect 49523 61886 49783 61914
rect 49915 61914 49943 62026
rect 50379 61914 50407 62026
rect 49915 61886 50175 61914
rect 49523 61774 49551 61886
rect 50147 61774 50175 61886
rect 50219 61886 50407 61914
rect 50539 61914 50567 62026
rect 51003 61914 51031 62026
rect 50539 61886 50727 61914
rect 50219 61774 50247 61886
rect 50699 61774 50727 61886
rect 50771 61886 51031 61914
rect 51163 61914 51191 62026
rect 51627 61914 51655 62026
rect 51163 61886 51423 61914
rect 50771 61774 50799 61886
rect 51395 61774 51423 61886
rect 51467 61886 51655 61914
rect 51787 61914 51815 62026
rect 52251 61914 52279 62026
rect 51787 61886 51975 61914
rect 51467 61774 51495 61886
rect 51947 61774 51975 61886
rect 52019 61886 52279 61914
rect 52411 61914 52439 62026
rect 52875 61914 52903 62026
rect 52411 61886 52671 61914
rect 52019 61774 52047 61886
rect 52643 61774 52671 61886
rect 52715 61886 52903 61914
rect 53035 61914 53063 62026
rect 53499 61914 53527 62026
rect 53035 61886 53223 61914
rect 52715 61774 52743 61886
rect 53195 61774 53223 61886
rect 53267 61886 53527 61914
rect 53659 61914 53687 62026
rect 54123 61914 54151 62026
rect 53659 61886 53919 61914
rect 53267 61774 53295 61886
rect 53891 61774 53919 61886
rect 53963 61886 54151 61914
rect 54283 61914 54311 62026
rect 54747 61914 54775 62026
rect 54283 61886 54471 61914
rect 53963 61774 53991 61886
rect 54443 61774 54471 61886
rect 54515 61886 54775 61914
rect 54907 61914 54935 62026
rect 55371 61914 55399 62026
rect 54907 61886 55167 61914
rect 54515 61774 54543 61886
rect 55139 61774 55167 61886
rect 55211 61886 55399 61914
rect 55531 61914 55559 62026
rect 55995 61914 56023 62026
rect 55531 61886 55719 61914
rect 55211 61774 55239 61886
rect 55691 61774 55719 61886
rect 55763 61886 56023 61914
rect 56155 61914 56183 62026
rect 56619 61914 56647 62026
rect 56155 61886 56415 61914
rect 55763 61774 55791 61886
rect 56387 61774 56415 61886
rect 56459 61886 56647 61914
rect 56779 61914 56807 62026
rect 57243 61914 57271 62026
rect 56779 61886 56967 61914
rect 56459 61774 56487 61886
rect 56939 61774 56967 61886
rect 57011 61886 57271 61914
rect 57403 61914 57431 62026
rect 57867 61914 57895 62026
rect 57403 61886 57663 61914
rect 57011 61774 57039 61886
rect 57635 61774 57663 61886
rect 57707 61886 57895 61914
rect 58027 61914 58055 62026
rect 58491 61914 58519 62026
rect 58027 61886 58215 61914
rect 57707 61774 57735 61886
rect 58187 61774 58215 61886
rect 58259 61886 58519 61914
rect 58651 61914 58679 62026
rect 59115 61914 59143 62026
rect 58651 61886 58911 61914
rect 58259 61774 58287 61886
rect 58883 61774 58911 61886
rect 58955 61886 59143 61914
rect 59275 61914 59303 62026
rect 59739 61914 59767 62026
rect 59275 61886 59463 61914
rect 58955 61774 58983 61886
rect 59435 61774 59463 61886
rect 59507 61886 59767 61914
rect 59899 61914 59927 62026
rect 60363 61914 60391 62026
rect 59899 61886 60159 61914
rect 59507 61774 59535 61886
rect 60131 61774 60159 61886
rect 60203 61886 60391 61914
rect 60523 61914 60551 62026
rect 60987 61914 61015 62026
rect 60523 61886 60711 61914
rect 60203 61774 60231 61886
rect 60683 61774 60711 61886
rect 60755 61886 61015 61914
rect 61147 61914 61175 62026
rect 61611 61914 61639 62026
rect 61147 61886 61407 61914
rect 60755 61774 60783 61886
rect 61379 61774 61407 61886
rect 61451 61886 61639 61914
rect 61771 61914 61799 62026
rect 62235 61914 62263 62026
rect 61771 61886 61959 61914
rect 61451 61774 61479 61886
rect 61931 61774 61959 61886
rect 62003 61886 62263 61914
rect 62395 61914 62423 62026
rect 62859 61914 62887 62026
rect 62395 61886 62655 61914
rect 62003 61774 62031 61886
rect 62627 61774 62655 61886
rect 62699 61886 62887 61914
rect 63019 61914 63047 62026
rect 63483 61914 63511 62026
rect 63019 61886 63207 61914
rect 62699 61774 62727 61886
rect 63179 61774 63207 61886
rect 63251 61886 63511 61914
rect 63643 61914 63671 62026
rect 64107 61914 64135 62026
rect 63643 61886 63903 61914
rect 63251 61774 63279 61886
rect 63875 61774 63903 61886
rect 63947 61886 64135 61914
rect 64267 61914 64295 62026
rect 64731 61914 64759 62026
rect 64267 61886 64455 61914
rect 63947 61774 63975 61886
rect 64427 61774 64455 61886
rect 64499 61886 64759 61914
rect 64891 61914 64919 62026
rect 65355 61914 65383 62026
rect 64891 61886 65151 61914
rect 64499 61774 64527 61886
rect 65123 61774 65151 61886
rect 65195 61886 65383 61914
rect 65515 61914 65543 62026
rect 65979 61914 66007 62026
rect 65515 61886 65703 61914
rect 65195 61774 65223 61886
rect 65675 61774 65703 61886
rect 65747 61886 66007 61914
rect 66139 61914 66167 62026
rect 66603 61914 66631 62026
rect 66139 61886 66399 61914
rect 65747 61774 65775 61886
rect 66371 61774 66399 61886
rect 66443 61886 66631 61914
rect 66763 61914 66791 62026
rect 67227 61914 67255 62026
rect 66763 61886 66951 61914
rect 66443 61774 66471 61886
rect 66923 61774 66951 61886
rect 66995 61886 67255 61914
rect 67387 61914 67415 62026
rect 67851 61914 67879 62026
rect 67387 61886 67647 61914
rect 66995 61774 67023 61886
rect 67619 61774 67647 61886
rect 67691 61886 67879 61914
rect 68011 61914 68039 62026
rect 68475 61914 68503 62026
rect 68011 61886 68199 61914
rect 67691 61774 67719 61886
rect 68171 61774 68199 61886
rect 68243 61886 68503 61914
rect 68635 61914 68663 62026
rect 69099 61914 69127 62026
rect 68635 61886 68895 61914
rect 68243 61774 68271 61886
rect 68867 61774 68895 61886
rect 68939 61886 69127 61914
rect 69259 61914 69287 62026
rect 69723 61914 69751 62026
rect 69259 61886 69447 61914
rect 68939 61774 68967 61886
rect 69419 61774 69447 61886
rect 69491 61886 69751 61914
rect 69883 61914 69911 62026
rect 70347 61914 70375 62026
rect 69883 61886 70143 61914
rect 69491 61774 69519 61886
rect 70115 61774 70143 61886
rect 70187 61886 70375 61914
rect 70507 61914 70535 62026
rect 70971 61914 70999 62026
rect 70507 61886 70695 61914
rect 70187 61774 70215 61886
rect 70667 61774 70695 61886
rect 70739 61886 70999 61914
rect 71131 61914 71159 62026
rect 71595 61914 71623 62026
rect 71131 61886 71391 61914
rect 70739 61774 70767 61886
rect 71363 61774 71391 61886
rect 71435 61886 71623 61914
rect 71755 61914 71783 62026
rect 72219 61914 72247 62026
rect 71755 61886 71943 61914
rect 71435 61774 71463 61886
rect 71915 61774 71943 61886
rect 71987 61886 72247 61914
rect 72379 61914 72407 62026
rect 72843 61914 72871 62026
rect 72379 61886 72639 61914
rect 71987 61774 72015 61886
rect 72611 61774 72639 61886
rect 72683 61886 72871 61914
rect 73003 61914 73031 62026
rect 73467 61914 73495 62026
rect 73003 61886 73191 61914
rect 72683 61774 72711 61886
rect 73163 61774 73191 61886
rect 73235 61886 73495 61914
rect 73627 61914 73655 62026
rect 74091 61914 74119 62026
rect 73627 61886 73887 61914
rect 73235 61774 73263 61886
rect 73859 61774 73887 61886
rect 73931 61886 74119 61914
rect 74251 61914 74279 62026
rect 74715 61914 74743 62026
rect 74251 61886 74439 61914
rect 73931 61774 73959 61886
rect 74411 61774 74439 61886
rect 74483 61886 74743 61914
rect 74875 61914 74903 62026
rect 75339 61914 75367 62026
rect 74875 61886 75135 61914
rect 74483 61774 74511 61886
rect 75107 61774 75135 61886
rect 75179 61886 75367 61914
rect 75499 61914 75527 62026
rect 75963 61914 75991 62026
rect 75499 61886 75687 61914
rect 75179 61774 75207 61886
rect 75659 61774 75687 61886
rect 75731 61886 75991 61914
rect 76123 61914 76151 62026
rect 76587 61914 76615 62026
rect 76123 61886 76383 61914
rect 75731 61774 75759 61886
rect 76355 61774 76383 61886
rect 76427 61886 76615 61914
rect 76747 61914 76775 62026
rect 77211 61914 77239 62026
rect 76747 61886 76935 61914
rect 76427 61774 76455 61886
rect 76907 61774 76935 61886
rect 76979 61886 77239 61914
rect 77371 61914 77399 62026
rect 77835 61914 77863 62026
rect 77371 61886 77631 61914
rect 76979 61774 77007 61886
rect 77603 61774 77631 61886
rect 77675 61886 77863 61914
rect 77995 61914 78023 62026
rect 78459 61914 78487 62026
rect 77995 61886 78183 61914
rect 77675 61774 77703 61886
rect 78155 61774 78183 61886
rect 78227 61886 78487 61914
rect 78619 61914 78647 62026
rect 79083 61914 79111 62026
rect 78619 61886 78879 61914
rect 78227 61774 78255 61886
rect 78851 61774 78879 61886
rect 78923 61886 79111 61914
rect 79243 61914 79271 62026
rect 79707 61914 79735 62026
rect 79243 61886 79431 61914
rect 78923 61774 78951 61886
rect 79403 61774 79431 61886
rect 79475 61886 79735 61914
rect 79867 61914 79895 62026
rect 80331 61914 80359 62026
rect 79867 61886 80127 61914
rect 79475 61774 79503 61886
rect 80099 61774 80127 61886
rect 80171 61886 80359 61914
rect 80491 61914 80519 62026
rect 80955 61914 80983 62026
rect 80491 61886 80679 61914
rect 80171 61774 80199 61886
rect 80651 61774 80679 61886
rect 80723 61886 80983 61914
rect 81115 61914 81143 62026
rect 81579 61914 81607 62026
rect 81115 61886 81375 61914
rect 80723 61774 80751 61886
rect 81347 61774 81375 61886
rect 81419 61886 81607 61914
rect 81739 61914 81767 62026
rect 82203 61914 82231 62026
rect 81739 61886 81927 61914
rect 81419 61774 81447 61886
rect 81899 61774 81927 61886
rect 81971 61886 82231 61914
rect 82363 61914 82391 62026
rect 82827 61914 82855 62026
rect 82363 61886 82623 61914
rect 81971 61774 81999 61886
rect 82595 61774 82623 61886
rect 82667 61886 82855 61914
rect 82987 61914 83015 62026
rect 83451 61914 83479 62026
rect 82987 61886 83175 61914
rect 82667 61774 82695 61886
rect 83147 61774 83175 61886
rect 83219 61886 83479 61914
rect 83611 61914 83639 62026
rect 84075 61914 84103 62026
rect 83611 61886 83871 61914
rect 83219 61774 83247 61886
rect 83843 61774 83871 61886
rect 83915 61886 84103 61914
rect 84235 61914 84263 62026
rect 84699 61914 84727 62026
rect 84235 61886 84423 61914
rect 83915 61774 83943 61886
rect 84395 61774 84423 61886
rect 84467 61886 84727 61914
rect 84859 61914 84887 62026
rect 85323 61914 85351 62026
rect 84859 61886 85119 61914
rect 84467 61774 84495 61886
rect 85091 61774 85119 61886
rect 85163 61886 85351 61914
rect 85483 61914 85511 62026
rect 85947 61914 85975 62026
rect 85483 61886 85671 61914
rect 85163 61774 85191 61886
rect 85643 61774 85671 61886
rect 85715 61886 85975 61914
rect 86107 61914 86135 62026
rect 86571 61914 86599 62026
rect 86107 61886 86367 61914
rect 85715 61774 85743 61886
rect 86339 61774 86367 61886
rect 86411 61886 86599 61914
rect 86731 61914 86759 62026
rect 87195 61914 87223 62026
rect 86731 61886 86919 61914
rect 86411 61774 86439 61886
rect 86891 61774 86919 61886
rect 86963 61886 87223 61914
rect 87355 61914 87383 62026
rect 87819 61914 87847 62026
rect 87355 61886 87615 61914
rect 86963 61774 86991 61886
rect 87587 61774 87615 61886
rect 87659 61886 87847 61914
rect 87979 61914 88007 62026
rect 88443 61914 88471 62026
rect 87979 61886 88167 61914
rect 87659 61774 87687 61886
rect 88139 61774 88167 61886
rect 88211 61886 88471 61914
rect 88603 61914 88631 62026
rect 89067 61914 89095 62026
rect 88603 61886 88863 61914
rect 88211 61774 88239 61886
rect 88835 61774 88863 61886
rect 88907 61886 89095 61914
rect 89227 61914 89255 62026
rect 89691 61914 89719 62026
rect 89227 61886 89415 61914
rect 88907 61774 88935 61886
rect 89387 61774 89415 61886
rect 89459 61886 89719 61914
rect 89851 61914 89879 62026
rect 90315 61914 90343 62026
rect 89851 61886 90111 61914
rect 89459 61774 89487 61886
rect 90083 61774 90111 61886
rect 90155 61886 90343 61914
rect 90475 61914 90503 62026
rect 90939 61914 90967 62026
rect 90475 61886 90663 61914
rect 90155 61774 90183 61886
rect 90635 61774 90663 61886
rect 90707 61886 90967 61914
rect 91099 61914 91127 62026
rect 91563 61914 91591 62026
rect 91099 61886 91359 61914
rect 90707 61774 90735 61886
rect 91331 61774 91359 61886
rect 91403 61886 91591 61914
rect 91723 61914 91751 62026
rect 92187 61914 92215 62026
rect 91723 61886 91911 61914
rect 91403 61774 91431 61886
rect 91883 61774 91911 61886
rect 91955 61886 92215 61914
rect 92347 61914 92375 62026
rect 92811 61914 92839 62026
rect 92347 61886 92607 61914
rect 91955 61774 91983 61886
rect 92579 61774 92607 61886
rect 92651 61886 92839 61914
rect 92971 61914 92999 62026
rect 93435 61914 93463 62026
rect 92971 61886 93159 61914
rect 92651 61774 92679 61886
rect 93131 61774 93159 61886
rect 93203 61886 93463 61914
rect 93595 61914 93623 62026
rect 94059 61914 94087 62026
rect 93595 61886 93855 61914
rect 93203 61774 93231 61886
rect 93827 61774 93855 61886
rect 93899 61886 94087 61914
rect 93899 61774 93927 61886
rect 94998 61078 95062 61130
rect 12124 60838 12188 60890
rect 94998 60838 95062 60890
rect 12124 60288 12188 60340
rect 94998 60288 95062 60340
rect 12124 60048 12188 60100
rect 94998 60048 95062 60100
rect 12124 59498 12188 59550
rect 94998 59498 95062 59550
rect 12124 59258 12188 59310
rect 94998 59258 95062 59310
rect 12124 58708 12188 58760
rect 94998 58708 95062 58760
rect 12124 58468 12188 58520
rect 94998 58468 95062 58520
rect 12124 57918 12188 57970
rect 94998 57918 95062 57970
rect 12124 57678 12188 57730
rect 94998 57678 95062 57730
rect 12124 57128 12188 57180
rect 94998 57128 95062 57180
rect 12124 56888 12188 56940
rect 94998 56888 95062 56940
rect 12124 56338 12188 56390
rect 94998 56338 95062 56390
rect 12124 56098 12188 56150
rect 94998 56098 95062 56150
rect 12124 55548 12188 55600
rect 94998 55548 95062 55600
rect 12124 55308 12188 55360
rect 94998 55308 95062 55360
rect 12124 54758 12188 54810
rect 94998 54758 95062 54810
rect 12124 54518 12188 54570
rect 94998 54518 95062 54570
rect 12124 53968 12188 54020
rect 94998 53968 95062 54020
rect 12124 53728 12188 53780
rect 94998 53728 95062 53780
rect 12124 53178 12188 53230
rect 94998 53178 95062 53230
rect 12124 52938 12188 52990
rect 94998 52938 95062 52990
rect 12124 52388 12188 52440
rect 94998 52388 95062 52440
rect 12124 52148 12188 52200
rect 94998 52148 95062 52200
rect 12124 51598 12188 51650
rect 94998 51598 95062 51650
rect 12124 51358 12188 51410
rect 94998 51358 95062 51410
rect 12124 50808 12188 50860
rect 94998 50808 95062 50860
rect 12124 50568 12188 50620
rect 94998 50568 95062 50620
rect 12124 50018 12188 50070
rect 94998 50018 95062 50070
rect 12124 49778 12188 49830
rect 94998 49778 95062 49830
rect 12124 49228 12188 49280
rect 94998 49228 95062 49280
rect 12124 48988 12188 49040
rect 94998 48988 95062 49040
rect 12124 48438 12188 48490
rect 94998 48438 95062 48490
rect 12124 48198 12188 48250
rect 94998 48198 95062 48250
rect 12124 47648 12188 47700
rect 94998 47648 95062 47700
rect 12124 47408 12188 47460
rect 94998 47408 95062 47460
rect 12124 46858 12188 46910
rect 94998 46858 95062 46910
rect 12124 46618 12188 46670
rect 94998 46618 95062 46670
rect 12124 46068 12188 46120
rect 94998 46068 95062 46120
rect 12124 45828 12188 45880
rect 94998 45828 95062 45880
rect 12124 45278 12188 45330
rect 94998 45278 95062 45330
rect 12124 45038 12188 45090
rect 94998 45038 95062 45090
rect 12124 44488 12188 44540
rect 94998 44488 95062 44540
rect 12124 44248 12188 44300
rect 94998 44248 95062 44300
rect 12124 43698 12188 43750
rect 94998 43698 95062 43750
rect 12124 43458 12188 43510
rect 94998 43458 95062 43510
rect 12124 42908 12188 42960
rect 94998 42908 95062 42960
rect 12124 42668 12188 42720
rect 94998 42668 95062 42720
rect 12124 42118 12188 42170
rect 94998 42118 95062 42170
rect 12124 41878 12188 41930
rect 94998 41878 95062 41930
rect 12124 41328 12188 41380
rect 94998 41328 95062 41380
rect 12124 41088 12188 41140
rect 94998 41088 95062 41140
rect 12124 40538 12188 40590
rect 94998 40538 95062 40590
rect 12124 40298 12188 40350
rect 94998 40298 95062 40350
rect 12124 39748 12188 39800
rect 94998 39748 95062 39800
rect 12124 39508 12188 39560
rect 94998 39508 95062 39560
rect 12124 38958 12188 39010
rect 94998 38958 95062 39010
rect 12124 38718 12188 38770
rect 94998 38718 95062 38770
rect 12124 38168 12188 38220
rect 94998 38168 95062 38220
rect 12124 37928 12188 37980
rect 94998 37928 95062 37980
rect 12124 37378 12188 37430
rect 94998 37378 95062 37430
rect 12124 37138 12188 37190
rect 94998 37138 95062 37190
rect 12124 36588 12188 36640
rect 94998 36588 95062 36640
rect 12124 36348 12188 36400
rect 94998 36348 95062 36400
rect 12124 35798 12188 35850
rect 94998 35798 95062 35850
rect 12124 35558 12188 35610
rect 94998 35558 95062 35610
rect 12124 35008 12188 35060
rect 94998 35008 95062 35060
rect 12124 34768 12188 34820
rect 94998 34768 95062 34820
rect 12124 34218 12188 34270
rect 94998 34218 95062 34270
rect 12124 33978 12188 34030
rect 94998 33978 95062 34030
rect 12124 33428 12188 33480
rect 94998 33428 95062 33480
rect 12124 33188 12188 33240
rect 94998 33188 95062 33240
rect 12124 32638 12188 32690
rect 94998 32638 95062 32690
rect 12124 32398 12188 32450
rect 94998 32398 95062 32450
rect 12124 31848 12188 31900
rect 94998 31848 95062 31900
rect 12124 31608 12188 31660
rect 94998 31608 95062 31660
rect 12124 31058 12188 31110
rect 94998 31058 95062 31110
rect 12124 30818 12188 30870
rect 94998 30818 95062 30870
rect 12124 30268 12188 30320
rect 94998 30268 95062 30320
rect 12124 30028 12188 30080
rect 94998 30028 95062 30080
rect 12124 29478 12188 29530
rect 94998 29478 95062 29530
rect 12124 29238 12188 29290
rect 94998 29238 95062 29290
rect 12124 28688 12188 28740
rect 94998 28688 95062 28740
rect 12124 28448 12188 28500
rect 94998 28448 95062 28500
rect 12124 27898 12188 27950
rect 94998 27898 95062 27950
rect 12124 27658 12188 27710
rect 94998 27658 95062 27710
rect 12124 27108 12188 27160
rect 94998 27108 95062 27160
rect 12124 26868 12188 26920
rect 94998 26868 95062 26920
rect 12124 26318 12188 26370
rect 94998 26318 95062 26370
rect 12124 26078 12188 26130
rect 94998 26078 95062 26130
rect 12124 25528 12188 25580
rect 94998 25528 95062 25580
rect 12124 25288 12188 25340
rect 94998 25288 95062 25340
rect 12124 24738 12188 24790
rect 94998 24738 95062 24790
rect 12124 24498 12188 24550
rect 94998 24498 95062 24550
rect 12124 23948 12188 24000
rect 94998 23948 95062 24000
rect 12124 23708 12188 23760
rect 94998 23708 95062 23760
rect 12124 23158 12188 23210
rect 94998 23158 95062 23210
rect 12124 22918 12188 22970
rect 94998 22918 95062 22970
rect 12124 22368 12188 22420
rect 94998 22368 95062 22420
rect 12124 22128 12188 22180
rect 94998 22128 95062 22180
rect 12124 21578 12188 21630
rect 94998 21578 95062 21630
rect 12124 21338 12188 21390
rect 94998 21338 95062 21390
rect 12124 20788 12188 20840
rect 94998 20788 95062 20840
rect 12124 20548 12188 20600
rect 94998 20548 95062 20600
rect 12124 19998 12188 20050
rect 94998 19998 95062 20050
rect 12124 19758 12188 19810
rect 94998 19758 95062 19810
rect 12124 19208 12188 19260
rect 94998 19208 95062 19260
rect 12124 18968 12188 19020
rect 94998 18968 95062 19020
rect 12124 18418 12188 18470
rect 94998 18418 95062 18470
rect 19 10424 47 18324
rect 99 10424 127 18324
rect 179 10424 207 18324
rect 259 10424 287 18324
rect 339 10424 367 18324
rect 419 10424 447 18324
rect 499 10424 527 18324
rect 12124 18178 12188 18230
rect 94998 18178 95062 18230
rect 12124 17628 12188 17680
rect 94998 17628 95062 17680
rect 12124 17388 12188 17440
rect 94998 17388 95062 17440
rect 12124 16838 12188 16890
rect 94998 16838 95062 16890
rect 12124 16598 12188 16650
rect 94998 16598 95062 16650
rect 12124 16048 12188 16100
rect 94998 16048 95062 16100
rect 12124 15808 12188 15860
rect 94998 15808 95062 15860
rect 12124 15258 12188 15310
rect 94998 15258 95062 15310
rect 12124 15018 12188 15070
rect 94998 15018 95062 15070
rect 12124 14468 12188 14520
rect 94998 14468 95062 14520
rect 12124 14228 12188 14280
rect 94998 14228 95062 14280
rect 12124 13678 12188 13730
rect 94998 13678 95062 13730
rect 12124 13438 12188 13490
rect 94998 13438 95062 13490
rect 12124 12888 12188 12940
rect 94998 12888 95062 12940
rect 12124 12648 12188 12700
rect 94998 12648 95062 12700
rect 12124 12098 12188 12150
rect 94998 12098 95062 12150
rect 12124 11858 12188 11910
rect 94998 11858 95062 11910
rect 12124 11308 12188 11360
rect 94998 11308 95062 11360
rect 12124 11068 12188 11120
rect 94998 11068 95062 11120
rect 12124 10518 12188 10570
rect 94998 10518 95062 10570
rect 106659 10424 106687 18324
rect 106739 10424 106767 18324
rect 106819 10424 106847 18324
rect 106899 10424 106927 18324
rect 106979 10424 107007 18324
rect 107059 10424 107087 18324
rect 107139 10424 107167 18324
rect 12124 10278 12188 10330
rect 13475 9522 13503 9634
rect 13099 9494 13503 9522
rect 13547 9522 13575 9634
rect 13739 9522 13767 9634
rect 13547 9494 13591 9522
rect 13099 9382 13127 9494
rect 13563 9382 13591 9494
rect 13723 9494 13767 9522
rect 13811 9522 13839 9634
rect 14723 9522 14751 9634
rect 13811 9494 14215 9522
rect 13723 9382 13751 9494
rect 14187 9382 14215 9494
rect 14347 9494 14751 9522
rect 14795 9522 14823 9634
rect 14987 9522 15015 9634
rect 14795 9494 14839 9522
rect 14347 9382 14375 9494
rect 14811 9382 14839 9494
rect 14971 9494 15015 9522
rect 15059 9522 15087 9634
rect 15971 9522 15999 9634
rect 15059 9494 15463 9522
rect 14971 9382 14999 9494
rect 15435 9382 15463 9494
rect 15595 9494 15999 9522
rect 16043 9522 16071 9634
rect 16235 9522 16263 9634
rect 16043 9494 16087 9522
rect 15595 9382 15623 9494
rect 16059 9382 16087 9494
rect 16219 9494 16263 9522
rect 16307 9522 16335 9634
rect 17219 9522 17247 9634
rect 16307 9494 16711 9522
rect 16219 9382 16247 9494
rect 16683 9382 16711 9494
rect 16843 9494 17247 9522
rect 17291 9522 17319 9634
rect 17483 9522 17511 9634
rect 17291 9494 17335 9522
rect 16843 9382 16871 9494
rect 17307 9382 17335 9494
rect 17467 9494 17511 9522
rect 17555 9522 17583 9634
rect 18467 9522 18495 9634
rect 17555 9494 17959 9522
rect 17467 9382 17495 9494
rect 17931 9382 17959 9494
rect 18091 9494 18495 9522
rect 18539 9522 18567 9634
rect 18731 9522 18759 9634
rect 18539 9494 18583 9522
rect 18091 9382 18119 9494
rect 18555 9382 18583 9494
rect 18715 9494 18759 9522
rect 18803 9522 18831 9634
rect 19715 9522 19743 9634
rect 18803 9494 19207 9522
rect 18715 9382 18743 9494
rect 19179 9382 19207 9494
rect 19339 9494 19743 9522
rect 19787 9522 19815 9634
rect 19979 9522 20007 9634
rect 19787 9494 19831 9522
rect 19339 9382 19367 9494
rect 19803 9382 19831 9494
rect 19963 9494 20007 9522
rect 20051 9522 20079 9634
rect 20963 9522 20991 9634
rect 20051 9494 20455 9522
rect 19963 9382 19991 9494
rect 20427 9382 20455 9494
rect 20587 9494 20991 9522
rect 21035 9522 21063 9634
rect 21227 9522 21255 9634
rect 21035 9494 21079 9522
rect 20587 9382 20615 9494
rect 21051 9382 21079 9494
rect 21211 9494 21255 9522
rect 21299 9522 21327 9634
rect 22211 9522 22239 9634
rect 21299 9494 21703 9522
rect 21211 9382 21239 9494
rect 21675 9382 21703 9494
rect 21835 9494 22239 9522
rect 22283 9522 22311 9634
rect 22475 9522 22503 9634
rect 22283 9494 22327 9522
rect 21835 9382 21863 9494
rect 22299 9382 22327 9494
rect 22459 9494 22503 9522
rect 22547 9522 22575 9634
rect 23459 9522 23487 9634
rect 22547 9494 22951 9522
rect 22459 9382 22487 9494
rect 22923 9382 22951 9494
rect 23083 9494 23487 9522
rect 23531 9522 23559 9634
rect 23723 9522 23751 9634
rect 23531 9494 23575 9522
rect 23083 9382 23111 9494
rect 23547 9382 23575 9494
rect 23707 9494 23751 9522
rect 23795 9522 23823 9634
rect 24707 9522 24735 9634
rect 23795 9494 24199 9522
rect 23707 9382 23735 9494
rect 24171 9382 24199 9494
rect 24331 9494 24735 9522
rect 24779 9522 24807 9634
rect 24971 9522 24999 9634
rect 24779 9494 24823 9522
rect 24331 9382 24359 9494
rect 24795 9382 24823 9494
rect 24955 9494 24999 9522
rect 25043 9522 25071 9634
rect 25955 9522 25983 9634
rect 25043 9494 25447 9522
rect 24955 9382 24983 9494
rect 25419 9382 25447 9494
rect 25579 9494 25983 9522
rect 26027 9522 26055 9634
rect 26219 9522 26247 9634
rect 26027 9494 26071 9522
rect 25579 9382 25607 9494
rect 26043 9382 26071 9494
rect 26203 9494 26247 9522
rect 26291 9522 26319 9634
rect 27203 9522 27231 9634
rect 26291 9494 26695 9522
rect 26203 9382 26231 9494
rect 26667 9382 26695 9494
rect 26827 9494 27231 9522
rect 27275 9522 27303 9634
rect 27467 9522 27495 9634
rect 27275 9494 27319 9522
rect 26827 9382 26855 9494
rect 27291 9382 27319 9494
rect 27451 9494 27495 9522
rect 27539 9522 27567 9634
rect 28451 9522 28479 9634
rect 27539 9494 27943 9522
rect 27451 9382 27479 9494
rect 27915 9382 27943 9494
rect 28075 9494 28479 9522
rect 28523 9522 28551 9634
rect 28715 9522 28743 9634
rect 28523 9494 28567 9522
rect 28075 9382 28103 9494
rect 28539 9382 28567 9494
rect 28699 9494 28743 9522
rect 28787 9522 28815 9634
rect 29699 9522 29727 9634
rect 28787 9494 29191 9522
rect 28699 9382 28727 9494
rect 29163 9382 29191 9494
rect 29323 9494 29727 9522
rect 29771 9522 29799 9634
rect 29963 9522 29991 9634
rect 29771 9494 29815 9522
rect 29323 9382 29351 9494
rect 29787 9382 29815 9494
rect 29947 9494 29991 9522
rect 30035 9522 30063 9634
rect 30947 9522 30975 9634
rect 30035 9494 30439 9522
rect 29947 9382 29975 9494
rect 30411 9382 30439 9494
rect 30571 9494 30975 9522
rect 31019 9522 31047 9634
rect 31211 9522 31239 9634
rect 31019 9494 31063 9522
rect 30571 9382 30599 9494
rect 31035 9382 31063 9494
rect 31195 9494 31239 9522
rect 31283 9522 31311 9634
rect 32195 9522 32223 9634
rect 31283 9494 31687 9522
rect 31195 9382 31223 9494
rect 31659 9382 31687 9494
rect 31819 9494 32223 9522
rect 32267 9522 32295 9634
rect 32459 9522 32487 9634
rect 32267 9494 32311 9522
rect 31819 9382 31847 9494
rect 32283 9382 32311 9494
rect 32443 9494 32487 9522
rect 32531 9522 32559 9634
rect 33443 9522 33471 9634
rect 32531 9494 32935 9522
rect 32443 9382 32471 9494
rect 32907 9382 32935 9494
rect 33067 9494 33471 9522
rect 33515 9522 33543 9634
rect 33707 9522 33735 9634
rect 33515 9494 33559 9522
rect 33067 9382 33095 9494
rect 33531 9382 33559 9494
rect 33691 9494 33735 9522
rect 33779 9522 33807 9634
rect 34691 9522 34719 9634
rect 33779 9494 34183 9522
rect 33691 9382 33719 9494
rect 34155 9382 34183 9494
rect 34315 9494 34719 9522
rect 34763 9522 34791 9634
rect 34955 9522 34983 9634
rect 34763 9494 34807 9522
rect 34315 9382 34343 9494
rect 34779 9382 34807 9494
rect 34939 9494 34983 9522
rect 35027 9522 35055 9634
rect 35939 9522 35967 9634
rect 35027 9494 35431 9522
rect 34939 9382 34967 9494
rect 35403 9382 35431 9494
rect 35563 9494 35967 9522
rect 36011 9522 36039 9634
rect 36203 9522 36231 9634
rect 36011 9494 36055 9522
rect 35563 9382 35591 9494
rect 36027 9382 36055 9494
rect 36187 9494 36231 9522
rect 36275 9522 36303 9634
rect 37187 9522 37215 9634
rect 36275 9494 36679 9522
rect 36187 9382 36215 9494
rect 36651 9382 36679 9494
rect 36811 9494 37215 9522
rect 37259 9522 37287 9634
rect 37451 9522 37479 9634
rect 37259 9494 37303 9522
rect 36811 9382 36839 9494
rect 37275 9382 37303 9494
rect 37435 9494 37479 9522
rect 37523 9522 37551 9634
rect 38435 9522 38463 9634
rect 37523 9494 37927 9522
rect 37435 9382 37463 9494
rect 37899 9382 37927 9494
rect 38059 9494 38463 9522
rect 38507 9522 38535 9634
rect 38699 9522 38727 9634
rect 38507 9494 38551 9522
rect 38059 9382 38087 9494
rect 38523 9382 38551 9494
rect 38683 9494 38727 9522
rect 38771 9522 38799 9634
rect 39683 9522 39711 9634
rect 38771 9494 39175 9522
rect 38683 9382 38711 9494
rect 39147 9382 39175 9494
rect 39307 9494 39711 9522
rect 39755 9522 39783 9634
rect 39947 9522 39975 9634
rect 39755 9494 39799 9522
rect 39307 9382 39335 9494
rect 39771 9382 39799 9494
rect 39931 9494 39975 9522
rect 40019 9522 40047 9634
rect 40931 9522 40959 9634
rect 40019 9494 40423 9522
rect 39931 9382 39959 9494
rect 40395 9382 40423 9494
rect 40555 9494 40959 9522
rect 41003 9522 41031 9634
rect 41195 9522 41223 9634
rect 41003 9494 41047 9522
rect 40555 9382 40583 9494
rect 41019 9382 41047 9494
rect 41179 9494 41223 9522
rect 41267 9522 41295 9634
rect 42179 9522 42207 9634
rect 41267 9494 41671 9522
rect 41179 9382 41207 9494
rect 41643 9382 41671 9494
rect 41803 9494 42207 9522
rect 42251 9522 42279 9634
rect 42443 9522 42471 9634
rect 42251 9494 42295 9522
rect 41803 9382 41831 9494
rect 42267 9382 42295 9494
rect 42427 9494 42471 9522
rect 42515 9522 42543 9634
rect 43427 9522 43455 9634
rect 42515 9494 42919 9522
rect 42427 9382 42455 9494
rect 42891 9382 42919 9494
rect 43051 9494 43455 9522
rect 43499 9522 43527 9634
rect 43691 9522 43719 9634
rect 43499 9494 43543 9522
rect 43051 9382 43079 9494
rect 43515 9382 43543 9494
rect 43675 9494 43719 9522
rect 43763 9522 43791 9634
rect 44675 9522 44703 9634
rect 43763 9494 44167 9522
rect 43675 9382 43703 9494
rect 44139 9382 44167 9494
rect 44299 9494 44703 9522
rect 44747 9522 44775 9634
rect 44939 9522 44967 9634
rect 44747 9494 44791 9522
rect 44299 9382 44327 9494
rect 44763 9382 44791 9494
rect 44923 9494 44967 9522
rect 45011 9522 45039 9634
rect 45923 9522 45951 9634
rect 45011 9494 45415 9522
rect 44923 9382 44951 9494
rect 45387 9382 45415 9494
rect 45547 9494 45951 9522
rect 45995 9522 46023 9634
rect 46187 9522 46215 9634
rect 45995 9494 46039 9522
rect 45547 9382 45575 9494
rect 46011 9382 46039 9494
rect 46171 9494 46215 9522
rect 46259 9522 46287 9634
rect 47171 9522 47199 9634
rect 46259 9494 46663 9522
rect 46171 9382 46199 9494
rect 46635 9382 46663 9494
rect 46795 9494 47199 9522
rect 47243 9522 47271 9634
rect 47435 9522 47463 9634
rect 47243 9494 47287 9522
rect 46795 9382 46823 9494
rect 47259 9382 47287 9494
rect 47419 9494 47463 9522
rect 47507 9522 47535 9634
rect 48419 9522 48447 9634
rect 47507 9494 47911 9522
rect 47419 9382 47447 9494
rect 47883 9382 47911 9494
rect 48043 9494 48447 9522
rect 48491 9522 48519 9634
rect 48683 9522 48711 9634
rect 48491 9494 48535 9522
rect 48043 9382 48071 9494
rect 48507 9382 48535 9494
rect 48667 9494 48711 9522
rect 48755 9522 48783 9634
rect 49667 9522 49695 9634
rect 48755 9494 49159 9522
rect 48667 9382 48695 9494
rect 49131 9382 49159 9494
rect 49291 9494 49695 9522
rect 49739 9522 49767 9634
rect 49931 9522 49959 9634
rect 49739 9494 49783 9522
rect 49291 9382 49319 9494
rect 49755 9382 49783 9494
rect 49915 9494 49959 9522
rect 50003 9522 50031 9634
rect 50915 9522 50943 9634
rect 50003 9494 50407 9522
rect 49915 9382 49943 9494
rect 50379 9382 50407 9494
rect 50539 9494 50943 9522
rect 50987 9522 51015 9634
rect 51179 9522 51207 9634
rect 50987 9494 51031 9522
rect 50539 9382 50567 9494
rect 51003 9382 51031 9494
rect 51163 9494 51207 9522
rect 51251 9522 51279 9634
rect 52163 9522 52191 9634
rect 51251 9494 51655 9522
rect 51163 9382 51191 9494
rect 51627 9382 51655 9494
rect 51787 9494 52191 9522
rect 52235 9522 52263 9634
rect 52427 9522 52455 9634
rect 52235 9494 52279 9522
rect 51787 9382 51815 9494
rect 52251 9382 52279 9494
rect 52411 9494 52455 9522
rect 52499 9522 52527 9634
rect 53411 9522 53439 9634
rect 52499 9494 52903 9522
rect 52411 9382 52439 9494
rect 52875 9382 52903 9494
rect 53035 9494 53439 9522
rect 53483 9522 53511 9634
rect 53675 9522 53703 9634
rect 53483 9494 53527 9522
rect 53035 9382 53063 9494
rect 53499 9382 53527 9494
rect 53659 9494 53703 9522
rect 53747 9522 53775 9634
rect 54659 9522 54687 9634
rect 53747 9494 54151 9522
rect 53659 9382 53687 9494
rect 54123 9382 54151 9494
rect 54283 9494 54687 9522
rect 54731 9522 54759 9634
rect 54923 9522 54951 9634
rect 54731 9494 54775 9522
rect 54283 9382 54311 9494
rect 54747 9382 54775 9494
rect 54907 9494 54951 9522
rect 54995 9522 55023 9634
rect 55907 9522 55935 9634
rect 54995 9494 55399 9522
rect 54907 9382 54935 9494
rect 55371 9382 55399 9494
rect 55531 9494 55935 9522
rect 55979 9522 56007 9634
rect 56171 9522 56199 9634
rect 55979 9494 56023 9522
rect 55531 9382 55559 9494
rect 55995 9382 56023 9494
rect 56155 9494 56199 9522
rect 56243 9522 56271 9634
rect 57155 9522 57183 9634
rect 56243 9494 56647 9522
rect 56155 9382 56183 9494
rect 56619 9382 56647 9494
rect 56779 9494 57183 9522
rect 57227 9522 57255 9634
rect 57419 9522 57447 9634
rect 57227 9494 57271 9522
rect 56779 9382 56807 9494
rect 57243 9382 57271 9494
rect 57403 9494 57447 9522
rect 57491 9522 57519 9634
rect 58403 9522 58431 9634
rect 57491 9494 57895 9522
rect 57403 9382 57431 9494
rect 57867 9382 57895 9494
rect 58027 9494 58431 9522
rect 58475 9522 58503 9634
rect 58667 9522 58695 9634
rect 58475 9494 58519 9522
rect 58027 9382 58055 9494
rect 58491 9382 58519 9494
rect 58651 9494 58695 9522
rect 58739 9522 58767 9634
rect 59651 9522 59679 9634
rect 58739 9494 59143 9522
rect 58651 9382 58679 9494
rect 59115 9382 59143 9494
rect 59275 9494 59679 9522
rect 59723 9522 59751 9634
rect 59915 9522 59943 9634
rect 59723 9494 59767 9522
rect 59275 9382 59303 9494
rect 59739 9382 59767 9494
rect 59899 9494 59943 9522
rect 59987 9522 60015 9634
rect 60899 9522 60927 9634
rect 59987 9494 60391 9522
rect 59899 9382 59927 9494
rect 60363 9382 60391 9494
rect 60523 9494 60927 9522
rect 60971 9522 60999 9634
rect 61163 9522 61191 9634
rect 60971 9494 61015 9522
rect 60523 9382 60551 9494
rect 60987 9382 61015 9494
rect 61147 9494 61191 9522
rect 61235 9522 61263 9634
rect 62147 9522 62175 9634
rect 61235 9494 61639 9522
rect 61147 9382 61175 9494
rect 61611 9382 61639 9494
rect 61771 9494 62175 9522
rect 62219 9522 62247 9634
rect 62411 9522 62439 9634
rect 62219 9494 62263 9522
rect 61771 9382 61799 9494
rect 62235 9382 62263 9494
rect 62395 9494 62439 9522
rect 62483 9522 62511 9634
rect 63395 9522 63423 9634
rect 62483 9494 62887 9522
rect 62395 9382 62423 9494
rect 62859 9382 62887 9494
rect 63019 9494 63423 9522
rect 63467 9522 63495 9634
rect 63659 9522 63687 9634
rect 63467 9494 63511 9522
rect 63019 9382 63047 9494
rect 63483 9382 63511 9494
rect 63643 9494 63687 9522
rect 63731 9522 63759 9634
rect 64643 9522 64671 9634
rect 63731 9494 64135 9522
rect 63643 9382 63671 9494
rect 64107 9382 64135 9494
rect 64267 9494 64671 9522
rect 64715 9522 64743 9634
rect 64907 9522 64935 9634
rect 64715 9494 64759 9522
rect 64267 9382 64295 9494
rect 64731 9382 64759 9494
rect 64891 9494 64935 9522
rect 64979 9522 65007 9634
rect 65891 9522 65919 9634
rect 64979 9494 65383 9522
rect 64891 9382 64919 9494
rect 65355 9382 65383 9494
rect 65515 9494 65919 9522
rect 65963 9522 65991 9634
rect 66155 9522 66183 9634
rect 65963 9494 66007 9522
rect 65515 9382 65543 9494
rect 65979 9382 66007 9494
rect 66139 9494 66183 9522
rect 66227 9522 66255 9634
rect 67139 9522 67167 9634
rect 66227 9494 66631 9522
rect 66139 9382 66167 9494
rect 66603 9382 66631 9494
rect 66763 9494 67167 9522
rect 67211 9522 67239 9634
rect 67403 9522 67431 9634
rect 67211 9494 67255 9522
rect 66763 9382 66791 9494
rect 67227 9382 67255 9494
rect 67387 9494 67431 9522
rect 67475 9522 67503 9634
rect 68387 9522 68415 9634
rect 67475 9494 67879 9522
rect 67387 9382 67415 9494
rect 67851 9382 67879 9494
rect 68011 9494 68415 9522
rect 68459 9522 68487 9634
rect 68651 9522 68679 9634
rect 68459 9494 68503 9522
rect 68011 9382 68039 9494
rect 68475 9382 68503 9494
rect 68635 9494 68679 9522
rect 68723 9522 68751 9634
rect 69635 9522 69663 9634
rect 68723 9494 69127 9522
rect 68635 9382 68663 9494
rect 69099 9382 69127 9494
rect 69259 9494 69663 9522
rect 69707 9522 69735 9634
rect 69899 9522 69927 9634
rect 69707 9494 69751 9522
rect 69259 9382 69287 9494
rect 69723 9382 69751 9494
rect 69883 9494 69927 9522
rect 69971 9522 69999 9634
rect 70883 9522 70911 9634
rect 69971 9494 70375 9522
rect 69883 9382 69911 9494
rect 70347 9382 70375 9494
rect 70507 9494 70911 9522
rect 70955 9522 70983 9634
rect 71147 9522 71175 9634
rect 70955 9494 70999 9522
rect 70507 9382 70535 9494
rect 70971 9382 70999 9494
rect 71131 9494 71175 9522
rect 71219 9522 71247 9634
rect 72131 9522 72159 9634
rect 71219 9494 71623 9522
rect 71131 9382 71159 9494
rect 71595 9382 71623 9494
rect 71755 9494 72159 9522
rect 72203 9522 72231 9634
rect 72395 9522 72423 9634
rect 72203 9494 72247 9522
rect 71755 9382 71783 9494
rect 72219 9382 72247 9494
rect 72379 9494 72423 9522
rect 72467 9522 72495 9634
rect 73379 9522 73407 9634
rect 72467 9494 72871 9522
rect 72379 9382 72407 9494
rect 72843 9382 72871 9494
rect 73003 9494 73407 9522
rect 73451 9522 73479 9634
rect 73643 9522 73671 9634
rect 73451 9494 73495 9522
rect 73003 9382 73031 9494
rect 73467 9382 73495 9494
rect 73627 9494 73671 9522
rect 73715 9522 73743 9634
rect 74627 9522 74655 9634
rect 73715 9494 74119 9522
rect 73627 9382 73655 9494
rect 74091 9382 74119 9494
rect 74251 9494 74655 9522
rect 74699 9522 74727 9634
rect 74891 9522 74919 9634
rect 74699 9494 74743 9522
rect 74251 9382 74279 9494
rect 74715 9382 74743 9494
rect 74875 9494 74919 9522
rect 74963 9522 74991 9634
rect 75875 9522 75903 9634
rect 74963 9494 75367 9522
rect 74875 9382 74903 9494
rect 75339 9382 75367 9494
rect 75499 9494 75903 9522
rect 75947 9522 75975 9634
rect 76139 9522 76167 9634
rect 75947 9494 75991 9522
rect 75499 9382 75527 9494
rect 75963 9382 75991 9494
rect 76123 9494 76167 9522
rect 76211 9522 76239 9634
rect 77123 9522 77151 9634
rect 76211 9494 76615 9522
rect 76123 9382 76151 9494
rect 76587 9382 76615 9494
rect 76747 9494 77151 9522
rect 77195 9522 77223 9634
rect 77387 9522 77415 9634
rect 77195 9494 77239 9522
rect 76747 9382 76775 9494
rect 77211 9382 77239 9494
rect 77371 9494 77415 9522
rect 77459 9522 77487 9634
rect 78371 9522 78399 9634
rect 77459 9494 77863 9522
rect 77371 9382 77399 9494
rect 77835 9382 77863 9494
rect 77995 9494 78399 9522
rect 78443 9522 78471 9634
rect 78635 9522 78663 9634
rect 78443 9494 78487 9522
rect 77995 9382 78023 9494
rect 78459 9382 78487 9494
rect 78619 9494 78663 9522
rect 78707 9522 78735 9634
rect 79619 9522 79647 9634
rect 78707 9494 79111 9522
rect 78619 9382 78647 9494
rect 79083 9382 79111 9494
rect 79243 9494 79647 9522
rect 79691 9522 79719 9634
rect 79883 9522 79911 9634
rect 79691 9494 79735 9522
rect 79243 9382 79271 9494
rect 79707 9382 79735 9494
rect 79867 9494 79911 9522
rect 79955 9522 79983 9634
rect 80867 9522 80895 9634
rect 79955 9494 80359 9522
rect 79867 9382 79895 9494
rect 80331 9382 80359 9494
rect 80491 9494 80895 9522
rect 80939 9522 80967 9634
rect 81131 9522 81159 9634
rect 80939 9494 80983 9522
rect 80491 9382 80519 9494
rect 80955 9382 80983 9494
rect 81115 9494 81159 9522
rect 81203 9522 81231 9634
rect 82115 9522 82143 9634
rect 81203 9494 81607 9522
rect 81115 9382 81143 9494
rect 81579 9382 81607 9494
rect 81739 9494 82143 9522
rect 82187 9522 82215 9634
rect 82379 9522 82407 9634
rect 82187 9494 82231 9522
rect 81739 9382 81767 9494
rect 82203 9382 82231 9494
rect 82363 9494 82407 9522
rect 82451 9522 82479 9634
rect 83363 9522 83391 9634
rect 82451 9494 82855 9522
rect 82363 9382 82391 9494
rect 82827 9382 82855 9494
rect 82987 9494 83391 9522
rect 83435 9522 83463 9634
rect 83627 9522 83655 9634
rect 83435 9494 83479 9522
rect 82987 9382 83015 9494
rect 83451 9382 83479 9494
rect 83611 9494 83655 9522
rect 83699 9522 83727 9634
rect 84611 9522 84639 9634
rect 83699 9494 84103 9522
rect 83611 9382 83639 9494
rect 84075 9382 84103 9494
rect 84235 9494 84639 9522
rect 84683 9522 84711 9634
rect 84875 9522 84903 9634
rect 84683 9494 84727 9522
rect 84235 9382 84263 9494
rect 84699 9382 84727 9494
rect 84859 9494 84903 9522
rect 84947 9522 84975 9634
rect 85859 9522 85887 9634
rect 84947 9494 85351 9522
rect 84859 9382 84887 9494
rect 85323 9382 85351 9494
rect 85483 9494 85887 9522
rect 85931 9522 85959 9634
rect 86123 9522 86151 9634
rect 85931 9494 85975 9522
rect 85483 9382 85511 9494
rect 85947 9382 85975 9494
rect 86107 9494 86151 9522
rect 86195 9522 86223 9634
rect 87107 9522 87135 9634
rect 86195 9494 86599 9522
rect 86107 9382 86135 9494
rect 86571 9382 86599 9494
rect 86731 9494 87135 9522
rect 87179 9522 87207 9634
rect 87371 9522 87399 9634
rect 87179 9494 87223 9522
rect 86731 9382 86759 9494
rect 87195 9382 87223 9494
rect 87355 9494 87399 9522
rect 87443 9522 87471 9634
rect 88355 9522 88383 9634
rect 87443 9494 87847 9522
rect 87355 9382 87383 9494
rect 87819 9382 87847 9494
rect 87979 9494 88383 9522
rect 88427 9522 88455 9634
rect 88619 9522 88647 9634
rect 88427 9494 88471 9522
rect 87979 9382 88007 9494
rect 88443 9382 88471 9494
rect 88603 9494 88647 9522
rect 88691 9522 88719 9634
rect 89603 9522 89631 9634
rect 88691 9494 89095 9522
rect 88603 9382 88631 9494
rect 89067 9382 89095 9494
rect 89227 9494 89631 9522
rect 89675 9522 89703 9634
rect 89867 9522 89895 9634
rect 89675 9494 89719 9522
rect 89227 9382 89255 9494
rect 89691 9382 89719 9494
rect 89851 9494 89895 9522
rect 89939 9522 89967 9634
rect 90851 9522 90879 9634
rect 89939 9494 90343 9522
rect 89851 9382 89879 9494
rect 90315 9382 90343 9494
rect 90475 9494 90879 9522
rect 90923 9522 90951 9634
rect 91115 9522 91143 9634
rect 90923 9494 90967 9522
rect 90475 9382 90503 9494
rect 90939 9382 90967 9494
rect 91099 9494 91143 9522
rect 91187 9522 91215 9634
rect 92099 9522 92127 9634
rect 91187 9494 91591 9522
rect 91099 9382 91127 9494
rect 91563 9382 91591 9494
rect 91723 9494 92127 9522
rect 92171 9522 92199 9634
rect 92363 9522 92391 9634
rect 92171 9494 92215 9522
rect 91723 9382 91751 9494
rect 92187 9382 92215 9494
rect 92347 9494 92391 9522
rect 92435 9522 92463 9634
rect 93347 9522 93375 9634
rect 92435 9494 92839 9522
rect 92347 9382 92375 9494
rect 92811 9382 92839 9494
rect 92971 9494 93375 9522
rect 93419 9522 93447 9634
rect 93419 9494 93463 9522
rect 92971 9382 92999 9494
rect 93435 9382 93463 9494
rect 13563 8504 13591 8628
rect 7170 7171 7234 7223
rect 7170 5681 7234 5733
rect 5242 4340 5288 4398
rect 7170 4343 7234 4395
rect 13761 3684 13807 3938
rect 16257 3684 16303 3938
rect 18753 3684 18799 3938
rect 21249 3684 21295 3938
rect 23745 3684 23791 3938
rect 26241 3684 26287 3938
rect 28737 3684 28783 3938
rect 31233 3684 31279 3938
rect 33729 3684 33775 3938
rect 36225 3684 36271 3938
rect 38721 3684 38767 3938
rect 41217 3684 41263 3938
rect 43713 3684 43759 3938
rect 46209 3684 46255 3938
rect 48705 3684 48751 3938
rect 51201 3684 51247 3938
rect 53697 3684 53743 3938
rect 56193 3684 56239 3938
rect 58689 3684 58735 3938
rect 61185 3684 61231 3938
rect 63681 3684 63727 3938
rect 66177 3684 66223 3938
rect 68673 3684 68719 3938
rect 71169 3684 71215 3938
rect 73665 3684 73711 3938
rect 76161 3684 76207 3938
rect 78657 3684 78703 3938
rect 81153 3684 81199 3938
rect 83649 3684 83695 3938
rect 86145 3684 86191 3938
rect 88641 3684 88687 3938
rect 91137 3684 91183 3938
rect 5118 2850 5164 2908
rect 7170 2853 7234 2905
rect 13912 1425 13972 1481
rect 16408 1425 16468 1481
rect 18904 1425 18964 1481
rect 21400 1425 21460 1481
rect 23896 1425 23956 1481
rect 26392 1425 26452 1481
rect 28888 1425 28948 1481
rect 31384 1425 31444 1481
rect 33880 1425 33940 1481
rect 36376 1425 36436 1481
rect 38872 1425 38932 1481
rect 41368 1425 41428 1481
rect 43864 1425 43924 1481
rect 46360 1425 46420 1481
rect 48856 1425 48916 1481
rect 51352 1425 51412 1481
rect 53848 1425 53908 1481
rect 56344 1425 56404 1481
rect 58840 1425 58900 1481
rect 61336 1425 61396 1481
rect 63832 1425 63892 1481
rect 66328 1425 66388 1481
rect 68824 1425 68884 1481
rect 71320 1425 71380 1481
rect 73816 1425 73876 1481
rect 76312 1425 76372 1481
rect 78808 1425 78868 1481
rect 81304 1425 81364 1481
rect 83800 1425 83860 1481
rect 86296 1425 86356 1481
rect 88792 1425 88852 1481
rect 91288 1425 91348 1481
<< metal2 >>
rect 93581 62880 93637 62928
rect 95213 61774 95241 69282
rect 95337 61774 95365 69282
rect 99071 64690 99099 67039
rect 99207 64566 99235 65701
rect 99343 64814 99371 68529
rect 99832 68505 99888 68553
rect 99832 67015 99888 67063
rect 99832 65677 99888 65725
rect 99071 64211 99099 64442
rect 99832 64187 99888 64235
rect 99198 61269 99226 61297
rect 94903 61097 95044 61125
rect 12142 60651 12170 60864
rect 94903 60843 95044 60871
rect 12142 60623 12283 60651
rect 12142 60527 12283 60555
rect 12142 60314 12170 60527
rect 94903 60307 95044 60335
rect 12142 59861 12170 60074
rect 94903 60053 95044 60081
rect 12142 59833 12283 59861
rect 12142 59737 12283 59765
rect 12142 59524 12170 59737
rect 94903 59517 95044 59545
rect 12142 59071 12170 59284
rect 94903 59263 95044 59291
rect 12142 59043 12283 59071
rect 12142 58947 12283 58975
rect 12142 58734 12170 58947
rect 94903 58727 95044 58755
rect 12142 58281 12170 58494
rect 94903 58473 95044 58501
rect 12142 58253 12283 58281
rect 12142 58157 12283 58185
rect 12142 57944 12170 58157
rect 94903 57937 95044 57965
rect 12142 57491 12170 57704
rect 94903 57683 95044 57711
rect 12142 57463 12283 57491
rect 12142 57367 12283 57395
rect 12142 57154 12170 57367
rect 94903 57147 95044 57175
rect 12142 56701 12170 56914
rect 94903 56893 95044 56921
rect 12142 56673 12283 56701
rect 12142 56577 12283 56605
rect 12142 56364 12170 56577
rect 94903 56357 95044 56385
rect 12142 55911 12170 56124
rect 94903 56103 95044 56131
rect 12142 55883 12283 55911
rect 12142 55787 12283 55815
rect 12142 55574 12170 55787
rect 94903 55567 95044 55595
rect 12142 55121 12170 55334
rect 94903 55313 95044 55341
rect 12142 55093 12283 55121
rect 12142 54997 12283 55025
rect 12142 54784 12170 54997
rect 94903 54777 95044 54805
rect 12142 54331 12170 54544
rect 94903 54523 95044 54551
rect 12142 54303 12283 54331
rect 12142 54207 12283 54235
rect 12142 53994 12170 54207
rect 94903 53987 95044 54015
rect 12142 53541 12170 53754
rect 94903 53733 95044 53761
rect 12142 53513 12283 53541
rect 12142 53417 12283 53445
rect 12142 53204 12170 53417
rect 94903 53197 95044 53225
rect 12142 52751 12170 52964
rect 94903 52943 95044 52971
rect 12142 52723 12283 52751
rect 12142 52627 12283 52655
rect 12142 52414 12170 52627
rect 94903 52407 95044 52435
rect 12142 51961 12170 52174
rect 94903 52153 95044 52181
rect 12142 51933 12283 51961
rect 12142 51837 12283 51865
rect 12142 51624 12170 51837
rect 94903 51617 95044 51645
rect 12142 51171 12170 51384
rect 94903 51363 95044 51391
rect 12142 51143 12283 51171
rect 12142 51047 12283 51075
rect 12142 50834 12170 51047
rect 94903 50827 95044 50855
rect 12142 50381 12170 50594
rect 94903 50573 95044 50601
rect 12142 50353 12283 50381
rect 12142 50257 12283 50285
rect 12142 50044 12170 50257
rect 94903 50037 95044 50065
rect 12142 49591 12170 49804
rect 94903 49783 95044 49811
rect 12142 49563 12283 49591
rect 12142 49467 12283 49495
rect 12142 49254 12170 49467
rect 94903 49247 95044 49275
rect 12142 48801 12170 49014
rect 94903 48993 95044 49021
rect 12142 48773 12283 48801
rect 12142 48677 12283 48705
rect 12142 48464 12170 48677
rect 94903 48457 95044 48485
rect 12142 48011 12170 48224
rect 94903 48203 95044 48231
rect 12142 47983 12283 48011
rect 12142 47887 12283 47915
rect 12142 47674 12170 47887
rect 94903 47667 95044 47695
rect 12142 47221 12170 47434
rect 94903 47413 95044 47441
rect 12142 47193 12283 47221
rect 12142 47097 12283 47125
rect 12142 46884 12170 47097
rect 94903 46877 95044 46905
rect 12142 46431 12170 46644
rect 94903 46623 95044 46651
rect 12142 46403 12283 46431
rect 12142 46307 12283 46335
rect 12142 46094 12170 46307
rect 94903 46087 95044 46115
rect 12142 45641 12170 45854
rect 94903 45833 95044 45861
rect 12142 45613 12283 45641
rect 12142 45517 12283 45545
rect 12142 45304 12170 45517
rect 94903 45297 95044 45325
rect 12142 44851 12170 45064
rect 94903 45043 95044 45071
rect 12142 44823 12283 44851
rect 12142 44727 12283 44755
rect 12142 44514 12170 44727
rect 94903 44507 95044 44535
rect 12142 44061 12170 44274
rect 94903 44253 95044 44281
rect 12142 44033 12283 44061
rect 12142 43937 12283 43965
rect 12142 43724 12170 43937
rect 94903 43717 95044 43745
rect 12142 43271 12170 43484
rect 94903 43463 95044 43491
rect 12142 43243 12283 43271
rect 12142 43147 12283 43175
rect 12142 42934 12170 43147
rect 94903 42927 95044 42955
rect 12142 42481 12170 42694
rect 94903 42673 95044 42701
rect 12142 42453 12283 42481
rect 12142 42357 12283 42385
rect 12142 42144 12170 42357
rect 94903 42137 95044 42165
rect 12142 41691 12170 41904
rect 94903 41883 95044 41911
rect 12142 41663 12283 41691
rect 12142 41567 12283 41595
rect 12142 41354 12170 41567
rect 94903 41347 95044 41375
rect 12142 40901 12170 41114
rect 94903 41093 95044 41121
rect 12142 40873 12283 40901
rect 12142 40777 12283 40805
rect 12142 40564 12170 40777
rect 94903 40557 95044 40585
rect 12142 40111 12170 40324
rect 94903 40303 95044 40331
rect 12142 40083 12283 40111
rect 12142 39987 12283 40015
rect 12142 39774 12170 39987
rect 94903 39767 95044 39795
rect 12142 39321 12170 39534
rect 94903 39513 95044 39541
rect 12142 39293 12283 39321
rect 12142 39197 12283 39225
rect 12142 38984 12170 39197
rect 94903 38977 95044 39005
rect 12142 38531 12170 38744
rect 94903 38723 95044 38751
rect 12142 38503 12283 38531
rect 12142 38407 12283 38435
rect 12142 38194 12170 38407
rect 94903 38187 95044 38215
rect 12142 37741 12170 37954
rect 94903 37933 95044 37961
rect 12142 37713 12283 37741
rect 12142 37617 12283 37645
rect 12142 37404 12170 37617
rect 94903 37397 95044 37425
rect 12142 36951 12170 37164
rect 94903 37143 95044 37171
rect 12142 36923 12283 36951
rect 12142 36827 12283 36855
rect 12142 36614 12170 36827
rect 94903 36607 95044 36635
rect 12142 36161 12170 36374
rect 94903 36353 95044 36381
rect 12142 36133 12283 36161
rect 12142 36037 12283 36065
rect 12142 35824 12170 36037
rect 94903 35817 95044 35845
rect 12142 35371 12170 35584
rect 94903 35563 95044 35591
rect 12142 35343 12283 35371
rect 12142 35247 12283 35275
rect 12142 35034 12170 35247
rect 94903 35027 95044 35055
rect 12142 34581 12170 34794
rect 94903 34773 95044 34801
rect 12142 34553 12283 34581
rect 12142 34457 12283 34485
rect 12142 34244 12170 34457
rect 94903 34237 95044 34265
rect 12142 33791 12170 34004
rect 94903 33983 95044 34011
rect 12142 33763 12283 33791
rect 12142 33667 12283 33695
rect 12142 33454 12170 33667
rect 94903 33447 95044 33475
rect 12142 33001 12170 33214
rect 94903 33193 95044 33221
rect 12142 32973 12283 33001
rect 12142 32877 12283 32905
rect 12142 32664 12170 32877
rect 94903 32657 95044 32685
rect 12142 32211 12170 32424
rect 94903 32403 95044 32431
rect 12142 32183 12283 32211
rect 12142 32087 12283 32115
rect 12142 31874 12170 32087
rect 94903 31867 95044 31895
rect 12142 31421 12170 31634
rect 94903 31613 95044 31641
rect 12142 31393 12283 31421
rect 12142 31297 12283 31325
rect 12142 31084 12170 31297
rect 94903 31077 95044 31105
rect 12142 30631 12170 30844
rect 94903 30823 95044 30851
rect 12142 30603 12283 30631
rect 12142 30507 12283 30535
rect 12142 30294 12170 30507
rect 94903 30287 95044 30315
rect 12142 29841 12170 30054
rect 94903 30033 95044 30061
rect 12142 29813 12283 29841
rect 12142 29717 12283 29745
rect 12142 29504 12170 29717
rect 94903 29497 95044 29525
rect 12142 29051 12170 29264
rect 94903 29243 95044 29271
rect 12142 29023 12283 29051
rect 12142 28927 12283 28955
rect 12142 28714 12170 28927
rect 94903 28707 95044 28735
rect 12142 28261 12170 28474
rect 94903 28453 95044 28481
rect 12142 28233 12283 28261
rect 12142 28137 12283 28165
rect 12142 27924 12170 28137
rect 94903 27917 95044 27945
rect 12142 27471 12170 27684
rect 94903 27663 95044 27691
rect 12142 27443 12283 27471
rect 12142 27347 12283 27375
rect 12142 27134 12170 27347
rect 94903 27127 95044 27155
rect 12142 26681 12170 26894
rect 94903 26873 95044 26901
rect 12142 26653 12283 26681
rect 12142 26557 12283 26585
rect 12142 26344 12170 26557
rect 94903 26337 95044 26365
rect 12142 25891 12170 26104
rect 94903 26083 95044 26111
rect 12142 25863 12283 25891
rect 12142 25767 12283 25795
rect 12142 25554 12170 25767
rect 94903 25547 95044 25575
rect 12142 25101 12170 25314
rect 94903 25293 95044 25321
rect 12142 25073 12283 25101
rect 12142 24977 12283 25005
rect 12142 24764 12170 24977
rect 94903 24757 95044 24785
rect 12142 24311 12170 24524
rect 94903 24503 95044 24531
rect 12142 24283 12283 24311
rect 12142 24187 12283 24215
rect 12142 23974 12170 24187
rect 94903 23967 95044 23995
rect 12142 23521 12170 23734
rect 94903 23713 95044 23741
rect 12142 23493 12283 23521
rect 12142 23397 12283 23425
rect 12142 23184 12170 23397
rect 94903 23177 95044 23205
rect 12142 22731 12170 22944
rect 94903 22923 95044 22951
rect 12142 22703 12283 22731
rect 12142 22607 12283 22635
rect 12142 22394 12170 22607
rect 94903 22387 95044 22415
rect 12142 21941 12170 22154
rect 94903 22133 95044 22161
rect 12142 21913 12283 21941
rect 12142 21817 12283 21845
rect 12142 21604 12170 21817
rect 94903 21597 95044 21625
rect 12142 21151 12170 21364
rect 94903 21343 95044 21371
rect 12142 21123 12283 21151
rect 12142 21027 12283 21055
rect 12142 20814 12170 21027
rect 94903 20807 95044 20835
rect 12142 20361 12170 20574
rect 94903 20553 95044 20581
rect 12142 20333 12283 20361
rect 12142 20237 12283 20265
rect 12142 20024 12170 20237
rect 94903 20017 95044 20045
rect 12142 19571 12170 19784
rect 94903 19763 95044 19791
rect 12142 19543 12283 19571
rect 12142 19447 12283 19475
rect 12142 19234 12170 19447
rect 94903 19227 95044 19255
rect 12142 18781 12170 18994
rect 94903 18973 95044 19001
rect 12142 18753 12283 18781
rect 12142 18657 12283 18685
rect 12142 18444 12170 18657
rect 94903 18437 95044 18465
rect 12142 17991 12170 18204
rect 94903 18183 95044 18211
rect 12142 17963 12283 17991
rect 12142 17867 12283 17895
rect 12142 17654 12170 17867
rect 94903 17647 95044 17675
rect 12142 17201 12170 17414
rect 94903 17393 95044 17421
rect 12142 17173 12283 17201
rect 12142 17077 12283 17105
rect 12142 16864 12170 17077
rect 94903 16857 95044 16885
rect 12142 16411 12170 16624
rect 94903 16603 95044 16631
rect 12142 16383 12283 16411
rect 12142 16287 12283 16315
rect 12142 16074 12170 16287
rect 94903 16067 95044 16095
rect 12142 15621 12170 15834
rect 94903 15813 95044 15841
rect 12142 15593 12283 15621
rect 12142 15497 12283 15525
rect 12142 15284 12170 15497
rect 94903 15277 95044 15305
rect 12142 14831 12170 15044
rect 94903 15023 95044 15051
rect 12142 14803 12283 14831
rect 12142 14707 12283 14735
rect 12142 14494 12170 14707
rect 94903 14487 95044 14515
rect 12142 14041 12170 14254
rect 94903 14233 95044 14261
rect 12142 14013 12283 14041
rect 12142 13917 12283 13945
rect 12142 13704 12170 13917
rect 94903 13697 95044 13725
rect 12142 13251 12170 13464
rect 94903 13443 95044 13471
rect 12142 13223 12283 13251
rect 12142 13127 12283 13155
rect 12142 12914 12170 13127
rect 94903 12907 95044 12935
rect 12142 12461 12170 12674
rect 94903 12653 95044 12681
rect 12142 12433 12283 12461
rect 12142 12337 12283 12365
rect 12142 12124 12170 12337
rect 94903 12117 95044 12145
rect 12142 11671 12170 11884
rect 94903 11863 95044 11891
rect 12142 11643 12283 11671
rect 12142 11547 12283 11575
rect 12142 11334 12170 11547
rect 94903 11327 95044 11355
rect 12142 10881 12170 11094
rect 94903 11073 95044 11101
rect 12142 10853 12283 10881
rect 12142 10757 12283 10785
rect 12142 10544 12170 10757
rect 94903 10537 95044 10565
rect 7960 10111 7988 10139
rect 12142 10091 12170 10304
rect 12142 10063 12283 10091
rect 7174 7173 7230 7221
rect 7467 6966 7495 7197
rect 7174 5683 7230 5731
rect 7174 4345 7230 4393
rect 7174 2855 7230 2903
rect 7467 2879 7495 6594
rect 7603 4369 7631 6718
rect 7739 5707 7767 6842
rect 11663 49 11691 9634
rect 11787 49 11815 9634
rect 11911 49 11939 9634
rect 13549 8480 13605 8528
rect 13643 305 13671 333
rect 33611 305 33639 333
rect 53579 305 53607 333
rect 73547 305 73575 333
<< metal3 >>
rect 100492 69149 100590 69247
rect 101604 69149 101702 69247
rect 99357 68499 99860 68559
rect 100492 67735 100590 67833
rect 101604 67735 101702 67833
rect 13989 67567 14087 67665
rect 16485 67567 16583 67665
rect 18981 67567 19079 67665
rect 21477 67567 21575 67665
rect 23973 67567 24071 67665
rect 26469 67567 26567 67665
rect 28965 67567 29063 67665
rect 31461 67567 31559 67665
rect 33957 67567 34055 67665
rect 36453 67567 36551 67665
rect 38949 67567 39047 67665
rect 41445 67567 41543 67665
rect 43941 67567 44039 67665
rect 46437 67567 46535 67665
rect 48933 67567 49031 67665
rect 51429 67567 51527 67665
rect 53925 67567 54023 67665
rect 56421 67567 56519 67665
rect 58917 67567 59015 67665
rect 61413 67567 61511 67665
rect 63909 67567 64007 67665
rect 66405 67567 66503 67665
rect 68901 67567 68999 67665
rect 71397 67567 71495 67665
rect 73893 67567 73991 67665
rect 76389 67567 76487 67665
rect 78885 67567 78983 67665
rect 81381 67567 81479 67665
rect 83877 67567 83975 67665
rect 86373 67567 86471 67665
rect 88869 67567 88967 67665
rect 91365 67567 91463 67665
rect 13989 67245 14087 67343
rect 16485 67245 16583 67343
rect 18981 67245 19079 67343
rect 21477 67245 21575 67343
rect 23973 67245 24071 67343
rect 26469 67245 26567 67343
rect 28965 67245 29063 67343
rect 31461 67245 31559 67343
rect 33957 67245 34055 67343
rect 36453 67245 36551 67343
rect 38949 67245 39047 67343
rect 41445 67245 41543 67343
rect 43941 67245 44039 67343
rect 46437 67245 46535 67343
rect 48933 67245 49031 67343
rect 51429 67245 51527 67343
rect 53925 67245 54023 67343
rect 56421 67245 56519 67343
rect 58917 67245 59015 67343
rect 61413 67245 61511 67343
rect 63909 67245 64007 67343
rect 66405 67245 66503 67343
rect 68901 67245 68999 67343
rect 71397 67245 71495 67343
rect 73893 67245 73991 67343
rect 76389 67245 76487 67343
rect 78885 67245 78983 67343
rect 81381 67245 81479 67343
rect 83877 67245 83975 67343
rect 86373 67245 86471 67343
rect 88869 67245 88967 67343
rect 91365 67245 91463 67343
rect 99085 67009 99860 67069
rect 13977 66407 14075 66505
rect 16473 66407 16571 66505
rect 18969 66407 19067 66505
rect 21465 66407 21563 66505
rect 23961 66407 24059 66505
rect 26457 66407 26555 66505
rect 28953 66407 29051 66505
rect 31449 66407 31547 66505
rect 33945 66407 34043 66505
rect 36441 66407 36539 66505
rect 38937 66407 39035 66505
rect 41433 66407 41531 66505
rect 43929 66407 44027 66505
rect 46425 66407 46523 66505
rect 48921 66407 49019 66505
rect 51417 66407 51515 66505
rect 53913 66407 54011 66505
rect 56409 66407 56507 66505
rect 58905 66407 59003 66505
rect 61401 66407 61499 66505
rect 63897 66407 63995 66505
rect 66393 66407 66491 66505
rect 68889 66407 68987 66505
rect 71385 66407 71483 66505
rect 73881 66407 73979 66505
rect 76377 66407 76475 66505
rect 78873 66407 78971 66505
rect 81369 66407 81467 66505
rect 83865 66407 83963 66505
rect 86361 66407 86459 66505
rect 88857 66407 88955 66505
rect 91353 66407 91451 66505
rect 100492 66321 100590 66419
rect 101604 66321 101702 66419
rect 14059 65633 14157 65731
rect 16555 65633 16653 65731
rect 19051 65633 19149 65731
rect 21547 65633 21645 65731
rect 24043 65633 24141 65731
rect 26539 65633 26637 65731
rect 29035 65633 29133 65731
rect 31531 65633 31629 65731
rect 34027 65633 34125 65731
rect 36523 65633 36621 65731
rect 39019 65633 39117 65731
rect 41515 65633 41613 65731
rect 44011 65633 44109 65731
rect 46507 65633 46605 65731
rect 49003 65633 49101 65731
rect 51499 65633 51597 65731
rect 53995 65633 54093 65731
rect 56491 65633 56589 65731
rect 58987 65633 59085 65731
rect 61483 65633 61581 65731
rect 63979 65633 64077 65731
rect 66475 65633 66573 65731
rect 68971 65633 69069 65731
rect 71467 65633 71565 65731
rect 73963 65633 74061 65731
rect 76459 65633 76557 65731
rect 78955 65633 79053 65731
rect 81451 65633 81549 65731
rect 83947 65633 84045 65731
rect 86443 65633 86541 65731
rect 88939 65633 89037 65731
rect 91435 65633 91533 65731
rect 99221 65671 99860 65731
rect 51908 65500 95227 65560
rect 100492 64907 100590 65005
rect 101604 64907 101702 65005
rect 93499 64784 99357 64844
rect 93499 64660 99085 64720
rect 93499 64536 99221 64596
rect 93499 64412 99085 64472
rect 99085 64181 99860 64241
rect 14232 63636 14330 63734
rect 15480 63636 15578 63734
rect 16728 63636 16826 63734
rect 17976 63636 18074 63734
rect 19224 63636 19322 63734
rect 20472 63636 20570 63734
rect 21720 63636 21818 63734
rect 22968 63636 23066 63734
rect 24216 63636 24314 63734
rect 25464 63636 25562 63734
rect 26712 63636 26810 63734
rect 27960 63636 28058 63734
rect 29208 63636 29306 63734
rect 30456 63636 30554 63734
rect 31704 63636 31802 63734
rect 32952 63636 33050 63734
rect 34200 63636 34298 63734
rect 35448 63636 35546 63734
rect 36696 63636 36794 63734
rect 37944 63636 38042 63734
rect 39192 63636 39290 63734
rect 40440 63636 40538 63734
rect 41688 63636 41786 63734
rect 42936 63636 43034 63734
rect 44184 63636 44282 63734
rect 45432 63636 45530 63734
rect 46680 63636 46778 63734
rect 47928 63636 48026 63734
rect 49176 63636 49274 63734
rect 50424 63636 50522 63734
rect 51672 63636 51770 63734
rect 52920 63636 53018 63734
rect 54168 63636 54266 63734
rect 55416 63636 55514 63734
rect 56664 63636 56762 63734
rect 57912 63636 58010 63734
rect 59160 63636 59258 63734
rect 60408 63636 60506 63734
rect 61656 63636 61754 63734
rect 62904 63636 63002 63734
rect 64152 63636 64250 63734
rect 65400 63636 65498 63734
rect 66648 63636 66746 63734
rect 67896 63636 67994 63734
rect 69144 63636 69242 63734
rect 70392 63636 70490 63734
rect 71640 63636 71738 63734
rect 72888 63636 72986 63734
rect 74136 63636 74234 63734
rect 75384 63636 75482 63734
rect 76632 63636 76730 63734
rect 77880 63636 77978 63734
rect 79128 63636 79226 63734
rect 80376 63636 80474 63734
rect 81624 63636 81722 63734
rect 82872 63636 82970 63734
rect 84120 63636 84218 63734
rect 85368 63636 85466 63734
rect 86616 63636 86714 63734
rect 87864 63636 87962 63734
rect 89112 63636 89210 63734
rect 90360 63636 90458 63734
rect 91608 63636 91706 63734
rect 92856 63636 92954 63734
rect 100492 63493 100590 63591
rect 101604 63493 101702 63591
rect 93609 62874 107270 62934
rect 53218 62725 95351 62785
rect 13801 62087 13899 62185
rect 14663 62087 14761 62185
rect 15049 62087 15147 62185
rect 15911 62087 16009 62185
rect 16297 62087 16395 62185
rect 17159 62087 17257 62185
rect 17545 62087 17643 62185
rect 18407 62087 18505 62185
rect 18793 62087 18891 62185
rect 19655 62087 19753 62185
rect 20041 62087 20139 62185
rect 20903 62087 21001 62185
rect 21289 62087 21387 62185
rect 22151 62087 22249 62185
rect 22537 62087 22635 62185
rect 23399 62087 23497 62185
rect 23785 62087 23883 62185
rect 24647 62087 24745 62185
rect 25033 62087 25131 62185
rect 25895 62087 25993 62185
rect 26281 62087 26379 62185
rect 27143 62087 27241 62185
rect 27529 62087 27627 62185
rect 28391 62087 28489 62185
rect 28777 62087 28875 62185
rect 29639 62087 29737 62185
rect 30025 62087 30123 62185
rect 30887 62087 30985 62185
rect 31273 62087 31371 62185
rect 32135 62087 32233 62185
rect 32521 62087 32619 62185
rect 33383 62087 33481 62185
rect 33769 62087 33867 62185
rect 34631 62087 34729 62185
rect 35017 62087 35115 62185
rect 35879 62087 35977 62185
rect 36265 62087 36363 62185
rect 37127 62087 37225 62185
rect 37513 62087 37611 62185
rect 38375 62087 38473 62185
rect 38761 62087 38859 62185
rect 39623 62087 39721 62185
rect 40009 62087 40107 62185
rect 40871 62087 40969 62185
rect 41257 62087 41355 62185
rect 42119 62087 42217 62185
rect 42505 62087 42603 62185
rect 43367 62087 43465 62185
rect 43753 62087 43851 62185
rect 44615 62087 44713 62185
rect 45001 62087 45099 62185
rect 45863 62087 45961 62185
rect 46249 62087 46347 62185
rect 47111 62087 47209 62185
rect 47497 62087 47595 62185
rect 48359 62087 48457 62185
rect 48745 62087 48843 62185
rect 49607 62087 49705 62185
rect 49993 62087 50091 62185
rect 50855 62087 50953 62185
rect 51241 62087 51339 62185
rect 52103 62087 52201 62185
rect 52489 62087 52587 62185
rect 53351 62087 53449 62185
rect 53737 62087 53835 62185
rect 54599 62087 54697 62185
rect 54985 62087 55083 62185
rect 55847 62087 55945 62185
rect 56233 62087 56331 62185
rect 57095 62087 57193 62185
rect 57481 62087 57579 62185
rect 58343 62087 58441 62185
rect 58729 62087 58827 62185
rect 59591 62087 59689 62185
rect 59977 62087 60075 62185
rect 60839 62087 60937 62185
rect 61225 62087 61323 62185
rect 62087 62087 62185 62185
rect 62473 62087 62571 62185
rect 63335 62087 63433 62185
rect 63721 62087 63819 62185
rect 64583 62087 64681 62185
rect 64969 62087 65067 62185
rect 65831 62087 65929 62185
rect 66217 62087 66315 62185
rect 67079 62087 67177 62185
rect 67465 62087 67563 62185
rect 68327 62087 68425 62185
rect 68713 62087 68811 62185
rect 69575 62087 69673 62185
rect 69961 62087 70059 62185
rect 70823 62087 70921 62185
rect 71209 62087 71307 62185
rect 72071 62087 72169 62185
rect 72457 62087 72555 62185
rect 73319 62087 73417 62185
rect 73705 62087 73803 62185
rect 74567 62087 74665 62185
rect 74953 62087 75051 62185
rect 75815 62087 75913 62185
rect 76201 62087 76299 62185
rect 77063 62087 77161 62185
rect 77449 62087 77547 62185
rect 78311 62087 78409 62185
rect 78697 62087 78795 62185
rect 79559 62087 79657 62185
rect 79945 62087 80043 62185
rect 80807 62087 80905 62185
rect 81193 62087 81291 62185
rect 82055 62087 82153 62185
rect 82441 62087 82539 62185
rect 83303 62087 83401 62185
rect 83689 62087 83787 62185
rect 84551 62087 84649 62185
rect 84937 62087 85035 62185
rect 85799 62087 85897 62185
rect 86185 62087 86283 62185
rect 87047 62087 87145 62185
rect 87433 62087 87531 62185
rect 88295 62087 88393 62185
rect 88681 62087 88779 62185
rect 89543 62087 89641 62185
rect 89929 62087 90027 62185
rect 90791 62087 90889 62185
rect 91177 62087 91275 62185
rect 92039 62087 92137 62185
rect 92425 62087 92523 62185
rect 93287 62087 93385 62185
rect 93673 62087 93771 62185
rect 13296 61496 13394 61594
rect 13920 61496 14018 61594
rect 14544 61496 14642 61594
rect 15168 61496 15266 61594
rect 15792 61496 15890 61594
rect 16416 61496 16514 61594
rect 17040 61496 17138 61594
rect 17664 61496 17762 61594
rect 18288 61496 18386 61594
rect 18912 61496 19010 61594
rect 19536 61496 19634 61594
rect 20160 61496 20258 61594
rect 20784 61496 20882 61594
rect 21408 61496 21506 61594
rect 22032 61496 22130 61594
rect 22656 61496 22754 61594
rect 23280 61496 23378 61594
rect 23904 61496 24002 61594
rect 24528 61496 24626 61594
rect 25152 61496 25250 61594
rect 25776 61496 25874 61594
rect 26400 61496 26498 61594
rect 27024 61496 27122 61594
rect 27648 61496 27746 61594
rect 28272 61496 28370 61594
rect 28896 61496 28994 61594
rect 29520 61496 29618 61594
rect 30144 61496 30242 61594
rect 30768 61496 30866 61594
rect 31392 61496 31490 61594
rect 32016 61496 32114 61594
rect 32640 61496 32738 61594
rect 33264 61496 33362 61594
rect 33888 61496 33986 61594
rect 34512 61496 34610 61594
rect 35136 61496 35234 61594
rect 35760 61496 35858 61594
rect 36384 61496 36482 61594
rect 37008 61496 37106 61594
rect 37632 61496 37730 61594
rect 38256 61496 38354 61594
rect 38880 61496 38978 61594
rect 39504 61496 39602 61594
rect 40128 61496 40226 61594
rect 40752 61496 40850 61594
rect 41376 61496 41474 61594
rect 42000 61496 42098 61594
rect 42624 61496 42722 61594
rect 43248 61496 43346 61594
rect 43872 61496 43970 61594
rect 44496 61496 44594 61594
rect 45120 61496 45218 61594
rect 45744 61496 45842 61594
rect 46368 61496 46466 61594
rect 46992 61496 47090 61594
rect 47616 61496 47714 61594
rect 48240 61496 48338 61594
rect 48864 61496 48962 61594
rect 49488 61496 49586 61594
rect 50112 61496 50210 61594
rect 50736 61496 50834 61594
rect 51360 61496 51458 61594
rect 51984 61496 52082 61594
rect 52608 61496 52706 61594
rect 53232 61496 53330 61594
rect 53856 61496 53954 61594
rect 54480 61496 54578 61594
rect 55104 61496 55202 61594
rect 55728 61496 55826 61594
rect 56352 61496 56450 61594
rect 56976 61496 57074 61594
rect 57600 61496 57698 61594
rect 58224 61496 58322 61594
rect 58848 61496 58946 61594
rect 59472 61496 59570 61594
rect 60096 61496 60194 61594
rect 60720 61496 60818 61594
rect 61344 61496 61442 61594
rect 61968 61496 62066 61594
rect 62592 61496 62690 61594
rect 63216 61496 63314 61594
rect 63840 61496 63938 61594
rect 64464 61496 64562 61594
rect 65088 61496 65186 61594
rect 65712 61496 65810 61594
rect 66336 61496 66434 61594
rect 66960 61496 67058 61594
rect 67584 61496 67682 61594
rect 68208 61496 68306 61594
rect 68832 61496 68930 61594
rect 69456 61496 69554 61594
rect 70080 61496 70178 61594
rect 70704 61496 70802 61594
rect 71328 61496 71426 61594
rect 71952 61496 72050 61594
rect 72576 61496 72674 61594
rect 73200 61496 73298 61594
rect 73824 61496 73922 61594
rect 74448 61496 74546 61594
rect 75072 61496 75170 61594
rect 75696 61496 75794 61594
rect 76320 61496 76418 61594
rect 76944 61496 77042 61594
rect 77568 61496 77666 61594
rect 78192 61496 78290 61594
rect 78816 61496 78914 61594
rect 79440 61496 79538 61594
rect 80064 61496 80162 61594
rect 80688 61496 80786 61594
rect 81312 61496 81410 61594
rect 81936 61496 82034 61594
rect 82560 61496 82658 61594
rect 83184 61496 83282 61594
rect 83808 61496 83906 61594
rect 84432 61496 84530 61594
rect 85056 61496 85154 61594
rect 85680 61496 85778 61594
rect 86304 61496 86402 61594
rect 86928 61496 87026 61594
rect 87552 61496 87650 61594
rect 88176 61496 88274 61594
rect 88800 61496 88898 61594
rect 89424 61496 89522 61594
rect 90048 61496 90146 61594
rect 90672 61496 90770 61594
rect 91296 61496 91394 61594
rect 91920 61496 92018 61594
rect 92544 61496 92642 61594
rect 93168 61496 93266 61594
rect 93792 61496 93890 61594
rect 12234 61282 12332 61380
rect 94854 61282 94952 61380
rect 95880 61132 95978 61230
rect 98571 61120 98669 61218
rect 99403 61126 99501 61224
rect 12600 60935 12698 61033
rect 94488 60935 94586 61033
rect 12600 60698 12698 60796
rect 94488 60698 94586 60796
rect 6025 60563 6123 60661
rect 6450 60563 6548 60661
rect 6882 60563 6980 60661
rect 7264 60540 7362 60638
rect 7660 60540 7758 60638
rect 99428 60540 99526 60638
rect 99824 60540 99922 60638
rect 100206 60563 100304 60661
rect 100638 60563 100736 60661
rect 101063 60563 101161 60661
rect 12600 60382 12698 60480
rect 94488 60382 94586 60480
rect 6025 60189 6123 60287
rect 6450 60131 6548 60229
rect 6882 60131 6980 60229
rect 7264 60145 7362 60243
rect 7660 60145 7758 60243
rect 12600 60145 12698 60243
rect 94488 60145 94586 60243
rect 99428 60145 99526 60243
rect 99824 60145 99922 60243
rect 100206 60131 100304 60229
rect 100638 60131 100736 60229
rect 101063 60189 101161 60287
rect 12600 59908 12698 60006
rect 94488 59908 94586 60006
rect 6025 59773 6123 59871
rect 6450 59773 6548 59871
rect 6882 59773 6980 59871
rect 7264 59750 7362 59848
rect 7660 59750 7758 59848
rect 99428 59750 99526 59848
rect 99824 59750 99922 59848
rect 100206 59773 100304 59871
rect 100638 59773 100736 59871
rect 101063 59773 101161 59871
rect 12600 59592 12698 59690
rect 94488 59592 94586 59690
rect 6025 59399 6123 59497
rect 6450 59341 6548 59439
rect 6882 59341 6980 59439
rect 7264 59355 7362 59453
rect 7660 59355 7758 59453
rect 12600 59355 12698 59453
rect 94488 59355 94586 59453
rect 99428 59355 99526 59453
rect 99824 59355 99922 59453
rect 100206 59341 100304 59439
rect 100638 59341 100736 59439
rect 101063 59399 101161 59497
rect 12600 59118 12698 59216
rect 94488 59118 94586 59216
rect 6025 58983 6123 59081
rect 6450 58983 6548 59081
rect 6882 58983 6980 59081
rect 7264 58960 7362 59058
rect 7660 58960 7758 59058
rect 99428 58960 99526 59058
rect 99824 58960 99922 59058
rect 100206 58983 100304 59081
rect 100638 58983 100736 59081
rect 101063 58983 101161 59081
rect 12600 58802 12698 58900
rect 94488 58802 94586 58900
rect 6025 58609 6123 58707
rect 6450 58551 6548 58649
rect 6882 58551 6980 58649
rect 7264 58565 7362 58663
rect 7660 58565 7758 58663
rect 12600 58565 12698 58663
rect 94488 58565 94586 58663
rect 99428 58565 99526 58663
rect 99824 58565 99922 58663
rect 100206 58551 100304 58649
rect 100638 58551 100736 58649
rect 101063 58609 101161 58707
rect 12600 58328 12698 58426
rect 94488 58328 94586 58426
rect 6025 58193 6123 58291
rect 6450 58193 6548 58291
rect 6882 58193 6980 58291
rect 7264 58170 7362 58268
rect 7660 58170 7758 58268
rect 99428 58170 99526 58268
rect 99824 58170 99922 58268
rect 100206 58193 100304 58291
rect 100638 58193 100736 58291
rect 101063 58193 101161 58291
rect 12600 58012 12698 58110
rect 94488 58012 94586 58110
rect 6025 57819 6123 57917
rect 6450 57761 6548 57859
rect 6882 57761 6980 57859
rect 7264 57775 7362 57873
rect 7660 57775 7758 57873
rect 12600 57775 12698 57873
rect 94488 57775 94586 57873
rect 99428 57775 99526 57873
rect 99824 57775 99922 57873
rect 100206 57761 100304 57859
rect 100638 57761 100736 57859
rect 101063 57819 101161 57917
rect 12600 57538 12698 57636
rect 94488 57538 94586 57636
rect 6025 57403 6123 57501
rect 6450 57403 6548 57501
rect 6882 57403 6980 57501
rect 7264 57380 7362 57478
rect 7660 57380 7758 57478
rect 99428 57380 99526 57478
rect 99824 57380 99922 57478
rect 100206 57403 100304 57501
rect 100638 57403 100736 57501
rect 101063 57403 101161 57501
rect 12600 57222 12698 57320
rect 94488 57222 94586 57320
rect 6025 57029 6123 57127
rect 6450 56971 6548 57069
rect 6882 56971 6980 57069
rect 7264 56985 7362 57083
rect 7660 56985 7758 57083
rect 12600 56985 12698 57083
rect 94488 56985 94586 57083
rect 99428 56985 99526 57083
rect 99824 56985 99922 57083
rect 100206 56971 100304 57069
rect 100638 56971 100736 57069
rect 101063 57029 101161 57127
rect 12600 56748 12698 56846
rect 94488 56748 94586 56846
rect 6025 56613 6123 56711
rect 6450 56613 6548 56711
rect 6882 56613 6980 56711
rect 7264 56590 7362 56688
rect 7660 56590 7758 56688
rect 99428 56590 99526 56688
rect 99824 56590 99922 56688
rect 100206 56613 100304 56711
rect 100638 56613 100736 56711
rect 101063 56613 101161 56711
rect 12600 56432 12698 56530
rect 94488 56432 94586 56530
rect 6025 56239 6123 56337
rect 6450 56181 6548 56279
rect 6882 56181 6980 56279
rect 7264 56195 7362 56293
rect 7660 56195 7758 56293
rect 12600 56195 12698 56293
rect 94488 56195 94586 56293
rect 99428 56195 99526 56293
rect 99824 56195 99922 56293
rect 100206 56181 100304 56279
rect 100638 56181 100736 56279
rect 101063 56239 101161 56337
rect 12600 55958 12698 56056
rect 94488 55958 94586 56056
rect 6025 55823 6123 55921
rect 6450 55823 6548 55921
rect 6882 55823 6980 55921
rect 7264 55800 7362 55898
rect 7660 55800 7758 55898
rect 99428 55800 99526 55898
rect 99824 55800 99922 55898
rect 100206 55823 100304 55921
rect 100638 55823 100736 55921
rect 101063 55823 101161 55921
rect 12600 55642 12698 55740
rect 94488 55642 94586 55740
rect 6025 55449 6123 55547
rect 6450 55391 6548 55489
rect 6882 55391 6980 55489
rect 7264 55405 7362 55503
rect 7660 55405 7758 55503
rect 12600 55405 12698 55503
rect 94488 55405 94586 55503
rect 99428 55405 99526 55503
rect 99824 55405 99922 55503
rect 100206 55391 100304 55489
rect 100638 55391 100736 55489
rect 101063 55449 101161 55547
rect 12600 55168 12698 55266
rect 94488 55168 94586 55266
rect 6025 55033 6123 55131
rect 6450 55033 6548 55131
rect 6882 55033 6980 55131
rect 7264 55010 7362 55108
rect 7660 55010 7758 55108
rect 99428 55010 99526 55108
rect 99824 55010 99922 55108
rect 100206 55033 100304 55131
rect 100638 55033 100736 55131
rect 101063 55033 101161 55131
rect 12600 54852 12698 54950
rect 94488 54852 94586 54950
rect 6025 54659 6123 54757
rect 6450 54601 6548 54699
rect 6882 54601 6980 54699
rect 7264 54615 7362 54713
rect 7660 54615 7758 54713
rect 12600 54615 12698 54713
rect 94488 54615 94586 54713
rect 99428 54615 99526 54713
rect 99824 54615 99922 54713
rect 100206 54601 100304 54699
rect 100638 54601 100736 54699
rect 101063 54659 101161 54757
rect 12600 54378 12698 54476
rect 94488 54378 94586 54476
rect 6025 54243 6123 54341
rect 6450 54243 6548 54341
rect 6882 54243 6980 54341
rect 7264 54220 7362 54318
rect 7660 54220 7758 54318
rect 99428 54220 99526 54318
rect 99824 54220 99922 54318
rect 100206 54243 100304 54341
rect 100638 54243 100736 54341
rect 101063 54243 101161 54341
rect 12600 54062 12698 54160
rect 94488 54062 94586 54160
rect 6025 53869 6123 53967
rect 6450 53811 6548 53909
rect 6882 53811 6980 53909
rect 7264 53825 7362 53923
rect 7660 53825 7758 53923
rect 12600 53825 12698 53923
rect 94488 53825 94586 53923
rect 99428 53825 99526 53923
rect 99824 53825 99922 53923
rect 100206 53811 100304 53909
rect 100638 53811 100736 53909
rect 101063 53869 101161 53967
rect 12600 53588 12698 53686
rect 94488 53588 94586 53686
rect 6025 53453 6123 53551
rect 6450 53453 6548 53551
rect 6882 53453 6980 53551
rect 7264 53430 7362 53528
rect 7660 53430 7758 53528
rect 99428 53430 99526 53528
rect 99824 53430 99922 53528
rect 100206 53453 100304 53551
rect 100638 53453 100736 53551
rect 101063 53453 101161 53551
rect 12600 53272 12698 53370
rect 94488 53272 94586 53370
rect 6025 53079 6123 53177
rect 6450 53021 6548 53119
rect 6882 53021 6980 53119
rect 7264 53035 7362 53133
rect 7660 53035 7758 53133
rect 12600 53035 12698 53133
rect 94488 53035 94586 53133
rect 99428 53035 99526 53133
rect 99824 53035 99922 53133
rect 100206 53021 100304 53119
rect 100638 53021 100736 53119
rect 101063 53079 101161 53177
rect 12600 52798 12698 52896
rect 94488 52798 94586 52896
rect 6025 52663 6123 52761
rect 6450 52663 6548 52761
rect 6882 52663 6980 52761
rect 7264 52640 7362 52738
rect 7660 52640 7758 52738
rect 99428 52640 99526 52738
rect 99824 52640 99922 52738
rect 100206 52663 100304 52761
rect 100638 52663 100736 52761
rect 101063 52663 101161 52761
rect 12600 52482 12698 52580
rect 94488 52482 94586 52580
rect 6025 52289 6123 52387
rect 6450 52231 6548 52329
rect 6882 52231 6980 52329
rect 7264 52245 7362 52343
rect 7660 52245 7758 52343
rect 12600 52245 12698 52343
rect 94488 52245 94586 52343
rect 99428 52245 99526 52343
rect 99824 52245 99922 52343
rect 100206 52231 100304 52329
rect 100638 52231 100736 52329
rect 101063 52289 101161 52387
rect 12600 52008 12698 52106
rect 94488 52008 94586 52106
rect 6025 51873 6123 51971
rect 6450 51873 6548 51971
rect 6882 51873 6980 51971
rect 7264 51850 7362 51948
rect 7660 51850 7758 51948
rect 99428 51850 99526 51948
rect 99824 51850 99922 51948
rect 100206 51873 100304 51971
rect 100638 51873 100736 51971
rect 101063 51873 101161 51971
rect 12600 51692 12698 51790
rect 94488 51692 94586 51790
rect 6025 51499 6123 51597
rect 6450 51441 6548 51539
rect 6882 51441 6980 51539
rect 7264 51455 7362 51553
rect 7660 51455 7758 51553
rect 12600 51455 12698 51553
rect 94488 51455 94586 51553
rect 99428 51455 99526 51553
rect 99824 51455 99922 51553
rect 100206 51441 100304 51539
rect 100638 51441 100736 51539
rect 101063 51499 101161 51597
rect 12600 51218 12698 51316
rect 94488 51218 94586 51316
rect 6025 51083 6123 51181
rect 6450 51083 6548 51181
rect 6882 51083 6980 51181
rect 7264 51060 7362 51158
rect 7660 51060 7758 51158
rect 99428 51060 99526 51158
rect 99824 51060 99922 51158
rect 100206 51083 100304 51181
rect 100638 51083 100736 51181
rect 101063 51083 101161 51181
rect 12600 50902 12698 51000
rect 94488 50902 94586 51000
rect 6025 50709 6123 50807
rect 6450 50651 6548 50749
rect 6882 50651 6980 50749
rect 7264 50665 7362 50763
rect 7660 50665 7758 50763
rect 12600 50665 12698 50763
rect 94488 50665 94586 50763
rect 99428 50665 99526 50763
rect 99824 50665 99922 50763
rect 100206 50651 100304 50749
rect 100638 50651 100736 50749
rect 101063 50709 101161 50807
rect 12600 50428 12698 50526
rect 94488 50428 94586 50526
rect 6025 50293 6123 50391
rect 6450 50293 6548 50391
rect 6882 50293 6980 50391
rect 7264 50270 7362 50368
rect 7660 50270 7758 50368
rect 99428 50270 99526 50368
rect 99824 50270 99922 50368
rect 100206 50293 100304 50391
rect 100638 50293 100736 50391
rect 101063 50293 101161 50391
rect 12600 50112 12698 50210
rect 94488 50112 94586 50210
rect 6025 49919 6123 50017
rect 6450 49861 6548 49959
rect 6882 49861 6980 49959
rect 7264 49875 7362 49973
rect 7660 49875 7758 49973
rect 12600 49875 12698 49973
rect 94488 49875 94586 49973
rect 99428 49875 99526 49973
rect 99824 49875 99922 49973
rect 100206 49861 100304 49959
rect 100638 49861 100736 49959
rect 101063 49919 101161 50017
rect 12600 49638 12698 49736
rect 94488 49638 94586 49736
rect 6025 49503 6123 49601
rect 6450 49503 6548 49601
rect 6882 49503 6980 49601
rect 7264 49480 7362 49578
rect 7660 49480 7758 49578
rect 99428 49480 99526 49578
rect 99824 49480 99922 49578
rect 100206 49503 100304 49601
rect 100638 49503 100736 49601
rect 101063 49503 101161 49601
rect 12600 49322 12698 49420
rect 94488 49322 94586 49420
rect 6025 49129 6123 49227
rect 6450 49071 6548 49169
rect 6882 49071 6980 49169
rect 7264 49085 7362 49183
rect 7660 49085 7758 49183
rect 12600 49085 12698 49183
rect 94488 49085 94586 49183
rect 99428 49085 99526 49183
rect 99824 49085 99922 49183
rect 100206 49071 100304 49169
rect 100638 49071 100736 49169
rect 101063 49129 101161 49227
rect 12600 48848 12698 48946
rect 94488 48848 94586 48946
rect 6025 48713 6123 48811
rect 6450 48713 6548 48811
rect 6882 48713 6980 48811
rect 7264 48690 7362 48788
rect 7660 48690 7758 48788
rect 99428 48690 99526 48788
rect 99824 48690 99922 48788
rect 100206 48713 100304 48811
rect 100638 48713 100736 48811
rect 101063 48713 101161 48811
rect 12600 48532 12698 48630
rect 94488 48532 94586 48630
rect 6025 48339 6123 48437
rect 6450 48281 6548 48379
rect 6882 48281 6980 48379
rect 7264 48295 7362 48393
rect 7660 48295 7758 48393
rect 12600 48295 12698 48393
rect 94488 48295 94586 48393
rect 99428 48295 99526 48393
rect 99824 48295 99922 48393
rect 100206 48281 100304 48379
rect 100638 48281 100736 48379
rect 101063 48339 101161 48437
rect 12600 48058 12698 48156
rect 94488 48058 94586 48156
rect 6025 47923 6123 48021
rect 6450 47923 6548 48021
rect 6882 47923 6980 48021
rect 7264 47900 7362 47998
rect 7660 47900 7758 47998
rect 99428 47900 99526 47998
rect 99824 47900 99922 47998
rect 100206 47923 100304 48021
rect 100638 47923 100736 48021
rect 101063 47923 101161 48021
rect 12600 47742 12698 47840
rect 94488 47742 94586 47840
rect 6025 47549 6123 47647
rect 6450 47491 6548 47589
rect 6882 47491 6980 47589
rect 7264 47505 7362 47603
rect 7660 47505 7758 47603
rect 12600 47505 12698 47603
rect 94488 47505 94586 47603
rect 99428 47505 99526 47603
rect 99824 47505 99922 47603
rect 100206 47491 100304 47589
rect 100638 47491 100736 47589
rect 101063 47549 101161 47647
rect 12600 47268 12698 47366
rect 94488 47268 94586 47366
rect 6025 47133 6123 47231
rect 6450 47133 6548 47231
rect 6882 47133 6980 47231
rect 7264 47110 7362 47208
rect 7660 47110 7758 47208
rect 99428 47110 99526 47208
rect 99824 47110 99922 47208
rect 100206 47133 100304 47231
rect 100638 47133 100736 47231
rect 101063 47133 101161 47231
rect 12600 46952 12698 47050
rect 94488 46952 94586 47050
rect 6025 46759 6123 46857
rect 6450 46701 6548 46799
rect 6882 46701 6980 46799
rect 7264 46715 7362 46813
rect 7660 46715 7758 46813
rect 12600 46715 12698 46813
rect 94488 46715 94586 46813
rect 99428 46715 99526 46813
rect 99824 46715 99922 46813
rect 100206 46701 100304 46799
rect 100638 46701 100736 46799
rect 101063 46759 101161 46857
rect 12600 46478 12698 46576
rect 94488 46478 94586 46576
rect 6025 46343 6123 46441
rect 6450 46343 6548 46441
rect 6882 46343 6980 46441
rect 7264 46320 7362 46418
rect 7660 46320 7758 46418
rect 99428 46320 99526 46418
rect 99824 46320 99922 46418
rect 100206 46343 100304 46441
rect 100638 46343 100736 46441
rect 101063 46343 101161 46441
rect 12600 46162 12698 46260
rect 94488 46162 94586 46260
rect 6025 45969 6123 46067
rect 6450 45911 6548 46009
rect 6882 45911 6980 46009
rect 7264 45925 7362 46023
rect 7660 45925 7758 46023
rect 12600 45925 12698 46023
rect 94488 45925 94586 46023
rect 99428 45925 99526 46023
rect 99824 45925 99922 46023
rect 100206 45911 100304 46009
rect 100638 45911 100736 46009
rect 101063 45969 101161 46067
rect 12600 45688 12698 45786
rect 94488 45688 94586 45786
rect 6025 45553 6123 45651
rect 6450 45553 6548 45651
rect 6882 45553 6980 45651
rect 7264 45530 7362 45628
rect 7660 45530 7758 45628
rect 99428 45530 99526 45628
rect 99824 45530 99922 45628
rect 100206 45553 100304 45651
rect 100638 45553 100736 45651
rect 101063 45553 101161 45651
rect 12600 45372 12698 45470
rect 94488 45372 94586 45470
rect 6025 45179 6123 45277
rect 6450 45121 6548 45219
rect 6882 45121 6980 45219
rect 7264 45135 7362 45233
rect 7660 45135 7758 45233
rect 12600 45135 12698 45233
rect 94488 45135 94586 45233
rect 99428 45135 99526 45233
rect 99824 45135 99922 45233
rect 100206 45121 100304 45219
rect 100638 45121 100736 45219
rect 101063 45179 101161 45277
rect 12600 44898 12698 44996
rect 94488 44898 94586 44996
rect 6025 44763 6123 44861
rect 6450 44763 6548 44861
rect 6882 44763 6980 44861
rect 7264 44740 7362 44838
rect 7660 44740 7758 44838
rect 99428 44740 99526 44838
rect 99824 44740 99922 44838
rect 100206 44763 100304 44861
rect 100638 44763 100736 44861
rect 101063 44763 101161 44861
rect 12600 44582 12698 44680
rect 94488 44582 94586 44680
rect 6025 44389 6123 44487
rect 6450 44331 6548 44429
rect 6882 44331 6980 44429
rect 7264 44345 7362 44443
rect 7660 44345 7758 44443
rect 12600 44345 12698 44443
rect 94488 44345 94586 44443
rect 99428 44345 99526 44443
rect 99824 44345 99922 44443
rect 100206 44331 100304 44429
rect 100638 44331 100736 44429
rect 101063 44389 101161 44487
rect 12600 44108 12698 44206
rect 94488 44108 94586 44206
rect 6025 43973 6123 44071
rect 6450 43973 6548 44071
rect 6882 43973 6980 44071
rect 7264 43950 7362 44048
rect 7660 43950 7758 44048
rect 99428 43950 99526 44048
rect 99824 43950 99922 44048
rect 100206 43973 100304 44071
rect 100638 43973 100736 44071
rect 101063 43973 101161 44071
rect 12600 43792 12698 43890
rect 94488 43792 94586 43890
rect 6025 43599 6123 43697
rect 6450 43541 6548 43639
rect 6882 43541 6980 43639
rect 7264 43555 7362 43653
rect 7660 43555 7758 43653
rect 12600 43555 12698 43653
rect 94488 43555 94586 43653
rect 99428 43555 99526 43653
rect 99824 43555 99922 43653
rect 100206 43541 100304 43639
rect 100638 43541 100736 43639
rect 101063 43599 101161 43697
rect 12600 43318 12698 43416
rect 94488 43318 94586 43416
rect 6025 43183 6123 43281
rect 6450 43183 6548 43281
rect 6882 43183 6980 43281
rect 7264 43160 7362 43258
rect 7660 43160 7758 43258
rect 99428 43160 99526 43258
rect 99824 43160 99922 43258
rect 100206 43183 100304 43281
rect 100638 43183 100736 43281
rect 101063 43183 101161 43281
rect 12600 43002 12698 43100
rect 94488 43002 94586 43100
rect 6025 42809 6123 42907
rect 6450 42751 6548 42849
rect 6882 42751 6980 42849
rect 7264 42765 7362 42863
rect 7660 42765 7758 42863
rect 12600 42765 12698 42863
rect 94488 42765 94586 42863
rect 99428 42765 99526 42863
rect 99824 42765 99922 42863
rect 100206 42751 100304 42849
rect 100638 42751 100736 42849
rect 101063 42809 101161 42907
rect 12600 42528 12698 42626
rect 94488 42528 94586 42626
rect 6025 42393 6123 42491
rect 6450 42393 6548 42491
rect 6882 42393 6980 42491
rect 7264 42370 7362 42468
rect 7660 42370 7758 42468
rect 99428 42370 99526 42468
rect 99824 42370 99922 42468
rect 100206 42393 100304 42491
rect 100638 42393 100736 42491
rect 101063 42393 101161 42491
rect 12600 42212 12698 42310
rect 94488 42212 94586 42310
rect 6025 42019 6123 42117
rect 6450 41961 6548 42059
rect 6882 41961 6980 42059
rect 7264 41975 7362 42073
rect 7660 41975 7758 42073
rect 12600 41975 12698 42073
rect 94488 41975 94586 42073
rect 99428 41975 99526 42073
rect 99824 41975 99922 42073
rect 100206 41961 100304 42059
rect 100638 41961 100736 42059
rect 101063 42019 101161 42117
rect 12600 41738 12698 41836
rect 94488 41738 94586 41836
rect 6025 41603 6123 41701
rect 6450 41603 6548 41701
rect 6882 41603 6980 41701
rect 7264 41580 7362 41678
rect 7660 41580 7758 41678
rect 99428 41580 99526 41678
rect 99824 41580 99922 41678
rect 100206 41603 100304 41701
rect 100638 41603 100736 41701
rect 101063 41603 101161 41701
rect 12600 41422 12698 41520
rect 94488 41422 94586 41520
rect 6025 41229 6123 41327
rect 6450 41171 6548 41269
rect 6882 41171 6980 41269
rect 7264 41185 7362 41283
rect 7660 41185 7758 41283
rect 12600 41185 12698 41283
rect 94488 41185 94586 41283
rect 99428 41185 99526 41283
rect 99824 41185 99922 41283
rect 100206 41171 100304 41269
rect 100638 41171 100736 41269
rect 101063 41229 101161 41327
rect 12600 40948 12698 41046
rect 94488 40948 94586 41046
rect 6025 40813 6123 40911
rect 6450 40813 6548 40911
rect 6882 40813 6980 40911
rect 7264 40790 7362 40888
rect 7660 40790 7758 40888
rect 99428 40790 99526 40888
rect 99824 40790 99922 40888
rect 100206 40813 100304 40911
rect 100638 40813 100736 40911
rect 101063 40813 101161 40911
rect 12600 40632 12698 40730
rect 94488 40632 94586 40730
rect 6025 40439 6123 40537
rect 6450 40381 6548 40479
rect 6882 40381 6980 40479
rect 7264 40395 7362 40493
rect 7660 40395 7758 40493
rect 12600 40395 12698 40493
rect 94488 40395 94586 40493
rect 99428 40395 99526 40493
rect 99824 40395 99922 40493
rect 100206 40381 100304 40479
rect 100638 40381 100736 40479
rect 101063 40439 101161 40537
rect 12600 40158 12698 40256
rect 94488 40158 94586 40256
rect 6025 40023 6123 40121
rect 6450 40023 6548 40121
rect 6882 40023 6980 40121
rect 7264 40000 7362 40098
rect 7660 40000 7758 40098
rect 99428 40000 99526 40098
rect 99824 40000 99922 40098
rect 100206 40023 100304 40121
rect 100638 40023 100736 40121
rect 101063 40023 101161 40121
rect 12600 39842 12698 39940
rect 94488 39842 94586 39940
rect 6025 39649 6123 39747
rect 6450 39591 6548 39689
rect 6882 39591 6980 39689
rect 7264 39605 7362 39703
rect 7660 39605 7758 39703
rect 12600 39605 12698 39703
rect 94488 39605 94586 39703
rect 99428 39605 99526 39703
rect 99824 39605 99922 39703
rect 100206 39591 100304 39689
rect 100638 39591 100736 39689
rect 101063 39649 101161 39747
rect 12600 39368 12698 39466
rect 94488 39368 94586 39466
rect 6025 39233 6123 39331
rect 6450 39233 6548 39331
rect 6882 39233 6980 39331
rect 7264 39210 7362 39308
rect 7660 39210 7758 39308
rect 99428 39210 99526 39308
rect 99824 39210 99922 39308
rect 100206 39233 100304 39331
rect 100638 39233 100736 39331
rect 101063 39233 101161 39331
rect 12600 39052 12698 39150
rect 94488 39052 94586 39150
rect 6025 38859 6123 38957
rect 6450 38801 6548 38899
rect 6882 38801 6980 38899
rect 7264 38815 7362 38913
rect 7660 38815 7758 38913
rect 12600 38815 12698 38913
rect 94488 38815 94586 38913
rect 99428 38815 99526 38913
rect 99824 38815 99922 38913
rect 100206 38801 100304 38899
rect 100638 38801 100736 38899
rect 101063 38859 101161 38957
rect 12600 38578 12698 38676
rect 94488 38578 94586 38676
rect 6025 38443 6123 38541
rect 6450 38443 6548 38541
rect 6882 38443 6980 38541
rect 7264 38420 7362 38518
rect 7660 38420 7758 38518
rect 99428 38420 99526 38518
rect 99824 38420 99922 38518
rect 100206 38443 100304 38541
rect 100638 38443 100736 38541
rect 101063 38443 101161 38541
rect 12600 38262 12698 38360
rect 94488 38262 94586 38360
rect 6025 38069 6123 38167
rect 6450 38011 6548 38109
rect 6882 38011 6980 38109
rect 7264 38025 7362 38123
rect 7660 38025 7758 38123
rect 12600 38025 12698 38123
rect 94488 38025 94586 38123
rect 99428 38025 99526 38123
rect 99824 38025 99922 38123
rect 100206 38011 100304 38109
rect 100638 38011 100736 38109
rect 101063 38069 101161 38167
rect 12600 37788 12698 37886
rect 94488 37788 94586 37886
rect 6025 37653 6123 37751
rect 6450 37653 6548 37751
rect 6882 37653 6980 37751
rect 7264 37630 7362 37728
rect 7660 37630 7758 37728
rect 99428 37630 99526 37728
rect 99824 37630 99922 37728
rect 100206 37653 100304 37751
rect 100638 37653 100736 37751
rect 101063 37653 101161 37751
rect 12600 37472 12698 37570
rect 94488 37472 94586 37570
rect 6025 37279 6123 37377
rect 6450 37221 6548 37319
rect 6882 37221 6980 37319
rect 7264 37235 7362 37333
rect 7660 37235 7758 37333
rect 12600 37235 12698 37333
rect 94488 37235 94586 37333
rect 99428 37235 99526 37333
rect 99824 37235 99922 37333
rect 100206 37221 100304 37319
rect 100638 37221 100736 37319
rect 101063 37279 101161 37377
rect 12600 36998 12698 37096
rect 94488 36998 94586 37096
rect 6025 36863 6123 36961
rect 6450 36863 6548 36961
rect 6882 36863 6980 36961
rect 7264 36840 7362 36938
rect 7660 36840 7758 36938
rect 99428 36840 99526 36938
rect 99824 36840 99922 36938
rect 100206 36863 100304 36961
rect 100638 36863 100736 36961
rect 101063 36863 101161 36961
rect 12600 36682 12698 36780
rect 94488 36682 94586 36780
rect 6025 36489 6123 36587
rect 6450 36431 6548 36529
rect 6882 36431 6980 36529
rect 7264 36445 7362 36543
rect 7660 36445 7758 36543
rect 12600 36445 12698 36543
rect 94488 36445 94586 36543
rect 99428 36445 99526 36543
rect 99824 36445 99922 36543
rect 100206 36431 100304 36529
rect 100638 36431 100736 36529
rect 101063 36489 101161 36587
rect 12600 36208 12698 36306
rect 94488 36208 94586 36306
rect 6025 36073 6123 36171
rect 6450 36073 6548 36171
rect 6882 36073 6980 36171
rect 7264 36050 7362 36148
rect 7660 36050 7758 36148
rect 99428 36050 99526 36148
rect 99824 36050 99922 36148
rect 100206 36073 100304 36171
rect 100638 36073 100736 36171
rect 101063 36073 101161 36171
rect 12600 35892 12698 35990
rect 94488 35892 94586 35990
rect 6025 35699 6123 35797
rect 6450 35641 6548 35739
rect 6882 35641 6980 35739
rect 7264 35655 7362 35753
rect 7660 35655 7758 35753
rect 8092 35640 8190 35738
rect 8517 35639 8615 35737
rect 9560 35655 9658 35753
rect 11208 35655 11306 35753
rect 12600 35655 12698 35753
rect 94488 35655 94586 35753
rect 95880 35655 95978 35753
rect 97528 35655 97626 35753
rect 98571 35639 98669 35737
rect 98996 35640 99094 35738
rect 99428 35655 99526 35753
rect 99824 35655 99922 35753
rect 100206 35641 100304 35739
rect 100638 35641 100736 35739
rect 101063 35699 101161 35797
rect 12600 35418 12698 35516
rect 94488 35418 94586 35516
rect 6025 35283 6123 35381
rect 6450 35283 6548 35381
rect 6882 35283 6980 35381
rect 7264 35260 7362 35358
rect 7660 35260 7758 35358
rect 99428 35260 99526 35358
rect 99824 35260 99922 35358
rect 100206 35283 100304 35381
rect 100638 35283 100736 35381
rect 101063 35283 101161 35381
rect 12600 35102 12698 35200
rect 94488 35102 94586 35200
rect 6025 34909 6123 35007
rect 6450 34851 6548 34949
rect 6882 34851 6980 34949
rect 7264 34865 7362 34963
rect 7660 34865 7758 34963
rect 12600 34865 12698 34963
rect 94488 34865 94586 34963
rect 99428 34865 99526 34963
rect 99824 34865 99922 34963
rect 100206 34851 100304 34949
rect 100638 34851 100736 34949
rect 101063 34909 101161 35007
rect 12600 34628 12698 34726
rect 94488 34628 94586 34726
rect 6025 34493 6123 34591
rect 6450 34493 6548 34591
rect 6882 34493 6980 34591
rect 7264 34470 7362 34568
rect 7660 34470 7758 34568
rect 99428 34470 99526 34568
rect 99824 34470 99922 34568
rect 100206 34493 100304 34591
rect 100638 34493 100736 34591
rect 101063 34493 101161 34591
rect 12600 34312 12698 34410
rect 94488 34312 94586 34410
rect 6025 34119 6123 34217
rect 6450 34061 6548 34159
rect 6882 34061 6980 34159
rect 7264 34075 7362 34173
rect 7660 34075 7758 34173
rect 12600 34075 12698 34173
rect 94488 34075 94586 34173
rect 99428 34075 99526 34173
rect 99824 34075 99922 34173
rect 100206 34061 100304 34159
rect 100638 34061 100736 34159
rect 101063 34119 101161 34217
rect 12600 33838 12698 33936
rect 94488 33838 94586 33936
rect 6025 33703 6123 33801
rect 6450 33703 6548 33801
rect 6882 33703 6980 33801
rect 7264 33680 7362 33778
rect 7660 33680 7758 33778
rect 99428 33680 99526 33778
rect 99824 33680 99922 33778
rect 100206 33703 100304 33801
rect 100638 33703 100736 33801
rect 101063 33703 101161 33801
rect 12600 33522 12698 33620
rect 94488 33522 94586 33620
rect 6025 33329 6123 33427
rect 6450 33271 6548 33369
rect 6882 33271 6980 33369
rect 7264 33285 7362 33383
rect 7660 33285 7758 33383
rect 12600 33285 12698 33383
rect 94488 33285 94586 33383
rect 99428 33285 99526 33383
rect 99824 33285 99922 33383
rect 100206 33271 100304 33369
rect 100638 33271 100736 33369
rect 101063 33329 101161 33427
rect 12600 33048 12698 33146
rect 94488 33048 94586 33146
rect 6025 32913 6123 33011
rect 6450 32913 6548 33011
rect 6882 32913 6980 33011
rect 7264 32890 7362 32988
rect 7660 32890 7758 32988
rect 99428 32890 99526 32988
rect 99824 32890 99922 32988
rect 100206 32913 100304 33011
rect 100638 32913 100736 33011
rect 101063 32913 101161 33011
rect 12600 32732 12698 32830
rect 94488 32732 94586 32830
rect 6025 32539 6123 32637
rect 6450 32481 6548 32579
rect 6882 32481 6980 32579
rect 7264 32495 7362 32593
rect 7660 32495 7758 32593
rect 12600 32495 12698 32593
rect 94488 32495 94586 32593
rect 99428 32495 99526 32593
rect 99824 32495 99922 32593
rect 100206 32481 100304 32579
rect 100638 32481 100736 32579
rect 101063 32539 101161 32637
rect 12600 32258 12698 32356
rect 94488 32258 94586 32356
rect 6025 32123 6123 32221
rect 6450 32123 6548 32221
rect 6882 32123 6980 32221
rect 7264 32100 7362 32198
rect 7660 32100 7758 32198
rect 99428 32100 99526 32198
rect 99824 32100 99922 32198
rect 100206 32123 100304 32221
rect 100638 32123 100736 32221
rect 101063 32123 101161 32221
rect 12600 31942 12698 32040
rect 94488 31942 94586 32040
rect 6025 31749 6123 31847
rect 6450 31691 6548 31789
rect 6882 31691 6980 31789
rect 7264 31705 7362 31803
rect 7660 31705 7758 31803
rect 12600 31705 12698 31803
rect 94488 31705 94586 31803
rect 99428 31705 99526 31803
rect 99824 31705 99922 31803
rect 100206 31691 100304 31789
rect 100638 31691 100736 31789
rect 101063 31749 101161 31847
rect 12600 31468 12698 31566
rect 94488 31468 94586 31566
rect 6025 31333 6123 31431
rect 6450 31333 6548 31431
rect 6882 31333 6980 31431
rect 7264 31310 7362 31408
rect 7660 31310 7758 31408
rect 99428 31310 99526 31408
rect 99824 31310 99922 31408
rect 100206 31333 100304 31431
rect 100638 31333 100736 31431
rect 101063 31333 101161 31431
rect 12600 31152 12698 31250
rect 94488 31152 94586 31250
rect 6025 30959 6123 31057
rect 6450 30901 6548 30999
rect 6882 30901 6980 30999
rect 7264 30915 7362 31013
rect 7660 30915 7758 31013
rect 12600 30915 12698 31013
rect 94488 30915 94586 31013
rect 99428 30915 99526 31013
rect 99824 30915 99922 31013
rect 100206 30901 100304 30999
rect 100638 30901 100736 30999
rect 101063 30959 101161 31057
rect 12600 30678 12698 30776
rect 94488 30678 94586 30776
rect 6025 30543 6123 30641
rect 6450 30543 6548 30641
rect 6882 30543 6980 30641
rect 7264 30520 7362 30618
rect 7660 30520 7758 30618
rect 99428 30520 99526 30618
rect 99824 30520 99922 30618
rect 100206 30543 100304 30641
rect 100638 30543 100736 30641
rect 101063 30543 101161 30641
rect 12600 30362 12698 30460
rect 94488 30362 94586 30460
rect 6025 30169 6123 30267
rect 6450 30111 6548 30209
rect 6882 30111 6980 30209
rect 7264 30125 7362 30223
rect 7660 30125 7758 30223
rect 12600 30125 12698 30223
rect 94488 30125 94586 30223
rect 99428 30125 99526 30223
rect 99824 30125 99922 30223
rect 100206 30111 100304 30209
rect 100638 30111 100736 30209
rect 101063 30169 101161 30267
rect 12600 29888 12698 29986
rect 94488 29888 94586 29986
rect 6025 29753 6123 29851
rect 6450 29753 6548 29851
rect 6882 29753 6980 29851
rect 7264 29730 7362 29828
rect 7660 29730 7758 29828
rect 99428 29730 99526 29828
rect 99824 29730 99922 29828
rect 100206 29753 100304 29851
rect 100638 29753 100736 29851
rect 101063 29753 101161 29851
rect 12600 29572 12698 29670
rect 94488 29572 94586 29670
rect 6025 29379 6123 29477
rect 6450 29321 6548 29419
rect 6882 29321 6980 29419
rect 7264 29335 7362 29433
rect 7660 29335 7758 29433
rect 12600 29335 12698 29433
rect 94488 29335 94586 29433
rect 99428 29335 99526 29433
rect 99824 29335 99922 29433
rect 100206 29321 100304 29419
rect 100638 29321 100736 29419
rect 101063 29379 101161 29477
rect 12600 29098 12698 29196
rect 94488 29098 94586 29196
rect 6025 28963 6123 29061
rect 6450 28963 6548 29061
rect 6882 28963 6980 29061
rect 7264 28940 7362 29038
rect 7660 28940 7758 29038
rect 99428 28940 99526 29038
rect 99824 28940 99922 29038
rect 100206 28963 100304 29061
rect 100638 28963 100736 29061
rect 101063 28963 101161 29061
rect 12600 28782 12698 28880
rect 94488 28782 94586 28880
rect 6025 28589 6123 28687
rect 6450 28531 6548 28629
rect 6882 28531 6980 28629
rect 7264 28545 7362 28643
rect 7660 28545 7758 28643
rect 12600 28545 12698 28643
rect 94488 28545 94586 28643
rect 99428 28545 99526 28643
rect 99824 28545 99922 28643
rect 100206 28531 100304 28629
rect 100638 28531 100736 28629
rect 101063 28589 101161 28687
rect 12600 28308 12698 28406
rect 94488 28308 94586 28406
rect 6025 28173 6123 28271
rect 6450 28173 6548 28271
rect 6882 28173 6980 28271
rect 7264 28150 7362 28248
rect 7660 28150 7758 28248
rect 99428 28150 99526 28248
rect 99824 28150 99922 28248
rect 100206 28173 100304 28271
rect 100638 28173 100736 28271
rect 101063 28173 101161 28271
rect 12600 27992 12698 28090
rect 94488 27992 94586 28090
rect 6025 27799 6123 27897
rect 6450 27741 6548 27839
rect 6882 27741 6980 27839
rect 7264 27755 7362 27853
rect 7660 27755 7758 27853
rect 12600 27755 12698 27853
rect 94488 27755 94586 27853
rect 99428 27755 99526 27853
rect 99824 27755 99922 27853
rect 100206 27741 100304 27839
rect 100638 27741 100736 27839
rect 101063 27799 101161 27897
rect 12600 27518 12698 27616
rect 94488 27518 94586 27616
rect 6025 27383 6123 27481
rect 6450 27383 6548 27481
rect 6882 27383 6980 27481
rect 7264 27360 7362 27458
rect 7660 27360 7758 27458
rect 99428 27360 99526 27458
rect 99824 27360 99922 27458
rect 100206 27383 100304 27481
rect 100638 27383 100736 27481
rect 101063 27383 101161 27481
rect 12600 27202 12698 27300
rect 94488 27202 94586 27300
rect 6025 27009 6123 27107
rect 6450 26951 6548 27049
rect 6882 26951 6980 27049
rect 7264 26965 7362 27063
rect 7660 26965 7758 27063
rect 12600 26965 12698 27063
rect 94488 26965 94586 27063
rect 99428 26965 99526 27063
rect 99824 26965 99922 27063
rect 100206 26951 100304 27049
rect 100638 26951 100736 27049
rect 101063 27009 101161 27107
rect 12600 26728 12698 26826
rect 94488 26728 94586 26826
rect 6025 26593 6123 26691
rect 6450 26593 6548 26691
rect 6882 26593 6980 26691
rect 7264 26570 7362 26668
rect 7660 26570 7758 26668
rect 99428 26570 99526 26668
rect 99824 26570 99922 26668
rect 100206 26593 100304 26691
rect 100638 26593 100736 26691
rect 101063 26593 101161 26691
rect 12600 26412 12698 26510
rect 94488 26412 94586 26510
rect 6025 26219 6123 26317
rect 6450 26161 6548 26259
rect 6882 26161 6980 26259
rect 7264 26175 7362 26273
rect 7660 26175 7758 26273
rect 12600 26175 12698 26273
rect 94488 26175 94586 26273
rect 99428 26175 99526 26273
rect 99824 26175 99922 26273
rect 100206 26161 100304 26259
rect 100638 26161 100736 26259
rect 101063 26219 101161 26317
rect 12600 25938 12698 26036
rect 94488 25938 94586 26036
rect 6025 25803 6123 25901
rect 6450 25803 6548 25901
rect 6882 25803 6980 25901
rect 7264 25780 7362 25878
rect 7660 25780 7758 25878
rect 99428 25780 99526 25878
rect 99824 25780 99922 25878
rect 100206 25803 100304 25901
rect 100638 25803 100736 25901
rect 101063 25803 101161 25901
rect 12600 25622 12698 25720
rect 94488 25622 94586 25720
rect 6025 25429 6123 25527
rect 6450 25371 6548 25469
rect 6882 25371 6980 25469
rect 7264 25385 7362 25483
rect 7660 25385 7758 25483
rect 12600 25385 12698 25483
rect 94488 25385 94586 25483
rect 99428 25385 99526 25483
rect 99824 25385 99922 25483
rect 100206 25371 100304 25469
rect 100638 25371 100736 25469
rect 101063 25429 101161 25527
rect 12600 25148 12698 25246
rect 94488 25148 94586 25246
rect 6025 25013 6123 25111
rect 6450 25013 6548 25111
rect 6882 25013 6980 25111
rect 7264 24990 7362 25088
rect 7660 24990 7758 25088
rect 99428 24990 99526 25088
rect 99824 24990 99922 25088
rect 100206 25013 100304 25111
rect 100638 25013 100736 25111
rect 101063 25013 101161 25111
rect 12600 24832 12698 24930
rect 94488 24832 94586 24930
rect 6025 24639 6123 24737
rect 6450 24581 6548 24679
rect 6882 24581 6980 24679
rect 7264 24595 7362 24693
rect 7660 24595 7758 24693
rect 12600 24595 12698 24693
rect 94488 24595 94586 24693
rect 99428 24595 99526 24693
rect 99824 24595 99922 24693
rect 100206 24581 100304 24679
rect 100638 24581 100736 24679
rect 101063 24639 101161 24737
rect 12600 24358 12698 24456
rect 94488 24358 94586 24456
rect 6025 24223 6123 24321
rect 6450 24223 6548 24321
rect 6882 24223 6980 24321
rect 7264 24200 7362 24298
rect 7660 24200 7758 24298
rect 99428 24200 99526 24298
rect 99824 24200 99922 24298
rect 100206 24223 100304 24321
rect 100638 24223 100736 24321
rect 101063 24223 101161 24321
rect 12600 24042 12698 24140
rect 94488 24042 94586 24140
rect 6025 23849 6123 23947
rect 6450 23791 6548 23889
rect 6882 23791 6980 23889
rect 7264 23805 7362 23903
rect 7660 23805 7758 23903
rect 12600 23805 12698 23903
rect 94488 23805 94586 23903
rect 99428 23805 99526 23903
rect 99824 23805 99922 23903
rect 100206 23791 100304 23889
rect 100638 23791 100736 23889
rect 101063 23849 101161 23947
rect 12600 23568 12698 23666
rect 94488 23568 94586 23666
rect 6025 23433 6123 23531
rect 6450 23433 6548 23531
rect 6882 23433 6980 23531
rect 7264 23410 7362 23508
rect 7660 23410 7758 23508
rect 99428 23410 99526 23508
rect 99824 23410 99922 23508
rect 100206 23433 100304 23531
rect 100638 23433 100736 23531
rect 101063 23433 101161 23531
rect 12600 23252 12698 23350
rect 94488 23252 94586 23350
rect 6025 23059 6123 23157
rect 6450 23001 6548 23099
rect 6882 23001 6980 23099
rect 7264 23015 7362 23113
rect 7660 23015 7758 23113
rect 12600 23015 12698 23113
rect 94488 23015 94586 23113
rect 99428 23015 99526 23113
rect 99824 23015 99922 23113
rect 100206 23001 100304 23099
rect 100638 23001 100736 23099
rect 101063 23059 101161 23157
rect 12600 22778 12698 22876
rect 94488 22778 94586 22876
rect 6025 22643 6123 22741
rect 6450 22643 6548 22741
rect 6882 22643 6980 22741
rect 7264 22620 7362 22718
rect 7660 22620 7758 22718
rect 99428 22620 99526 22718
rect 99824 22620 99922 22718
rect 100206 22643 100304 22741
rect 100638 22643 100736 22741
rect 101063 22643 101161 22741
rect 12600 22462 12698 22560
rect 94488 22462 94586 22560
rect 6025 22269 6123 22367
rect 6450 22211 6548 22309
rect 6882 22211 6980 22309
rect 7264 22225 7362 22323
rect 7660 22225 7758 22323
rect 12600 22225 12698 22323
rect 94488 22225 94586 22323
rect 99428 22225 99526 22323
rect 99824 22225 99922 22323
rect 100206 22211 100304 22309
rect 100638 22211 100736 22309
rect 101063 22269 101161 22367
rect 12600 21988 12698 22086
rect 94488 21988 94586 22086
rect 6025 21853 6123 21951
rect 6450 21853 6548 21951
rect 6882 21853 6980 21951
rect 7264 21830 7362 21928
rect 7660 21830 7758 21928
rect 99428 21830 99526 21928
rect 99824 21830 99922 21928
rect 100206 21853 100304 21951
rect 100638 21853 100736 21951
rect 101063 21853 101161 21951
rect 12600 21672 12698 21770
rect 94488 21672 94586 21770
rect 6025 21479 6123 21577
rect 6450 21421 6548 21519
rect 6882 21421 6980 21519
rect 7264 21435 7362 21533
rect 7660 21435 7758 21533
rect 12600 21435 12698 21533
rect 94488 21435 94586 21533
rect 99428 21435 99526 21533
rect 99824 21435 99922 21533
rect 100206 21421 100304 21519
rect 100638 21421 100736 21519
rect 101063 21479 101161 21577
rect 12600 21198 12698 21296
rect 94488 21198 94586 21296
rect 6025 21063 6123 21161
rect 6450 21063 6548 21161
rect 6882 21063 6980 21161
rect 7264 21040 7362 21138
rect 7660 21040 7758 21138
rect 99428 21040 99526 21138
rect 99824 21040 99922 21138
rect 100206 21063 100304 21161
rect 100638 21063 100736 21161
rect 101063 21063 101161 21161
rect 12600 20882 12698 20980
rect 94488 20882 94586 20980
rect 6025 20689 6123 20787
rect 6450 20631 6548 20729
rect 6882 20631 6980 20729
rect 7264 20645 7362 20743
rect 7660 20645 7758 20743
rect 12600 20645 12698 20743
rect 94488 20645 94586 20743
rect 99428 20645 99526 20743
rect 99824 20645 99922 20743
rect 100206 20631 100304 20729
rect 100638 20631 100736 20729
rect 101063 20689 101161 20787
rect 12600 20408 12698 20506
rect 94488 20408 94586 20506
rect 6025 20273 6123 20371
rect 6450 20273 6548 20371
rect 6882 20273 6980 20371
rect 7264 20250 7362 20348
rect 7660 20250 7758 20348
rect 99428 20250 99526 20348
rect 99824 20250 99922 20348
rect 100206 20273 100304 20371
rect 100638 20273 100736 20371
rect 101063 20273 101161 20371
rect 12600 20092 12698 20190
rect 94488 20092 94586 20190
rect 6025 19899 6123 19997
rect 6450 19841 6548 19939
rect 6882 19841 6980 19939
rect 7264 19855 7362 19953
rect 7660 19855 7758 19953
rect 12600 19855 12698 19953
rect 94488 19855 94586 19953
rect 99428 19855 99526 19953
rect 99824 19855 99922 19953
rect 100206 19841 100304 19939
rect 100638 19841 100736 19939
rect 101063 19899 101161 19997
rect 12600 19618 12698 19716
rect 94488 19618 94586 19716
rect 6025 19483 6123 19581
rect 6450 19483 6548 19581
rect 6882 19483 6980 19581
rect 7264 19460 7362 19558
rect 7660 19460 7758 19558
rect 99428 19460 99526 19558
rect 99824 19460 99922 19558
rect 100206 19483 100304 19581
rect 100638 19483 100736 19581
rect 101063 19483 101161 19581
rect 12600 19302 12698 19400
rect 94488 19302 94586 19400
rect 6025 19109 6123 19207
rect 6450 19051 6548 19149
rect 6882 19051 6980 19149
rect 7264 19065 7362 19163
rect 7660 19065 7758 19163
rect 12600 19065 12698 19163
rect 94488 19065 94586 19163
rect 99428 19065 99526 19163
rect 99824 19065 99922 19163
rect 100206 19051 100304 19149
rect 100638 19051 100736 19149
rect 101063 19109 101161 19207
rect 12600 18828 12698 18926
rect 94488 18828 94586 18926
rect 6025 18693 6123 18791
rect 6450 18693 6548 18791
rect 6882 18693 6980 18791
rect 7264 18670 7362 18768
rect 7660 18670 7758 18768
rect 99428 18670 99526 18768
rect 99824 18670 99922 18768
rect 100206 18693 100304 18791
rect 100638 18693 100736 18791
rect 101063 18693 101161 18791
rect 12600 18512 12698 18610
rect 94488 18512 94586 18610
rect 6025 18319 6123 18417
rect 6450 18261 6548 18359
rect 6882 18261 6980 18359
rect 7264 18275 7362 18373
rect 7660 18275 7758 18373
rect 12600 18275 12698 18373
rect 94488 18275 94586 18373
rect 99428 18275 99526 18373
rect 99824 18275 99922 18373
rect 100206 18261 100304 18359
rect 100638 18261 100736 18359
rect 101063 18319 101161 18417
rect 12600 18038 12698 18136
rect 94488 18038 94586 18136
rect 2611 17903 2709 18001
rect 3036 17903 3134 18001
rect 3468 17903 3566 18001
rect 3850 17880 3948 17978
rect 4246 17880 4344 17978
rect 6025 17903 6123 18001
rect 6450 17903 6548 18001
rect 6882 17903 6980 18001
rect 7264 17880 7362 17978
rect 7660 17880 7758 17978
rect 99428 17880 99526 17978
rect 99824 17880 99922 17978
rect 100206 17903 100304 18001
rect 100638 17903 100736 18001
rect 101063 17903 101161 18001
rect 102842 17880 102940 17978
rect 103238 17880 103336 17978
rect 103620 17903 103718 18001
rect 104052 17903 104150 18001
rect 104477 17903 104575 18001
rect 12600 17722 12698 17820
rect 94488 17722 94586 17820
rect 6025 17529 6123 17627
rect 6450 17471 6548 17569
rect 6882 17471 6980 17569
rect 7264 17485 7362 17583
rect 7660 17485 7758 17583
rect 12600 17485 12698 17583
rect 94488 17485 94586 17583
rect 99428 17485 99526 17583
rect 99824 17485 99922 17583
rect 100206 17471 100304 17569
rect 100638 17471 100736 17569
rect 101063 17529 101161 17627
rect 12600 17248 12698 17346
rect 94488 17248 94586 17346
rect 2611 17113 2709 17211
rect 3036 17113 3134 17211
rect 3468 17113 3566 17211
rect 3850 17090 3948 17188
rect 4246 17090 4344 17188
rect 6025 17113 6123 17211
rect 6450 17113 6548 17211
rect 6882 17113 6980 17211
rect 7264 17090 7362 17188
rect 7660 17090 7758 17188
rect 99428 17090 99526 17188
rect 99824 17090 99922 17188
rect 100206 17113 100304 17211
rect 100638 17113 100736 17211
rect 101063 17113 101161 17211
rect 102842 17090 102940 17188
rect 103238 17090 103336 17188
rect 103620 17113 103718 17211
rect 104052 17113 104150 17211
rect 104477 17113 104575 17211
rect 12600 16932 12698 17030
rect 94488 16932 94586 17030
rect 6025 16739 6123 16837
rect 6450 16681 6548 16779
rect 6882 16681 6980 16779
rect 7264 16695 7362 16793
rect 7660 16695 7758 16793
rect 12600 16695 12698 16793
rect 94488 16695 94586 16793
rect 99428 16695 99526 16793
rect 99824 16695 99922 16793
rect 100206 16681 100304 16779
rect 100638 16681 100736 16779
rect 101063 16739 101161 16837
rect 12600 16458 12698 16556
rect 94488 16458 94586 16556
rect 2611 16323 2709 16421
rect 3036 16323 3134 16421
rect 3468 16323 3566 16421
rect 3850 16300 3948 16398
rect 4246 16300 4344 16398
rect 6025 16323 6123 16421
rect 6450 16323 6548 16421
rect 6882 16323 6980 16421
rect 7264 16300 7362 16398
rect 7660 16300 7758 16398
rect 99428 16300 99526 16398
rect 99824 16300 99922 16398
rect 100206 16323 100304 16421
rect 100638 16323 100736 16421
rect 101063 16323 101161 16421
rect 102842 16300 102940 16398
rect 103238 16300 103336 16398
rect 103620 16323 103718 16421
rect 104052 16323 104150 16421
rect 104477 16323 104575 16421
rect 12600 16142 12698 16240
rect 94488 16142 94586 16240
rect 6025 15949 6123 16047
rect 6450 15891 6548 15989
rect 6882 15891 6980 15989
rect 7264 15905 7362 16003
rect 7660 15905 7758 16003
rect 12600 15905 12698 16003
rect 94488 15905 94586 16003
rect 99428 15905 99526 16003
rect 99824 15905 99922 16003
rect 100206 15891 100304 15989
rect 100638 15891 100736 15989
rect 101063 15949 101161 16047
rect 12600 15668 12698 15766
rect 94488 15668 94586 15766
rect 1156 15510 1254 15608
rect 1552 15510 1650 15608
rect 2611 15533 2709 15631
rect 3036 15533 3134 15631
rect 3468 15533 3566 15631
rect 3850 15510 3948 15608
rect 4246 15510 4344 15608
rect 6025 15533 6123 15631
rect 6450 15533 6548 15631
rect 6882 15533 6980 15631
rect 7264 15510 7362 15608
rect 7660 15510 7758 15608
rect 99428 15510 99526 15608
rect 99824 15510 99922 15608
rect 100206 15533 100304 15631
rect 100638 15533 100736 15631
rect 101063 15533 101161 15631
rect 102842 15510 102940 15608
rect 103238 15510 103336 15608
rect 103620 15533 103718 15631
rect 104052 15533 104150 15631
rect 104477 15533 104575 15631
rect 105536 15510 105634 15608
rect 105932 15510 106030 15608
rect 12600 15352 12698 15450
rect 94488 15352 94586 15450
rect 6025 15159 6123 15257
rect 6450 15101 6548 15199
rect 6882 15101 6980 15199
rect 7264 15115 7362 15213
rect 7660 15115 7758 15213
rect 12600 15115 12698 15213
rect 94488 15115 94586 15213
rect 99428 15115 99526 15213
rect 99824 15115 99922 15213
rect 100206 15101 100304 15199
rect 100638 15101 100736 15199
rect 101063 15159 101161 15257
rect 12600 14878 12698 14976
rect 94488 14878 94586 14976
rect 6025 14743 6123 14841
rect 6450 14743 6548 14841
rect 6882 14743 6980 14841
rect 7264 14720 7362 14818
rect 7660 14720 7758 14818
rect 99428 14720 99526 14818
rect 99824 14720 99922 14818
rect 100206 14743 100304 14841
rect 100638 14743 100736 14841
rect 101063 14743 101161 14841
rect 12600 14562 12698 14660
rect 94488 14562 94586 14660
rect 6025 14369 6123 14467
rect 6450 14311 6548 14409
rect 6882 14311 6980 14409
rect 7264 14325 7362 14423
rect 7660 14325 7758 14423
rect 12600 14325 12698 14423
rect 94488 14325 94586 14423
rect 99428 14325 99526 14423
rect 99824 14325 99922 14423
rect 100206 14311 100304 14409
rect 100638 14311 100736 14409
rect 101063 14369 101161 14467
rect 12600 14088 12698 14186
rect 94488 14088 94586 14186
rect 3046 13937 3144 14035
rect 3471 13937 3569 14035
rect 3850 13930 3948 14028
rect 4246 13930 4344 14028
rect 6025 13953 6123 14051
rect 6450 13953 6548 14051
rect 6882 13953 6980 14051
rect 7264 13930 7362 14028
rect 7660 13930 7758 14028
rect 99428 13930 99526 14028
rect 99824 13930 99922 14028
rect 100206 13953 100304 14051
rect 100638 13953 100736 14051
rect 101063 13953 101161 14051
rect 102842 13930 102940 14028
rect 103238 13930 103336 14028
rect 103617 13937 103715 14035
rect 104042 13937 104140 14035
rect 12600 13772 12698 13870
rect 94488 13772 94586 13870
rect 6025 13579 6123 13677
rect 6450 13521 6548 13619
rect 6882 13521 6980 13619
rect 7264 13535 7362 13633
rect 7660 13535 7758 13633
rect 12600 13535 12698 13633
rect 94488 13535 94586 13633
rect 99428 13535 99526 13633
rect 99824 13535 99922 13633
rect 100206 13521 100304 13619
rect 100638 13521 100736 13619
rect 101063 13579 101161 13677
rect 12600 13298 12698 13396
rect 94488 13298 94586 13396
rect 1752 13140 1850 13238
rect 2148 13140 2246 13238
rect 3046 13147 3144 13245
rect 3471 13147 3569 13245
rect 3850 13140 3948 13238
rect 4246 13140 4344 13238
rect 6025 13163 6123 13261
rect 6450 13163 6548 13261
rect 6882 13163 6980 13261
rect 7264 13140 7362 13238
rect 7660 13140 7758 13238
rect 99428 13140 99526 13238
rect 99824 13140 99922 13238
rect 100206 13163 100304 13261
rect 100638 13163 100736 13261
rect 101063 13163 101161 13261
rect 102842 13140 102940 13238
rect 103238 13140 103336 13238
rect 103617 13147 103715 13245
rect 104042 13147 104140 13245
rect 104940 13140 105038 13238
rect 105336 13140 105434 13238
rect 12600 12982 12698 13080
rect 94488 12982 94586 13080
rect 6025 12789 6123 12887
rect 6450 12731 6548 12829
rect 6882 12731 6980 12829
rect 7264 12745 7362 12843
rect 7660 12745 7758 12843
rect 12600 12745 12698 12843
rect 94488 12745 94586 12843
rect 99428 12745 99526 12843
rect 99824 12745 99922 12843
rect 100206 12731 100304 12829
rect 100638 12731 100736 12829
rect 101063 12789 101161 12887
rect 12600 12508 12698 12606
rect 94488 12508 94586 12606
rect 6025 12373 6123 12471
rect 6450 12373 6548 12471
rect 6882 12373 6980 12471
rect 7264 12350 7362 12448
rect 7660 12350 7758 12448
rect 99428 12350 99526 12448
rect 99824 12350 99922 12448
rect 100206 12373 100304 12471
rect 100638 12373 100736 12471
rect 101063 12373 101161 12471
rect 12600 12192 12698 12290
rect 94488 12192 94586 12290
rect 6025 11999 6123 12097
rect 6450 11941 6548 12039
rect 6882 11941 6980 12039
rect 7264 11955 7362 12053
rect 7660 11955 7758 12053
rect 12600 11955 12698 12053
rect 94488 11955 94586 12053
rect 99428 11955 99526 12053
rect 99824 11955 99922 12053
rect 100206 11941 100304 12039
rect 100638 11941 100736 12039
rect 101063 11999 101161 12097
rect 12600 11718 12698 11816
rect 94488 11718 94586 11816
rect 3046 11567 3144 11665
rect 3471 11567 3569 11665
rect 3850 11560 3948 11658
rect 4246 11560 4344 11658
rect 6025 11583 6123 11681
rect 6450 11583 6548 11681
rect 6882 11583 6980 11681
rect 7264 11560 7362 11658
rect 7660 11560 7758 11658
rect 99428 11560 99526 11658
rect 99824 11560 99922 11658
rect 100206 11583 100304 11681
rect 100638 11583 100736 11681
rect 101063 11583 101161 11681
rect 102842 11560 102940 11658
rect 103238 11560 103336 11658
rect 103617 11567 103715 11665
rect 104042 11567 104140 11665
rect 12600 11402 12698 11500
rect 94488 11402 94586 11500
rect 6025 11209 6123 11307
rect 6450 11151 6548 11249
rect 6882 11151 6980 11249
rect 7264 11165 7362 11263
rect 7660 11165 7758 11263
rect 12600 11165 12698 11263
rect 94488 11165 94586 11263
rect 99428 11165 99526 11263
rect 99824 11165 99922 11263
rect 100206 11151 100304 11249
rect 100638 11151 100736 11249
rect 101063 11209 101161 11307
rect 12600 10928 12698 11026
rect 94488 10928 94586 11026
rect 1752 10770 1850 10868
rect 2148 10770 2246 10868
rect 3046 10777 3144 10875
rect 3471 10777 3569 10875
rect 3850 10770 3948 10868
rect 4246 10770 4344 10868
rect 6025 10793 6123 10891
rect 6450 10793 6548 10891
rect 6882 10793 6980 10891
rect 7264 10770 7362 10868
rect 7660 10770 7758 10868
rect 99428 10770 99526 10868
rect 99824 10770 99922 10868
rect 100206 10793 100304 10891
rect 100638 10793 100736 10891
rect 101063 10793 101161 10891
rect 102842 10770 102940 10868
rect 103238 10770 103336 10868
rect 103617 10777 103715 10875
rect 104042 10777 104140 10875
rect 104940 10770 105038 10868
rect 105336 10770 105434 10868
rect 12600 10612 12698 10710
rect 94488 10612 94586 10710
rect 12600 10375 12698 10473
rect 94488 10375 94586 10473
rect 7685 10184 7783 10282
rect 8517 10190 8615 10288
rect 11208 10178 11306 10276
rect 12234 10248 12332 10346
rect 94854 10248 94952 10346
rect 13296 9814 13394 9912
rect 13920 9814 14018 9912
rect 14544 9814 14642 9912
rect 15168 9814 15266 9912
rect 15792 9814 15890 9912
rect 16416 9814 16514 9912
rect 17040 9814 17138 9912
rect 17664 9814 17762 9912
rect 18288 9814 18386 9912
rect 18912 9814 19010 9912
rect 19536 9814 19634 9912
rect 20160 9814 20258 9912
rect 20784 9814 20882 9912
rect 21408 9814 21506 9912
rect 22032 9814 22130 9912
rect 22656 9814 22754 9912
rect 23280 9814 23378 9912
rect 23904 9814 24002 9912
rect 24528 9814 24626 9912
rect 25152 9814 25250 9912
rect 25776 9814 25874 9912
rect 26400 9814 26498 9912
rect 27024 9814 27122 9912
rect 27648 9814 27746 9912
rect 28272 9814 28370 9912
rect 28896 9814 28994 9912
rect 29520 9814 29618 9912
rect 30144 9814 30242 9912
rect 30768 9814 30866 9912
rect 31392 9814 31490 9912
rect 32016 9814 32114 9912
rect 32640 9814 32738 9912
rect 33264 9814 33362 9912
rect 33888 9814 33986 9912
rect 34512 9814 34610 9912
rect 35136 9814 35234 9912
rect 35760 9814 35858 9912
rect 36384 9814 36482 9912
rect 37008 9814 37106 9912
rect 37632 9814 37730 9912
rect 38256 9814 38354 9912
rect 38880 9814 38978 9912
rect 39504 9814 39602 9912
rect 40128 9814 40226 9912
rect 40752 9814 40850 9912
rect 41376 9814 41474 9912
rect 42000 9814 42098 9912
rect 42624 9814 42722 9912
rect 43248 9814 43346 9912
rect 43872 9814 43970 9912
rect 44496 9814 44594 9912
rect 45120 9814 45218 9912
rect 45744 9814 45842 9912
rect 46368 9814 46466 9912
rect 46992 9814 47090 9912
rect 47616 9814 47714 9912
rect 48240 9814 48338 9912
rect 48864 9814 48962 9912
rect 49488 9814 49586 9912
rect 50112 9814 50210 9912
rect 50736 9814 50834 9912
rect 51360 9814 51458 9912
rect 51984 9814 52082 9912
rect 52608 9814 52706 9912
rect 53232 9814 53330 9912
rect 53856 9814 53954 9912
rect 54480 9814 54578 9912
rect 55104 9814 55202 9912
rect 55728 9814 55826 9912
rect 56352 9814 56450 9912
rect 56976 9814 57074 9912
rect 57600 9814 57698 9912
rect 58224 9814 58322 9912
rect 58848 9814 58946 9912
rect 59472 9814 59570 9912
rect 60096 9814 60194 9912
rect 60720 9814 60818 9912
rect 61344 9814 61442 9912
rect 61968 9814 62066 9912
rect 62592 9814 62690 9912
rect 63216 9814 63314 9912
rect 63840 9814 63938 9912
rect 64464 9814 64562 9912
rect 65088 9814 65186 9912
rect 65712 9814 65810 9912
rect 66336 9814 66434 9912
rect 66960 9814 67058 9912
rect 67584 9814 67682 9912
rect 68208 9814 68306 9912
rect 68832 9814 68930 9912
rect 69456 9814 69554 9912
rect 70080 9814 70178 9912
rect 70704 9814 70802 9912
rect 71328 9814 71426 9912
rect 71952 9814 72050 9912
rect 72576 9814 72674 9912
rect 73200 9814 73298 9912
rect 73824 9814 73922 9912
rect 74448 9814 74546 9912
rect 75072 9814 75170 9912
rect 75696 9814 75794 9912
rect 76320 9814 76418 9912
rect 76944 9814 77042 9912
rect 77568 9814 77666 9912
rect 78192 9814 78290 9912
rect 78816 9814 78914 9912
rect 79440 9814 79538 9912
rect 80064 9814 80162 9912
rect 80688 9814 80786 9912
rect 81312 9814 81410 9912
rect 81936 9814 82034 9912
rect 82560 9814 82658 9912
rect 83184 9814 83282 9912
rect 83808 9814 83906 9912
rect 84432 9814 84530 9912
rect 85056 9814 85154 9912
rect 85680 9814 85778 9912
rect 86304 9814 86402 9912
rect 86928 9814 87026 9912
rect 87552 9814 87650 9912
rect 88176 9814 88274 9912
rect 88800 9814 88898 9912
rect 89424 9814 89522 9912
rect 90048 9814 90146 9912
rect 90672 9814 90770 9912
rect 91296 9814 91394 9912
rect 91920 9814 92018 9912
rect 92544 9814 92642 9912
rect 93168 9814 93266 9912
rect 93792 9814 93890 9912
rect 13415 9223 13513 9321
rect 13801 9223 13899 9321
rect 14663 9223 14761 9321
rect 15049 9223 15147 9321
rect 15911 9223 16009 9321
rect 16297 9223 16395 9321
rect 17159 9223 17257 9321
rect 17545 9223 17643 9321
rect 18407 9223 18505 9321
rect 18793 9223 18891 9321
rect 19655 9223 19753 9321
rect 20041 9223 20139 9321
rect 20903 9223 21001 9321
rect 21289 9223 21387 9321
rect 22151 9223 22249 9321
rect 22537 9223 22635 9321
rect 23399 9223 23497 9321
rect 23785 9223 23883 9321
rect 24647 9223 24745 9321
rect 25033 9223 25131 9321
rect 25895 9223 25993 9321
rect 26281 9223 26379 9321
rect 27143 9223 27241 9321
rect 27529 9223 27627 9321
rect 28391 9223 28489 9321
rect 28777 9223 28875 9321
rect 29639 9223 29737 9321
rect 30025 9223 30123 9321
rect 30887 9223 30985 9321
rect 31273 9223 31371 9321
rect 32135 9223 32233 9321
rect 32521 9223 32619 9321
rect 33383 9223 33481 9321
rect 33769 9223 33867 9321
rect 34631 9223 34729 9321
rect 35017 9223 35115 9321
rect 35879 9223 35977 9321
rect 36265 9223 36363 9321
rect 37127 9223 37225 9321
rect 37513 9223 37611 9321
rect 38375 9223 38473 9321
rect 38761 9223 38859 9321
rect 39623 9223 39721 9321
rect 40009 9223 40107 9321
rect 40871 9223 40969 9321
rect 41257 9223 41355 9321
rect 42119 9223 42217 9321
rect 42505 9223 42603 9321
rect 43367 9223 43465 9321
rect 43753 9223 43851 9321
rect 44615 9223 44713 9321
rect 45001 9223 45099 9321
rect 45863 9223 45961 9321
rect 46249 9223 46347 9321
rect 47111 9223 47209 9321
rect 47497 9223 47595 9321
rect 48359 9223 48457 9321
rect 48745 9223 48843 9321
rect 49607 9223 49705 9321
rect 49993 9223 50091 9321
rect 50855 9223 50953 9321
rect 51241 9223 51339 9321
rect 52103 9223 52201 9321
rect 52489 9223 52587 9321
rect 53351 9223 53449 9321
rect 53737 9223 53835 9321
rect 54599 9223 54697 9321
rect 54985 9223 55083 9321
rect 55847 9223 55945 9321
rect 56233 9223 56331 9321
rect 57095 9223 57193 9321
rect 57481 9223 57579 9321
rect 58343 9223 58441 9321
rect 58729 9223 58827 9321
rect 59591 9223 59689 9321
rect 59977 9223 60075 9321
rect 60839 9223 60937 9321
rect 61225 9223 61323 9321
rect 62087 9223 62185 9321
rect 62473 9223 62571 9321
rect 63335 9223 63433 9321
rect 63721 9223 63819 9321
rect 64583 9223 64681 9321
rect 64969 9223 65067 9321
rect 65831 9223 65929 9321
rect 66217 9223 66315 9321
rect 67079 9223 67177 9321
rect 67465 9223 67563 9321
rect 68327 9223 68425 9321
rect 68713 9223 68811 9321
rect 69575 9223 69673 9321
rect 69961 9223 70059 9321
rect 70823 9223 70921 9321
rect 71209 9223 71307 9321
rect 72071 9223 72169 9321
rect 72457 9223 72555 9321
rect 73319 9223 73417 9321
rect 73705 9223 73803 9321
rect 74567 9223 74665 9321
rect 74953 9223 75051 9321
rect 75815 9223 75913 9321
rect 76201 9223 76299 9321
rect 77063 9223 77161 9321
rect 77449 9223 77547 9321
rect 78311 9223 78409 9321
rect 78697 9223 78795 9321
rect 79559 9223 79657 9321
rect 79945 9223 80043 9321
rect 80807 9223 80905 9321
rect 81193 9223 81291 9321
rect 82055 9223 82153 9321
rect 82441 9223 82539 9321
rect 83303 9223 83401 9321
rect 83689 9223 83787 9321
rect 84551 9223 84649 9321
rect 84937 9223 85035 9321
rect 85799 9223 85897 9321
rect 86185 9223 86283 9321
rect 87047 9223 87145 9321
rect 87433 9223 87531 9321
rect 88295 9223 88393 9321
rect 88681 9223 88779 9321
rect 89543 9223 89641 9321
rect 89929 9223 90027 9321
rect 90791 9223 90889 9321
rect 91177 9223 91275 9321
rect 92039 9223 92137 9321
rect 92425 9223 92523 9321
rect 93287 9223 93385 9321
rect 11677 8623 52906 8683
rect 0 8474 13577 8534
rect 5360 7817 5458 7915
rect 6472 7817 6570 7915
rect 14232 7674 14330 7772
rect 15480 7674 15578 7772
rect 16728 7674 16826 7772
rect 17976 7674 18074 7772
rect 19224 7674 19322 7772
rect 20472 7674 20570 7772
rect 21720 7674 21818 7772
rect 22968 7674 23066 7772
rect 24216 7674 24314 7772
rect 25464 7674 25562 7772
rect 26712 7674 26810 7772
rect 27960 7674 28058 7772
rect 29208 7674 29306 7772
rect 30456 7674 30554 7772
rect 31704 7674 31802 7772
rect 32952 7674 33050 7772
rect 34200 7674 34298 7772
rect 35448 7674 35546 7772
rect 36696 7674 36794 7772
rect 37944 7674 38042 7772
rect 39192 7674 39290 7772
rect 40440 7674 40538 7772
rect 41688 7674 41786 7772
rect 42936 7674 43034 7772
rect 44184 7674 44282 7772
rect 45432 7674 45530 7772
rect 46680 7674 46778 7772
rect 47928 7674 48026 7772
rect 49176 7674 49274 7772
rect 50424 7674 50522 7772
rect 51672 7674 51770 7772
rect 52920 7674 53018 7772
rect 54168 7674 54266 7772
rect 55416 7674 55514 7772
rect 56664 7674 56762 7772
rect 57912 7674 58010 7772
rect 59160 7674 59258 7772
rect 60408 7674 60506 7772
rect 61656 7674 61754 7772
rect 62904 7674 63002 7772
rect 64152 7674 64250 7772
rect 65400 7674 65498 7772
rect 66648 7674 66746 7772
rect 67896 7674 67994 7772
rect 69144 7674 69242 7772
rect 70392 7674 70490 7772
rect 71640 7674 71738 7772
rect 72888 7674 72986 7772
rect 74136 7674 74234 7772
rect 75384 7674 75482 7772
rect 76632 7674 76730 7772
rect 77880 7674 77978 7772
rect 79128 7674 79226 7772
rect 80376 7674 80474 7772
rect 81624 7674 81722 7772
rect 82872 7674 82970 7772
rect 84120 7674 84218 7772
rect 85368 7674 85466 7772
rect 86616 7674 86714 7772
rect 87864 7674 87962 7772
rect 89112 7674 89210 7772
rect 90360 7674 90458 7772
rect 91608 7674 91706 7772
rect 92856 7674 92954 7772
rect 7202 7167 7481 7227
rect 7481 6936 12313 6996
rect 7753 6812 12313 6872
rect 7617 6688 12313 6748
rect 7481 6564 12313 6624
rect 5360 6403 5458 6501
rect 6472 6403 6570 6501
rect 11801 5848 51908 5908
rect 7202 5677 7753 5737
rect 14059 5677 14157 5775
rect 16555 5677 16653 5775
rect 19051 5677 19149 5775
rect 21547 5677 21645 5775
rect 24043 5677 24141 5775
rect 26539 5677 26637 5775
rect 29035 5677 29133 5775
rect 31531 5677 31629 5775
rect 34027 5677 34125 5775
rect 36523 5677 36621 5775
rect 39019 5677 39117 5775
rect 41515 5677 41613 5775
rect 44011 5677 44109 5775
rect 46507 5677 46605 5775
rect 49003 5677 49101 5775
rect 51499 5677 51597 5775
rect 53995 5677 54093 5775
rect 56491 5677 56589 5775
rect 58987 5677 59085 5775
rect 61483 5677 61581 5775
rect 63979 5677 64077 5775
rect 66475 5677 66573 5775
rect 68971 5677 69069 5775
rect 71467 5677 71565 5775
rect 73963 5677 74061 5775
rect 76459 5677 76557 5775
rect 78955 5677 79053 5775
rect 81451 5677 81549 5775
rect 83947 5677 84045 5775
rect 86443 5677 86541 5775
rect 88939 5677 89037 5775
rect 91435 5677 91533 5775
rect 5360 4989 5458 5087
rect 6472 4989 6570 5087
rect 13977 4903 14075 5001
rect 16473 4903 16571 5001
rect 18969 4903 19067 5001
rect 21465 4903 21563 5001
rect 23961 4903 24059 5001
rect 26457 4903 26555 5001
rect 28953 4903 29051 5001
rect 31449 4903 31547 5001
rect 33945 4903 34043 5001
rect 36441 4903 36539 5001
rect 38937 4903 39035 5001
rect 41433 4903 41531 5001
rect 43929 4903 44027 5001
rect 46425 4903 46523 5001
rect 48921 4903 49019 5001
rect 51417 4903 51515 5001
rect 53913 4903 54011 5001
rect 56409 4903 56507 5001
rect 58905 4903 59003 5001
rect 61401 4903 61499 5001
rect 63897 4903 63995 5001
rect 66393 4903 66491 5001
rect 68889 4903 68987 5001
rect 71385 4903 71483 5001
rect 73881 4903 73979 5001
rect 76377 4903 76475 5001
rect 78873 4903 78971 5001
rect 81369 4903 81467 5001
rect 83865 4903 83963 5001
rect 86361 4903 86459 5001
rect 88857 4903 88955 5001
rect 91353 4903 91451 5001
rect 7202 4339 7617 4399
rect 13989 4065 14087 4163
rect 16485 4065 16583 4163
rect 18981 4065 19079 4163
rect 21477 4065 21575 4163
rect 23973 4065 24071 4163
rect 26469 4065 26567 4163
rect 28965 4065 29063 4163
rect 31461 4065 31559 4163
rect 33957 4065 34055 4163
rect 36453 4065 36551 4163
rect 38949 4065 39047 4163
rect 41445 4065 41543 4163
rect 43941 4065 44039 4163
rect 46437 4065 46535 4163
rect 48933 4065 49031 4163
rect 51429 4065 51527 4163
rect 53925 4065 54023 4163
rect 56421 4065 56519 4163
rect 58917 4065 59015 4163
rect 61413 4065 61511 4163
rect 63909 4065 64007 4163
rect 66405 4065 66503 4163
rect 68901 4065 68999 4163
rect 71397 4065 71495 4163
rect 73893 4065 73991 4163
rect 76389 4065 76487 4163
rect 78885 4065 78983 4163
rect 81381 4065 81479 4163
rect 83877 4065 83975 4163
rect 86373 4065 86471 4163
rect 88869 4065 88967 4163
rect 91365 4065 91463 4163
rect 13989 3743 14087 3841
rect 16485 3743 16583 3841
rect 18981 3743 19079 3841
rect 21477 3743 21575 3841
rect 23973 3743 24071 3841
rect 26469 3743 26567 3841
rect 28965 3743 29063 3841
rect 31461 3743 31559 3841
rect 33957 3743 34055 3841
rect 36453 3743 36551 3841
rect 38949 3743 39047 3841
rect 41445 3743 41543 3841
rect 43941 3743 44039 3841
rect 46437 3743 46535 3841
rect 48933 3743 49031 3841
rect 51429 3743 51527 3841
rect 53925 3743 54023 3841
rect 56421 3743 56519 3841
rect 58917 3743 59015 3841
rect 61413 3743 61511 3841
rect 63909 3743 64007 3841
rect 66405 3743 66503 3841
rect 68901 3743 68999 3841
rect 71397 3743 71495 3841
rect 73893 3743 73991 3841
rect 76389 3743 76487 3841
rect 78885 3743 78983 3841
rect 81381 3743 81479 3841
rect 83877 3743 83975 3841
rect 86373 3743 86471 3841
rect 88869 3743 88967 3841
rect 91365 3743 91463 3841
rect 5360 3575 5458 3673
rect 6472 3575 6570 3673
rect 13875 2950 13973 3048
rect 16371 2950 16469 3048
rect 18867 2950 18965 3048
rect 21363 2950 21461 3048
rect 23859 2950 23957 3048
rect 26355 2950 26453 3048
rect 28851 2950 28949 3048
rect 31347 2950 31445 3048
rect 33843 2950 33941 3048
rect 36339 2950 36437 3048
rect 38835 2950 38933 3048
rect 41331 2950 41429 3048
rect 43827 2950 43925 3048
rect 46323 2950 46421 3048
rect 48819 2950 48917 3048
rect 51315 2950 51413 3048
rect 53811 2950 53909 3048
rect 56307 2950 56405 3048
rect 58803 2950 58901 3048
rect 61299 2950 61397 3048
rect 63795 2950 63893 3048
rect 66291 2950 66389 3048
rect 68787 2950 68885 3048
rect 71283 2950 71381 3048
rect 73779 2950 73877 3048
rect 76275 2950 76373 3048
rect 78771 2950 78869 3048
rect 81267 2950 81365 3048
rect 83763 2950 83861 3048
rect 86259 2950 86357 3048
rect 88755 2950 88853 3048
rect 91251 2950 91349 3048
rect 7202 2849 7481 2909
rect 13864 2513 13962 2611
rect 16360 2513 16458 2611
rect 18856 2513 18954 2611
rect 21352 2513 21450 2611
rect 23848 2513 23946 2611
rect 26344 2513 26442 2611
rect 28840 2513 28938 2611
rect 31336 2513 31434 2611
rect 33832 2513 33930 2611
rect 36328 2513 36426 2611
rect 38824 2513 38922 2611
rect 41320 2513 41418 2611
rect 43816 2513 43914 2611
rect 46312 2513 46410 2611
rect 48808 2513 48906 2611
rect 51304 2513 51402 2611
rect 53800 2513 53898 2611
rect 56296 2513 56394 2611
rect 58792 2513 58890 2611
rect 61288 2513 61386 2611
rect 63784 2513 63882 2611
rect 66280 2513 66378 2611
rect 68776 2513 68874 2611
rect 71272 2513 71370 2611
rect 73768 2513 73866 2611
rect 76264 2513 76362 2611
rect 78760 2513 78858 2611
rect 81256 2513 81354 2611
rect 83752 2513 83850 2611
rect 86248 2513 86346 2611
rect 88744 2513 88842 2611
rect 91240 2513 91338 2611
rect 5360 2161 5458 2259
rect 6472 2161 6570 2259
rect 13985 2181 14083 2279
rect 16481 2181 16579 2279
rect 18977 2181 19075 2279
rect 21473 2181 21571 2279
rect 23969 2181 24067 2279
rect 26465 2181 26563 2279
rect 28961 2181 29059 2279
rect 31457 2181 31555 2279
rect 33953 2181 34051 2279
rect 36449 2181 36547 2279
rect 38945 2181 39043 2279
rect 41441 2181 41539 2279
rect 43937 2181 44035 2279
rect 46433 2181 46531 2279
rect 48929 2181 49027 2279
rect 51425 2181 51523 2279
rect 53921 2181 54019 2279
rect 56417 2181 56515 2279
rect 58913 2181 59011 2279
rect 61409 2181 61507 2279
rect 63905 2181 64003 2279
rect 66401 2181 66499 2279
rect 68897 2181 68995 2279
rect 71393 2181 71491 2279
rect 73889 2181 73987 2279
rect 76385 2181 76483 2279
rect 78881 2181 78979 2279
rect 81377 2181 81475 2279
rect 83873 2181 83971 2279
rect 86369 2181 86467 2279
rect 88865 2181 88963 2279
rect 91361 2181 91459 2279
rect 13870 1979 13968 2077
rect 16366 1979 16464 2077
rect 18862 1979 18960 2077
rect 21358 1979 21456 2077
rect 23854 1979 23952 2077
rect 26350 1979 26448 2077
rect 28846 1979 28944 2077
rect 31342 1979 31440 2077
rect 33838 1979 33936 2077
rect 36334 1979 36432 2077
rect 38830 1979 38928 2077
rect 41326 1979 41424 2077
rect 43822 1979 43920 2077
rect 46318 1979 46416 2077
rect 48814 1979 48912 2077
rect 51310 1979 51408 2077
rect 53806 1979 53904 2077
rect 56302 1979 56400 2077
rect 58798 1979 58896 2077
rect 61294 1979 61392 2077
rect 63790 1979 63888 2077
rect 66286 1979 66384 2077
rect 68782 1979 68880 2077
rect 71278 1979 71376 2077
rect 73774 1979 73872 2077
rect 76270 1979 76368 2077
rect 78766 1979 78864 2077
rect 81262 1979 81360 2077
rect 83758 1979 83856 2077
rect 86254 1979 86352 2077
rect 88750 1979 88848 2077
rect 91246 1979 91344 2077
rect 13884 1563 13982 1661
rect 16380 1563 16478 1661
rect 18876 1563 18974 1661
rect 21372 1563 21470 1661
rect 23868 1563 23966 1661
rect 26364 1563 26462 1661
rect 28860 1563 28958 1661
rect 31356 1563 31454 1661
rect 33852 1563 33950 1661
rect 36348 1563 36446 1661
rect 38844 1563 38942 1661
rect 41340 1563 41438 1661
rect 43836 1563 43934 1661
rect 46332 1563 46430 1661
rect 48828 1563 48926 1661
rect 51324 1563 51422 1661
rect 53820 1563 53918 1661
rect 56316 1563 56414 1661
rect 58812 1563 58910 1661
rect 61308 1563 61406 1661
rect 63804 1563 63902 1661
rect 66300 1563 66398 1661
rect 68796 1563 68894 1661
rect 71292 1563 71390 1661
rect 73788 1563 73886 1661
rect 76284 1563 76382 1661
rect 78780 1563 78878 1661
rect 81276 1563 81374 1661
rect 83772 1563 83870 1661
rect 86268 1563 86366 1661
rect 88764 1563 88862 1661
rect 91260 1563 91358 1661
rect 12234 1120 12332 1218
rect 93480 1120 93578 1218
rect 11925 537 52906 597
rect 12234 0 12332 98
rect 93480 0 93578 98
use sky130_sram_2kbyte_1rw1r_32x512_8_port_address  sky130_sram_2kbyte_1rw1r_32x512_8_port_address_0
timestamp 1626065694
transform 1 0 0 0 1 10424
box 0 -490 12011 50620
use sky130_sram_2kbyte_1rw1r_32x512_8_port_address_0  sky130_sram_2kbyte_1rw1r_32x512_8_port_address_0_0
timestamp 1626065694
transform -1 0 107186 0 1 10424
box 0 -60 12011 51050
use sky130_sram_2kbyte_1rw1r_32x512_8_hierarchical_predecode2x4_0  sky130_sram_2kbyte_1rw1r_32x512_8_hierarchical_predecode2x4_0_1
timestamp 1626065694
transform -1 0 102059 0 -1 69198
box 0 -49 2390 5705
use sky130_sram_2kbyte_1rw1r_32x512_8_hierarchical_predecode2x4_0  sky130_sram_2kbyte_1rw1r_32x512_8_hierarchical_predecode2x4_0_0
timestamp 1626065694
transform 1 0 5003 0 1 2210
box 0 -49 2390 5705
use sky130_sram_2kbyte_1rw1r_32x512_8_port_data_0  sky130_sram_2kbyte_1rw1r_32x512_8_port_data_0_0
timestamp 1626065694
transform 1 0 12283 0 1 61774
box 0 238 81870 5950
use sky130_sram_2kbyte_1rw1r_32x512_8_port_data  sky130_sram_2kbyte_1rw1r_32x512_8_port_data_0
timestamp 1626065694
transform 1 0 12283 0 -1 9634
box -49 238 81295 9634
use sky130_sram_2kbyte_1rw1r_32x512_8_replica_bitcell_array  sky130_sram_2kbyte_1rw1r_32x512_8_replica_bitcell_array_0
timestamp 1626065694
transform 1 0 12283 0 1 9634
box -49 0 82669 52140
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_30
timestamp 1626065694
transform 1 0 93576 0 1 62867
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_29
timestamp 1626065694
transform 1 0 99052 0 1 64174
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_28
timestamp 1626065694
transform 1 0 99827 0 1 64174
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_27
timestamp 1626065694
transform 1 0 99052 0 1 64405
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_26
timestamp 1626065694
transform 1 0 99052 0 1 67002
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_25
timestamp 1626065694
transform 1 0 99827 0 1 67002
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_24
timestamp 1626065694
transform 1 0 99052 0 1 64653
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_23
timestamp 1626065694
transform 1 0 99188 0 1 65664
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_22
timestamp 1626065694
transform 1 0 99827 0 1 65664
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_21
timestamp 1626065694
transform 1 0 99188 0 1 64529
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_20
timestamp 1626065694
transform 1 0 99324 0 1 68492
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_19
timestamp 1626065694
transform 1 0 99827 0 1 68492
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_18
timestamp 1626065694
transform 1 0 99324 0 1 64777
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_17
timestamp 1626065694
transform 1 0 95318 0 1 62718
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_16
timestamp 1626065694
transform 1 0 95194 0 1 65493
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_15
timestamp 1626065694
transform 1 0 13544 0 1 8467
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_14
timestamp 1626065694
transform 1 0 7448 0 1 2842
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_13
timestamp 1626065694
transform 1 0 7169 0 1 2842
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_12
timestamp 1626065694
transform 1 0 7448 0 1 6557
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_11
timestamp 1626065694
transform 1 0 7448 0 1 7160
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_10
timestamp 1626065694
transform 1 0 7169 0 1 7160
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_9
timestamp 1626065694
transform 1 0 7448 0 1 6929
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_8
timestamp 1626065694
transform 1 0 7584 0 1 4332
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_7
timestamp 1626065694
transform 1 0 7169 0 1 4332
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_6
timestamp 1626065694
transform 1 0 7584 0 1 6681
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_5
timestamp 1626065694
transform 1 0 7720 0 1 5670
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_4
timestamp 1626065694
transform 1 0 7169 0 1 5670
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_3
timestamp 1626065694
transform 1 0 7720 0 1 6805
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_2
timestamp 1626065694
transform 1 0 11644 0 1 8616
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_1
timestamp 1626065694
transform 1 0 11892 0 1 530
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_0
timestamp 1626065694
transform 1 0 11768 0 1 5841
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_267
timestamp 1626065694
transform 1 0 93577 0 1 62872
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_266
timestamp 1626065694
transform 1 0 94998 0 1 52142
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_265
timestamp 1626065694
transform 1 0 94998 0 1 52382
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_264
timestamp 1626065694
transform 1 0 94998 0 1 52932
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_263
timestamp 1626065694
transform 1 0 94998 0 1 53172
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_262
timestamp 1626065694
transform 1 0 94998 0 1 53722
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_261
timestamp 1626065694
transform 1 0 94998 0 1 53962
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_260
timestamp 1626065694
transform 1 0 94998 0 1 54512
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_259
timestamp 1626065694
transform 1 0 94998 0 1 54752
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_258
timestamp 1626065694
transform 1 0 94998 0 1 55302
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_257
timestamp 1626065694
transform 1 0 94998 0 1 55542
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_256
timestamp 1626065694
transform 1 0 94998 0 1 56092
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_255
timestamp 1626065694
transform 1 0 94998 0 1 56332
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_254
timestamp 1626065694
transform 1 0 94998 0 1 56882
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_253
timestamp 1626065694
transform 1 0 94998 0 1 57122
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_252
timestamp 1626065694
transform 1 0 94998 0 1 57672
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_251
timestamp 1626065694
transform 1 0 94998 0 1 57912
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_250
timestamp 1626065694
transform 1 0 94998 0 1 58462
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_249
timestamp 1626065694
transform 1 0 94998 0 1 58702
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_248
timestamp 1626065694
transform 1 0 94998 0 1 59252
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_247
timestamp 1626065694
transform 1 0 94998 0 1 59492
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_246
timestamp 1626065694
transform 1 0 94998 0 1 60042
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_245
timestamp 1626065694
transform 1 0 94998 0 1 60282
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_244
timestamp 1626065694
transform 1 0 94998 0 1 60832
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_243
timestamp 1626065694
transform 1 0 94998 0 1 61072
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_242
timestamp 1626065694
transform 1 0 99828 0 1 64179
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_241
timestamp 1626065694
transform 1 0 99828 0 1 67007
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_240
timestamp 1626065694
transform 1 0 99828 0 1 65669
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_239
timestamp 1626065694
transform 1 0 99828 0 1 68497
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_238
timestamp 1626065694
transform 1 0 94998 0 1 48432
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_237
timestamp 1626065694
transform 1 0 94998 0 1 48982
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_236
timestamp 1626065694
transform 1 0 94998 0 1 49222
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_235
timestamp 1626065694
transform 1 0 94998 0 1 49772
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_234
timestamp 1626065694
transform 1 0 94998 0 1 50012
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_233
timestamp 1626065694
transform 1 0 94998 0 1 50562
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_232
timestamp 1626065694
transform 1 0 94998 0 1 50802
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_231
timestamp 1626065694
transform 1 0 94998 0 1 51352
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_230
timestamp 1626065694
transform 1 0 94998 0 1 51592
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_229
timestamp 1626065694
transform 1 0 94998 0 1 34762
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_228
timestamp 1626065694
transform 1 0 94998 0 1 35002
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_227
timestamp 1626065694
transform 1 0 94998 0 1 35552
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_226
timestamp 1626065694
transform 1 0 94998 0 1 35792
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_225
timestamp 1626065694
transform 1 0 94998 0 1 36342
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_224
timestamp 1626065694
transform 1 0 94998 0 1 36582
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_223
timestamp 1626065694
transform 1 0 94998 0 1 37132
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_222
timestamp 1626065694
transform 1 0 94998 0 1 37372
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_221
timestamp 1626065694
transform 1 0 94998 0 1 37922
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_220
timestamp 1626065694
transform 1 0 94998 0 1 38162
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_219
timestamp 1626065694
transform 1 0 94998 0 1 38712
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_218
timestamp 1626065694
transform 1 0 94998 0 1 38952
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_217
timestamp 1626065694
transform 1 0 94998 0 1 39502
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_216
timestamp 1626065694
transform 1 0 94998 0 1 39742
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_215
timestamp 1626065694
transform 1 0 94998 0 1 40292
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_214
timestamp 1626065694
transform 1 0 94998 0 1 40532
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_213
timestamp 1626065694
transform 1 0 94998 0 1 41082
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_212
timestamp 1626065694
transform 1 0 94998 0 1 41322
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_211
timestamp 1626065694
transform 1 0 94998 0 1 41872
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_210
timestamp 1626065694
transform 1 0 94998 0 1 42112
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_209
timestamp 1626065694
transform 1 0 94998 0 1 42662
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_208
timestamp 1626065694
transform 1 0 94998 0 1 42902
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_207
timestamp 1626065694
transform 1 0 94998 0 1 43452
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_206
timestamp 1626065694
transform 1 0 94998 0 1 43692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_205
timestamp 1626065694
transform 1 0 94998 0 1 44242
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_204
timestamp 1626065694
transform 1 0 94998 0 1 44482
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_203
timestamp 1626065694
transform 1 0 94998 0 1 45032
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_202
timestamp 1626065694
transform 1 0 94998 0 1 45272
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_201
timestamp 1626065694
transform 1 0 94998 0 1 45822
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_200
timestamp 1626065694
transform 1 0 94998 0 1 46062
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_199
timestamp 1626065694
transform 1 0 94998 0 1 46612
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_198
timestamp 1626065694
transform 1 0 94998 0 1 46852
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_197
timestamp 1626065694
transform 1 0 94998 0 1 47402
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_196
timestamp 1626065694
transform 1 0 94998 0 1 47642
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_195
timestamp 1626065694
transform 1 0 94998 0 1 48192
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_194
timestamp 1626065694
transform 1 0 12124 0 1 52142
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_193
timestamp 1626065694
transform 1 0 12124 0 1 52382
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_192
timestamp 1626065694
transform 1 0 12124 0 1 52932
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_191
timestamp 1626065694
transform 1 0 12124 0 1 53172
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_190
timestamp 1626065694
transform 1 0 12124 0 1 53722
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_189
timestamp 1626065694
transform 1 0 12124 0 1 53962
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_188
timestamp 1626065694
transform 1 0 12124 0 1 54512
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_187
timestamp 1626065694
transform 1 0 12124 0 1 54752
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_186
timestamp 1626065694
transform 1 0 12124 0 1 55302
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_185
timestamp 1626065694
transform 1 0 12124 0 1 55542
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_184
timestamp 1626065694
transform 1 0 12124 0 1 56092
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_183
timestamp 1626065694
transform 1 0 12124 0 1 56332
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_182
timestamp 1626065694
transform 1 0 12124 0 1 56882
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_181
timestamp 1626065694
transform 1 0 12124 0 1 57122
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_180
timestamp 1626065694
transform 1 0 12124 0 1 57672
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_179
timestamp 1626065694
transform 1 0 12124 0 1 57912
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_178
timestamp 1626065694
transform 1 0 12124 0 1 58462
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_177
timestamp 1626065694
transform 1 0 12124 0 1 58702
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_176
timestamp 1626065694
transform 1 0 12124 0 1 59252
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_175
timestamp 1626065694
transform 1 0 12124 0 1 59492
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_174
timestamp 1626065694
transform 1 0 12124 0 1 60042
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_173
timestamp 1626065694
transform 1 0 12124 0 1 60282
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_172
timestamp 1626065694
transform 1 0 12124 0 1 60832
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_171
timestamp 1626065694
transform 1 0 12124 0 1 48982
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_170
timestamp 1626065694
transform 1 0 12124 0 1 49222
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_169
timestamp 1626065694
transform 1 0 12124 0 1 49772
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_168
timestamp 1626065694
transform 1 0 12124 0 1 50012
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_167
timestamp 1626065694
transform 1 0 12124 0 1 50562
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_166
timestamp 1626065694
transform 1 0 12124 0 1 50802
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_165
timestamp 1626065694
transform 1 0 12124 0 1 51352
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_164
timestamp 1626065694
transform 1 0 12124 0 1 51592
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_163
timestamp 1626065694
transform 1 0 12124 0 1 39742
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_162
timestamp 1626065694
transform 1 0 12124 0 1 40292
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_161
timestamp 1626065694
transform 1 0 12124 0 1 40532
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_160
timestamp 1626065694
transform 1 0 12124 0 1 41082
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_159
timestamp 1626065694
transform 1 0 12124 0 1 41322
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_158
timestamp 1626065694
transform 1 0 12124 0 1 41872
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_157
timestamp 1626065694
transform 1 0 12124 0 1 42112
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_156
timestamp 1626065694
transform 1 0 12124 0 1 42662
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_155
timestamp 1626065694
transform 1 0 12124 0 1 42902
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_154
timestamp 1626065694
transform 1 0 12124 0 1 43452
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_153
timestamp 1626065694
transform 1 0 12124 0 1 43692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_152
timestamp 1626065694
transform 1 0 12124 0 1 44242
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_151
timestamp 1626065694
transform 1 0 12124 0 1 44482
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_150
timestamp 1626065694
transform 1 0 12124 0 1 45032
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_149
timestamp 1626065694
transform 1 0 12124 0 1 45272
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_148
timestamp 1626065694
transform 1 0 12124 0 1 45822
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_147
timestamp 1626065694
transform 1 0 12124 0 1 46062
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_146
timestamp 1626065694
transform 1 0 12124 0 1 46612
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_145
timestamp 1626065694
transform 1 0 12124 0 1 46852
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_144
timestamp 1626065694
transform 1 0 12124 0 1 47402
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_143
timestamp 1626065694
transform 1 0 12124 0 1 47642
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_142
timestamp 1626065694
transform 1 0 12124 0 1 48192
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_141
timestamp 1626065694
transform 1 0 12124 0 1 48432
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_140
timestamp 1626065694
transform 1 0 12124 0 1 34762
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_139
timestamp 1626065694
transform 1 0 12124 0 1 35002
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_138
timestamp 1626065694
transform 1 0 12124 0 1 35552
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_137
timestamp 1626065694
transform 1 0 12124 0 1 35792
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_136
timestamp 1626065694
transform 1 0 12124 0 1 36342
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_135
timestamp 1626065694
transform 1 0 12124 0 1 36582
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_134
timestamp 1626065694
transform 1 0 12124 0 1 37132
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_133
timestamp 1626065694
transform 1 0 12124 0 1 37372
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_132
timestamp 1626065694
transform 1 0 12124 0 1 37922
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_131
timestamp 1626065694
transform 1 0 12124 0 1 38162
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_130
timestamp 1626065694
transform 1 0 12124 0 1 38712
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_129
timestamp 1626065694
transform 1 0 12124 0 1 38952
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_128
timestamp 1626065694
transform 1 0 12124 0 1 39502
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_127
timestamp 1626065694
transform 1 0 12124 0 1 17382
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_126
timestamp 1626065694
transform 1 0 12124 0 1 17622
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_125
timestamp 1626065694
transform 1 0 12124 0 1 18172
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_124
timestamp 1626065694
transform 1 0 12124 0 1 18412
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_123
timestamp 1626065694
transform 1 0 12124 0 1 18962
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_122
timestamp 1626065694
transform 1 0 12124 0 1 19202
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_121
timestamp 1626065694
transform 1 0 12124 0 1 19752
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_120
timestamp 1626065694
transform 1 0 12124 0 1 19992
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_119
timestamp 1626065694
transform 1 0 12124 0 1 20542
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_118
timestamp 1626065694
transform 1 0 12124 0 1 20782
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_117
timestamp 1626065694
transform 1 0 12124 0 1 21332
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_116
timestamp 1626065694
transform 1 0 12124 0 1 21572
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_115
timestamp 1626065694
transform 1 0 12124 0 1 22122
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_114
timestamp 1626065694
transform 1 0 12124 0 1 22362
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_113
timestamp 1626065694
transform 1 0 12124 0 1 22912
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_112
timestamp 1626065694
transform 1 0 12124 0 1 23152
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_111
timestamp 1626065694
transform 1 0 12124 0 1 23702
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_110
timestamp 1626065694
transform 1 0 12124 0 1 23942
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_109
timestamp 1626065694
transform 1 0 12124 0 1 24492
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_108
timestamp 1626065694
transform 1 0 12124 0 1 24732
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_107
timestamp 1626065694
transform 1 0 12124 0 1 25282
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_106
timestamp 1626065694
transform 1 0 12124 0 1 25522
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_105
timestamp 1626065694
transform 1 0 12124 0 1 26072
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_104
timestamp 1626065694
transform 1 0 12124 0 1 26312
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_103
timestamp 1626065694
transform 1 0 12124 0 1 26862
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_102
timestamp 1626065694
transform 1 0 12124 0 1 27102
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_101
timestamp 1626065694
transform 1 0 12124 0 1 27652
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_100
timestamp 1626065694
transform 1 0 12124 0 1 27892
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_99
timestamp 1626065694
transform 1 0 12124 0 1 28442
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_98
timestamp 1626065694
transform 1 0 12124 0 1 28682
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_97
timestamp 1626065694
transform 1 0 12124 0 1 29232
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_96
timestamp 1626065694
transform 1 0 12124 0 1 29472
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_95
timestamp 1626065694
transform 1 0 12124 0 1 30022
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_94
timestamp 1626065694
transform 1 0 12124 0 1 30262
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_93
timestamp 1626065694
transform 1 0 12124 0 1 30812
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_92
timestamp 1626065694
transform 1 0 12124 0 1 31052
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_91
timestamp 1626065694
transform 1 0 12124 0 1 31602
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_90
timestamp 1626065694
transform 1 0 12124 0 1 31842
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_89
timestamp 1626065694
transform 1 0 12124 0 1 32392
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_88
timestamp 1626065694
transform 1 0 12124 0 1 32632
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_87
timestamp 1626065694
transform 1 0 12124 0 1 33182
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_86
timestamp 1626065694
transform 1 0 12124 0 1 33422
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_85
timestamp 1626065694
transform 1 0 12124 0 1 33972
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_84
timestamp 1626065694
transform 1 0 12124 0 1 34212
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_83
timestamp 1626065694
transform 1 0 12124 0 1 16832
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_82
timestamp 1626065694
transform 1 0 12124 0 1 13672
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_81
timestamp 1626065694
transform 1 0 12124 0 1 14222
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_80
timestamp 1626065694
transform 1 0 12124 0 1 14462
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_79
timestamp 1626065694
transform 1 0 12124 0 1 15012
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_78
timestamp 1626065694
transform 1 0 12124 0 1 15252
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_77
timestamp 1626065694
transform 1 0 12124 0 1 15802
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_76
timestamp 1626065694
transform 1 0 12124 0 1 16042
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_75
timestamp 1626065694
transform 1 0 12124 0 1 16592
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_74
timestamp 1626065694
transform 1 0 13545 0 1 8472
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_73
timestamp 1626065694
transform 1 0 12124 0 1 10512
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_72
timestamp 1626065694
transform 1 0 12124 0 1 11062
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_71
timestamp 1626065694
transform 1 0 12124 0 1 11302
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_70
timestamp 1626065694
transform 1 0 12124 0 1 10272
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_69
timestamp 1626065694
transform 1 0 7170 0 1 2847
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_68
timestamp 1626065694
transform 1 0 7170 0 1 7165
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_67
timestamp 1626065694
transform 1 0 7170 0 1 4337
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_66
timestamp 1626065694
transform 1 0 7170 0 1 5675
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_65
timestamp 1626065694
transform 1 0 12124 0 1 11852
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_64
timestamp 1626065694
transform 1 0 12124 0 1 12092
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_63
timestamp 1626065694
transform 1 0 12124 0 1 12642
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_62
timestamp 1626065694
transform 1 0 12124 0 1 12882
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_61
timestamp 1626065694
transform 1 0 12124 0 1 13432
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_60
timestamp 1626065694
transform 1 0 94998 0 1 17622
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_59
timestamp 1626065694
transform 1 0 94998 0 1 18172
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_58
timestamp 1626065694
transform 1 0 94998 0 1 18412
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_57
timestamp 1626065694
transform 1 0 94998 0 1 18962
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_56
timestamp 1626065694
transform 1 0 94998 0 1 19202
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_55
timestamp 1626065694
transform 1 0 94998 0 1 19752
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_54
timestamp 1626065694
transform 1 0 94998 0 1 19992
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_53
timestamp 1626065694
transform 1 0 94998 0 1 20542
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_52
timestamp 1626065694
transform 1 0 94998 0 1 20782
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_51
timestamp 1626065694
transform 1 0 94998 0 1 21332
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_50
timestamp 1626065694
transform 1 0 94998 0 1 21572
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_49
timestamp 1626065694
transform 1 0 94998 0 1 22122
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_48
timestamp 1626065694
transform 1 0 94998 0 1 22362
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_47
timestamp 1626065694
transform 1 0 94998 0 1 22912
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_46
timestamp 1626065694
transform 1 0 94998 0 1 23152
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_45
timestamp 1626065694
transform 1 0 94998 0 1 23702
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_44
timestamp 1626065694
transform 1 0 94998 0 1 23942
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_43
timestamp 1626065694
transform 1 0 94998 0 1 24492
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_42
timestamp 1626065694
transform 1 0 94998 0 1 24732
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_41
timestamp 1626065694
transform 1 0 94998 0 1 25282
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_40
timestamp 1626065694
transform 1 0 94998 0 1 25522
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_39
timestamp 1626065694
transform 1 0 94998 0 1 26072
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_38
timestamp 1626065694
transform 1 0 94998 0 1 26312
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_37
timestamp 1626065694
transform 1 0 94998 0 1 26862
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_36
timestamp 1626065694
transform 1 0 94998 0 1 27102
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_35
timestamp 1626065694
transform 1 0 94998 0 1 27652
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_34
timestamp 1626065694
transform 1 0 94998 0 1 27892
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_33
timestamp 1626065694
transform 1 0 94998 0 1 28442
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_32
timestamp 1626065694
transform 1 0 94998 0 1 28682
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_31
timestamp 1626065694
transform 1 0 94998 0 1 29232
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_30
timestamp 1626065694
transform 1 0 94998 0 1 29472
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_29
timestamp 1626065694
transform 1 0 94998 0 1 30022
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_28
timestamp 1626065694
transform 1 0 94998 0 1 30262
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_27
timestamp 1626065694
transform 1 0 94998 0 1 30812
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_26
timestamp 1626065694
transform 1 0 94998 0 1 31052
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_25
timestamp 1626065694
transform 1 0 94998 0 1 31602
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_24
timestamp 1626065694
transform 1 0 94998 0 1 31842
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_23
timestamp 1626065694
transform 1 0 94998 0 1 32392
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_22
timestamp 1626065694
transform 1 0 94998 0 1 32632
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_21
timestamp 1626065694
transform 1 0 94998 0 1 33182
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_20
timestamp 1626065694
transform 1 0 94998 0 1 33422
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_19
timestamp 1626065694
transform 1 0 94998 0 1 33972
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_18
timestamp 1626065694
transform 1 0 94998 0 1 34212
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_17
timestamp 1626065694
transform 1 0 94998 0 1 17382
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_16
timestamp 1626065694
transform 1 0 94998 0 1 11062
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_15
timestamp 1626065694
transform 1 0 94998 0 1 11302
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_14
timestamp 1626065694
transform 1 0 94998 0 1 11852
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_13
timestamp 1626065694
transform 1 0 94998 0 1 12092
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_12
timestamp 1626065694
transform 1 0 94998 0 1 12642
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_11
timestamp 1626065694
transform 1 0 94998 0 1 12882
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_10
timestamp 1626065694
transform 1 0 94998 0 1 13432
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_9
timestamp 1626065694
transform 1 0 94998 0 1 13672
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_8
timestamp 1626065694
transform 1 0 94998 0 1 14222
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_7
timestamp 1626065694
transform 1 0 94998 0 1 14462
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_6
timestamp 1626065694
transform 1 0 94998 0 1 15012
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_5
timestamp 1626065694
transform 1 0 94998 0 1 15252
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_4
timestamp 1626065694
transform 1 0 94998 0 1 15802
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_3
timestamp 1626065694
transform 1 0 94998 0 1 16042
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_2
timestamp 1626065694
transform 1 0 94998 0 1 16592
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_1
timestamp 1626065694
transform 1 0 94998 0 1 16832
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_0
timestamp 1626065694
transform 1 0 94998 0 1 10512
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_265
timestamp 1626065694
transform 1 0 95001 0 1 52141
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_264
timestamp 1626065694
transform 1 0 95001 0 1 52381
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_263
timestamp 1626065694
transform 1 0 95001 0 1 52931
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_262
timestamp 1626065694
transform 1 0 95001 0 1 53171
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_261
timestamp 1626065694
transform 1 0 95001 0 1 53721
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_260
timestamp 1626065694
transform 1 0 95001 0 1 53961
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_259
timestamp 1626065694
transform 1 0 95001 0 1 54511
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_258
timestamp 1626065694
transform 1 0 95001 0 1 54751
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_257
timestamp 1626065694
transform 1 0 95001 0 1 55301
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_256
timestamp 1626065694
transform 1 0 95001 0 1 55541
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_255
timestamp 1626065694
transform 1 0 95001 0 1 56091
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_254
timestamp 1626065694
transform 1 0 95001 0 1 56331
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_253
timestamp 1626065694
transform 1 0 95001 0 1 56881
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_252
timestamp 1626065694
transform 1 0 95001 0 1 57121
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_251
timestamp 1626065694
transform 1 0 95001 0 1 57671
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_250
timestamp 1626065694
transform 1 0 95001 0 1 57911
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_249
timestamp 1626065694
transform 1 0 95001 0 1 58461
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_248
timestamp 1626065694
transform 1 0 95001 0 1 58701
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_247
timestamp 1626065694
transform 1 0 95001 0 1 59251
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_246
timestamp 1626065694
transform 1 0 95001 0 1 59491
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_245
timestamp 1626065694
transform 1 0 95001 0 1 60041
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_244
timestamp 1626065694
transform 1 0 95001 0 1 60281
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_243
timestamp 1626065694
transform 1 0 95001 0 1 60831
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_242
timestamp 1626065694
transform 1 0 95001 0 1 61071
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_241
timestamp 1626065694
transform 1 0 99831 0 1 64178
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_240
timestamp 1626065694
transform 1 0 99831 0 1 67006
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_239
timestamp 1626065694
transform 1 0 99831 0 1 65668
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_238
timestamp 1626065694
transform 1 0 99831 0 1 68496
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_237
timestamp 1626065694
transform 1 0 95001 0 1 48431
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_236
timestamp 1626065694
transform 1 0 95001 0 1 48981
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_235
timestamp 1626065694
transform 1 0 95001 0 1 49221
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_234
timestamp 1626065694
transform 1 0 95001 0 1 49771
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_233
timestamp 1626065694
transform 1 0 95001 0 1 50011
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_232
timestamp 1626065694
transform 1 0 95001 0 1 50561
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_231
timestamp 1626065694
transform 1 0 95001 0 1 50801
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_230
timestamp 1626065694
transform 1 0 95001 0 1 51351
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_229
timestamp 1626065694
transform 1 0 95001 0 1 51591
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_228
timestamp 1626065694
transform 1 0 95001 0 1 34761
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_227
timestamp 1626065694
transform 1 0 95001 0 1 35001
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_226
timestamp 1626065694
transform 1 0 95001 0 1 35551
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_225
timestamp 1626065694
transform 1 0 95001 0 1 35791
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_224
timestamp 1626065694
transform 1 0 95001 0 1 36341
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_223
timestamp 1626065694
transform 1 0 95001 0 1 36581
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_222
timestamp 1626065694
transform 1 0 95001 0 1 37131
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_221
timestamp 1626065694
transform 1 0 95001 0 1 37371
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_220
timestamp 1626065694
transform 1 0 95001 0 1 37921
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_219
timestamp 1626065694
transform 1 0 95001 0 1 38161
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_218
timestamp 1626065694
transform 1 0 95001 0 1 38711
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_217
timestamp 1626065694
transform 1 0 95001 0 1 38951
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_216
timestamp 1626065694
transform 1 0 95001 0 1 39501
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_215
timestamp 1626065694
transform 1 0 95001 0 1 39741
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_214
timestamp 1626065694
transform 1 0 95001 0 1 40291
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_213
timestamp 1626065694
transform 1 0 95001 0 1 40531
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_212
timestamp 1626065694
transform 1 0 95001 0 1 41081
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_211
timestamp 1626065694
transform 1 0 95001 0 1 41321
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_210
timestamp 1626065694
transform 1 0 95001 0 1 41871
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_209
timestamp 1626065694
transform 1 0 95001 0 1 42111
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_208
timestamp 1626065694
transform 1 0 95001 0 1 42661
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_207
timestamp 1626065694
transform 1 0 95001 0 1 42901
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_206
timestamp 1626065694
transform 1 0 95001 0 1 43451
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_205
timestamp 1626065694
transform 1 0 95001 0 1 43691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_204
timestamp 1626065694
transform 1 0 95001 0 1 44241
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_203
timestamp 1626065694
transform 1 0 95001 0 1 44481
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_202
timestamp 1626065694
transform 1 0 95001 0 1 45031
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_201
timestamp 1626065694
transform 1 0 95001 0 1 45271
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_200
timestamp 1626065694
transform 1 0 95001 0 1 45821
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_199
timestamp 1626065694
transform 1 0 95001 0 1 46061
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_198
timestamp 1626065694
transform 1 0 95001 0 1 46611
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_197
timestamp 1626065694
transform 1 0 95001 0 1 46851
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_196
timestamp 1626065694
transform 1 0 95001 0 1 47401
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_195
timestamp 1626065694
transform 1 0 95001 0 1 47641
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_194
timestamp 1626065694
transform 1 0 95001 0 1 48191
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_193
timestamp 1626065694
transform 1 0 12127 0 1 52141
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_192
timestamp 1626065694
transform 1 0 12127 0 1 52381
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_191
timestamp 1626065694
transform 1 0 12127 0 1 52931
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_190
timestamp 1626065694
transform 1 0 12127 0 1 53171
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_189
timestamp 1626065694
transform 1 0 12127 0 1 53721
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_188
timestamp 1626065694
transform 1 0 12127 0 1 53961
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_187
timestamp 1626065694
transform 1 0 12127 0 1 54511
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_186
timestamp 1626065694
transform 1 0 12127 0 1 54751
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_185
timestamp 1626065694
transform 1 0 12127 0 1 55301
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_184
timestamp 1626065694
transform 1 0 12127 0 1 55541
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_183
timestamp 1626065694
transform 1 0 12127 0 1 56091
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_182
timestamp 1626065694
transform 1 0 12127 0 1 56331
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_181
timestamp 1626065694
transform 1 0 12127 0 1 56881
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_180
timestamp 1626065694
transform 1 0 12127 0 1 57121
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_179
timestamp 1626065694
transform 1 0 12127 0 1 57671
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_178
timestamp 1626065694
transform 1 0 12127 0 1 57911
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_177
timestamp 1626065694
transform 1 0 12127 0 1 58461
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_176
timestamp 1626065694
transform 1 0 12127 0 1 58701
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_175
timestamp 1626065694
transform 1 0 12127 0 1 59251
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_174
timestamp 1626065694
transform 1 0 12127 0 1 59491
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_173
timestamp 1626065694
transform 1 0 12127 0 1 60041
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_172
timestamp 1626065694
transform 1 0 12127 0 1 60281
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_171
timestamp 1626065694
transform 1 0 12127 0 1 60831
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_170
timestamp 1626065694
transform 1 0 12127 0 1 48981
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_169
timestamp 1626065694
transform 1 0 12127 0 1 49221
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_168
timestamp 1626065694
transform 1 0 12127 0 1 49771
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_167
timestamp 1626065694
transform 1 0 12127 0 1 50011
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_166
timestamp 1626065694
transform 1 0 12127 0 1 50561
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_165
timestamp 1626065694
transform 1 0 12127 0 1 50801
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_164
timestamp 1626065694
transform 1 0 12127 0 1 51351
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_163
timestamp 1626065694
transform 1 0 12127 0 1 51591
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_162
timestamp 1626065694
transform 1 0 12127 0 1 39741
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_161
timestamp 1626065694
transform 1 0 12127 0 1 40291
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_160
timestamp 1626065694
transform 1 0 12127 0 1 40531
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_159
timestamp 1626065694
transform 1 0 12127 0 1 41081
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_158
timestamp 1626065694
transform 1 0 12127 0 1 41321
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_157
timestamp 1626065694
transform 1 0 12127 0 1 41871
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_156
timestamp 1626065694
transform 1 0 12127 0 1 42111
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_155
timestamp 1626065694
transform 1 0 12127 0 1 42661
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_154
timestamp 1626065694
transform 1 0 12127 0 1 42901
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_153
timestamp 1626065694
transform 1 0 12127 0 1 43451
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_152
timestamp 1626065694
transform 1 0 12127 0 1 43691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_151
timestamp 1626065694
transform 1 0 12127 0 1 44241
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_150
timestamp 1626065694
transform 1 0 12127 0 1 44481
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_149
timestamp 1626065694
transform 1 0 12127 0 1 45031
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_148
timestamp 1626065694
transform 1 0 12127 0 1 45271
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_147
timestamp 1626065694
transform 1 0 12127 0 1 45821
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_146
timestamp 1626065694
transform 1 0 12127 0 1 46061
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_145
timestamp 1626065694
transform 1 0 12127 0 1 46611
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_144
timestamp 1626065694
transform 1 0 12127 0 1 46851
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_143
timestamp 1626065694
transform 1 0 12127 0 1 47401
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_142
timestamp 1626065694
transform 1 0 12127 0 1 47641
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_141
timestamp 1626065694
transform 1 0 12127 0 1 48191
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_140
timestamp 1626065694
transform 1 0 12127 0 1 48431
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_139
timestamp 1626065694
transform 1 0 12127 0 1 34761
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_138
timestamp 1626065694
transform 1 0 12127 0 1 35001
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_137
timestamp 1626065694
transform 1 0 12127 0 1 35551
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_136
timestamp 1626065694
transform 1 0 12127 0 1 35791
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_135
timestamp 1626065694
transform 1 0 12127 0 1 36341
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_134
timestamp 1626065694
transform 1 0 12127 0 1 36581
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_133
timestamp 1626065694
transform 1 0 12127 0 1 37131
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_132
timestamp 1626065694
transform 1 0 12127 0 1 37371
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_131
timestamp 1626065694
transform 1 0 12127 0 1 37921
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_130
timestamp 1626065694
transform 1 0 12127 0 1 38161
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_129
timestamp 1626065694
transform 1 0 12127 0 1 38711
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_128
timestamp 1626065694
transform 1 0 12127 0 1 38951
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_127
timestamp 1626065694
transform 1 0 12127 0 1 39501
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_126
timestamp 1626065694
transform 1 0 12127 0 1 17381
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_125
timestamp 1626065694
transform 1 0 12127 0 1 17621
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_124
timestamp 1626065694
transform 1 0 12127 0 1 18171
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_123
timestamp 1626065694
transform 1 0 12127 0 1 18411
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_122
timestamp 1626065694
transform 1 0 12127 0 1 18961
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_121
timestamp 1626065694
transform 1 0 12127 0 1 19201
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_120
timestamp 1626065694
transform 1 0 12127 0 1 19751
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_119
timestamp 1626065694
transform 1 0 12127 0 1 19991
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_118
timestamp 1626065694
transform 1 0 12127 0 1 20541
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_117
timestamp 1626065694
transform 1 0 12127 0 1 20781
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_116
timestamp 1626065694
transform 1 0 12127 0 1 21331
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_115
timestamp 1626065694
transform 1 0 12127 0 1 21571
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_114
timestamp 1626065694
transform 1 0 12127 0 1 22121
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_113
timestamp 1626065694
transform 1 0 12127 0 1 22361
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_112
timestamp 1626065694
transform 1 0 12127 0 1 22911
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_111
timestamp 1626065694
transform 1 0 12127 0 1 23151
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_110
timestamp 1626065694
transform 1 0 12127 0 1 23701
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_109
timestamp 1626065694
transform 1 0 12127 0 1 23941
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_108
timestamp 1626065694
transform 1 0 12127 0 1 24491
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_107
timestamp 1626065694
transform 1 0 12127 0 1 24731
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_106
timestamp 1626065694
transform 1 0 12127 0 1 25281
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_105
timestamp 1626065694
transform 1 0 12127 0 1 25521
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_104
timestamp 1626065694
transform 1 0 12127 0 1 26071
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_103
timestamp 1626065694
transform 1 0 12127 0 1 26311
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_102
timestamp 1626065694
transform 1 0 12127 0 1 26861
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_101
timestamp 1626065694
transform 1 0 12127 0 1 27101
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_100
timestamp 1626065694
transform 1 0 12127 0 1 27651
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_99
timestamp 1626065694
transform 1 0 12127 0 1 27891
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_98
timestamp 1626065694
transform 1 0 12127 0 1 28441
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_97
timestamp 1626065694
transform 1 0 12127 0 1 28681
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_96
timestamp 1626065694
transform 1 0 12127 0 1 29231
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_95
timestamp 1626065694
transform 1 0 12127 0 1 29471
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_94
timestamp 1626065694
transform 1 0 12127 0 1 30021
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_93
timestamp 1626065694
transform 1 0 12127 0 1 30261
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_92
timestamp 1626065694
transform 1 0 12127 0 1 30811
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_91
timestamp 1626065694
transform 1 0 12127 0 1 31051
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_90
timestamp 1626065694
transform 1 0 12127 0 1 31601
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_89
timestamp 1626065694
transform 1 0 12127 0 1 31841
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_88
timestamp 1626065694
transform 1 0 12127 0 1 32391
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_87
timestamp 1626065694
transform 1 0 12127 0 1 32631
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_86
timestamp 1626065694
transform 1 0 12127 0 1 33181
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_85
timestamp 1626065694
transform 1 0 12127 0 1 33421
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_84
timestamp 1626065694
transform 1 0 12127 0 1 33971
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_83
timestamp 1626065694
transform 1 0 12127 0 1 34211
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_82
timestamp 1626065694
transform 1 0 12127 0 1 16831
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_81
timestamp 1626065694
transform 1 0 12127 0 1 13671
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_80
timestamp 1626065694
transform 1 0 12127 0 1 14221
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_79
timestamp 1626065694
transform 1 0 12127 0 1 14461
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_78
timestamp 1626065694
transform 1 0 12127 0 1 15011
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_77
timestamp 1626065694
transform 1 0 12127 0 1 15251
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_76
timestamp 1626065694
transform 1 0 12127 0 1 15801
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_75
timestamp 1626065694
transform 1 0 12127 0 1 16041
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_74
timestamp 1626065694
transform 1 0 12127 0 1 16591
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_73
timestamp 1626065694
transform 1 0 12127 0 1 10511
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_72
timestamp 1626065694
transform 1 0 12127 0 1 11061
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_71
timestamp 1626065694
transform 1 0 12127 0 1 11301
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_70
timestamp 1626065694
transform 1 0 12127 0 1 10271
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_69
timestamp 1626065694
transform 1 0 7173 0 1 2846
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_68
timestamp 1626065694
transform 1 0 7173 0 1 7164
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_67
timestamp 1626065694
transform 1 0 7173 0 1 4336
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_66
timestamp 1626065694
transform 1 0 7173 0 1 5674
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_65
timestamp 1626065694
transform 1 0 12127 0 1 11851
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_64
timestamp 1626065694
transform 1 0 12127 0 1 12091
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_63
timestamp 1626065694
transform 1 0 12127 0 1 12641
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_62
timestamp 1626065694
transform 1 0 12127 0 1 12881
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_61
timestamp 1626065694
transform 1 0 12127 0 1 13431
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_60
timestamp 1626065694
transform 1 0 95001 0 1 17621
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_59
timestamp 1626065694
transform 1 0 95001 0 1 18171
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_58
timestamp 1626065694
transform 1 0 95001 0 1 18411
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_57
timestamp 1626065694
transform 1 0 95001 0 1 18961
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_56
timestamp 1626065694
transform 1 0 95001 0 1 19201
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_55
timestamp 1626065694
transform 1 0 95001 0 1 19751
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_54
timestamp 1626065694
transform 1 0 95001 0 1 19991
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_53
timestamp 1626065694
transform 1 0 95001 0 1 20541
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_52
timestamp 1626065694
transform 1 0 95001 0 1 20781
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_51
timestamp 1626065694
transform 1 0 95001 0 1 21331
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_50
timestamp 1626065694
transform 1 0 95001 0 1 21571
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_49
timestamp 1626065694
transform 1 0 95001 0 1 22121
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_48
timestamp 1626065694
transform 1 0 95001 0 1 22361
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_47
timestamp 1626065694
transform 1 0 95001 0 1 22911
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_46
timestamp 1626065694
transform 1 0 95001 0 1 23151
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_45
timestamp 1626065694
transform 1 0 95001 0 1 23701
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_44
timestamp 1626065694
transform 1 0 95001 0 1 23941
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_43
timestamp 1626065694
transform 1 0 95001 0 1 24491
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_42
timestamp 1626065694
transform 1 0 95001 0 1 24731
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_41
timestamp 1626065694
transform 1 0 95001 0 1 25281
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_40
timestamp 1626065694
transform 1 0 95001 0 1 25521
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_39
timestamp 1626065694
transform 1 0 95001 0 1 26071
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_38
timestamp 1626065694
transform 1 0 95001 0 1 26311
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_37
timestamp 1626065694
transform 1 0 95001 0 1 26861
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_36
timestamp 1626065694
transform 1 0 95001 0 1 27101
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_35
timestamp 1626065694
transform 1 0 95001 0 1 27651
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_34
timestamp 1626065694
transform 1 0 95001 0 1 27891
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_33
timestamp 1626065694
transform 1 0 95001 0 1 28441
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_32
timestamp 1626065694
transform 1 0 95001 0 1 28681
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_31
timestamp 1626065694
transform 1 0 95001 0 1 29231
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_30
timestamp 1626065694
transform 1 0 95001 0 1 29471
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_29
timestamp 1626065694
transform 1 0 95001 0 1 30021
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_28
timestamp 1626065694
transform 1 0 95001 0 1 30261
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_27
timestamp 1626065694
transform 1 0 95001 0 1 30811
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_26
timestamp 1626065694
transform 1 0 95001 0 1 31051
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_25
timestamp 1626065694
transform 1 0 95001 0 1 31601
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_24
timestamp 1626065694
transform 1 0 95001 0 1 31841
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_23
timestamp 1626065694
transform 1 0 95001 0 1 32391
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_22
timestamp 1626065694
transform 1 0 95001 0 1 32631
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_21
timestamp 1626065694
transform 1 0 95001 0 1 33181
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_20
timestamp 1626065694
transform 1 0 95001 0 1 33421
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_19
timestamp 1626065694
transform 1 0 95001 0 1 33971
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_18
timestamp 1626065694
transform 1 0 95001 0 1 34211
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_17
timestamp 1626065694
transform 1 0 95001 0 1 17381
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_16
timestamp 1626065694
transform 1 0 95001 0 1 11061
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_15
timestamp 1626065694
transform 1 0 95001 0 1 11301
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_14
timestamp 1626065694
transform 1 0 95001 0 1 11851
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_13
timestamp 1626065694
transform 1 0 95001 0 1 12091
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_12
timestamp 1626065694
transform 1 0 95001 0 1 12641
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_11
timestamp 1626065694
transform 1 0 95001 0 1 12881
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_10
timestamp 1626065694
transform 1 0 95001 0 1 13431
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_9
timestamp 1626065694
transform 1 0 95001 0 1 13671
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_8
timestamp 1626065694
transform 1 0 95001 0 1 14221
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_7
timestamp 1626065694
transform 1 0 95001 0 1 14461
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_6
timestamp 1626065694
transform 1 0 95001 0 1 15011
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_5
timestamp 1626065694
transform 1 0 95001 0 1 15251
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_4
timestamp 1626065694
transform 1 0 95001 0 1 15801
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_3
timestamp 1626065694
transform 1 0 95001 0 1 16041
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_2
timestamp 1626065694
transform 1 0 95001 0 1 16591
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1
timestamp 1626065694
transform 1 0 95001 0 1 16831
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_0
timestamp 1626065694
transform 1 0 95001 0 1 10511
box 0 0 58 66
<< labels >>
rlabel metal3 s 93609 62874 107270 62934 4 rbl_bl_1_1
rlabel metal3 s 93287 62087 93385 62185 4 vdd
rlabel metal3 s 100492 64907 100590 65005 4 vdd
rlabel metal3 s 93673 62087 93771 62185 4 vdd
rlabel metal3 s 93168 61496 93266 61594 4 vdd
rlabel metal3 s 99403 61126 99501 61224 4 vdd
rlabel metal3 s 95880 61132 95978 61230 4 vdd
rlabel metal3 s 100492 67735 100590 67833 4 vdd
rlabel metal3 s 101604 64907 101702 65005 4 vdd
rlabel metal3 s 101604 67735 101702 67833 4 vdd
rlabel metal3 s 99428 60540 99526 60638 4 vdd
rlabel metal3 s 100638 60563 100736 60661 4 vdd
rlabel metal3 s 100206 60563 100304 60661 4 vdd
rlabel metal3 s 98571 61120 98669 61218 4 vdd
rlabel metal3 s 93792 61496 93890 61594 4 vdd
rlabel metal3 s 101604 66321 101702 66419 4 gnd
rlabel metal3 s 101604 69149 101702 69247 4 gnd
rlabel metal3 s 100492 69149 100590 69247 4 gnd
rlabel metal3 s 94854 61282 94952 61380 4 gnd
rlabel metal3 s 101604 63493 101702 63591 4 gnd
rlabel metal3 s 92856 63636 92954 63734 4 gnd
rlabel metal3 s 100492 63493 100590 63591 4 gnd
rlabel metal3 s 94488 60698 94586 60796 4 gnd
rlabel metal3 s 94488 60935 94586 61033 4 gnd
rlabel metal3 s 99824 60540 99922 60638 4 gnd
rlabel metal3 s 101063 60563 101161 60661 4 gnd
rlabel metal3 s 100492 66321 100590 66419 4 gnd
rlabel metal3 s 79945 62087 80043 62185 4 vdd
rlabel metal3 s 92039 62087 92137 62185 4 vdd
rlabel metal3 s 88176 61496 88274 61594 4 vdd
rlabel metal3 s 80688 61496 80786 61594 4 vdd
rlabel metal3 s 82055 62087 82153 62185 4 vdd
rlabel metal3 s 90791 62087 90889 62185 4 vdd
rlabel metal3 s 82441 62087 82539 62185 4 vdd
rlabel metal3 s 84432 61496 84530 61594 4 vdd
rlabel metal3 s 86361 66407 86459 66505 4 vdd
rlabel metal3 s 88681 62087 88779 62185 4 vdd
rlabel metal3 s 81381 67245 81479 67343 4 vdd
rlabel metal3 s 86373 67245 86471 67343 4 vdd
rlabel metal3 s 80064 61496 80162 61594 4 vdd
rlabel metal3 s 89424 61496 89522 61594 4 vdd
rlabel metal3 s 81312 61496 81410 61594 4 vdd
rlabel metal3 s 81936 61496 82034 61594 4 vdd
rlabel metal3 s 88295 62087 88393 62185 4 vdd
rlabel metal3 s 92425 62087 92523 62185 4 vdd
rlabel metal3 s 85799 62087 85897 62185 4 vdd
rlabel metal3 s 88857 66407 88955 66505 4 vdd
rlabel metal3 s 91353 66407 91451 66505 4 vdd
rlabel metal3 s 83877 67245 83975 67343 4 vdd
rlabel metal3 s 90048 61496 90146 61594 4 vdd
rlabel metal3 s 81369 66407 81467 66505 4 vdd
rlabel metal3 s 89543 62087 89641 62185 4 vdd
rlabel metal3 s 83865 66407 83963 66505 4 vdd
rlabel metal3 s 88869 67245 88967 67343 4 vdd
rlabel metal3 s 85056 61496 85154 61594 4 vdd
rlabel metal3 s 87433 62087 87531 62185 4 vdd
rlabel metal3 s 89929 62087 90027 62185 4 vdd
rlabel metal3 s 83303 62087 83401 62185 4 vdd
rlabel metal3 s 83184 61496 83282 61594 4 vdd
rlabel metal3 s 84937 62087 85035 62185 4 vdd
rlabel metal3 s 83689 62087 83787 62185 4 vdd
rlabel metal3 s 84551 62087 84649 62185 4 vdd
rlabel metal3 s 86928 61496 87026 61594 4 vdd
rlabel metal3 s 88800 61496 88898 61594 4 vdd
rlabel metal3 s 91920 61496 92018 61594 4 vdd
rlabel metal3 s 90672 61496 90770 61594 4 vdd
rlabel metal3 s 86185 62087 86283 62185 4 vdd
rlabel metal3 s 80376 63636 80474 63734 4 gnd
rlabel metal3 s 91177 62087 91275 62185 4 vdd
rlabel metal3 s 81381 67567 81479 67665 4 gnd
rlabel metal3 s 91608 63636 91706 63734 4 gnd
rlabel metal3 s 82560 61496 82658 61594 4 vdd
rlabel metal3 s 86373 67567 86471 67665 4 gnd
rlabel metal3 s 90360 63636 90458 63734 4 gnd
rlabel metal3 s 85368 63636 85466 63734 4 gnd
rlabel metal3 s 86443 65633 86541 65731 4 gnd
rlabel metal3 s 81193 62087 81291 62185 4 vdd
rlabel metal3 s 87047 62087 87145 62185 4 vdd
rlabel metal3 s 84120 63636 84218 63734 4 gnd
rlabel metal3 s 81624 63636 81722 63734 4 gnd
rlabel metal3 s 86304 61496 86402 61594 4 vdd
rlabel metal3 s 80807 62087 80905 62185 4 vdd
rlabel metal3 s 81451 65633 81549 65731 4 gnd
rlabel metal3 s 87552 61496 87650 61594 4 vdd
rlabel metal3 s 87864 63636 87962 63734 4 gnd
rlabel metal3 s 88869 67567 88967 67665 4 gnd
rlabel metal3 s 91296 61496 91394 61594 4 vdd
rlabel metal3 s 83877 67567 83975 67665 4 gnd
rlabel metal3 s 91365 67567 91463 67665 4 gnd
rlabel metal3 s 88939 65633 89037 65731 4 gnd
rlabel metal3 s 85680 61496 85778 61594 4 vdd
rlabel metal3 s 89112 63636 89210 63734 4 gnd
rlabel metal3 s 82872 63636 82970 63734 4 gnd
rlabel metal3 s 91435 65633 91533 65731 4 gnd
rlabel metal3 s 83808 61496 83906 61594 4 vdd
rlabel metal3 s 86616 63636 86714 63734 4 gnd
rlabel metal3 s 83947 65633 84045 65731 4 gnd
rlabel metal3 s 91365 67245 91463 67343 4 vdd
rlabel metal3 s 92544 61496 92642 61594 4 vdd
rlabel metal3 s 99428 59355 99526 59453 4 vdd
rlabel metal3 s 100206 57761 100304 57859 4 vdd
rlabel metal3 s 100638 56613 100736 56711 4 vdd
rlabel metal3 s 99428 58565 99526 58663 4 vdd
rlabel metal3 s 100638 59773 100736 59871 4 vdd
rlabel metal3 s 99428 56985 99526 57083 4 vdd
rlabel metal3 s 100638 56971 100736 57069 4 vdd
rlabel metal3 s 100638 57761 100736 57859 4 vdd
rlabel metal3 s 99428 57380 99526 57478 4 vdd
rlabel metal3 s 100206 58551 100304 58649 4 vdd
rlabel metal3 s 100638 58551 100736 58649 4 vdd
rlabel metal3 s 100206 57403 100304 57501 4 vdd
rlabel metal3 s 100206 58983 100304 59081 4 vdd
rlabel metal3 s 99824 57775 99922 57873 4 gnd
rlabel metal3 s 100206 58193 100304 58291 4 vdd
rlabel metal3 s 99428 58170 99526 58268 4 vdd
rlabel metal3 s 99824 60145 99922 60243 4 gnd
rlabel metal3 s 100206 56613 100304 56711 4 vdd
rlabel metal3 s 99428 60145 99526 60243 4 vdd
rlabel metal3 s 99428 57775 99526 57873 4 vdd
rlabel metal3 s 100206 60131 100304 60229 4 vdd
rlabel metal3 s 99824 56985 99922 57083 4 gnd
rlabel metal3 s 99824 56590 99922 56688 4 gnd
rlabel metal3 s 100638 59341 100736 59439 4 vdd
rlabel metal3 s 101063 59773 101161 59871 4 gnd
rlabel metal3 s 99824 56195 99922 56293 4 gnd
rlabel metal3 s 99428 58960 99526 59058 4 vdd
rlabel metal3 s 100638 58193 100736 58291 4 vdd
rlabel metal3 s 99824 59750 99922 59848 4 gnd
rlabel metal3 s 99824 57380 99922 57478 4 gnd
rlabel metal3 s 101063 60189 101161 60287 4 gnd
rlabel metal3 s 101063 56613 101161 56711 4 gnd
rlabel metal3 s 99428 59750 99526 59848 4 vdd
rlabel metal3 s 101063 58609 101161 58707 4 gnd
rlabel metal3 s 99824 58960 99922 59058 4 gnd
rlabel metal3 s 100638 60131 100736 60229 4 vdd
rlabel metal3 s 100206 56971 100304 57069 4 vdd
rlabel metal3 s 101063 58983 101161 59081 4 gnd
rlabel metal3 s 101063 56239 101161 56337 4 gnd
rlabel metal3 s 101063 59399 101161 59497 4 gnd
rlabel metal3 s 101063 57403 101161 57501 4 gnd
rlabel metal3 s 99824 58565 99922 58663 4 gnd
rlabel metal3 s 100206 59773 100304 59871 4 vdd
rlabel metal3 s 100206 59341 100304 59439 4 vdd
rlabel metal3 s 101063 57819 101161 57917 4 gnd
rlabel metal3 s 99824 59355 99922 59453 4 gnd
rlabel metal3 s 100638 57403 100736 57501 4 vdd
rlabel metal3 s 101063 58193 101161 58291 4 gnd
rlabel metal3 s 99824 58170 99922 58268 4 gnd
rlabel metal3 s 99428 56590 99526 56688 4 vdd
rlabel metal3 s 99428 56195 99526 56293 4 vdd
rlabel metal3 s 101063 57029 101161 57127 4 gnd
rlabel metal3 s 100638 58983 100736 59081 4 vdd
rlabel metal3 s 94488 59355 94586 59453 4 gnd
rlabel metal3 s 94488 57222 94586 57320 4 gnd
rlabel metal3 s 94488 58012 94586 58110 4 gnd
rlabel metal3 s 94488 58565 94586 58663 4 gnd
rlabel metal3 s 94488 58802 94586 58900 4 gnd
rlabel metal3 s 94488 56432 94586 56530 4 gnd
rlabel metal3 s 94488 59592 94586 59690 4 gnd
rlabel metal3 s 94488 56195 94586 56293 4 gnd
rlabel metal3 s 94488 60145 94586 60243 4 gnd
rlabel metal3 s 94488 56985 94586 57083 4 gnd
rlabel metal3 s 94488 58328 94586 58426 4 gnd
rlabel metal3 s 94488 57775 94586 57873 4 gnd
rlabel metal3 s 94488 57538 94586 57636 4 gnd
rlabel metal3 s 94488 59908 94586 60006 4 gnd
rlabel metal3 s 94488 59118 94586 59216 4 gnd
rlabel metal3 s 94488 56748 94586 56846 4 gnd
rlabel metal3 s 94488 60382 94586 60480 4 gnd
rlabel metal3 s 94488 53272 94586 53370 4 gnd
rlabel metal3 s 94488 55958 94586 56056 4 gnd
rlabel metal3 s 94488 55405 94586 55503 4 gnd
rlabel metal3 s 94488 54852 94586 54950 4 gnd
rlabel metal3 s 94488 52798 94586 52896 4 gnd
rlabel metal3 s 94488 52482 94586 52580 4 gnd
rlabel metal3 s 94488 54062 94586 54160 4 gnd
rlabel metal3 s 94488 52245 94586 52343 4 gnd
rlabel metal3 s 94488 55642 94586 55740 4 gnd
rlabel metal3 s 94488 54378 94586 54476 4 gnd
rlabel metal3 s 94488 54615 94586 54713 4 gnd
rlabel metal3 s 94488 52008 94586 52106 4 gnd
rlabel metal3 s 94488 53035 94586 53133 4 gnd
rlabel metal3 s 94488 53825 94586 53923 4 gnd
rlabel metal3 s 94488 55168 94586 55266 4 gnd
rlabel metal3 s 94488 53588 94586 53686 4 gnd
rlabel metal3 s 101063 54659 101161 54757 4 gnd
rlabel metal3 s 99824 55010 99922 55108 4 gnd
rlabel metal3 s 99428 54615 99526 54713 4 vdd
rlabel metal3 s 100206 52663 100304 52761 4 vdd
rlabel metal3 s 100638 53811 100736 53909 4 vdd
rlabel metal3 s 100638 55823 100736 55921 4 vdd
rlabel metal3 s 99428 53035 99526 53133 4 vdd
rlabel metal3 s 100206 55823 100304 55921 4 vdd
rlabel metal3 s 99824 53035 99922 53133 4 gnd
rlabel metal3 s 99428 55405 99526 55503 4 vdd
rlabel metal3 s 101063 52289 101161 52387 4 gnd
rlabel metal3 s 100638 55033 100736 55131 4 vdd
rlabel metal3 s 100206 55391 100304 55489 4 vdd
rlabel metal3 s 101063 54243 101161 54341 4 gnd
rlabel metal3 s 100638 54243 100736 54341 4 vdd
rlabel metal3 s 100638 56181 100736 56279 4 vdd
rlabel metal3 s 101063 51873 101161 51971 4 gnd
rlabel metal3 s 101063 55449 101161 55547 4 gnd
rlabel metal3 s 99428 53825 99526 53923 4 vdd
rlabel metal3 s 99428 55010 99526 55108 4 vdd
rlabel metal3 s 100638 53453 100736 53551 4 vdd
rlabel metal3 s 99824 54615 99922 54713 4 gnd
rlabel metal3 s 100638 54601 100736 54699 4 vdd
rlabel metal3 s 100206 53021 100304 53119 4 vdd
rlabel metal3 s 100638 55391 100736 55489 4 vdd
rlabel metal3 s 100206 51873 100304 51971 4 vdd
rlabel metal3 s 99824 55800 99922 55898 4 gnd
rlabel metal3 s 100638 51873 100736 51971 4 vdd
rlabel metal3 s 100206 55033 100304 55131 4 vdd
rlabel metal3 s 100638 52231 100736 52329 4 vdd
rlabel metal3 s 99428 52640 99526 52738 4 vdd
rlabel metal3 s 99824 55405 99922 55503 4 gnd
rlabel metal3 s 99824 53430 99922 53528 4 gnd
rlabel metal3 s 100206 54601 100304 54699 4 vdd
rlabel metal3 s 101063 55823 101161 55921 4 gnd
rlabel metal3 s 100206 56181 100304 56279 4 vdd
rlabel metal3 s 99428 52245 99526 52343 4 vdd
rlabel metal3 s 99428 54220 99526 54318 4 vdd
rlabel metal3 s 99824 52640 99922 52738 4 gnd
rlabel metal3 s 101063 53869 101161 53967 4 gnd
rlabel metal3 s 101063 55033 101161 55131 4 gnd
rlabel metal3 s 101063 53079 101161 53177 4 gnd
rlabel metal3 s 99428 53430 99526 53528 4 vdd
rlabel metal3 s 101063 53453 101161 53551 4 gnd
rlabel metal3 s 100206 52231 100304 52329 4 vdd
rlabel metal3 s 99824 52245 99922 52343 4 gnd
rlabel metal3 s 99824 54220 99922 54318 4 gnd
rlabel metal3 s 100206 53811 100304 53909 4 vdd
rlabel metal3 s 100638 52663 100736 52761 4 vdd
rlabel metal3 s 99824 53825 99922 53923 4 gnd
rlabel metal3 s 100206 53453 100304 53551 4 vdd
rlabel metal3 s 100638 53021 100736 53119 4 vdd
rlabel metal3 s 101063 52663 101161 52761 4 gnd
rlabel metal3 s 99428 55800 99526 55898 4 vdd
rlabel metal3 s 100206 54243 100304 54341 4 vdd
rlabel metal3 s 76632 63636 76730 63734 4 gnd
rlabel metal3 s 79440 61496 79538 61594 4 vdd
rlabel metal3 s 72888 63636 72986 63734 4 gnd
rlabel metal3 s 71397 67245 71495 67343 4 vdd
rlabel metal3 s 78885 67567 78983 67665 4 gnd
rlabel metal3 s 75696 61496 75794 61594 4 vdd
rlabel metal3 s 77880 63636 77978 63734 4 gnd
rlabel metal3 s 78885 67245 78983 67343 4 vdd
rlabel metal3 s 73893 67567 73991 67665 4 gnd
rlabel metal3 s 74953 62087 75051 62185 4 vdd
rlabel metal3 s 67584 61496 67682 61594 4 vdd
rlabel metal3 s 71385 66407 71483 66505 4 vdd
rlabel metal3 s 76389 67567 76487 67665 4 gnd
rlabel metal3 s 78955 65633 79053 65731 4 gnd
rlabel metal3 s 75072 61496 75170 61594 4 vdd
rlabel metal3 s 66960 61496 67058 61594 4 vdd
rlabel metal3 s 67079 62087 67177 62185 4 vdd
rlabel metal3 s 68901 67567 68999 67665 4 gnd
rlabel metal3 s 78311 62087 78409 62185 4 vdd
rlabel metal3 s 72071 62087 72169 62185 4 vdd
rlabel metal3 s 68208 61496 68306 61594 4 vdd
rlabel metal3 s 76320 61496 76418 61594 4 vdd
rlabel metal3 s 66648 63636 66746 63734 4 gnd
rlabel metal3 s 67465 62087 67563 62185 4 vdd
rlabel metal3 s 78873 66407 78971 66505 4 vdd
rlabel metal3 s 73319 62087 73417 62185 4 vdd
rlabel metal3 s 68901 67245 68999 67343 4 vdd
rlabel metal3 s 69575 62087 69673 62185 4 vdd
rlabel metal3 s 71397 67567 71495 67665 4 gnd
rlabel metal3 s 73200 61496 73298 61594 4 vdd
rlabel metal3 s 73963 65633 74061 65731 4 gnd
rlabel metal3 s 69456 61496 69554 61594 4 vdd
rlabel metal3 s 73881 66407 73979 66505 4 vdd
rlabel metal3 s 77063 62087 77161 62185 4 vdd
rlabel metal3 s 72576 61496 72674 61594 4 vdd
rlabel metal3 s 69144 63636 69242 63734 4 gnd
rlabel metal3 s 79559 62087 79657 62185 4 vdd
rlabel metal3 s 78816 61496 78914 61594 4 vdd
rlabel metal3 s 67896 63636 67994 63734 4 gnd
rlabel metal3 s 74567 62087 74665 62185 4 vdd
rlabel metal3 s 71467 65633 71565 65731 4 gnd
rlabel metal3 s 70080 61496 70178 61594 4 vdd
rlabel metal3 s 74448 61496 74546 61594 4 vdd
rlabel metal3 s 70823 62087 70921 62185 4 vdd
rlabel metal3 s 68832 61496 68930 61594 4 vdd
rlabel metal3 s 75384 63636 75482 63734 4 gnd
rlabel metal3 s 78697 62087 78795 62185 4 vdd
rlabel metal3 s 76201 62087 76299 62185 4 vdd
rlabel metal3 s 76944 61496 77042 61594 4 vdd
rlabel metal3 s 73824 61496 73922 61594 4 vdd
rlabel metal3 s 76459 65633 76557 65731 4 gnd
rlabel metal3 s 70392 63636 70490 63734 4 gnd
rlabel metal3 s 71328 61496 71426 61594 4 vdd
rlabel metal3 s 79128 63636 79226 63734 4 gnd
rlabel metal3 s 75815 62087 75913 62185 4 vdd
rlabel metal3 s 77449 62087 77547 62185 4 vdd
rlabel metal3 s 69961 62087 70059 62185 4 vdd
rlabel metal3 s 68713 62087 68811 62185 4 vdd
rlabel metal3 s 73705 62087 73803 62185 4 vdd
rlabel metal3 s 68889 66407 68987 66505 4 vdd
rlabel metal3 s 76377 66407 76475 66505 4 vdd
rlabel metal3 s 71952 61496 72050 61594 4 vdd
rlabel metal3 s 70704 61496 70802 61594 4 vdd
rlabel metal3 s 71640 63636 71738 63734 4 gnd
rlabel metal3 s 71209 62087 71307 62185 4 vdd
rlabel metal3 s 78192 61496 78290 61594 4 vdd
rlabel metal3 s 68327 62087 68425 62185 4 vdd
rlabel metal3 s 77568 61496 77666 61594 4 vdd
rlabel metal3 s 72457 62087 72555 62185 4 vdd
rlabel metal3 s 74136 63636 74234 63734 4 gnd
rlabel metal3 s 73893 67245 73991 67343 4 vdd
rlabel metal3 s 76389 67245 76487 67343 4 vdd
rlabel metal3 s 68971 65633 69069 65731 4 gnd
rlabel metal3 s 59591 62087 59689 62185 4 vdd
rlabel metal3 s 53995 65633 54093 65731 4 gnd
rlabel metal3 s 58905 66407 59003 66505 4 vdd
rlabel metal3 s 61401 66407 61499 66505 4 vdd
rlabel metal3 s 58224 61496 58322 61594 4 vdd
rlabel metal3 s 55847 62087 55945 62185 4 vdd
rlabel metal3 s 54599 62087 54697 62185 4 vdd
rlabel metal3 s 53913 66407 54011 66505 4 vdd
rlabel metal3 s 61413 67567 61511 67665 4 gnd
rlabel metal3 s 58343 62087 58441 62185 4 vdd
rlabel metal3 s 58917 67245 59015 67343 4 vdd
rlabel metal3 s 63897 66407 63995 66505 4 vdd
rlabel metal3 s 61413 67245 61511 67343 4 vdd
rlabel metal3 s 66405 67567 66503 67665 4 gnd
rlabel metal3 s 63840 61496 63938 61594 4 vdd
rlabel metal3 s 61656 63636 61754 63734 4 gnd
rlabel metal3 s 54480 61496 54578 61594 4 vdd
rlabel metal3 s 55104 61496 55202 61594 4 vdd
rlabel metal3 s 62087 62087 62185 62185 4 vdd
rlabel metal3 s 63335 62087 63433 62185 4 vdd
rlabel metal3 s 63909 67245 64007 67343 4 vdd
rlabel metal3 s 53737 62087 53835 62185 4 vdd
rlabel metal3 s 61225 62087 61323 62185 4 vdd
rlabel metal3 s 54985 62087 55083 62185 4 vdd
rlabel metal3 s 64464 61496 64562 61594 4 vdd
rlabel metal3 s 60720 61496 60818 61594 4 vdd
rlabel metal3 s 53925 67245 54023 67343 4 vdd
rlabel metal3 s 66217 62087 66315 62185 4 vdd
rlabel metal3 s 60839 62087 60937 62185 4 vdd
rlabel metal3 s 56233 62087 56331 62185 4 vdd
rlabel metal3 s 57912 63636 58010 63734 4 gnd
rlabel metal3 s 63909 67567 64007 67665 4 gnd
rlabel metal3 s 53925 67567 54023 67665 4 gnd
rlabel metal3 s 64969 62087 65067 62185 4 vdd
rlabel metal3 s 58917 67567 59015 67665 4 gnd
rlabel metal3 s 61968 61496 62066 61594 4 vdd
rlabel metal3 s 58729 62087 58827 62185 4 vdd
rlabel metal3 s 57600 61496 57698 61594 4 vdd
rlabel metal3 s 56421 67245 56519 67343 4 vdd
rlabel metal3 s 66405 67245 66503 67343 4 vdd
rlabel metal3 s 55728 61496 55826 61594 4 vdd
rlabel metal3 s 57095 62087 57193 62185 4 vdd
rlabel metal3 s 63216 61496 63314 61594 4 vdd
rlabel metal3 s 58848 61496 58946 61594 4 vdd
rlabel metal3 s 59977 62087 60075 62185 4 vdd
rlabel metal3 s 54168 63636 54266 63734 4 gnd
rlabel metal3 s 64583 62087 64681 62185 4 vdd
rlabel metal3 s 62473 62087 62571 62185 4 vdd
rlabel metal3 s 53856 61496 53954 61594 4 vdd
rlabel metal3 s 60408 63636 60506 63734 4 gnd
rlabel metal3 s 65712 61496 65810 61594 4 vdd
rlabel metal3 s 62592 61496 62690 61594 4 vdd
rlabel metal3 s 60096 61496 60194 61594 4 vdd
rlabel metal3 s 65088 61496 65186 61594 4 vdd
rlabel metal3 s 56664 63636 56762 63734 4 gnd
rlabel metal3 s 56409 66407 56507 66505 4 vdd
rlabel metal3 s 62904 63636 63002 63734 4 gnd
rlabel metal3 s 55416 63636 55514 63734 4 gnd
rlabel metal3 s 56976 61496 57074 61594 4 vdd
rlabel metal3 s 61483 65633 61581 65731 4 gnd
rlabel metal3 s 57481 62087 57579 62185 4 vdd
rlabel metal3 s 59472 61496 59570 61594 4 vdd
rlabel metal3 s 64152 63636 64250 63734 4 gnd
rlabel metal3 s 66336 61496 66434 61594 4 vdd
rlabel metal3 s 59160 63636 59258 63734 4 gnd
rlabel metal3 s 58987 65633 59085 65731 4 gnd
rlabel metal3 s 56491 65633 56589 65731 4 gnd
rlabel metal3 s 66393 66407 66491 66505 4 vdd
rlabel metal3 s 56421 67567 56519 67665 4 gnd
rlabel metal3 s 66475 65633 66573 65731 4 gnd
rlabel metal3 s 56352 61496 56450 61594 4 vdd
rlabel metal3 s 63979 65633 64077 65731 4 gnd
rlabel metal3 s 63721 62087 63819 62185 4 vdd
rlabel metal3 s 61344 61496 61442 61594 4 vdd
rlabel metal3 s 65831 62087 65929 62185 4 vdd
rlabel metal3 s 65400 63636 65498 63734 4 gnd
rlabel metal3 s 99824 51060 99922 51158 4 gnd
rlabel metal3 s 99824 49480 99922 49578 4 gnd
rlabel metal3 s 99428 47900 99526 47998 4 vdd
rlabel metal3 s 99824 48690 99922 48788 4 gnd
rlabel metal3 s 100206 48281 100304 48379 4 vdd
rlabel metal3 s 100206 49071 100304 49169 4 vdd
rlabel metal3 s 101063 51499 101161 51597 4 gnd
rlabel metal3 s 101063 51083 101161 51181 4 gnd
rlabel metal3 s 100638 48713 100736 48811 4 vdd
rlabel metal3 s 100638 47923 100736 48021 4 vdd
rlabel metal3 s 99428 51455 99526 51553 4 vdd
rlabel metal3 s 100638 48281 100736 48379 4 vdd
rlabel metal3 s 100638 49071 100736 49169 4 vdd
rlabel metal3 s 100638 51441 100736 51539 4 vdd
rlabel metal3 s 101063 48713 101161 48811 4 gnd
rlabel metal3 s 100638 49503 100736 49601 4 vdd
rlabel metal3 s 100638 50651 100736 50749 4 vdd
rlabel metal3 s 100638 51083 100736 51181 4 vdd
rlabel metal3 s 100206 50651 100304 50749 4 vdd
rlabel metal3 s 100206 51441 100304 51539 4 vdd
rlabel metal3 s 99428 50270 99526 50368 4 vdd
rlabel metal3 s 100206 47923 100304 48021 4 vdd
rlabel metal3 s 100206 48713 100304 48811 4 vdd
rlabel metal3 s 99428 48295 99526 48393 4 vdd
rlabel metal3 s 101063 48339 101161 48437 4 gnd
rlabel metal3 s 99428 51060 99526 51158 4 vdd
rlabel metal3 s 101063 49919 101161 50017 4 gnd
rlabel metal3 s 99824 51455 99922 51553 4 gnd
rlabel metal3 s 99428 51850 99526 51948 4 vdd
rlabel metal3 s 101063 50293 101161 50391 4 gnd
rlabel metal3 s 100638 50293 100736 50391 4 vdd
rlabel metal3 s 100206 49861 100304 49959 4 vdd
rlabel metal3 s 100206 50293 100304 50391 4 vdd
rlabel metal3 s 99428 49875 99526 49973 4 vdd
rlabel metal3 s 100206 49503 100304 49601 4 vdd
rlabel metal3 s 101063 49129 101161 49227 4 gnd
rlabel metal3 s 99428 50665 99526 50763 4 vdd
rlabel metal3 s 101063 49503 101161 49601 4 gnd
rlabel metal3 s 99824 50270 99922 50368 4 gnd
rlabel metal3 s 99824 48295 99922 48393 4 gnd
rlabel metal3 s 101063 47923 101161 48021 4 gnd
rlabel metal3 s 100638 49861 100736 49959 4 vdd
rlabel metal3 s 100206 51083 100304 51181 4 vdd
rlabel metal3 s 99824 49085 99922 49183 4 gnd
rlabel metal3 s 99824 51850 99922 51948 4 gnd
rlabel metal3 s 99824 49875 99922 49973 4 gnd
rlabel metal3 s 99428 48690 99526 48788 4 vdd
rlabel metal3 s 101063 50709 101161 50807 4 gnd
rlabel metal3 s 99428 49085 99526 49183 4 vdd
rlabel metal3 s 99824 50665 99922 50763 4 gnd
rlabel metal3 s 99824 47900 99922 47998 4 gnd
rlabel metal3 s 99428 49480 99526 49578 4 vdd
rlabel metal3 s 101063 47549 101161 47647 4 gnd
rlabel metal3 s 94488 48295 94586 48393 4 gnd
rlabel metal3 s 94488 48058 94586 48156 4 gnd
rlabel metal3 s 94488 49085 94586 49183 4 gnd
rlabel metal3 s 94488 51218 94586 51316 4 gnd
rlabel metal3 s 94488 49322 94586 49420 4 gnd
rlabel metal3 s 94488 49638 94586 49736 4 gnd
rlabel metal3 s 94488 49875 94586 49973 4 gnd
rlabel metal3 s 94488 50902 94586 51000 4 gnd
rlabel metal3 s 94488 47742 94586 47840 4 gnd
rlabel metal3 s 94488 50665 94586 50763 4 gnd
rlabel metal3 s 94488 50428 94586 50526 4 gnd
rlabel metal3 s 94488 51455 94586 51553 4 gnd
rlabel metal3 s 94488 48848 94586 48946 4 gnd
rlabel metal3 s 94488 48532 94586 48630 4 gnd
rlabel metal3 s 94488 50112 94586 50210 4 gnd
rlabel metal3 s 94488 51692 94586 51790 4 gnd
rlabel metal3 s 94488 43555 94586 43653 4 gnd
rlabel metal3 s 94488 46478 94586 46576 4 gnd
rlabel metal3 s 94488 45688 94586 45786 4 gnd
rlabel metal3 s 94488 46952 94586 47050 4 gnd
rlabel metal3 s 94488 43318 94586 43416 4 gnd
rlabel metal3 s 94488 46162 94586 46260 4 gnd
rlabel metal3 s 94488 45135 94586 45233 4 gnd
rlabel metal3 s 94488 44108 94586 44206 4 gnd
rlabel metal3 s 94488 45372 94586 45470 4 gnd
rlabel metal3 s 94488 46715 94586 46813 4 gnd
rlabel metal3 s 94488 47505 94586 47603 4 gnd
rlabel metal3 s 94488 47268 94586 47366 4 gnd
rlabel metal3 s 94488 43792 94586 43890 4 gnd
rlabel metal3 s 94488 45925 94586 46023 4 gnd
rlabel metal3 s 94488 44345 94586 44443 4 gnd
rlabel metal3 s 94488 44898 94586 44996 4 gnd
rlabel metal3 s 94488 44582 94586 44680 4 gnd
rlabel metal3 s 101063 46759 101161 46857 4 gnd
rlabel metal3 s 101063 43973 101161 44071 4 gnd
rlabel metal3 s 100638 43973 100736 44071 4 vdd
rlabel metal3 s 101063 45179 101161 45277 4 gnd
rlabel metal3 s 100638 44763 100736 44861 4 vdd
rlabel metal3 s 99824 47505 99922 47603 4 gnd
rlabel metal3 s 101063 44763 101161 44861 4 gnd
rlabel metal3 s 100638 46701 100736 46799 4 vdd
rlabel metal3 s 99824 43950 99922 44048 4 gnd
rlabel metal3 s 100206 47133 100304 47231 4 vdd
rlabel metal3 s 100206 45911 100304 46009 4 vdd
rlabel metal3 s 100206 44763 100304 44861 4 vdd
rlabel metal3 s 100206 44331 100304 44429 4 vdd
rlabel metal3 s 99428 45925 99526 46023 4 vdd
rlabel metal3 s 100638 44331 100736 44429 4 vdd
rlabel metal3 s 100206 46701 100304 46799 4 vdd
rlabel metal3 s 99428 44345 99526 44443 4 vdd
rlabel metal3 s 99428 46320 99526 46418 4 vdd
rlabel metal3 s 99428 47505 99526 47603 4 vdd
rlabel metal3 s 100206 47491 100304 47589 4 vdd
rlabel metal3 s 100638 47491 100736 47589 4 vdd
rlabel metal3 s 101063 45553 101161 45651 4 gnd
rlabel metal3 s 99428 47110 99526 47208 4 vdd
rlabel metal3 s 99428 45135 99526 45233 4 vdd
rlabel metal3 s 100206 45121 100304 45219 4 vdd
rlabel metal3 s 99824 45925 99922 46023 4 gnd
rlabel metal3 s 99824 46320 99922 46418 4 gnd
rlabel metal3 s 99824 44345 99922 44443 4 gnd
rlabel metal3 s 101063 43599 101161 43697 4 gnd
rlabel metal3 s 100638 46343 100736 46441 4 vdd
rlabel metal3 s 100206 43973 100304 44071 4 vdd
rlabel metal3 s 101063 46343 101161 46441 4 gnd
rlabel metal3 s 99428 46715 99526 46813 4 vdd
rlabel metal3 s 101063 47133 101161 47231 4 gnd
rlabel metal3 s 100638 45121 100736 45219 4 vdd
rlabel metal3 s 99824 44740 99922 44838 4 gnd
rlabel metal3 s 99428 43950 99526 44048 4 vdd
rlabel metal3 s 99428 43555 99526 43653 4 vdd
rlabel metal3 s 100206 45553 100304 45651 4 vdd
rlabel metal3 s 100206 43541 100304 43639 4 vdd
rlabel metal3 s 99824 43555 99922 43653 4 gnd
rlabel metal3 s 99824 46715 99922 46813 4 gnd
rlabel metal3 s 100638 45911 100736 46009 4 vdd
rlabel metal3 s 100638 47133 100736 47231 4 vdd
rlabel metal3 s 99428 44740 99526 44838 4 vdd
rlabel metal3 s 99824 45135 99922 45233 4 gnd
rlabel metal3 s 99428 45530 99526 45628 4 vdd
rlabel metal3 s 100638 45553 100736 45651 4 vdd
rlabel metal3 s 99824 45530 99922 45628 4 gnd
rlabel metal3 s 101063 44389 101161 44487 4 gnd
rlabel metal3 s 99824 47110 99922 47208 4 gnd
rlabel metal3 s 101063 45969 101161 46067 4 gnd
rlabel metal3 s 100638 43541 100736 43639 4 vdd
rlabel metal3 s 100206 46343 100304 46441 4 vdd
rlabel metal3 s 101063 39233 101161 39331 4 gnd
rlabel metal3 s 100206 40023 100304 40121 4 vdd
rlabel metal3 s 100206 40381 100304 40479 4 vdd
rlabel metal3 s 101063 41229 101161 41327 4 gnd
rlabel metal3 s 99428 40000 99526 40098 4 vdd
rlabel metal3 s 99824 39210 99922 39308 4 gnd
rlabel metal3 s 99428 41580 99526 41678 4 vdd
rlabel metal3 s 99824 42370 99922 42468 4 gnd
rlabel metal3 s 99824 41580 99922 41678 4 gnd
rlabel metal3 s 99824 40395 99922 40493 4 gnd
rlabel metal3 s 100638 41171 100736 41269 4 vdd
rlabel metal3 s 100206 39591 100304 39689 4 vdd
rlabel metal3 s 100206 41961 100304 42059 4 vdd
rlabel metal3 s 100638 42751 100736 42849 4 vdd
rlabel metal3 s 100638 39233 100736 39331 4 vdd
rlabel metal3 s 99428 42370 99526 42468 4 vdd
rlabel metal3 s 100638 43183 100736 43281 4 vdd
rlabel metal3 s 100206 42393 100304 42491 4 vdd
rlabel metal3 s 101063 41603 101161 41701 4 gnd
rlabel metal3 s 101063 43183 101161 43281 4 gnd
rlabel metal3 s 99428 40790 99526 40888 4 vdd
rlabel metal3 s 99824 43160 99922 43258 4 gnd
rlabel metal3 s 101063 40023 101161 40121 4 gnd
rlabel metal3 s 99428 39210 99526 39308 4 vdd
rlabel metal3 s 100206 40813 100304 40911 4 vdd
rlabel metal3 s 100638 41603 100736 41701 4 vdd
rlabel metal3 s 100638 39591 100736 39689 4 vdd
rlabel metal3 s 99428 40395 99526 40493 4 vdd
rlabel metal3 s 99824 41185 99922 41283 4 gnd
rlabel metal3 s 99428 41185 99526 41283 4 vdd
rlabel metal3 s 99824 41975 99922 42073 4 gnd
rlabel metal3 s 99428 41975 99526 42073 4 vdd
rlabel metal3 s 100206 41603 100304 41701 4 vdd
rlabel metal3 s 100206 42751 100304 42849 4 vdd
rlabel metal3 s 99428 42765 99526 42863 4 vdd
rlabel metal3 s 99428 43160 99526 43258 4 vdd
rlabel metal3 s 101063 39649 101161 39747 4 gnd
rlabel metal3 s 99428 39605 99526 39703 4 vdd
rlabel metal3 s 101063 40813 101161 40911 4 gnd
rlabel metal3 s 101063 42019 101161 42117 4 gnd
rlabel metal3 s 99824 42765 99922 42863 4 gnd
rlabel metal3 s 100206 43183 100304 43281 4 vdd
rlabel metal3 s 100206 39233 100304 39331 4 vdd
rlabel metal3 s 100638 40813 100736 40911 4 vdd
rlabel metal3 s 100638 42393 100736 42491 4 vdd
rlabel metal3 s 99824 39605 99922 39703 4 gnd
rlabel metal3 s 101063 42809 101161 42907 4 gnd
rlabel metal3 s 99824 40000 99922 40098 4 gnd
rlabel metal3 s 99824 40790 99922 40888 4 gnd
rlabel metal3 s 100638 40381 100736 40479 4 vdd
rlabel metal3 s 101063 42393 101161 42491 4 gnd
rlabel metal3 s 100206 41171 100304 41269 4 vdd
rlabel metal3 s 100638 40023 100736 40121 4 vdd
rlabel metal3 s 101063 40439 101161 40537 4 gnd
rlabel metal3 s 100638 41961 100736 42059 4 vdd
rlabel metal3 s 94488 40158 94586 40256 4 gnd
rlabel metal3 s 94488 39842 94586 39940 4 gnd
rlabel metal3 s 94488 42212 94586 42310 4 gnd
rlabel metal3 s 94488 39052 94586 39150 4 gnd
rlabel metal3 s 94488 42765 94586 42863 4 gnd
rlabel metal3 s 94488 39605 94586 39703 4 gnd
rlabel metal3 s 94488 40632 94586 40730 4 gnd
rlabel metal3 s 94488 42528 94586 42626 4 gnd
rlabel metal3 s 94488 41975 94586 42073 4 gnd
rlabel metal3 s 94488 43002 94586 43100 4 gnd
rlabel metal3 s 94488 40948 94586 41046 4 gnd
rlabel metal3 s 94488 40395 94586 40493 4 gnd
rlabel metal3 s 94488 41738 94586 41836 4 gnd
rlabel metal3 s 94488 41422 94586 41520 4 gnd
rlabel metal3 s 94488 39368 94586 39466 4 gnd
rlabel metal3 s 94488 41185 94586 41283 4 gnd
rlabel metal3 s 94488 34865 94586 34963 4 gnd
rlabel metal3 s 94488 34628 94586 34726 4 gnd
rlabel metal3 s 94488 36682 94586 36780 4 gnd
rlabel metal3 s 98571 35639 98669 35737 4 vdd
rlabel metal3 s 94488 38262 94586 38360 4 gnd
rlabel metal3 s 94488 38815 94586 38913 4 gnd
rlabel metal3 s 94488 38578 94586 38676 4 gnd
rlabel metal3 s 94488 35892 94586 35990 4 gnd
rlabel metal3 s 94488 35655 94586 35753 4 gnd
rlabel metal3 s 94488 37788 94586 37886 4 gnd
rlabel metal3 s 97528 35655 97626 35753 4 gnd
rlabel metal3 s 94488 35418 94586 35516 4 gnd
rlabel metal3 s 94488 36208 94586 36306 4 gnd
rlabel metal3 s 94488 38025 94586 38123 4 gnd
rlabel metal3 s 94488 36998 94586 37096 4 gnd
rlabel metal3 s 94488 37472 94586 37570 4 gnd
rlabel metal3 s 94488 35102 94586 35200 4 gnd
rlabel metal3 s 94488 36445 94586 36543 4 gnd
rlabel metal3 s 95880 35655 95978 35753 4 vdd
rlabel metal3 s 98996 35640 99094 35738 4 gnd
rlabel metal3 s 94488 37235 94586 37333 4 gnd
rlabel metal3 s 100638 36863 100736 36961 4 vdd
rlabel metal3 s 101063 36073 101161 36171 4 gnd
rlabel metal3 s 99428 38815 99526 38913 4 vdd
rlabel metal3 s 99824 35655 99922 35753 4 gnd
rlabel metal3 s 100206 36863 100304 36961 4 vdd
rlabel metal3 s 101063 38069 101161 38167 4 gnd
rlabel metal3 s 100206 38011 100304 38109 4 vdd
rlabel metal3 s 100206 37653 100304 37751 4 vdd
rlabel metal3 s 100638 36073 100736 36171 4 vdd
rlabel metal3 s 99428 38420 99526 38518 4 vdd
rlabel metal3 s 99428 36840 99526 36938 4 vdd
rlabel metal3 s 100638 36431 100736 36529 4 vdd
rlabel metal3 s 99428 36445 99526 36543 4 vdd
rlabel metal3 s 100206 34851 100304 34949 4 vdd
rlabel metal3 s 99428 34865 99526 34963 4 vdd
rlabel metal3 s 99824 37630 99922 37728 4 gnd
rlabel metal3 s 101063 36489 101161 36587 4 gnd
rlabel metal3 s 99824 38815 99922 38913 4 gnd
rlabel metal3 s 99824 36445 99922 36543 4 gnd
rlabel metal3 s 100638 34851 100736 34949 4 vdd
rlabel metal3 s 100206 36431 100304 36529 4 vdd
rlabel metal3 s 100638 35641 100736 35739 4 vdd
rlabel metal3 s 100638 38011 100736 38109 4 vdd
rlabel metal3 s 100206 38443 100304 38541 4 vdd
rlabel metal3 s 100638 37221 100736 37319 4 vdd
rlabel metal3 s 99824 37235 99922 37333 4 gnd
rlabel metal3 s 100638 38801 100736 38899 4 vdd
rlabel metal3 s 101063 35283 101161 35381 4 gnd
rlabel metal3 s 99824 36840 99922 36938 4 gnd
rlabel metal3 s 99428 36050 99526 36148 4 vdd
rlabel metal3 s 99824 38420 99922 38518 4 gnd
rlabel metal3 s 100206 36073 100304 36171 4 vdd
rlabel metal3 s 99824 34865 99922 34963 4 gnd
rlabel metal3 s 99428 37630 99526 37728 4 vdd
rlabel metal3 s 100638 38443 100736 38541 4 vdd
rlabel metal3 s 100638 35283 100736 35381 4 vdd
rlabel metal3 s 99824 35260 99922 35358 4 gnd
rlabel metal3 s 99824 38025 99922 38123 4 gnd
rlabel metal3 s 101063 35699 101161 35797 4 gnd
rlabel metal3 s 101063 38443 101161 38541 4 gnd
rlabel metal3 s 101063 34909 101161 35007 4 gnd
rlabel metal3 s 100638 37653 100736 37751 4 vdd
rlabel metal3 s 99428 35655 99526 35753 4 vdd
rlabel metal3 s 101063 37279 101161 37377 4 gnd
rlabel metal3 s 100206 38801 100304 38899 4 vdd
rlabel metal3 s 101063 36863 101161 36961 4 gnd
rlabel metal3 s 99428 38025 99526 38123 4 vdd
rlabel metal3 s 99428 37235 99526 37333 4 vdd
rlabel metal3 s 101063 37653 101161 37751 4 gnd
rlabel metal3 s 100206 35641 100304 35739 4 vdd
rlabel metal3 s 101063 38859 101161 38957 4 gnd
rlabel metal3 s 100206 35283 100304 35381 4 vdd
rlabel metal3 s 99428 35260 99526 35358 4 vdd
rlabel metal3 s 100206 37221 100304 37319 4 vdd
rlabel metal3 s 99824 36050 99922 36148 4 gnd
rlabel metal3 s 45001 62087 45099 62185 4 vdd
rlabel metal3 s 42119 62087 42217 62185 4 vdd
rlabel metal3 s 51984 61496 52082 61594 4 vdd
rlabel metal3 s 41445 67245 41543 67343 4 vdd
rlabel metal3 s 52608 61496 52706 61594 4 vdd
rlabel metal3 s 51417 66407 51515 66505 4 vdd
rlabel metal3 s 51429 67245 51527 67343 4 vdd
rlabel metal3 s 40752 61496 40850 61594 4 vdd
rlabel metal3 s 53232 61496 53330 61594 4 vdd
rlabel metal3 s 46992 61496 47090 61594 4 vdd
rlabel metal3 s 44184 63636 44282 63734 4 gnd
rlabel metal3 s 50855 62087 50953 62185 4 vdd
rlabel metal3 s 46249 62087 46347 62185 4 vdd
rlabel metal3 s 52920 63636 53018 63734 4 gnd
rlabel metal3 s 51429 67567 51527 67665 4 gnd
rlabel metal3 s 44496 61496 44594 61594 4 vdd
rlabel metal3 s 47497 62087 47595 62185 4 vdd
rlabel metal3 s 47616 61496 47714 61594 4 vdd
rlabel metal3 s 42505 62087 42603 62185 4 vdd
rlabel metal3 s 52489 62087 52587 62185 4 vdd
rlabel metal3 s 51499 65633 51597 65731 4 gnd
rlabel metal3 s 51672 63636 51770 63734 4 gnd
rlabel metal3 s 41433 66407 41531 66505 4 vdd
rlabel metal3 s 48864 61496 48962 61594 4 vdd
rlabel metal3 s 45120 61496 45218 61594 4 vdd
rlabel metal3 s 50424 63636 50522 63734 4 gnd
rlabel metal3 s 40871 62087 40969 62185 4 vdd
rlabel metal3 s 45744 61496 45842 61594 4 vdd
rlabel metal3 s 49607 62087 49705 62185 4 vdd
rlabel metal3 s 42936 63636 43034 63734 4 gnd
rlabel metal3 s 52103 62087 52201 62185 4 vdd
rlabel metal3 s 43872 61496 43970 61594 4 vdd
rlabel metal3 s 48933 67567 49031 67665 4 gnd
rlabel metal3 s 46680 63636 46778 63734 4 gnd
rlabel metal3 s 50736 61496 50834 61594 4 vdd
rlabel metal3 s 41688 63636 41786 63734 4 gnd
rlabel metal3 s 44011 65633 44109 65731 4 gnd
rlabel metal3 s 43248 61496 43346 61594 4 vdd
rlabel metal3 s 49993 62087 50091 62185 4 vdd
rlabel metal3 s 48240 61496 48338 61594 4 vdd
rlabel metal3 s 41445 67567 41543 67665 4 gnd
rlabel metal3 s 43929 66407 44027 66505 4 vdd
rlabel metal3 s 48933 67245 49031 67343 4 vdd
rlabel metal3 s 42624 61496 42722 61594 4 vdd
rlabel metal3 s 53351 62087 53449 62185 4 vdd
rlabel metal3 s 46507 65633 46605 65731 4 gnd
rlabel metal3 s 43367 62087 43465 62185 4 vdd
rlabel metal3 s 45432 63636 45530 63734 4 gnd
rlabel metal3 s 47111 62087 47209 62185 4 vdd
rlabel metal3 s 42000 61496 42098 61594 4 vdd
rlabel metal3 s 49176 63636 49274 63734 4 gnd
rlabel metal3 s 48921 66407 49019 66505 4 vdd
rlabel metal3 s 49003 65633 49101 65731 4 gnd
rlabel metal3 s 50112 61496 50210 61594 4 vdd
rlabel metal3 s 43753 62087 43851 62185 4 vdd
rlabel metal3 s 44615 62087 44713 62185 4 vdd
rlabel metal3 s 49488 61496 49586 61594 4 vdd
rlabel metal3 s 46437 67245 46535 67343 4 vdd
rlabel metal3 s 48359 62087 48457 62185 4 vdd
rlabel metal3 s 46425 66407 46523 66505 4 vdd
rlabel metal3 s 41515 65633 41613 65731 4 gnd
rlabel metal3 s 41257 62087 41355 62185 4 vdd
rlabel metal3 s 51360 61496 51458 61594 4 vdd
rlabel metal3 s 46437 67567 46535 67665 4 gnd
rlabel metal3 s 46368 61496 46466 61594 4 vdd
rlabel metal3 s 41376 61496 41474 61594 4 vdd
rlabel metal3 s 43941 67245 44039 67343 4 vdd
rlabel metal3 s 45863 62087 45961 62185 4 vdd
rlabel metal3 s 51241 62087 51339 62185 4 vdd
rlabel metal3 s 47928 63636 48026 63734 4 gnd
rlabel metal3 s 48745 62087 48843 62185 4 vdd
rlabel metal3 s 43941 67567 44039 67665 4 gnd
rlabel metal3 s 36453 67245 36551 67343 4 vdd
rlabel metal3 s 31273 62087 31371 62185 4 vdd
rlabel metal3 s 36523 65633 36621 65731 4 gnd
rlabel metal3 s 38949 67567 39047 67665 4 gnd
rlabel metal3 s 36384 61496 36482 61594 4 vdd
rlabel metal3 s 28272 61496 28370 61594 4 vdd
rlabel metal3 s 36441 66407 36539 66505 4 vdd
rlabel metal3 s 27960 63636 28058 63734 4 gnd
rlabel metal3 s 28953 66407 29051 66505 4 vdd
rlabel metal3 s 31392 61496 31490 61594 4 vdd
rlabel metal3 s 34512 61496 34610 61594 4 vdd
rlabel metal3 s 35136 61496 35234 61594 4 vdd
rlabel metal3 s 37008 61496 37106 61594 4 vdd
rlabel metal3 s 29208 63636 29306 63734 4 gnd
rlabel metal3 s 28896 61496 28994 61594 4 vdd
rlabel metal3 s 39019 65633 39117 65731 4 gnd
rlabel metal3 s 30025 62087 30123 62185 4 vdd
rlabel metal3 s 27648 61496 27746 61594 4 vdd
rlabel metal3 s 33957 67245 34055 67343 4 vdd
rlabel metal3 s 35448 63636 35546 63734 4 gnd
rlabel metal3 s 38949 67245 39047 67343 4 vdd
rlabel metal3 s 29639 62087 29737 62185 4 vdd
rlabel metal3 s 38761 62087 38859 62185 4 vdd
rlabel metal3 s 27529 62087 27627 62185 4 vdd
rlabel metal3 s 38256 61496 38354 61594 4 vdd
rlabel metal3 s 32952 63636 33050 63734 4 gnd
rlabel metal3 s 28965 67567 29063 67665 4 gnd
rlabel metal3 s 35760 61496 35858 61594 4 vdd
rlabel metal3 s 33957 67567 34055 67665 4 gnd
rlabel metal3 s 33945 66407 34043 66505 4 vdd
rlabel metal3 s 35017 62087 35115 62185 4 vdd
rlabel metal3 s 30768 61496 30866 61594 4 vdd
rlabel metal3 s 39504 61496 39602 61594 4 vdd
rlabel metal3 s 40128 61496 40226 61594 4 vdd
rlabel metal3 s 33383 62087 33481 62185 4 vdd
rlabel metal3 s 37944 63636 38042 63734 4 gnd
rlabel metal3 s 38937 66407 39035 66505 4 vdd
rlabel metal3 s 37513 62087 37611 62185 4 vdd
rlabel metal3 s 39192 63636 39290 63734 4 gnd
rlabel metal3 s 33888 61496 33986 61594 4 vdd
rlabel metal3 s 33769 62087 33867 62185 4 vdd
rlabel metal3 s 40009 62087 40107 62185 4 vdd
rlabel metal3 s 30144 61496 30242 61594 4 vdd
rlabel metal3 s 30456 63636 30554 63734 4 gnd
rlabel metal3 s 35879 62087 35977 62185 4 vdd
rlabel metal3 s 33264 61496 33362 61594 4 vdd
rlabel metal3 s 32016 61496 32114 61594 4 vdd
rlabel metal3 s 31531 65633 31629 65731 4 gnd
rlabel metal3 s 34027 65633 34125 65731 4 gnd
rlabel metal3 s 31461 67245 31559 67343 4 vdd
rlabel metal3 s 32135 62087 32233 62185 4 vdd
rlabel metal3 s 31449 66407 31547 66505 4 vdd
rlabel metal3 s 38375 62087 38473 62185 4 vdd
rlabel metal3 s 34631 62087 34729 62185 4 vdd
rlabel metal3 s 28965 67245 29063 67343 4 vdd
rlabel metal3 s 29035 65633 29133 65731 4 gnd
rlabel metal3 s 36696 63636 36794 63734 4 gnd
rlabel metal3 s 30887 62087 30985 62185 4 vdd
rlabel metal3 s 36265 62087 36363 62185 4 vdd
rlabel metal3 s 28777 62087 28875 62185 4 vdd
rlabel metal3 s 38880 61496 38978 61594 4 vdd
rlabel metal3 s 29520 61496 29618 61594 4 vdd
rlabel metal3 s 39623 62087 39721 62185 4 vdd
rlabel metal3 s 37632 61496 37730 61594 4 vdd
rlabel metal3 s 28391 62087 28489 62185 4 vdd
rlabel metal3 s 31461 67567 31559 67665 4 gnd
rlabel metal3 s 34200 63636 34298 63734 4 gnd
rlabel metal3 s 32640 61496 32738 61594 4 vdd
rlabel metal3 s 32521 62087 32619 62185 4 vdd
rlabel metal3 s 40440 63636 40538 63734 4 gnd
rlabel metal3 s 36453 67567 36551 67665 4 gnd
rlabel metal3 s 37127 62087 37225 62185 4 vdd
rlabel metal3 s 31704 63636 31802 63734 4 gnd
rlabel metal3 s 27024 61496 27122 61594 4 vdd
rlabel metal3 s 17976 63636 18074 63734 4 gnd
rlabel metal3 s 20041 62087 20139 62185 4 vdd
rlabel metal3 s 15792 61496 15890 61594 4 vdd
rlabel metal3 s 16485 67567 16583 67665 4 gnd
rlabel metal3 s 26539 65633 26637 65731 4 gnd
rlabel metal3 s 22032 61496 22130 61594 4 vdd
rlabel metal3 s 26712 63636 26810 63734 4 gnd
rlabel metal3 s 24647 62087 24745 62185 4 vdd
rlabel metal3 s 16485 67245 16583 67343 4 vdd
rlabel metal3 s 19536 61496 19634 61594 4 vdd
rlabel metal3 s 18288 61496 18386 61594 4 vdd
rlabel metal3 s 25152 61496 25250 61594 4 vdd
rlabel metal3 s 18912 61496 19010 61594 4 vdd
rlabel metal3 s 15168 61496 15266 61594 4 vdd
rlabel metal3 s 23399 62087 23497 62185 4 vdd
rlabel metal3 s 21289 62087 21387 62185 4 vdd
rlabel metal3 s 21408 61496 21506 61594 4 vdd
rlabel metal3 s 26469 67245 26567 67343 4 vdd
rlabel metal3 s 16473 66407 16571 66505 4 vdd
rlabel metal3 s 24216 63636 24314 63734 4 gnd
rlabel metal3 s 26281 62087 26379 62185 4 vdd
rlabel metal3 s 16555 65633 16653 65731 4 gnd
rlabel metal3 s 23973 67567 24071 67665 4 gnd
rlabel metal3 s 26400 61496 26498 61594 4 vdd
rlabel metal3 s 19224 63636 19322 63734 4 gnd
rlabel metal3 s 20472 63636 20570 63734 4 gnd
rlabel metal3 s 23280 61496 23378 61594 4 vdd
rlabel metal3 s 18793 62087 18891 62185 4 vdd
rlabel metal3 s 26457 66407 26555 66505 4 vdd
rlabel metal3 s 14663 62087 14761 62185 4 vdd
rlabel metal3 s 18969 66407 19067 66505 4 vdd
rlabel metal3 s 21477 67245 21575 67343 4 vdd
rlabel metal3 s 15049 62087 15147 62185 4 vdd
rlabel metal3 s 17040 61496 17138 61594 4 vdd
rlabel metal3 s 21720 63636 21818 63734 4 gnd
rlabel metal3 s 25776 61496 25874 61594 4 vdd
rlabel metal3 s 15480 63636 15578 63734 4 gnd
rlabel metal3 s 22151 62087 22249 62185 4 vdd
rlabel metal3 s 21547 65633 21645 65731 4 gnd
rlabel metal3 s 19655 62087 19753 62185 4 vdd
rlabel metal3 s 24528 61496 24626 61594 4 vdd
rlabel metal3 s 25033 62087 25131 62185 4 vdd
rlabel metal3 s 16416 61496 16514 61594 4 vdd
rlabel metal3 s 21465 66407 21563 66505 4 vdd
rlabel metal3 s 19051 65633 19149 65731 4 gnd
rlabel metal3 s 20784 61496 20882 61594 4 vdd
rlabel metal3 s 16728 63636 16826 63734 4 gnd
rlabel metal3 s 25895 62087 25993 62185 4 vdd
rlabel metal3 s 18981 67245 19079 67343 4 vdd
rlabel metal3 s 24043 65633 24141 65731 4 gnd
rlabel metal3 s 15911 62087 16009 62185 4 vdd
rlabel metal3 s 23785 62087 23883 62185 4 vdd
rlabel metal3 s 18981 67567 19079 67665 4 gnd
rlabel metal3 s 17159 62087 17257 62185 4 vdd
rlabel metal3 s 23904 61496 24002 61594 4 vdd
rlabel metal3 s 25464 63636 25562 63734 4 gnd
rlabel metal3 s 21477 67567 21575 67665 4 gnd
rlabel metal3 s 23973 67245 24071 67343 4 vdd
rlabel metal3 s 22968 63636 23066 63734 4 gnd
rlabel metal3 s 22656 61496 22754 61594 4 vdd
rlabel metal3 s 17664 61496 17762 61594 4 vdd
rlabel metal3 s 16297 62087 16395 62185 4 vdd
rlabel metal3 s 18407 62087 18505 62185 4 vdd
rlabel metal3 s 22537 62087 22635 62185 4 vdd
rlabel metal3 s 14544 61496 14642 61594 4 vdd
rlabel metal3 s 20160 61496 20258 61594 4 vdd
rlabel metal3 s 26469 67567 26567 67665 4 gnd
rlabel metal3 s 27143 62087 27241 62185 4 vdd
rlabel metal3 s 17545 62087 17643 62185 4 vdd
rlabel metal3 s 20903 62087 21001 62185 4 vdd
rlabel metal3 s 23961 66407 24059 66505 4 vdd
rlabel metal3 s 7660 60540 7758 60638 4 vdd
rlabel metal3 s 13989 67567 14087 67665 4 gnd
rlabel metal3 s 6882 60563 6980 60661 4 vdd
rlabel metal3 s 13801 62087 13899 62185 4 vdd
rlabel metal3 s 13920 61496 14018 61594 4 vdd
rlabel metal3 s 12600 60935 12698 61033 4 gnd
rlabel metal3 s 12600 60698 12698 60796 4 gnd
rlabel metal3 s 13296 61496 13394 61594 4 vdd
rlabel metal3 s 12234 61282 12332 61380 4 gnd
rlabel metal3 s 13989 67245 14087 67343 4 vdd
rlabel metal3 s 13977 66407 14075 66505 4 vdd
rlabel metal3 s 14059 65633 14157 65731 4 gnd
rlabel metal3 s 6450 60563 6548 60661 4 vdd
rlabel metal3 s 14232 63636 14330 63734 4 gnd
rlabel metal3 s 6025 60563 6123 60661 4 gnd
rlabel metal3 s 7264 60540 7362 60638 4 gnd
rlabel metal3 s 12600 59355 12698 59453 4 gnd
rlabel metal3 s 12600 56748 12698 56846 4 gnd
rlabel metal3 s 12600 59908 12698 60006 4 gnd
rlabel metal3 s 12600 60145 12698 60243 4 gnd
rlabel metal3 s 12600 58565 12698 58663 4 gnd
rlabel metal3 s 12600 56195 12698 56293 4 gnd
rlabel metal3 s 12600 60382 12698 60480 4 gnd
rlabel metal3 s 12600 58012 12698 58110 4 gnd
rlabel metal3 s 12600 58328 12698 58426 4 gnd
rlabel metal3 s 12600 56985 12698 57083 4 gnd
rlabel metal3 s 12600 59592 12698 59690 4 gnd
rlabel metal3 s 12600 57775 12698 57873 4 gnd
rlabel metal3 s 12600 56432 12698 56530 4 gnd
rlabel metal3 s 12600 57538 12698 57636 4 gnd
rlabel metal3 s 12600 59118 12698 59216 4 gnd
rlabel metal3 s 12600 58802 12698 58900 4 gnd
rlabel metal3 s 12600 57222 12698 57320 4 gnd
rlabel metal3 s 6025 57819 6123 57917 4 gnd
rlabel metal3 s 6882 56971 6980 57069 4 vdd
rlabel metal3 s 6025 58609 6123 58707 4 gnd
rlabel metal3 s 7660 57380 7758 57478 4 vdd
rlabel metal3 s 7264 58960 7362 59058 4 gnd
rlabel metal3 s 7264 59355 7362 59453 4 gnd
rlabel metal3 s 6025 56239 6123 56337 4 gnd
rlabel metal3 s 6450 59341 6548 59439 4 vdd
rlabel metal3 s 6450 56971 6548 57069 4 vdd
rlabel metal3 s 6882 57761 6980 57859 4 vdd
rlabel metal3 s 7660 59750 7758 59848 4 vdd
rlabel metal3 s 6025 59399 6123 59497 4 gnd
rlabel metal3 s 6882 58983 6980 59081 4 vdd
rlabel metal3 s 6450 58551 6548 58649 4 vdd
rlabel metal3 s 7660 60145 7758 60243 4 vdd
rlabel metal3 s 7660 58565 7758 58663 4 vdd
rlabel metal3 s 6450 59773 6548 59871 4 vdd
rlabel metal3 s 7264 59750 7362 59848 4 gnd
rlabel metal3 s 6882 58193 6980 58291 4 vdd
rlabel metal3 s 7660 58170 7758 58268 4 vdd
rlabel metal3 s 6025 59773 6123 59871 4 gnd
rlabel metal3 s 7264 56985 7362 57083 4 gnd
rlabel metal3 s 6450 60131 6548 60229 4 vdd
rlabel metal3 s 6882 56613 6980 56711 4 vdd
rlabel metal3 s 6025 60189 6123 60287 4 gnd
rlabel metal3 s 7660 58960 7758 59058 4 vdd
rlabel metal3 s 6025 56613 6123 56711 4 gnd
rlabel metal3 s 7660 59355 7758 59453 4 vdd
rlabel metal3 s 6025 57403 6123 57501 4 gnd
rlabel metal3 s 7660 56590 7758 56688 4 vdd
rlabel metal3 s 7264 58565 7362 58663 4 gnd
rlabel metal3 s 6882 59341 6980 59439 4 vdd
rlabel metal3 s 6450 58983 6548 59081 4 vdd
rlabel metal3 s 7660 56195 7758 56293 4 vdd
rlabel metal3 s 6450 56613 6548 56711 4 vdd
rlabel metal3 s 7660 56985 7758 57083 4 vdd
rlabel metal3 s 6025 58193 6123 58291 4 gnd
rlabel metal3 s 6882 58551 6980 58649 4 vdd
rlabel metal3 s 7264 57380 7362 57478 4 gnd
rlabel metal3 s 6450 57761 6548 57859 4 vdd
rlabel metal3 s 7264 58170 7362 58268 4 gnd
rlabel metal3 s 7264 56590 7362 56688 4 gnd
rlabel metal3 s 6025 57029 6123 57127 4 gnd
rlabel metal3 s 7264 60145 7362 60243 4 gnd
rlabel metal3 s 7264 56195 7362 56293 4 gnd
rlabel metal3 s 6882 60131 6980 60229 4 vdd
rlabel metal3 s 6450 58193 6548 58291 4 vdd
rlabel metal3 s 6882 57403 6980 57501 4 vdd
rlabel metal3 s 7660 57775 7758 57873 4 vdd
rlabel metal3 s 6450 57403 6548 57501 4 vdd
rlabel metal3 s 6025 58983 6123 59081 4 gnd
rlabel metal3 s 7264 57775 7362 57873 4 gnd
rlabel metal3 s 6882 59773 6980 59871 4 vdd
rlabel metal3 s 7264 53430 7362 53528 4 gnd
rlabel metal3 s 6450 52231 6548 52329 4 vdd
rlabel metal3 s 6450 51873 6548 51971 4 vdd
rlabel metal3 s 7660 53035 7758 53133 4 vdd
rlabel metal3 s 6450 55391 6548 55489 4 vdd
rlabel metal3 s 6025 51873 6123 51971 4 gnd
rlabel metal3 s 6882 52663 6980 52761 4 vdd
rlabel metal3 s 6882 54601 6980 54699 4 vdd
rlabel metal3 s 6882 56181 6980 56279 4 vdd
rlabel metal3 s 6025 55449 6123 55547 4 gnd
rlabel metal3 s 7264 53035 7362 53133 4 gnd
rlabel metal3 s 7264 52245 7362 52343 4 gnd
rlabel metal3 s 7264 55010 7362 55108 4 gnd
rlabel metal3 s 6882 53021 6980 53119 4 vdd
rlabel metal3 s 7660 52245 7758 52343 4 vdd
rlabel metal3 s 6882 53453 6980 53551 4 vdd
rlabel metal3 s 6882 52231 6980 52329 4 vdd
rlabel metal3 s 7264 53825 7362 53923 4 gnd
rlabel metal3 s 7264 55800 7362 55898 4 gnd
rlabel metal3 s 6025 53453 6123 53551 4 gnd
rlabel metal3 s 7660 54615 7758 54713 4 vdd
rlabel metal3 s 7660 55010 7758 55108 4 vdd
rlabel metal3 s 6450 53021 6548 53119 4 vdd
rlabel metal3 s 6025 55033 6123 55131 4 gnd
rlabel metal3 s 6025 54243 6123 54341 4 gnd
rlabel metal3 s 6450 56181 6548 56279 4 vdd
rlabel metal3 s 7264 55405 7362 55503 4 gnd
rlabel metal3 s 6450 54601 6548 54699 4 vdd
rlabel metal3 s 6025 54659 6123 54757 4 gnd
rlabel metal3 s 6025 55823 6123 55921 4 gnd
rlabel metal3 s 6882 51873 6980 51971 4 vdd
rlabel metal3 s 6025 53869 6123 53967 4 gnd
rlabel metal3 s 6882 55391 6980 55489 4 vdd
rlabel metal3 s 6025 52663 6123 52761 4 gnd
rlabel metal3 s 6450 53453 6548 53551 4 vdd
rlabel metal3 s 7264 54220 7362 54318 4 gnd
rlabel metal3 s 6450 52663 6548 52761 4 vdd
rlabel metal3 s 6025 53079 6123 53177 4 gnd
rlabel metal3 s 7660 53825 7758 53923 4 vdd
rlabel metal3 s 6450 55823 6548 55921 4 vdd
rlabel metal3 s 6450 53811 6548 53909 4 vdd
rlabel metal3 s 7660 53430 7758 53528 4 vdd
rlabel metal3 s 6882 53811 6980 53909 4 vdd
rlabel metal3 s 7264 54615 7362 54713 4 gnd
rlabel metal3 s 7660 55800 7758 55898 4 vdd
rlabel metal3 s 6882 55033 6980 55131 4 vdd
rlabel metal3 s 7660 55405 7758 55503 4 vdd
rlabel metal3 s 6450 54243 6548 54341 4 vdd
rlabel metal3 s 6025 52289 6123 52387 4 gnd
rlabel metal3 s 7660 52640 7758 52738 4 vdd
rlabel metal3 s 6450 55033 6548 55131 4 vdd
rlabel metal3 s 7660 54220 7758 54318 4 vdd
rlabel metal3 s 6882 55823 6980 55921 4 vdd
rlabel metal3 s 6882 54243 6980 54341 4 vdd
rlabel metal3 s 7264 52640 7362 52738 4 gnd
rlabel metal3 s 12600 54062 12698 54160 4 gnd
rlabel metal3 s 12600 53588 12698 53686 4 gnd
rlabel metal3 s 12600 55642 12698 55740 4 gnd
rlabel metal3 s 12600 52798 12698 52896 4 gnd
rlabel metal3 s 12600 54852 12698 54950 4 gnd
rlabel metal3 s 12600 53825 12698 53923 4 gnd
rlabel metal3 s 12600 55405 12698 55503 4 gnd
rlabel metal3 s 12600 55958 12698 56056 4 gnd
rlabel metal3 s 12600 52008 12698 52106 4 gnd
rlabel metal3 s 12600 52245 12698 52343 4 gnd
rlabel metal3 s 12600 53272 12698 53370 4 gnd
rlabel metal3 s 12600 55168 12698 55266 4 gnd
rlabel metal3 s 12600 52482 12698 52580 4 gnd
rlabel metal3 s 12600 53035 12698 53133 4 gnd
rlabel metal3 s 12600 54378 12698 54476 4 gnd
rlabel metal3 s 12600 54615 12698 54713 4 gnd
rlabel metal3 s 12600 47742 12698 47840 4 gnd
rlabel metal3 s 12600 50665 12698 50763 4 gnd
rlabel metal3 s 12600 51455 12698 51553 4 gnd
rlabel metal3 s 12600 48532 12698 48630 4 gnd
rlabel metal3 s 12600 48848 12698 48946 4 gnd
rlabel metal3 s 12600 51218 12698 51316 4 gnd
rlabel metal3 s 12600 48295 12698 48393 4 gnd
rlabel metal3 s 12600 50902 12698 51000 4 gnd
rlabel metal3 s 12600 49085 12698 49183 4 gnd
rlabel metal3 s 12600 50428 12698 50526 4 gnd
rlabel metal3 s 12600 51692 12698 51790 4 gnd
rlabel metal3 s 12600 49875 12698 49973 4 gnd
rlabel metal3 s 12600 50112 12698 50210 4 gnd
rlabel metal3 s 12600 49322 12698 49420 4 gnd
rlabel metal3 s 12600 49638 12698 49736 4 gnd
rlabel metal3 s 12600 48058 12698 48156 4 gnd
rlabel metal3 s 7660 51850 7758 51948 4 vdd
rlabel metal3 s 6882 47923 6980 48021 4 vdd
rlabel metal3 s 6450 48281 6548 48379 4 vdd
rlabel metal3 s 6882 50651 6980 50749 4 vdd
rlabel metal3 s 7264 48690 7362 48788 4 gnd
rlabel metal3 s 6025 47549 6123 47647 4 gnd
rlabel metal3 s 7660 51455 7758 51553 4 vdd
rlabel metal3 s 7660 50665 7758 50763 4 vdd
rlabel metal3 s 7660 49085 7758 49183 4 vdd
rlabel metal3 s 7264 47900 7362 47998 4 gnd
rlabel metal3 s 6882 51083 6980 51181 4 vdd
rlabel metal3 s 7660 49875 7758 49973 4 vdd
rlabel metal3 s 6025 50709 6123 50807 4 gnd
rlabel metal3 s 7660 48690 7758 48788 4 vdd
rlabel metal3 s 6882 48281 6980 48379 4 vdd
rlabel metal3 s 6882 49503 6980 49601 4 vdd
rlabel metal3 s 6450 47923 6548 48021 4 vdd
rlabel metal3 s 6025 47923 6123 48021 4 gnd
rlabel metal3 s 6450 48713 6548 48811 4 vdd
rlabel metal3 s 7660 48295 7758 48393 4 vdd
rlabel metal3 s 7264 50270 7362 50368 4 gnd
rlabel metal3 s 7660 51060 7758 51158 4 vdd
rlabel metal3 s 6025 48339 6123 48437 4 gnd
rlabel metal3 s 7264 51455 7362 51553 4 gnd
rlabel metal3 s 7264 51850 7362 51948 4 gnd
rlabel metal3 s 6025 50293 6123 50391 4 gnd
rlabel metal3 s 6882 48713 6980 48811 4 vdd
rlabel metal3 s 6025 49503 6123 49601 4 gnd
rlabel metal3 s 7264 50665 7362 50763 4 gnd
rlabel metal3 s 6450 49503 6548 49601 4 vdd
rlabel metal3 s 6450 50293 6548 50391 4 vdd
rlabel metal3 s 6025 49129 6123 49227 4 gnd
rlabel metal3 s 6025 51083 6123 51181 4 gnd
rlabel metal3 s 7660 50270 7758 50368 4 vdd
rlabel metal3 s 6450 51083 6548 51181 4 vdd
rlabel metal3 s 6882 49071 6980 49169 4 vdd
rlabel metal3 s 7264 49085 7362 49183 4 gnd
rlabel metal3 s 7264 49480 7362 49578 4 gnd
rlabel metal3 s 6882 50293 6980 50391 4 vdd
rlabel metal3 s 7264 48295 7362 48393 4 gnd
rlabel metal3 s 6882 49861 6980 49959 4 vdd
rlabel metal3 s 6450 51441 6548 51539 4 vdd
rlabel metal3 s 7660 47900 7758 47998 4 vdd
rlabel metal3 s 6450 49861 6548 49959 4 vdd
rlabel metal3 s 7264 51060 7362 51158 4 gnd
rlabel metal3 s 7264 49875 7362 49973 4 gnd
rlabel metal3 s 6882 51441 6980 51539 4 vdd
rlabel metal3 s 6450 50651 6548 50749 4 vdd
rlabel metal3 s 6025 49919 6123 50017 4 gnd
rlabel metal3 s 6025 48713 6123 48811 4 gnd
rlabel metal3 s 6450 49071 6548 49169 4 vdd
rlabel metal3 s 7660 49480 7758 49578 4 vdd
rlabel metal3 s 6025 51499 6123 51597 4 gnd
rlabel metal3 s 6882 45553 6980 45651 4 vdd
rlabel metal3 s 7264 44345 7362 44443 4 gnd
rlabel metal3 s 6882 44763 6980 44861 4 vdd
rlabel metal3 s 7264 43950 7362 44048 4 gnd
rlabel metal3 s 6025 43973 6123 44071 4 gnd
rlabel metal3 s 6025 46343 6123 46441 4 gnd
rlabel metal3 s 7660 47505 7758 47603 4 vdd
rlabel metal3 s 6025 45969 6123 46067 4 gnd
rlabel metal3 s 7264 45530 7362 45628 4 gnd
rlabel metal3 s 6450 46701 6548 46799 4 vdd
rlabel metal3 s 6882 45911 6980 46009 4 vdd
rlabel metal3 s 6025 47133 6123 47231 4 gnd
rlabel metal3 s 7264 44740 7362 44838 4 gnd
rlabel metal3 s 7264 45135 7362 45233 4 gnd
rlabel metal3 s 6450 47491 6548 47589 4 vdd
rlabel metal3 s 6450 43541 6548 43639 4 vdd
rlabel metal3 s 7660 46320 7758 46418 4 vdd
rlabel metal3 s 7660 44740 7758 44838 4 vdd
rlabel metal3 s 7264 46320 7362 46418 4 gnd
rlabel metal3 s 6882 43541 6980 43639 4 vdd
rlabel metal3 s 6450 45553 6548 45651 4 vdd
rlabel metal3 s 6025 45553 6123 45651 4 gnd
rlabel metal3 s 6882 47133 6980 47231 4 vdd
rlabel metal3 s 7660 44345 7758 44443 4 vdd
rlabel metal3 s 6025 43599 6123 43697 4 gnd
rlabel metal3 s 6025 44763 6123 44861 4 gnd
rlabel metal3 s 7660 45530 7758 45628 4 vdd
rlabel metal3 s 7660 47110 7758 47208 4 vdd
rlabel metal3 s 6450 43973 6548 44071 4 vdd
rlabel metal3 s 6882 43973 6980 44071 4 vdd
rlabel metal3 s 6450 44331 6548 44429 4 vdd
rlabel metal3 s 6882 46343 6980 46441 4 vdd
rlabel metal3 s 7264 46715 7362 46813 4 gnd
rlabel metal3 s 7660 43555 7758 43653 4 vdd
rlabel metal3 s 6882 45121 6980 45219 4 vdd
rlabel metal3 s 6882 47491 6980 47589 4 vdd
rlabel metal3 s 6025 44389 6123 44487 4 gnd
rlabel metal3 s 6450 46343 6548 46441 4 vdd
rlabel metal3 s 6450 45911 6548 46009 4 vdd
rlabel metal3 s 6025 46759 6123 46857 4 gnd
rlabel metal3 s 6450 47133 6548 47231 4 vdd
rlabel metal3 s 7660 46715 7758 46813 4 vdd
rlabel metal3 s 7264 47505 7362 47603 4 gnd
rlabel metal3 s 7264 47110 7362 47208 4 gnd
rlabel metal3 s 7264 45925 7362 46023 4 gnd
rlabel metal3 s 6450 44763 6548 44861 4 vdd
rlabel metal3 s 6882 44331 6980 44429 4 vdd
rlabel metal3 s 7660 43950 7758 44048 4 vdd
rlabel metal3 s 7264 43555 7362 43653 4 gnd
rlabel metal3 s 6025 45179 6123 45277 4 gnd
rlabel metal3 s 7660 45135 7758 45233 4 vdd
rlabel metal3 s 6450 45121 6548 45219 4 vdd
rlabel metal3 s 7660 45925 7758 46023 4 vdd
rlabel metal3 s 6882 46701 6980 46799 4 vdd
rlabel metal3 s 12600 47505 12698 47603 4 gnd
rlabel metal3 s 12600 44898 12698 44996 4 gnd
rlabel metal3 s 12600 46952 12698 47050 4 gnd
rlabel metal3 s 12600 46162 12698 46260 4 gnd
rlabel metal3 s 12600 44582 12698 44680 4 gnd
rlabel metal3 s 12600 45372 12698 45470 4 gnd
rlabel metal3 s 12600 46478 12698 46576 4 gnd
rlabel metal3 s 12600 43555 12698 43653 4 gnd
rlabel metal3 s 12600 46715 12698 46813 4 gnd
rlabel metal3 s 12600 45135 12698 45233 4 gnd
rlabel metal3 s 12600 43318 12698 43416 4 gnd
rlabel metal3 s 12600 45925 12698 46023 4 gnd
rlabel metal3 s 12600 45688 12698 45786 4 gnd
rlabel metal3 s 12600 44108 12698 44206 4 gnd
rlabel metal3 s 12600 43792 12698 43890 4 gnd
rlabel metal3 s 12600 47268 12698 47366 4 gnd
rlabel metal3 s 12600 44345 12698 44443 4 gnd
rlabel metal3 s 12600 40158 12698 40256 4 gnd
rlabel metal3 s 12600 41185 12698 41283 4 gnd
rlabel metal3 s 12600 42212 12698 42310 4 gnd
rlabel metal3 s 12600 41422 12698 41520 4 gnd
rlabel metal3 s 12600 39052 12698 39150 4 gnd
rlabel metal3 s 12600 40395 12698 40493 4 gnd
rlabel metal3 s 12600 42765 12698 42863 4 gnd
rlabel metal3 s 12600 40948 12698 41046 4 gnd
rlabel metal3 s 12600 39605 12698 39703 4 gnd
rlabel metal3 s 12600 41975 12698 42073 4 gnd
rlabel metal3 s 12600 42528 12698 42626 4 gnd
rlabel metal3 s 12600 39368 12698 39466 4 gnd
rlabel metal3 s 12600 40632 12698 40730 4 gnd
rlabel metal3 s 12600 41738 12698 41836 4 gnd
rlabel metal3 s 12600 39842 12698 39940 4 gnd
rlabel metal3 s 12600 43002 12698 43100 4 gnd
rlabel metal3 s 6882 41603 6980 41701 4 vdd
rlabel metal3 s 7264 41975 7362 42073 4 gnd
rlabel metal3 s 6025 39649 6123 39747 4 gnd
rlabel metal3 s 6025 41603 6123 41701 4 gnd
rlabel metal3 s 7660 41185 7758 41283 4 vdd
rlabel metal3 s 6450 42393 6548 42491 4 vdd
rlabel metal3 s 7660 40790 7758 40888 4 vdd
rlabel metal3 s 7264 42370 7362 42468 4 gnd
rlabel metal3 s 6025 40023 6123 40121 4 gnd
rlabel metal3 s 6450 42751 6548 42849 4 vdd
rlabel metal3 s 7264 40395 7362 40493 4 gnd
rlabel metal3 s 6450 41171 6548 41269 4 vdd
rlabel metal3 s 6882 40023 6980 40121 4 vdd
rlabel metal3 s 6450 39591 6548 39689 4 vdd
rlabel metal3 s 7660 43160 7758 43258 4 vdd
rlabel metal3 s 6882 39233 6980 39331 4 vdd
rlabel metal3 s 6025 41229 6123 41327 4 gnd
rlabel metal3 s 7264 42765 7362 42863 4 gnd
rlabel metal3 s 7660 42370 7758 42468 4 vdd
rlabel metal3 s 6882 39591 6980 39689 4 vdd
rlabel metal3 s 6025 42809 6123 42907 4 gnd
rlabel metal3 s 6882 42393 6980 42491 4 vdd
rlabel metal3 s 6025 42019 6123 42117 4 gnd
rlabel metal3 s 6025 40439 6123 40537 4 gnd
rlabel metal3 s 7660 39210 7758 39308 4 vdd
rlabel metal3 s 6450 39233 6548 39331 4 vdd
rlabel metal3 s 6882 40813 6980 40911 4 vdd
rlabel metal3 s 7660 41975 7758 42073 4 vdd
rlabel metal3 s 7264 39605 7362 39703 4 gnd
rlabel metal3 s 7264 40000 7362 40098 4 gnd
rlabel metal3 s 6450 41961 6548 42059 4 vdd
rlabel metal3 s 6025 42393 6123 42491 4 gnd
rlabel metal3 s 6882 40381 6980 40479 4 vdd
rlabel metal3 s 6882 41171 6980 41269 4 vdd
rlabel metal3 s 6882 42751 6980 42849 4 vdd
rlabel metal3 s 7660 42765 7758 42863 4 vdd
rlabel metal3 s 7264 39210 7362 39308 4 gnd
rlabel metal3 s 6450 41603 6548 41701 4 vdd
rlabel metal3 s 7660 39605 7758 39703 4 vdd
rlabel metal3 s 6882 41961 6980 42059 4 vdd
rlabel metal3 s 6450 40813 6548 40911 4 vdd
rlabel metal3 s 6882 43183 6980 43281 4 vdd
rlabel metal3 s 7660 41580 7758 41678 4 vdd
rlabel metal3 s 7264 43160 7362 43258 4 gnd
rlabel metal3 s 7264 40790 7362 40888 4 gnd
rlabel metal3 s 6025 40813 6123 40911 4 gnd
rlabel metal3 s 7660 40395 7758 40493 4 vdd
rlabel metal3 s 7264 41580 7362 41678 4 gnd
rlabel metal3 s 7264 41185 7362 41283 4 gnd
rlabel metal3 s 7660 40000 7758 40098 4 vdd
rlabel metal3 s 6450 40023 6548 40121 4 vdd
rlabel metal3 s 6025 39233 6123 39331 4 gnd
rlabel metal3 s 6450 40381 6548 40479 4 vdd
rlabel metal3 s 6450 43183 6548 43281 4 vdd
rlabel metal3 s 6025 43183 6123 43281 4 gnd
rlabel metal3 s 6882 35641 6980 35739 4 vdd
rlabel metal3 s 7660 38420 7758 38518 4 vdd
rlabel metal3 s 6450 36431 6548 36529 4 vdd
rlabel metal3 s 6450 36863 6548 36961 4 vdd
rlabel metal3 s 6450 38443 6548 38541 4 vdd
rlabel metal3 s 6025 38443 6123 38541 4 gnd
rlabel metal3 s 7660 38815 7758 38913 4 vdd
rlabel metal3 s 6025 38069 6123 38167 4 gnd
rlabel metal3 s 6882 38801 6980 38899 4 vdd
rlabel metal3 s 7660 35655 7758 35753 4 vdd
rlabel metal3 s 7660 35260 7758 35358 4 vdd
rlabel metal3 s 7660 34865 7758 34963 4 vdd
rlabel metal3 s 6025 34909 6123 35007 4 gnd
rlabel metal3 s 7264 36050 7362 36148 4 gnd
rlabel metal3 s 6450 37653 6548 37751 4 vdd
rlabel metal3 s 6025 35283 6123 35381 4 gnd
rlabel metal3 s 6450 36073 6548 36171 4 vdd
rlabel metal3 s 6025 36863 6123 36961 4 gnd
rlabel metal3 s 6025 35699 6123 35797 4 gnd
rlabel metal3 s 6450 35641 6548 35739 4 vdd
rlabel metal3 s 6025 38859 6123 38957 4 gnd
rlabel metal3 s 7264 35260 7362 35358 4 gnd
rlabel metal3 s 7264 37630 7362 37728 4 gnd
rlabel metal3 s 7660 36050 7758 36148 4 vdd
rlabel metal3 s 7660 37235 7758 37333 4 vdd
rlabel metal3 s 6025 36073 6123 36171 4 gnd
rlabel metal3 s 7264 34865 7362 34963 4 gnd
rlabel metal3 s 7660 36445 7758 36543 4 vdd
rlabel metal3 s 7660 36840 7758 36938 4 vdd
rlabel metal3 s 6450 38801 6548 38899 4 vdd
rlabel metal3 s 6882 36431 6980 36529 4 vdd
rlabel metal3 s 6025 36489 6123 36587 4 gnd
rlabel metal3 s 6450 34851 6548 34949 4 vdd
rlabel metal3 s 7264 38025 7362 38123 4 gnd
rlabel metal3 s 7264 36840 7362 36938 4 gnd
rlabel metal3 s 6882 38011 6980 38109 4 vdd
rlabel metal3 s 7264 38815 7362 38913 4 gnd
rlabel metal3 s 6450 35283 6548 35381 4 vdd
rlabel metal3 s 6025 37653 6123 37751 4 gnd
rlabel metal3 s 6882 34851 6980 34949 4 vdd
rlabel metal3 s 6882 36863 6980 36961 4 vdd
rlabel metal3 s 7264 38420 7362 38518 4 gnd
rlabel metal3 s 7264 37235 7362 37333 4 gnd
rlabel metal3 s 7660 37630 7758 37728 4 vdd
rlabel metal3 s 6882 36073 6980 36171 4 vdd
rlabel metal3 s 7660 38025 7758 38123 4 vdd
rlabel metal3 s 7264 35655 7362 35753 4 gnd
rlabel metal3 s 6025 37279 6123 37377 4 gnd
rlabel metal3 s 7264 36445 7362 36543 4 gnd
rlabel metal3 s 6450 38011 6548 38109 4 vdd
rlabel metal3 s 6882 38443 6980 38541 4 vdd
rlabel metal3 s 6882 37653 6980 37751 4 vdd
rlabel metal3 s 6450 37221 6548 37319 4 vdd
rlabel metal3 s 6882 35283 6980 35381 4 vdd
rlabel metal3 s 6882 37221 6980 37319 4 vdd
rlabel metal3 s 12600 38815 12698 38913 4 gnd
rlabel metal3 s 12600 38025 12698 38123 4 gnd
rlabel metal3 s 12600 38578 12698 38676 4 gnd
rlabel metal3 s 12600 35892 12698 35990 4 gnd
rlabel metal3 s 11208 35655 11306 35753 4 vdd
rlabel metal3 s 9560 35655 9658 35753 4 gnd
rlabel metal3 s 12600 36998 12698 37096 4 gnd
rlabel metal3 s 12600 38262 12698 38360 4 gnd
rlabel metal3 s 8092 35640 8190 35738 4 gnd
rlabel metal3 s 12600 35655 12698 35753 4 gnd
rlabel metal3 s 12600 37235 12698 37333 4 gnd
rlabel metal3 s 12600 34865 12698 34963 4 gnd
rlabel metal3 s 12600 37788 12698 37886 4 gnd
rlabel metal3 s 12600 37472 12698 37570 4 gnd
rlabel metal3 s 12600 34628 12698 34726 4 gnd
rlabel metal3 s 12600 36445 12698 36543 4 gnd
rlabel metal3 s 12600 36208 12698 36306 4 gnd
rlabel metal3 s 12600 35102 12698 35200 4 gnd
rlabel metal3 s 8517 35639 8615 35737 4 vdd
rlabel metal3 s 12600 36682 12698 36780 4 gnd
rlabel metal3 s 12600 35418 12698 35516 4 gnd
rlabel metal3 s 12600 33285 12698 33383 4 gnd
rlabel metal3 s 12600 30915 12698 31013 4 gnd
rlabel metal3 s 12600 30678 12698 30776 4 gnd
rlabel metal3 s 12600 33838 12698 33936 4 gnd
rlabel metal3 s 12600 31705 12698 31803 4 gnd
rlabel metal3 s 12600 31942 12698 32040 4 gnd
rlabel metal3 s 12600 32495 12698 32593 4 gnd
rlabel metal3 s 12600 31152 12698 31250 4 gnd
rlabel metal3 s 12600 34312 12698 34410 4 gnd
rlabel metal3 s 12600 34075 12698 34173 4 gnd
rlabel metal3 s 12600 30362 12698 30460 4 gnd
rlabel metal3 s 12600 33522 12698 33620 4 gnd
rlabel metal3 s 12600 32732 12698 32830 4 gnd
rlabel metal3 s 12600 32258 12698 32356 4 gnd
rlabel metal3 s 12600 33048 12698 33146 4 gnd
rlabel metal3 s 12600 31468 12698 31566 4 gnd
rlabel metal3 s 6450 32481 6548 32579 4 vdd
rlabel metal3 s 7264 31705 7362 31803 4 gnd
rlabel metal3 s 6025 34119 6123 34217 4 gnd
rlabel metal3 s 7264 30520 7362 30618 4 gnd
rlabel metal3 s 6025 30543 6123 30641 4 gnd
rlabel metal3 s 6882 34061 6980 34159 4 vdd
rlabel metal3 s 6450 32913 6548 33011 4 vdd
rlabel metal3 s 7660 32495 7758 32593 4 vdd
rlabel metal3 s 6025 32123 6123 32221 4 gnd
rlabel metal3 s 6882 31333 6980 31431 4 vdd
rlabel metal3 s 6025 30959 6123 31057 4 gnd
rlabel metal3 s 7660 31705 7758 31803 4 vdd
rlabel metal3 s 6025 33329 6123 33427 4 gnd
rlabel metal3 s 7660 32100 7758 32198 4 vdd
rlabel metal3 s 6450 33703 6548 33801 4 vdd
rlabel metal3 s 7660 34470 7758 34568 4 vdd
rlabel metal3 s 7660 30915 7758 31013 4 vdd
rlabel metal3 s 7660 34075 7758 34173 4 vdd
rlabel metal3 s 7660 30520 7758 30618 4 vdd
rlabel metal3 s 6882 34493 6980 34591 4 vdd
rlabel metal3 s 6025 31333 6123 31431 4 gnd
rlabel metal3 s 6025 31749 6123 31847 4 gnd
rlabel metal3 s 6882 30901 6980 30999 4 vdd
rlabel metal3 s 6450 30901 6548 30999 4 vdd
rlabel metal3 s 7660 33680 7758 33778 4 vdd
rlabel metal3 s 6450 33271 6548 33369 4 vdd
rlabel metal3 s 7660 33285 7758 33383 4 vdd
rlabel metal3 s 7264 33285 7362 33383 4 gnd
rlabel metal3 s 7660 31310 7758 31408 4 vdd
rlabel metal3 s 7264 30915 7362 31013 4 gnd
rlabel metal3 s 6025 34493 6123 34591 4 gnd
rlabel metal3 s 7264 34470 7362 34568 4 gnd
rlabel metal3 s 6450 32123 6548 32221 4 vdd
rlabel metal3 s 7660 32890 7758 32988 4 vdd
rlabel metal3 s 7264 34075 7362 34173 4 gnd
rlabel metal3 s 6882 32123 6980 32221 4 vdd
rlabel metal3 s 6882 33703 6980 33801 4 vdd
rlabel metal3 s 7264 32890 7362 32988 4 gnd
rlabel metal3 s 6450 31691 6548 31789 4 vdd
rlabel metal3 s 7264 32495 7362 32593 4 gnd
rlabel metal3 s 6882 31691 6980 31789 4 vdd
rlabel metal3 s 6025 32913 6123 33011 4 gnd
rlabel metal3 s 7264 32100 7362 32198 4 gnd
rlabel metal3 s 6450 31333 6548 31431 4 vdd
rlabel metal3 s 6025 33703 6123 33801 4 gnd
rlabel metal3 s 6025 32539 6123 32637 4 gnd
rlabel metal3 s 6450 34493 6548 34591 4 vdd
rlabel metal3 s 6882 32481 6980 32579 4 vdd
rlabel metal3 s 7264 31310 7362 31408 4 gnd
rlabel metal3 s 6882 33271 6980 33369 4 vdd
rlabel metal3 s 6450 30543 6548 30641 4 vdd
rlabel metal3 s 6882 32913 6980 33011 4 vdd
rlabel metal3 s 6450 34061 6548 34159 4 vdd
rlabel metal3 s 6882 30543 6980 30641 4 vdd
rlabel metal3 s 7264 33680 7362 33778 4 gnd
rlabel metal3 s 7264 26175 7362 26273 4 gnd
rlabel metal3 s 6882 28963 6980 29061 4 vdd
rlabel metal3 s 6450 26161 6548 26259 4 vdd
rlabel metal3 s 6025 28963 6123 29061 4 gnd
rlabel metal3 s 6882 26593 6980 26691 4 vdd
rlabel metal3 s 6025 29753 6123 29851 4 gnd
rlabel metal3 s 6450 27741 6548 27839 4 vdd
rlabel metal3 s 7660 26175 7758 26273 4 vdd
rlabel metal3 s 7264 28150 7362 28248 4 gnd
rlabel metal3 s 6882 27741 6980 27839 4 vdd
rlabel metal3 s 6450 26593 6548 26691 4 vdd
rlabel metal3 s 7660 30125 7758 30223 4 vdd
rlabel metal3 s 6450 28531 6548 28629 4 vdd
rlabel metal3 s 7264 29335 7362 29433 4 gnd
rlabel metal3 s 7264 27755 7362 27853 4 gnd
rlabel metal3 s 7660 29335 7758 29433 4 vdd
rlabel metal3 s 7264 30125 7362 30223 4 gnd
rlabel metal3 s 6450 30111 6548 30209 4 vdd
rlabel metal3 s 6882 28173 6980 28271 4 vdd
rlabel metal3 s 6882 29753 6980 29851 4 vdd
rlabel metal3 s 7660 28545 7758 28643 4 vdd
rlabel metal3 s 6882 29321 6980 29419 4 vdd
rlabel metal3 s 6025 26593 6123 26691 4 gnd
rlabel metal3 s 7660 26965 7758 27063 4 vdd
rlabel metal3 s 7660 26570 7758 26668 4 vdd
rlabel metal3 s 6450 28173 6548 28271 4 vdd
rlabel metal3 s 7264 29730 7362 29828 4 gnd
rlabel metal3 s 6025 30169 6123 30267 4 gnd
rlabel metal3 s 6882 26161 6980 26259 4 vdd
rlabel metal3 s 7264 27360 7362 27458 4 gnd
rlabel metal3 s 7660 29730 7758 29828 4 vdd
rlabel metal3 s 7660 27360 7758 27458 4 vdd
rlabel metal3 s 6025 28173 6123 28271 4 gnd
rlabel metal3 s 7660 27755 7758 27853 4 vdd
rlabel metal3 s 6025 29379 6123 29477 4 gnd
rlabel metal3 s 6882 27383 6980 27481 4 vdd
rlabel metal3 s 6025 27799 6123 27897 4 gnd
rlabel metal3 s 7264 26965 7362 27063 4 gnd
rlabel metal3 s 6882 30111 6980 30209 4 vdd
rlabel metal3 s 6450 26951 6548 27049 4 vdd
rlabel metal3 s 6025 27383 6123 27481 4 gnd
rlabel metal3 s 7264 28940 7362 29038 4 gnd
rlabel metal3 s 7264 26570 7362 26668 4 gnd
rlabel metal3 s 6025 28589 6123 28687 4 gnd
rlabel metal3 s 6450 29753 6548 29851 4 vdd
rlabel metal3 s 6025 27009 6123 27107 4 gnd
rlabel metal3 s 7264 28545 7362 28643 4 gnd
rlabel metal3 s 6882 26951 6980 27049 4 vdd
rlabel metal3 s 6025 26219 6123 26317 4 gnd
rlabel metal3 s 6882 28531 6980 28629 4 vdd
rlabel metal3 s 6450 27383 6548 27481 4 vdd
rlabel metal3 s 7660 28940 7758 29038 4 vdd
rlabel metal3 s 6450 28963 6548 29061 4 vdd
rlabel metal3 s 7660 28150 7758 28248 4 vdd
rlabel metal3 s 6450 29321 6548 29419 4 vdd
rlabel metal3 s 12600 29888 12698 29986 4 gnd
rlabel metal3 s 12600 26175 12698 26273 4 gnd
rlabel metal3 s 12600 27202 12698 27300 4 gnd
rlabel metal3 s 12600 28545 12698 28643 4 gnd
rlabel metal3 s 12600 26412 12698 26510 4 gnd
rlabel metal3 s 12600 26965 12698 27063 4 gnd
rlabel metal3 s 12600 29098 12698 29196 4 gnd
rlabel metal3 s 12600 27992 12698 28090 4 gnd
rlabel metal3 s 12600 29335 12698 29433 4 gnd
rlabel metal3 s 12600 28782 12698 28880 4 gnd
rlabel metal3 s 12600 27518 12698 27616 4 gnd
rlabel metal3 s 12600 26728 12698 26826 4 gnd
rlabel metal3 s 12600 27755 12698 27853 4 gnd
rlabel metal3 s 12600 28308 12698 28406 4 gnd
rlabel metal3 s 12600 29572 12698 29670 4 gnd
rlabel metal3 s 12600 25938 12698 26036 4 gnd
rlabel metal3 s 12600 30125 12698 30223 4 gnd
rlabel metal3 s 12600 24595 12698 24693 4 gnd
rlabel metal3 s 12600 25148 12698 25246 4 gnd
rlabel metal3 s 12600 25622 12698 25720 4 gnd
rlabel metal3 s 12600 22462 12698 22560 4 gnd
rlabel metal3 s 12600 24832 12698 24930 4 gnd
rlabel metal3 s 12600 25385 12698 25483 4 gnd
rlabel metal3 s 12600 23252 12698 23350 4 gnd
rlabel metal3 s 12600 21672 12698 21770 4 gnd
rlabel metal3 s 12600 23568 12698 23666 4 gnd
rlabel metal3 s 12600 24042 12698 24140 4 gnd
rlabel metal3 s 12600 22778 12698 22876 4 gnd
rlabel metal3 s 12600 21988 12698 22086 4 gnd
rlabel metal3 s 12600 23015 12698 23113 4 gnd
rlabel metal3 s 12600 22225 12698 22323 4 gnd
rlabel metal3 s 12600 23805 12698 23903 4 gnd
rlabel metal3 s 12600 24358 12698 24456 4 gnd
rlabel metal3 s 7660 22225 7758 22323 4 vdd
rlabel metal3 s 7660 25780 7758 25878 4 vdd
rlabel metal3 s 6450 24223 6548 24321 4 vdd
rlabel metal3 s 6882 25371 6980 25469 4 vdd
rlabel metal3 s 7660 24990 7758 25088 4 vdd
rlabel metal3 s 6882 24581 6980 24679 4 vdd
rlabel metal3 s 6025 25429 6123 25527 4 gnd
rlabel metal3 s 6450 25803 6548 25901 4 vdd
rlabel metal3 s 7264 24595 7362 24693 4 gnd
rlabel metal3 s 6025 25803 6123 25901 4 gnd
rlabel metal3 s 6882 25013 6980 25111 4 vdd
rlabel metal3 s 7660 25385 7758 25483 4 vdd
rlabel metal3 s 6025 22643 6123 22741 4 gnd
rlabel metal3 s 6450 23791 6548 23889 4 vdd
rlabel metal3 s 6450 23001 6548 23099 4 vdd
rlabel metal3 s 7264 21830 7362 21928 4 gnd
rlabel metal3 s 6025 24639 6123 24737 4 gnd
rlabel metal3 s 6882 22643 6980 22741 4 vdd
rlabel metal3 s 6882 23433 6980 23531 4 vdd
rlabel metal3 s 6025 23849 6123 23947 4 gnd
rlabel metal3 s 7660 21830 7758 21928 4 vdd
rlabel metal3 s 7660 23805 7758 23903 4 vdd
rlabel metal3 s 7264 24200 7362 24298 4 gnd
rlabel metal3 s 6450 21853 6548 21951 4 vdd
rlabel metal3 s 6450 25013 6548 25111 4 vdd
rlabel metal3 s 7264 22620 7362 22718 4 gnd
rlabel metal3 s 6882 25803 6980 25901 4 vdd
rlabel metal3 s 7264 23805 7362 23903 4 gnd
rlabel metal3 s 7264 23410 7362 23508 4 gnd
rlabel metal3 s 7660 24595 7758 24693 4 vdd
rlabel metal3 s 6450 22211 6548 22309 4 vdd
rlabel metal3 s 6450 25371 6548 25469 4 vdd
rlabel metal3 s 6025 23433 6123 23531 4 gnd
rlabel metal3 s 6882 21853 6980 21951 4 vdd
rlabel metal3 s 6882 23001 6980 23099 4 vdd
rlabel metal3 s 6882 23791 6980 23889 4 vdd
rlabel metal3 s 6025 23059 6123 23157 4 gnd
rlabel metal3 s 6882 24223 6980 24321 4 vdd
rlabel metal3 s 6882 22211 6980 22309 4 vdd
rlabel metal3 s 6450 24581 6548 24679 4 vdd
rlabel metal3 s 6025 24223 6123 24321 4 gnd
rlabel metal3 s 7264 25780 7362 25878 4 gnd
rlabel metal3 s 7264 24990 7362 25088 4 gnd
rlabel metal3 s 7660 24200 7758 24298 4 vdd
rlabel metal3 s 7264 25385 7362 25483 4 gnd
rlabel metal3 s 6025 21853 6123 21951 4 gnd
rlabel metal3 s 7660 23015 7758 23113 4 vdd
rlabel metal3 s 7264 23015 7362 23113 4 gnd
rlabel metal3 s 6450 23433 6548 23531 4 vdd
rlabel metal3 s 6450 22643 6548 22741 4 vdd
rlabel metal3 s 7660 23410 7758 23508 4 vdd
rlabel metal3 s 6025 22269 6123 22367 4 gnd
rlabel metal3 s 6025 25013 6123 25111 4 gnd
rlabel metal3 s 7660 22620 7758 22718 4 vdd
rlabel metal3 s 7264 22225 7362 22323 4 gnd
rlabel metal3 s 7660 21435 7758 21533 4 vdd
rlabel metal3 s 6025 17903 6123 18001 4 gnd
rlabel metal3 s 6450 21421 6548 21519 4 vdd
rlabel metal3 s 7264 20645 7362 20743 4 gnd
rlabel metal3 s 6882 17903 6980 18001 4 vdd
rlabel metal3 s 6882 21063 6980 21161 4 vdd
rlabel metal3 s 6025 21479 6123 21577 4 gnd
rlabel metal3 s 4246 17880 4344 17978 4 vdd
rlabel metal3 s 7264 18670 7362 18768 4 gnd
rlabel metal3 s 6882 19051 6980 19149 4 vdd
rlabel metal3 s 3468 17903 3566 18001 4 vdd
rlabel metal3 s 7660 20645 7758 20743 4 vdd
rlabel metal3 s 6025 18693 6123 18791 4 gnd
rlabel metal3 s 6025 17529 6123 17627 4 gnd
rlabel metal3 s 6025 18319 6123 18417 4 gnd
rlabel metal3 s 6882 18693 6980 18791 4 vdd
rlabel metal3 s 7660 18275 7758 18373 4 vdd
rlabel metal3 s 7264 18275 7362 18373 4 gnd
rlabel metal3 s 7264 21435 7362 21533 4 gnd
rlabel metal3 s 7264 20250 7362 20348 4 gnd
rlabel metal3 s 7660 20250 7758 20348 4 vdd
rlabel metal3 s 7660 19855 7758 19953 4 vdd
rlabel metal3 s 6450 20631 6548 20729 4 vdd
rlabel metal3 s 6025 19899 6123 19997 4 gnd
rlabel metal3 s 6025 19483 6123 19581 4 gnd
rlabel metal3 s 7660 17485 7758 17583 4 vdd
rlabel metal3 s 7264 17880 7362 17978 4 gnd
rlabel metal3 s 7660 18670 7758 18768 4 vdd
rlabel metal3 s 7660 19065 7758 19163 4 vdd
rlabel metal3 s 6450 18693 6548 18791 4 vdd
rlabel metal3 s 6882 20273 6980 20371 4 vdd
rlabel metal3 s 7264 19855 7362 19953 4 gnd
rlabel metal3 s 6025 21063 6123 21161 4 gnd
rlabel metal3 s 6450 21063 6548 21161 4 vdd
rlabel metal3 s 6025 20689 6123 20787 4 gnd
rlabel metal3 s 7264 19460 7362 19558 4 gnd
rlabel metal3 s 6450 19051 6548 19149 4 vdd
rlabel metal3 s 7264 19065 7362 19163 4 gnd
rlabel metal3 s 6450 19483 6548 19581 4 vdd
rlabel metal3 s 6450 17471 6548 17569 4 vdd
rlabel metal3 s 7660 19460 7758 19558 4 vdd
rlabel metal3 s 6882 17471 6980 17569 4 vdd
rlabel metal3 s 7264 21040 7362 21138 4 gnd
rlabel metal3 s 2611 17903 2709 18001 4 gnd
rlabel metal3 s 7264 17485 7362 17583 4 gnd
rlabel metal3 s 6882 20631 6980 20729 4 vdd
rlabel metal3 s 6882 18261 6980 18359 4 vdd
rlabel metal3 s 7660 21040 7758 21138 4 vdd
rlabel metal3 s 6882 19483 6980 19581 4 vdd
rlabel metal3 s 6450 19841 6548 19939 4 vdd
rlabel metal3 s 6025 20273 6123 20371 4 gnd
rlabel metal3 s 3036 17903 3134 18001 4 vdd
rlabel metal3 s 6882 19841 6980 19939 4 vdd
rlabel metal3 s 6450 18261 6548 18359 4 vdd
rlabel metal3 s 3850 17880 3948 17978 4 gnd
rlabel metal3 s 6882 21421 6980 21519 4 vdd
rlabel metal3 s 6025 19109 6123 19207 4 gnd
rlabel metal3 s 6450 20273 6548 20371 4 vdd
rlabel metal3 s 6450 17903 6548 18001 4 vdd
rlabel metal3 s 7660 17880 7758 17978 4 vdd
rlabel metal3 s 12600 19065 12698 19163 4 gnd
rlabel metal3 s 12600 18828 12698 18926 4 gnd
rlabel metal3 s 12600 20645 12698 20743 4 gnd
rlabel metal3 s 12600 21198 12698 21296 4 gnd
rlabel metal3 s 12600 18275 12698 18373 4 gnd
rlabel metal3 s 12600 19302 12698 19400 4 gnd
rlabel metal3 s 12600 18512 12698 18610 4 gnd
rlabel metal3 s 12600 21435 12698 21533 4 gnd
rlabel metal3 s 12600 20092 12698 20190 4 gnd
rlabel metal3 s 12600 20408 12698 20506 4 gnd
rlabel metal3 s 12600 19618 12698 19716 4 gnd
rlabel metal3 s 12600 17485 12698 17583 4 gnd
rlabel metal3 s 12600 20882 12698 20980 4 gnd
rlabel metal3 s 12600 19855 12698 19953 4 gnd
rlabel metal3 s 12600 18038 12698 18136 4 gnd
rlabel metal3 s 12600 17722 12698 17820 4 gnd
rlabel metal3 s 15792 9814 15890 9912 4 vdd
rlabel metal3 s 20784 9814 20882 9912 4 vdd
rlabel metal3 s 26400 9814 26498 9912 4 vdd
rlabel metal3 s 18793 9223 18891 9321 4 vdd
rlabel metal3 s 18407 9223 18505 9321 4 vdd
rlabel metal3 s 18912 9814 19010 9912 4 vdd
rlabel metal3 s 23280 9814 23378 9912 4 vdd
rlabel metal3 s 19655 9223 19753 9321 4 vdd
rlabel metal3 s 25776 9814 25874 9912 4 vdd
rlabel metal3 s 15049 9223 15147 9321 4 vdd
rlabel metal3 s 16416 9814 16514 9912 4 vdd
rlabel metal3 s 17664 9814 17762 9912 4 vdd
rlabel metal3 s 16297 9223 16395 9321 4 vdd
rlabel metal3 s 21289 9223 21387 9321 4 vdd
rlabel metal3 s 25152 9814 25250 9912 4 vdd
rlabel metal3 s 22032 9814 22130 9912 4 vdd
rlabel metal3 s 22151 9223 22249 9321 4 vdd
rlabel metal3 s 14663 9223 14761 9321 4 vdd
rlabel metal3 s 20041 9223 20139 9321 4 vdd
rlabel metal3 s 25033 9223 25131 9321 4 vdd
rlabel metal3 s 23785 9223 23883 9321 4 vdd
rlabel metal3 s 20160 9814 20258 9912 4 vdd
rlabel metal3 s 21408 9814 21506 9912 4 vdd
rlabel metal3 s 19536 9814 19634 9912 4 vdd
rlabel metal3 s 22656 9814 22754 9912 4 vdd
rlabel metal3 s 14544 9814 14642 9912 4 vdd
rlabel metal3 s 20903 9223 21001 9321 4 vdd
rlabel metal3 s 17545 9223 17643 9321 4 vdd
rlabel metal3 s 23904 9814 24002 9912 4 vdd
rlabel metal3 s 24528 9814 24626 9912 4 vdd
rlabel metal3 s 15168 9814 15266 9912 4 vdd
rlabel metal3 s 24647 9223 24745 9321 4 vdd
rlabel metal3 s 22537 9223 22635 9321 4 vdd
rlabel metal3 s 15911 9223 16009 9321 4 vdd
rlabel metal3 s 27143 9223 27241 9321 4 vdd
rlabel metal3 s 17040 9814 17138 9912 4 vdd
rlabel metal3 s 18288 9814 18386 9912 4 vdd
rlabel metal3 s 23399 9223 23497 9321 4 vdd
rlabel metal3 s 27024 9814 27122 9912 4 vdd
rlabel metal3 s 26281 9223 26379 9321 4 vdd
rlabel metal3 s 17159 9223 17257 9321 4 vdd
rlabel metal3 s 25895 9223 25993 9321 4 vdd
rlabel metal3 s 12600 13535 12698 13633 4 gnd
rlabel metal3 s 12600 16458 12698 16556 4 gnd
rlabel metal3 s 12600 14088 12698 14186 4 gnd
rlabel metal3 s 12600 12982 12698 13080 4 gnd
rlabel metal3 s 12600 13298 12698 13396 4 gnd
rlabel metal3 s 12600 14562 12698 14660 4 gnd
rlabel metal3 s 12600 16142 12698 16240 4 gnd
rlabel metal3 s 12600 17248 12698 17346 4 gnd
rlabel metal3 s 12600 15352 12698 15450 4 gnd
rlabel metal3 s 12600 16695 12698 16793 4 gnd
rlabel metal3 s 12600 13772 12698 13870 4 gnd
rlabel metal3 s 12600 15905 12698 16003 4 gnd
rlabel metal3 s 12600 15668 12698 15766 4 gnd
rlabel metal3 s 12600 16932 12698 17030 4 gnd
rlabel metal3 s 12600 14878 12698 14976 4 gnd
rlabel metal3 s 12600 14325 12698 14423 4 gnd
rlabel metal3 s 12600 15115 12698 15213 4 gnd
rlabel metal3 s 7264 13930 7362 14028 4 gnd
rlabel metal3 s 6450 14311 6548 14409 4 vdd
rlabel metal3 s 6882 13953 6980 14051 4 vdd
rlabel metal3 s 4246 15510 4344 15608 4 vdd
rlabel metal3 s 7660 13535 7758 13633 4 vdd
rlabel metal3 s 6025 15159 6123 15257 4 gnd
rlabel metal3 s 6450 16681 6548 16779 4 vdd
rlabel metal3 s 3036 16323 3134 16421 4 vdd
rlabel metal3 s 6882 16681 6980 16779 4 vdd
rlabel metal3 s 6025 15949 6123 16047 4 gnd
rlabel metal3 s 6025 13163 6123 13261 4 gnd
rlabel metal3 s 6025 15533 6123 15631 4 gnd
rlabel metal3 s 6025 13579 6123 13677 4 gnd
rlabel metal3 s 6450 15533 6548 15631 4 vdd
rlabel metal3 s 7264 15115 7362 15213 4 gnd
rlabel metal3 s 6882 15101 6980 15199 4 vdd
rlabel metal3 s 7264 13140 7362 13238 4 gnd
rlabel metal3 s 7660 14325 7758 14423 4 vdd
rlabel metal3 s 6025 17113 6123 17211 4 gnd
rlabel metal3 s 6450 15891 6548 15989 4 vdd
rlabel metal3 s 7660 14720 7758 14818 4 vdd
rlabel metal3 s 1752 13140 1850 13238 4 gnd
rlabel metal3 s 4246 13930 4344 14028 4 vdd
rlabel metal3 s 2611 16323 2709 16421 4 gnd
rlabel metal3 s 7660 16300 7758 16398 4 vdd
rlabel metal3 s 7264 14720 7362 14818 4 gnd
rlabel metal3 s 2611 15533 2709 15631 4 gnd
rlabel metal3 s 3850 13140 3948 13238 4 gnd
rlabel metal3 s 6450 14743 6548 14841 4 vdd
rlabel metal3 s 7264 14325 7362 14423 4 gnd
rlabel metal3 s 3850 15510 3948 15608 4 gnd
rlabel metal3 s 4246 16300 4344 16398 4 vdd
rlabel metal3 s 7660 13930 7758 14028 4 vdd
rlabel metal3 s 2611 17113 2709 17211 4 gnd
rlabel metal3 s 7660 13140 7758 13238 4 vdd
rlabel metal3 s 4246 13140 4344 13238 4 vdd
rlabel metal3 s 7660 17090 7758 17188 4 vdd
rlabel metal3 s 6025 14743 6123 14841 4 gnd
rlabel metal3 s 6450 13163 6548 13261 4 vdd
rlabel metal3 s 3046 13937 3144 14035 4 gnd
rlabel metal3 s 7264 17090 7362 17188 4 gnd
rlabel metal3 s 2148 13140 2246 13238 4 vdd
rlabel metal3 s 6882 14743 6980 14841 4 vdd
rlabel metal3 s 6882 16323 6980 16421 4 vdd
rlabel metal3 s 7264 13535 7362 13633 4 gnd
rlabel metal3 s 6025 16739 6123 16837 4 gnd
rlabel metal3 s 7660 16695 7758 16793 4 vdd
rlabel metal3 s 6882 17113 6980 17211 4 vdd
rlabel metal3 s 6882 13163 6980 13261 4 vdd
rlabel metal3 s 6025 16323 6123 16421 4 gnd
rlabel metal3 s 3036 17113 3134 17211 4 vdd
rlabel metal3 s 7660 15905 7758 16003 4 vdd
rlabel metal3 s 3471 13147 3569 13245 4 vdd
rlabel metal3 s 3471 13937 3569 14035 4 vdd
rlabel metal3 s 6450 17113 6548 17211 4 vdd
rlabel metal3 s 6025 13953 6123 14051 4 gnd
rlabel metal3 s 6882 14311 6980 14409 4 vdd
rlabel metal3 s 6450 13953 6548 14051 4 vdd
rlabel metal3 s 3036 15533 3134 15631 4 vdd
rlabel metal3 s 7264 16695 7362 16793 4 gnd
rlabel metal3 s 6450 13521 6548 13619 4 vdd
rlabel metal3 s 1552 15510 1650 15608 4 vdd
rlabel metal3 s 1156 15510 1254 15608 4 gnd
rlabel metal3 s 7264 15510 7362 15608 4 gnd
rlabel metal3 s 6450 15101 6548 15199 4 vdd
rlabel metal3 s 3850 17090 3948 17188 4 gnd
rlabel metal3 s 3468 17113 3566 17211 4 vdd
rlabel metal3 s 3468 15533 3566 15631 4 vdd
rlabel metal3 s 6025 14369 6123 14467 4 gnd
rlabel metal3 s 3468 16323 3566 16421 4 vdd
rlabel metal3 s 4246 17090 4344 17188 4 vdd
rlabel metal3 s 3046 13147 3144 13245 4 gnd
rlabel metal3 s 6882 15891 6980 15989 4 vdd
rlabel metal3 s 6450 16323 6548 16421 4 vdd
rlabel metal3 s 6882 15533 6980 15631 4 vdd
rlabel metal3 s 3850 13930 3948 14028 4 gnd
rlabel metal3 s 7264 16300 7362 16398 4 gnd
rlabel metal3 s 7660 15510 7758 15608 4 vdd
rlabel metal3 s 6882 13521 6980 13619 4 vdd
rlabel metal3 s 7660 15115 7758 15213 4 vdd
rlabel metal3 s 7264 15905 7362 16003 4 gnd
rlabel metal3 s 3850 16300 3948 16398 4 gnd
rlabel metal3 s 7264 11955 7362 12053 4 gnd
rlabel metal3 s 3046 10777 3144 10875 4 gnd
rlabel metal3 s 7264 11165 7362 11263 4 gnd
rlabel metal3 s 4246 11560 4344 11658 4 vdd
rlabel metal3 s 6025 11209 6123 11307 4 gnd
rlabel metal3 s 7264 12350 7362 12448 4 gnd
rlabel metal3 s 7264 10770 7362 10868 4 gnd
rlabel metal3 s 6450 11941 6548 12039 4 vdd
rlabel metal3 s 1752 10770 1850 10868 4 gnd
rlabel metal3 s 7264 12745 7362 12843 4 gnd
rlabel metal3 s 7660 11560 7758 11658 4 vdd
rlabel metal3 s 2148 10770 2246 10868 4 vdd
rlabel metal3 s 6882 12373 6980 12471 4 vdd
rlabel metal3 s 6882 11941 6980 12039 4 vdd
rlabel metal3 s 7264 11560 7362 11658 4 gnd
rlabel metal3 s 7660 12350 7758 12448 4 vdd
rlabel metal3 s 6025 11583 6123 11681 4 gnd
rlabel metal3 s 7660 11165 7758 11263 4 vdd
rlabel metal3 s 6450 11151 6548 11249 4 vdd
rlabel metal3 s 6882 11151 6980 11249 4 vdd
rlabel metal3 s 3850 11560 3948 11658 4 gnd
rlabel metal3 s 6450 12731 6548 12829 4 vdd
rlabel metal3 s 7660 12745 7758 12843 4 vdd
rlabel metal3 s 6882 12731 6980 12829 4 vdd
rlabel metal3 s 3046 11567 3144 11665 4 gnd
rlabel metal3 s 6025 11999 6123 12097 4 gnd
rlabel metal3 s 4246 10770 4344 10868 4 vdd
rlabel metal3 s 6450 10793 6548 10891 4 vdd
rlabel metal3 s 6025 12373 6123 12471 4 gnd
rlabel metal3 s 6025 10793 6123 10891 4 gnd
rlabel metal3 s 6450 12373 6548 12471 4 vdd
rlabel metal3 s 6450 11583 6548 11681 4 vdd
rlabel metal3 s 7685 10184 7783 10282 4 vdd
rlabel metal3 s 6882 11583 6980 11681 4 vdd
rlabel metal3 s 3850 10770 3948 10868 4 gnd
rlabel metal3 s 6882 10793 6980 10891 4 vdd
rlabel metal3 s 3471 11567 3569 11665 4 vdd
rlabel metal3 s 3471 10777 3569 10875 4 vdd
rlabel metal3 s 6025 12789 6123 12887 4 gnd
rlabel metal3 s 7660 10770 7758 10868 4 vdd
rlabel metal3 s 7660 11955 7758 12053 4 vdd
rlabel metal3 s 13296 9814 13394 9912 4 vdd
rlabel metal3 s 12600 12508 12698 12606 4 gnd
rlabel metal3 s 12600 10375 12698 10473 4 gnd
rlabel metal3 s 12234 10248 12332 10346 4 gnd
rlabel metal3 s 11208 10178 11306 10276 4 vdd
rlabel metal3 s 13801 9223 13899 9321 4 vdd
rlabel metal3 s 12600 11165 12698 11263 4 gnd
rlabel metal3 s 12600 12192 12698 12290 4 gnd
rlabel metal3 s 12600 11718 12698 11816 4 gnd
rlabel metal3 s 12600 10612 12698 10710 4 gnd
rlabel metal3 s 12600 10928 12698 11026 4 gnd
rlabel metal3 s 8517 10190 8615 10288 4 vdd
rlabel metal3 s 13415 9223 13513 9321 4 vdd
rlabel metal3 s 12600 12745 12698 12843 4 gnd
rlabel metal3 s 13920 9814 14018 9912 4 vdd
rlabel metal3 s 12600 11402 12698 11500 4 gnd
rlabel metal3 s 12600 11955 12698 12053 4 gnd
rlabel metal3 s 6472 4989 6570 5087 4 gnd
rlabel metal3 s 13989 3743 14087 3841 4 gnd
rlabel metal3 s 6472 2161 6570 2259 4 gnd
rlabel metal3 s 13989 4065 14087 4163 4 vdd
rlabel metal3 s 5360 6403 5458 6501 4 vdd
rlabel metal3 s 0 8474 13577 8534 4 rbl_bl_0_0
rlabel metal3 s 6472 3575 6570 3673 4 vdd
rlabel metal3 s 13884 1563 13982 1661 4 vdd
rlabel metal3 s 12234 1120 12332 1218 4 vdd
rlabel metal3 s 6472 7817 6570 7915 4 gnd
rlabel metal3 s 14059 5677 14157 5775 4 gnd
rlabel metal3 s 5360 3575 5458 3673 4 vdd
rlabel metal3 s 14232 7674 14330 7772 4 gnd
rlabel metal3 s 5360 7817 5458 7915 4 gnd
rlabel metal3 s 13985 2181 14083 2279 4 gnd
rlabel metal3 s 5360 2161 5458 2259 4 gnd
rlabel metal3 s 12234 0 12332 98 4 gnd
rlabel metal3 s 13875 2950 13973 3048 4 gnd
rlabel metal3 s 5360 4989 5458 5087 4 gnd
rlabel metal3 s 13864 2513 13962 2611 4 vdd
rlabel metal3 s 13870 1979 13968 2077 4 gnd
rlabel metal3 s 13977 4903 14075 5001 4 vdd
rlabel metal3 s 6472 6403 6570 6501 4 vdd
rlabel metal3 s 18876 1563 18974 1661 4 vdd
rlabel metal3 s 18867 2950 18965 3048 4 gnd
rlabel metal3 s 21473 2181 21571 2279 4 gnd
rlabel metal3 s 18862 1979 18960 2077 4 gnd
rlabel metal3 s 21372 1563 21470 1661 4 vdd
rlabel metal3 s 16481 2181 16579 2279 4 gnd
rlabel metal3 s 26469 3743 26567 3841 4 gnd
rlabel metal3 s 21547 5677 21645 5775 4 gnd
rlabel metal3 s 25464 7674 25562 7772 4 gnd
rlabel metal3 s 17976 7674 18074 7772 4 gnd
rlabel metal3 s 21358 1979 21456 2077 4 gnd
rlabel metal3 s 19224 7674 19322 7772 4 gnd
rlabel metal3 s 22968 7674 23066 7772 4 gnd
rlabel metal3 s 16366 1979 16464 2077 4 gnd
rlabel metal3 s 21477 4065 21575 4163 4 vdd
rlabel metal3 s 16473 4903 16571 5001 4 vdd
rlabel metal3 s 20472 7674 20570 7772 4 gnd
rlabel metal3 s 26469 4065 26567 4163 4 vdd
rlabel metal3 s 16555 5677 16653 5775 4 gnd
rlabel metal3 s 26465 2181 26563 2279 4 gnd
rlabel metal3 s 23854 1979 23952 2077 4 gnd
rlabel metal3 s 24216 7674 24314 7772 4 gnd
rlabel metal3 s 26350 1979 26448 2077 4 gnd
rlabel metal3 s 18981 3743 19079 3841 4 gnd
rlabel metal3 s 26712 7674 26810 7772 4 gnd
rlabel metal3 s 23969 2181 24067 2279 4 gnd
rlabel metal3 s 18981 4065 19079 4163 4 vdd
rlabel metal3 s 16380 1563 16478 1661 4 vdd
rlabel metal3 s 16485 4065 16583 4163 4 vdd
rlabel metal3 s 23848 2513 23946 2611 4 vdd
rlabel metal3 s 16485 3743 16583 3841 4 gnd
rlabel metal3 s 26344 2513 26442 2611 4 vdd
rlabel metal3 s 16360 2513 16458 2611 4 vdd
rlabel metal3 s 18856 2513 18954 2611 4 vdd
rlabel metal3 s 26539 5677 26637 5775 4 gnd
rlabel metal3 s 16371 2950 16469 3048 4 gnd
rlabel metal3 s 26457 4903 26555 5001 4 vdd
rlabel metal3 s 21363 2950 21461 3048 4 gnd
rlabel metal3 s 23868 1563 23966 1661 4 vdd
rlabel metal3 s 23973 4065 24071 4163 4 vdd
rlabel metal3 s 26364 1563 26462 1661 4 vdd
rlabel metal3 s 16728 7674 16826 7772 4 gnd
rlabel metal3 s 18969 4903 19067 5001 4 vdd
rlabel metal3 s 21477 3743 21575 3841 4 gnd
rlabel metal3 s 24043 5677 24141 5775 4 gnd
rlabel metal3 s 21720 7674 21818 7772 4 gnd
rlabel metal3 s 23973 3743 24071 3841 4 gnd
rlabel metal3 s 23859 2950 23957 3048 4 gnd
rlabel metal3 s 21352 2513 21450 2611 4 vdd
rlabel metal3 s 18977 2181 19075 2279 4 gnd
rlabel metal3 s 15480 7674 15578 7772 4 gnd
rlabel metal3 s 26355 2950 26453 3048 4 gnd
rlabel metal3 s 19051 5677 19149 5775 4 gnd
rlabel metal3 s 21465 4903 21563 5001 4 vdd
rlabel metal3 s 23961 4903 24059 5001 4 vdd
rlabel metal3 s 48240 9814 48338 9912 4 vdd
rlabel metal3 s 43367 9223 43465 9321 4 vdd
rlabel metal3 s 49488 9814 49586 9912 4 vdd
rlabel metal3 s 48745 9223 48843 9321 4 vdd
rlabel metal3 s 42000 9814 42098 9912 4 vdd
rlabel metal3 s 42505 9223 42603 9321 4 vdd
rlabel metal3 s 50855 9223 50953 9321 4 vdd
rlabel metal3 s 49607 9223 49705 9321 4 vdd
rlabel metal3 s 45863 9223 45961 9321 4 vdd
rlabel metal3 s 52489 9223 52587 9321 4 vdd
rlabel metal3 s 47497 9223 47595 9321 4 vdd
rlabel metal3 s 50112 9814 50210 9912 4 vdd
rlabel metal3 s 41376 9814 41474 9912 4 vdd
rlabel metal3 s 42119 9223 42217 9321 4 vdd
rlabel metal3 s 51984 9814 52082 9912 4 vdd
rlabel metal3 s 52608 9814 52706 9912 4 vdd
rlabel metal3 s 51241 9223 51339 9321 4 vdd
rlabel metal3 s 43872 9814 43970 9912 4 vdd
rlabel metal3 s 45744 9814 45842 9912 4 vdd
rlabel metal3 s 46992 9814 47090 9912 4 vdd
rlabel metal3 s 46368 9814 46466 9912 4 vdd
rlabel metal3 s 49993 9223 50091 9321 4 vdd
rlabel metal3 s 42624 9814 42722 9912 4 vdd
rlabel metal3 s 44496 9814 44594 9912 4 vdd
rlabel metal3 s 47616 9814 47714 9912 4 vdd
rlabel metal3 s 40871 9223 40969 9321 4 vdd
rlabel metal3 s 43248 9814 43346 9912 4 vdd
rlabel metal3 s 51360 9814 51458 9912 4 vdd
rlabel metal3 s 53232 9814 53330 9912 4 vdd
rlabel metal3 s 53351 9223 53449 9321 4 vdd
rlabel metal3 s 45120 9814 45218 9912 4 vdd
rlabel metal3 s 52103 9223 52201 9321 4 vdd
rlabel metal3 s 40752 9814 40850 9912 4 vdd
rlabel metal3 s 43753 9223 43851 9321 4 vdd
rlabel metal3 s 48359 9223 48457 9321 4 vdd
rlabel metal3 s 48864 9814 48962 9912 4 vdd
rlabel metal3 s 45001 9223 45099 9321 4 vdd
rlabel metal3 s 47111 9223 47209 9321 4 vdd
rlabel metal3 s 50736 9814 50834 9912 4 vdd
rlabel metal3 s 41257 9223 41355 9321 4 vdd
rlabel metal3 s 46249 9223 46347 9321 4 vdd
rlabel metal3 s 44615 9223 44713 9321 4 vdd
rlabel metal3 s 37513 9223 37611 9321 4 vdd
rlabel metal3 s 37632 9814 37730 9912 4 vdd
rlabel metal3 s 36384 9814 36482 9912 4 vdd
rlabel metal3 s 29520 9814 29618 9912 4 vdd
rlabel metal3 s 38880 9814 38978 9912 4 vdd
rlabel metal3 s 34512 9814 34610 9912 4 vdd
rlabel metal3 s 32640 9814 32738 9912 4 vdd
rlabel metal3 s 35017 9223 35115 9321 4 vdd
rlabel metal3 s 37008 9814 37106 9912 4 vdd
rlabel metal3 s 28272 9814 28370 9912 4 vdd
rlabel metal3 s 32521 9223 32619 9321 4 vdd
rlabel metal3 s 40128 9814 40226 9912 4 vdd
rlabel metal3 s 35136 9814 35234 9912 4 vdd
rlabel metal3 s 30144 9814 30242 9912 4 vdd
rlabel metal3 s 28391 9223 28489 9321 4 vdd
rlabel metal3 s 27648 9814 27746 9912 4 vdd
rlabel metal3 s 40009 9223 40107 9321 4 vdd
rlabel metal3 s 27529 9223 27627 9321 4 vdd
rlabel metal3 s 30025 9223 30123 9321 4 vdd
rlabel metal3 s 34631 9223 34729 9321 4 vdd
rlabel metal3 s 31392 9814 31490 9912 4 vdd
rlabel metal3 s 28896 9814 28994 9912 4 vdd
rlabel metal3 s 30768 9814 30866 9912 4 vdd
rlabel metal3 s 29639 9223 29737 9321 4 vdd
rlabel metal3 s 35760 9814 35858 9912 4 vdd
rlabel metal3 s 36265 9223 36363 9321 4 vdd
rlabel metal3 s 31273 9223 31371 9321 4 vdd
rlabel metal3 s 33888 9814 33986 9912 4 vdd
rlabel metal3 s 32016 9814 32114 9912 4 vdd
rlabel metal3 s 38761 9223 38859 9321 4 vdd
rlabel metal3 s 33264 9814 33362 9912 4 vdd
rlabel metal3 s 32135 9223 32233 9321 4 vdd
rlabel metal3 s 39623 9223 39721 9321 4 vdd
rlabel metal3 s 38256 9814 38354 9912 4 vdd
rlabel metal3 s 39504 9814 39602 9912 4 vdd
rlabel metal3 s 35879 9223 35977 9321 4 vdd
rlabel metal3 s 38375 9223 38473 9321 4 vdd
rlabel metal3 s 37127 9223 37225 9321 4 vdd
rlabel metal3 s 33383 9223 33481 9321 4 vdd
rlabel metal3 s 28777 9223 28875 9321 4 vdd
rlabel metal3 s 30887 9223 30985 9321 4 vdd
rlabel metal3 s 33769 9223 33867 9321 4 vdd
rlabel metal3 s 38949 4065 39047 4163 4 vdd
rlabel metal3 s 38937 4903 39035 5001 4 vdd
rlabel metal3 s 38949 3743 39047 3841 4 gnd
rlabel metal3 s 28953 4903 29051 5001 4 vdd
rlabel metal3 s 36441 4903 36539 5001 4 vdd
rlabel metal3 s 31461 4065 31559 4163 4 vdd
rlabel metal3 s 39192 7674 39290 7772 4 gnd
rlabel metal3 s 36696 7674 36794 7772 4 gnd
rlabel metal3 s 38824 2513 38922 2611 4 vdd
rlabel metal3 s 36339 2950 36437 3048 4 gnd
rlabel metal3 s 36453 4065 36551 4163 4 vdd
rlabel metal3 s 31336 2513 31434 2611 4 vdd
rlabel metal3 s 30456 7674 30554 7772 4 gnd
rlabel metal3 s 33852 1563 33950 1661 4 vdd
rlabel metal3 s 36453 3743 36551 3841 4 gnd
rlabel metal3 s 28840 2513 28938 2611 4 vdd
rlabel metal3 s 31356 1563 31454 1661 4 vdd
rlabel metal3 s 40440 7674 40538 7772 4 gnd
rlabel metal3 s 29035 5677 29133 5775 4 gnd
rlabel metal3 s 27960 7674 28058 7772 4 gnd
rlabel metal3 s 33945 4903 34043 5001 4 vdd
rlabel metal3 s 37944 7674 38042 7772 4 gnd
rlabel metal3 s 38830 1979 38928 2077 4 gnd
rlabel metal3 s 34200 7674 34298 7772 4 gnd
rlabel metal3 s 31531 5677 31629 5775 4 gnd
rlabel metal3 s 28860 1563 28958 1661 4 vdd
rlabel metal3 s 36328 2513 36426 2611 4 vdd
rlabel metal3 s 28846 1979 28944 2077 4 gnd
rlabel metal3 s 31704 7674 31802 7772 4 gnd
rlabel metal3 s 33957 3743 34055 3841 4 gnd
rlabel metal3 s 35448 7674 35546 7772 4 gnd
rlabel metal3 s 28851 2950 28949 3048 4 gnd
rlabel metal3 s 38835 2950 38933 3048 4 gnd
rlabel metal3 s 34027 5677 34125 5775 4 gnd
rlabel metal3 s 33957 4065 34055 4163 4 vdd
rlabel metal3 s 28965 4065 29063 4163 4 vdd
rlabel metal3 s 33843 2950 33941 3048 4 gnd
rlabel metal3 s 31347 2950 31445 3048 4 gnd
rlabel metal3 s 31342 1979 31440 2077 4 gnd
rlabel metal3 s 28961 2181 29059 2279 4 gnd
rlabel metal3 s 32952 7674 33050 7772 4 gnd
rlabel metal3 s 39019 5677 39117 5775 4 gnd
rlabel metal3 s 36449 2181 36547 2279 4 gnd
rlabel metal3 s 33838 1979 33936 2077 4 gnd
rlabel metal3 s 38844 1563 38942 1661 4 vdd
rlabel metal3 s 31449 4903 31547 5001 4 vdd
rlabel metal3 s 36348 1563 36446 1661 4 vdd
rlabel metal3 s 28965 3743 29063 3841 4 gnd
rlabel metal3 s 31457 2181 31555 2279 4 gnd
rlabel metal3 s 36523 5677 36621 5775 4 gnd
rlabel metal3 s 38945 2181 39043 2279 4 gnd
rlabel metal3 s 33953 2181 34051 2279 4 gnd
rlabel metal3 s 36334 1979 36432 2077 4 gnd
rlabel metal3 s 29208 7674 29306 7772 4 gnd
rlabel metal3 s 33832 2513 33930 2611 4 vdd
rlabel metal3 s 31461 3743 31559 3841 4 gnd
rlabel metal3 s 49003 5677 49101 5775 4 gnd
rlabel metal3 s 43816 2513 43914 2611 4 vdd
rlabel metal3 s 52920 7674 53018 7772 4 gnd
rlabel metal3 s 51417 4903 51515 5001 4 vdd
rlabel metal3 s 50424 7674 50522 7772 4 gnd
rlabel metal3 s 46433 2181 46531 2279 4 gnd
rlabel metal3 s 51429 4065 51527 4163 4 vdd
rlabel metal3 s 43827 2950 43925 3048 4 gnd
rlabel metal3 s 48933 4065 49031 4163 4 vdd
rlabel metal3 s 51324 1563 51422 1661 4 vdd
rlabel metal3 s 43822 1979 43920 2077 4 gnd
rlabel metal3 s 44011 5677 44109 5775 4 gnd
rlabel metal3 s 46323 2950 46421 3048 4 gnd
rlabel metal3 s 51304 2513 51402 2611 4 vdd
rlabel metal3 s 51672 7674 51770 7772 4 gnd
rlabel metal3 s 43937 2181 44035 2279 4 gnd
rlabel metal3 s 48814 1979 48912 2077 4 gnd
rlabel metal3 s 51315 2950 51413 3048 4 gnd
rlabel metal3 s 43941 3743 44039 3841 4 gnd
rlabel metal3 s 49176 7674 49274 7772 4 gnd
rlabel metal3 s 48819 2950 48917 3048 4 gnd
rlabel metal3 s 45432 7674 45530 7772 4 gnd
rlabel metal3 s 48808 2513 48906 2611 4 vdd
rlabel metal3 s 41688 7674 41786 7772 4 gnd
rlabel metal3 s 41433 4903 41531 5001 4 vdd
rlabel metal3 s 46425 4903 46523 5001 4 vdd
rlabel metal3 s 51429 3743 51527 3841 4 gnd
rlabel metal3 s 51499 5677 51597 5775 4 gnd
rlabel metal3 s 48933 3743 49031 3841 4 gnd
rlabel metal3 s 46437 3743 46535 3841 4 gnd
rlabel metal3 s 41340 1563 41438 1661 4 vdd
rlabel metal3 s 51310 1979 51408 2077 4 gnd
rlabel metal3 s 46507 5677 46605 5775 4 gnd
rlabel metal3 s 41445 3743 41543 3841 4 gnd
rlabel metal3 s 41445 4065 41543 4163 4 vdd
rlabel metal3 s 41515 5677 41613 5775 4 gnd
rlabel metal3 s 44184 7674 44282 7772 4 gnd
rlabel metal3 s 41326 1979 41424 2077 4 gnd
rlabel metal3 s 46318 1979 46416 2077 4 gnd
rlabel metal3 s 42936 7674 43034 7772 4 gnd
rlabel metal3 s 41331 2950 41429 3048 4 gnd
rlabel metal3 s 48929 2181 49027 2279 4 gnd
rlabel metal3 s 46312 2513 46410 2611 4 vdd
rlabel metal3 s 41441 2181 41539 2279 4 gnd
rlabel metal3 s 43836 1563 43934 1661 4 vdd
rlabel metal3 s 46332 1563 46430 1661 4 vdd
rlabel metal3 s 43929 4903 44027 5001 4 vdd
rlabel metal3 s 48921 4903 49019 5001 4 vdd
rlabel metal3 s 51425 2181 51523 2279 4 gnd
rlabel metal3 s 47928 7674 48026 7772 4 gnd
rlabel metal3 s 46437 4065 46535 4163 4 vdd
rlabel metal3 s 46680 7674 46778 7772 4 gnd
rlabel metal3 s 41320 2513 41418 2611 4 vdd
rlabel metal3 s 48828 1563 48926 1661 4 vdd
rlabel metal3 s 43941 4065 44039 4163 4 vdd
rlabel metal3 s 100638 32481 100736 32579 4 vdd
rlabel metal3 s 100206 33271 100304 33369 4 vdd
rlabel metal3 s 99824 33285 99922 33383 4 gnd
rlabel metal3 s 99824 32890 99922 32988 4 gnd
rlabel metal3 s 99428 34470 99526 34568 4 vdd
rlabel metal3 s 100638 33703 100736 33801 4 vdd
rlabel metal3 s 99824 34470 99922 34568 4 gnd
rlabel metal3 s 101063 32913 101161 33011 4 gnd
rlabel metal3 s 101063 32539 101161 32637 4 gnd
rlabel metal3 s 100206 31333 100304 31431 4 vdd
rlabel metal3 s 99428 33680 99526 33778 4 vdd
rlabel metal3 s 99428 32890 99526 32988 4 vdd
rlabel metal3 s 100638 33271 100736 33369 4 vdd
rlabel metal3 s 99824 32100 99922 32198 4 gnd
rlabel metal3 s 100206 33703 100304 33801 4 vdd
rlabel metal3 s 100206 32481 100304 32579 4 vdd
rlabel metal3 s 99428 30915 99526 31013 4 vdd
rlabel metal3 s 99428 33285 99526 33383 4 vdd
rlabel metal3 s 100206 32913 100304 33011 4 vdd
rlabel metal3 s 99824 30520 99922 30618 4 gnd
rlabel metal3 s 99824 34075 99922 34173 4 gnd
rlabel metal3 s 100206 30901 100304 30999 4 vdd
rlabel metal3 s 101063 33329 101161 33427 4 gnd
rlabel metal3 s 99428 34075 99526 34173 4 vdd
rlabel metal3 s 101063 30959 101161 31057 4 gnd
rlabel metal3 s 100638 30901 100736 30999 4 vdd
rlabel metal3 s 99428 30520 99526 30618 4 vdd
rlabel metal3 s 100206 32123 100304 32221 4 vdd
rlabel metal3 s 100638 34493 100736 34591 4 vdd
rlabel metal3 s 100638 30543 100736 30641 4 vdd
rlabel metal3 s 100638 34061 100736 34159 4 vdd
rlabel metal3 s 100638 32913 100736 33011 4 vdd
rlabel metal3 s 99824 31705 99922 31803 4 gnd
rlabel metal3 s 100206 30543 100304 30641 4 vdd
rlabel metal3 s 99428 31310 99526 31408 4 vdd
rlabel metal3 s 99824 30915 99922 31013 4 gnd
rlabel metal3 s 100206 34061 100304 34159 4 vdd
rlabel metal3 s 99428 31705 99526 31803 4 vdd
rlabel metal3 s 101063 31749 101161 31847 4 gnd
rlabel metal3 s 101063 30543 101161 30641 4 gnd
rlabel metal3 s 101063 34493 101161 34591 4 gnd
rlabel metal3 s 100638 31333 100736 31431 4 vdd
rlabel metal3 s 101063 32123 101161 32221 4 gnd
rlabel metal3 s 100638 32123 100736 32221 4 vdd
rlabel metal3 s 101063 33703 101161 33801 4 gnd
rlabel metal3 s 101063 31333 101161 31431 4 gnd
rlabel metal3 s 100206 31691 100304 31789 4 vdd
rlabel metal3 s 101063 34119 101161 34217 4 gnd
rlabel metal3 s 99428 32495 99526 32593 4 vdd
rlabel metal3 s 99824 31310 99922 31408 4 gnd
rlabel metal3 s 99824 33680 99922 33778 4 gnd
rlabel metal3 s 99428 32100 99526 32198 4 vdd
rlabel metal3 s 100638 31691 100736 31789 4 vdd
rlabel metal3 s 100206 34493 100304 34591 4 vdd
rlabel metal3 s 99824 32495 99922 32593 4 gnd
rlabel metal3 s 94488 33522 94586 33620 4 gnd
rlabel metal3 s 94488 33048 94586 33146 4 gnd
rlabel metal3 s 94488 33285 94586 33383 4 gnd
rlabel metal3 s 94488 32732 94586 32830 4 gnd
rlabel metal3 s 94488 34075 94586 34173 4 gnd
rlabel metal3 s 94488 32495 94586 32593 4 gnd
rlabel metal3 s 94488 33838 94586 33936 4 gnd
rlabel metal3 s 94488 31705 94586 31803 4 gnd
rlabel metal3 s 94488 31152 94586 31250 4 gnd
rlabel metal3 s 94488 30915 94586 31013 4 gnd
rlabel metal3 s 94488 32258 94586 32356 4 gnd
rlabel metal3 s 94488 31468 94586 31566 4 gnd
rlabel metal3 s 94488 30678 94586 30776 4 gnd
rlabel metal3 s 94488 34312 94586 34410 4 gnd
rlabel metal3 s 94488 30362 94586 30460 4 gnd
rlabel metal3 s 94488 31942 94586 32040 4 gnd
rlabel metal3 s 94488 28782 94586 28880 4 gnd
rlabel metal3 s 94488 29098 94586 29196 4 gnd
rlabel metal3 s 94488 30125 94586 30223 4 gnd
rlabel metal3 s 94488 29572 94586 29670 4 gnd
rlabel metal3 s 94488 27518 94586 27616 4 gnd
rlabel metal3 s 94488 26965 94586 27063 4 gnd
rlabel metal3 s 94488 29335 94586 29433 4 gnd
rlabel metal3 s 94488 27755 94586 27853 4 gnd
rlabel metal3 s 94488 27992 94586 28090 4 gnd
rlabel metal3 s 94488 28545 94586 28643 4 gnd
rlabel metal3 s 94488 29888 94586 29986 4 gnd
rlabel metal3 s 94488 25938 94586 26036 4 gnd
rlabel metal3 s 94488 26175 94586 26273 4 gnd
rlabel metal3 s 94488 26412 94586 26510 4 gnd
rlabel metal3 s 94488 27202 94586 27300 4 gnd
rlabel metal3 s 94488 26728 94586 26826 4 gnd
rlabel metal3 s 94488 28308 94586 28406 4 gnd
rlabel metal3 s 99428 28940 99526 29038 4 vdd
rlabel metal3 s 100638 27383 100736 27481 4 vdd
rlabel metal3 s 101063 26593 101161 26691 4 gnd
rlabel metal3 s 99824 26965 99922 27063 4 gnd
rlabel metal3 s 99824 30125 99922 30223 4 gnd
rlabel metal3 s 100206 28173 100304 28271 4 vdd
rlabel metal3 s 100206 28963 100304 29061 4 vdd
rlabel metal3 s 101063 29379 101161 29477 4 gnd
rlabel metal3 s 100206 29753 100304 29851 4 vdd
rlabel metal3 s 100638 26951 100736 27049 4 vdd
rlabel metal3 s 101063 28173 101161 28271 4 gnd
rlabel metal3 s 100638 27741 100736 27839 4 vdd
rlabel metal3 s 99824 27360 99922 27458 4 gnd
rlabel metal3 s 99824 28150 99922 28248 4 gnd
rlabel metal3 s 101063 26219 101161 26317 4 gnd
rlabel metal3 s 100638 26593 100736 26691 4 vdd
rlabel metal3 s 100638 28963 100736 29061 4 vdd
rlabel metal3 s 100206 26593 100304 26691 4 vdd
rlabel metal3 s 99428 28545 99526 28643 4 vdd
rlabel metal3 s 99824 29730 99922 29828 4 gnd
rlabel metal3 s 99428 26965 99526 27063 4 vdd
rlabel metal3 s 100206 26951 100304 27049 4 vdd
rlabel metal3 s 100638 29321 100736 29419 4 vdd
rlabel metal3 s 99428 26175 99526 26273 4 vdd
rlabel metal3 s 100206 27383 100304 27481 4 vdd
rlabel metal3 s 99428 29335 99526 29433 4 vdd
rlabel metal3 s 100638 28173 100736 28271 4 vdd
rlabel metal3 s 100638 30111 100736 30209 4 vdd
rlabel metal3 s 99428 27360 99526 27458 4 vdd
rlabel metal3 s 99824 26570 99922 26668 4 gnd
rlabel metal3 s 101063 27009 101161 27107 4 gnd
rlabel metal3 s 100638 29753 100736 29851 4 vdd
rlabel metal3 s 100638 28531 100736 28629 4 vdd
rlabel metal3 s 99824 27755 99922 27853 4 gnd
rlabel metal3 s 99428 26570 99526 26668 4 vdd
rlabel metal3 s 101063 27799 101161 27897 4 gnd
rlabel metal3 s 101063 29753 101161 29851 4 gnd
rlabel metal3 s 99428 30125 99526 30223 4 vdd
rlabel metal3 s 101063 28589 101161 28687 4 gnd
rlabel metal3 s 100206 28531 100304 28629 4 vdd
rlabel metal3 s 100206 26161 100304 26259 4 vdd
rlabel metal3 s 101063 28963 101161 29061 4 gnd
rlabel metal3 s 99824 28940 99922 29038 4 gnd
rlabel metal3 s 99824 29335 99922 29433 4 gnd
rlabel metal3 s 100206 30111 100304 30209 4 vdd
rlabel metal3 s 99428 27755 99526 27853 4 vdd
rlabel metal3 s 100206 29321 100304 29419 4 vdd
rlabel metal3 s 100206 27741 100304 27839 4 vdd
rlabel metal3 s 99428 28150 99526 28248 4 vdd
rlabel metal3 s 101063 30169 101161 30267 4 gnd
rlabel metal3 s 101063 27383 101161 27481 4 gnd
rlabel metal3 s 99428 29730 99526 29828 4 vdd
rlabel metal3 s 100638 26161 100736 26259 4 vdd
rlabel metal3 s 99824 28545 99922 28643 4 gnd
rlabel metal3 s 99824 26175 99922 26273 4 gnd
rlabel metal3 s 99428 21830 99526 21928 4 vdd
rlabel metal3 s 99824 23015 99922 23113 4 gnd
rlabel metal3 s 100206 22643 100304 22741 4 vdd
rlabel metal3 s 99428 23805 99526 23903 4 vdd
rlabel metal3 s 101063 23433 101161 23531 4 gnd
rlabel metal3 s 100206 23791 100304 23889 4 vdd
rlabel metal3 s 100206 23001 100304 23099 4 vdd
rlabel metal3 s 99428 24990 99526 25088 4 vdd
rlabel metal3 s 101063 25429 101161 25527 4 gnd
rlabel metal3 s 100638 23791 100736 23889 4 vdd
rlabel metal3 s 100638 21853 100736 21951 4 vdd
rlabel metal3 s 100638 22211 100736 22309 4 vdd
rlabel metal3 s 101063 22269 101161 22367 4 gnd
rlabel metal3 s 100206 21853 100304 21951 4 vdd
rlabel metal3 s 99824 24200 99922 24298 4 gnd
rlabel metal3 s 100638 23001 100736 23099 4 vdd
rlabel metal3 s 99428 23015 99526 23113 4 vdd
rlabel metal3 s 99824 25385 99922 25483 4 gnd
rlabel metal3 s 100638 25803 100736 25901 4 vdd
rlabel metal3 s 99824 23805 99922 23903 4 gnd
rlabel metal3 s 99824 23410 99922 23508 4 gnd
rlabel metal3 s 100206 23433 100304 23531 4 vdd
rlabel metal3 s 100206 25013 100304 25111 4 vdd
rlabel metal3 s 100206 24581 100304 24679 4 vdd
rlabel metal3 s 99428 22225 99526 22323 4 vdd
rlabel metal3 s 100638 25371 100736 25469 4 vdd
rlabel metal3 s 101063 23059 101161 23157 4 gnd
rlabel metal3 s 101063 23849 101161 23947 4 gnd
rlabel metal3 s 99824 24595 99922 24693 4 gnd
rlabel metal3 s 99824 24990 99922 25088 4 gnd
rlabel metal3 s 101063 25013 101161 25111 4 gnd
rlabel metal3 s 101063 21853 101161 21951 4 gnd
rlabel metal3 s 99428 22620 99526 22718 4 vdd
rlabel metal3 s 100638 22643 100736 22741 4 vdd
rlabel metal3 s 99824 25780 99922 25878 4 gnd
rlabel metal3 s 100638 24223 100736 24321 4 vdd
rlabel metal3 s 99428 24200 99526 24298 4 vdd
rlabel metal3 s 100206 24223 100304 24321 4 vdd
rlabel metal3 s 99428 23410 99526 23508 4 vdd
rlabel metal3 s 99428 25385 99526 25483 4 vdd
rlabel metal3 s 99428 25780 99526 25878 4 vdd
rlabel metal3 s 99824 21830 99922 21928 4 gnd
rlabel metal3 s 101063 25803 101161 25901 4 gnd
rlabel metal3 s 100638 24581 100736 24679 4 vdd
rlabel metal3 s 99824 22620 99922 22718 4 gnd
rlabel metal3 s 100638 23433 100736 23531 4 vdd
rlabel metal3 s 101063 22643 101161 22741 4 gnd
rlabel metal3 s 100206 25803 100304 25901 4 vdd
rlabel metal3 s 100206 25371 100304 25469 4 vdd
rlabel metal3 s 100638 25013 100736 25111 4 vdd
rlabel metal3 s 100206 22211 100304 22309 4 vdd
rlabel metal3 s 99428 24595 99526 24693 4 vdd
rlabel metal3 s 101063 24223 101161 24321 4 gnd
rlabel metal3 s 99824 22225 99922 22323 4 gnd
rlabel metal3 s 101063 24639 101161 24737 4 gnd
rlabel metal3 s 94488 24595 94586 24693 4 gnd
rlabel metal3 s 94488 24042 94586 24140 4 gnd
rlabel metal3 s 94488 22225 94586 22323 4 gnd
rlabel metal3 s 94488 23252 94586 23350 4 gnd
rlabel metal3 s 94488 24832 94586 24930 4 gnd
rlabel metal3 s 94488 23568 94586 23666 4 gnd
rlabel metal3 s 94488 25148 94586 25246 4 gnd
rlabel metal3 s 94488 25622 94586 25720 4 gnd
rlabel metal3 s 94488 23805 94586 23903 4 gnd
rlabel metal3 s 94488 22778 94586 22876 4 gnd
rlabel metal3 s 94488 25385 94586 25483 4 gnd
rlabel metal3 s 94488 21672 94586 21770 4 gnd
rlabel metal3 s 94488 23015 94586 23113 4 gnd
rlabel metal3 s 94488 22462 94586 22560 4 gnd
rlabel metal3 s 94488 21988 94586 22086 4 gnd
rlabel metal3 s 94488 24358 94586 24456 4 gnd
rlabel metal3 s 94488 19065 94586 19163 4 gnd
rlabel metal3 s 94488 19855 94586 19953 4 gnd
rlabel metal3 s 94488 19302 94586 19400 4 gnd
rlabel metal3 s 94488 21198 94586 21296 4 gnd
rlabel metal3 s 94488 18275 94586 18373 4 gnd
rlabel metal3 s 94488 17722 94586 17820 4 gnd
rlabel metal3 s 94488 20882 94586 20980 4 gnd
rlabel metal3 s 94488 20092 94586 20190 4 gnd
rlabel metal3 s 94488 18038 94586 18136 4 gnd
rlabel metal3 s 94488 21435 94586 21533 4 gnd
rlabel metal3 s 94488 19618 94586 19716 4 gnd
rlabel metal3 s 94488 18828 94586 18926 4 gnd
rlabel metal3 s 94488 18512 94586 18610 4 gnd
rlabel metal3 s 94488 17485 94586 17583 4 gnd
rlabel metal3 s 94488 20408 94586 20506 4 gnd
rlabel metal3 s 94488 20645 94586 20743 4 gnd
rlabel metal3 s 99428 17880 99526 17978 4 vdd
rlabel metal3 s 103620 17903 103718 18001 4 vdd
rlabel metal3 s 100206 18261 100304 18359 4 vdd
rlabel metal3 s 100206 20631 100304 20729 4 vdd
rlabel metal3 s 100206 20273 100304 20371 4 vdd
rlabel metal3 s 99428 18670 99526 18768 4 vdd
rlabel metal3 s 99824 18670 99922 18768 4 gnd
rlabel metal3 s 100206 19483 100304 19581 4 vdd
rlabel metal3 s 99824 21040 99922 21138 4 gnd
rlabel metal3 s 99824 20645 99922 20743 4 gnd
rlabel metal3 s 99428 20250 99526 20348 4 vdd
rlabel metal3 s 100638 18261 100736 18359 4 vdd
rlabel metal3 s 101063 19899 101161 19997 4 gnd
rlabel metal3 s 99428 20645 99526 20743 4 vdd
rlabel metal3 s 100638 18693 100736 18791 4 vdd
rlabel metal3 s 100638 19483 100736 19581 4 vdd
rlabel metal3 s 100206 17903 100304 18001 4 vdd
rlabel metal3 s 100638 19841 100736 19939 4 vdd
rlabel metal3 s 101063 17903 101161 18001 4 gnd
rlabel metal3 s 99428 19855 99526 19953 4 vdd
rlabel metal3 s 100206 21063 100304 21161 4 vdd
rlabel metal3 s 99428 19460 99526 19558 4 vdd
rlabel metal3 s 101063 19483 101161 19581 4 gnd
rlabel metal3 s 100206 19051 100304 19149 4 vdd
rlabel metal3 s 100206 17471 100304 17569 4 vdd
rlabel metal3 s 104052 17903 104150 18001 4 vdd
rlabel metal3 s 100638 20631 100736 20729 4 vdd
rlabel metal3 s 99824 17880 99922 17978 4 gnd
rlabel metal3 s 102842 17880 102940 17978 4 vdd
rlabel metal3 s 99824 19065 99922 19163 4 gnd
rlabel metal3 s 100206 21421 100304 21519 4 vdd
rlabel metal3 s 100638 19051 100736 19149 4 vdd
rlabel metal3 s 100638 17903 100736 18001 4 vdd
rlabel metal3 s 99428 19065 99526 19163 4 vdd
rlabel metal3 s 100206 18693 100304 18791 4 vdd
rlabel metal3 s 99824 19460 99922 19558 4 gnd
rlabel metal3 s 104477 17903 104575 18001 4 gnd
rlabel metal3 s 100638 21421 100736 21519 4 vdd
rlabel metal3 s 101063 21063 101161 21161 4 gnd
rlabel metal3 s 99824 20250 99922 20348 4 gnd
rlabel metal3 s 99824 17485 99922 17583 4 gnd
rlabel metal3 s 99428 18275 99526 18373 4 vdd
rlabel metal3 s 101063 18693 101161 18791 4 gnd
rlabel metal3 s 100638 21063 100736 21161 4 vdd
rlabel metal3 s 99824 21435 99922 21533 4 gnd
rlabel metal3 s 100638 20273 100736 20371 4 vdd
rlabel metal3 s 100206 19841 100304 19939 4 vdd
rlabel metal3 s 101063 21479 101161 21577 4 gnd
rlabel metal3 s 101063 20689 101161 20787 4 gnd
rlabel metal3 s 101063 17529 101161 17627 4 gnd
rlabel metal3 s 99428 17485 99526 17583 4 vdd
rlabel metal3 s 101063 19109 101161 19207 4 gnd
rlabel metal3 s 103238 17880 103336 17978 4 gnd
rlabel metal3 s 101063 20273 101161 20371 4 gnd
rlabel metal3 s 99428 21435 99526 21533 4 vdd
rlabel metal3 s 100638 17471 100736 17569 4 vdd
rlabel metal3 s 99428 21040 99526 21138 4 vdd
rlabel metal3 s 101063 18319 101161 18417 4 gnd
rlabel metal3 s 99824 18275 99922 18373 4 gnd
rlabel metal3 s 99824 19855 99922 19953 4 gnd
rlabel metal3 s 70080 9814 70178 9912 4 vdd
rlabel metal3 s 67465 9223 67563 9321 4 vdd
rlabel metal3 s 73705 9223 73803 9321 4 vdd
rlabel metal3 s 67584 9814 67682 9912 4 vdd
rlabel metal3 s 74567 9223 74665 9321 4 vdd
rlabel metal3 s 72576 9814 72674 9912 4 vdd
rlabel metal3 s 69961 9223 70059 9321 4 vdd
rlabel metal3 s 74448 9814 74546 9912 4 vdd
rlabel metal3 s 68327 9223 68425 9321 4 vdd
rlabel metal3 s 72071 9223 72169 9321 4 vdd
rlabel metal3 s 71952 9814 72050 9912 4 vdd
rlabel metal3 s 77449 9223 77547 9321 4 vdd
rlabel metal3 s 75696 9814 75794 9912 4 vdd
rlabel metal3 s 66960 9814 67058 9912 4 vdd
rlabel metal3 s 79559 9223 79657 9321 4 vdd
rlabel metal3 s 76320 9814 76418 9912 4 vdd
rlabel metal3 s 76201 9223 76299 9321 4 vdd
rlabel metal3 s 73200 9814 73298 9912 4 vdd
rlabel metal3 s 78192 9814 78290 9912 4 vdd
rlabel metal3 s 78816 9814 78914 9912 4 vdd
rlabel metal3 s 69456 9814 69554 9912 4 vdd
rlabel metal3 s 78697 9223 78795 9321 4 vdd
rlabel metal3 s 70704 9814 70802 9912 4 vdd
rlabel metal3 s 67079 9223 67177 9321 4 vdd
rlabel metal3 s 78311 9223 78409 9321 4 vdd
rlabel metal3 s 70823 9223 70921 9321 4 vdd
rlabel metal3 s 75815 9223 75913 9321 4 vdd
rlabel metal3 s 68713 9223 68811 9321 4 vdd
rlabel metal3 s 77063 9223 77161 9321 4 vdd
rlabel metal3 s 73319 9223 73417 9321 4 vdd
rlabel metal3 s 73824 9814 73922 9912 4 vdd
rlabel metal3 s 79440 9814 79538 9912 4 vdd
rlabel metal3 s 72457 9223 72555 9321 4 vdd
rlabel metal3 s 74953 9223 75051 9321 4 vdd
rlabel metal3 s 77568 9814 77666 9912 4 vdd
rlabel metal3 s 71209 9223 71307 9321 4 vdd
rlabel metal3 s 75072 9814 75170 9912 4 vdd
rlabel metal3 s 71328 9814 71426 9912 4 vdd
rlabel metal3 s 69575 9223 69673 9321 4 vdd
rlabel metal3 s 76944 9814 77042 9912 4 vdd
rlabel metal3 s 68208 9814 68306 9912 4 vdd
rlabel metal3 s 68832 9814 68930 9912 4 vdd
rlabel metal3 s 62592 9814 62690 9912 4 vdd
rlabel metal3 s 58729 9223 58827 9321 4 vdd
rlabel metal3 s 66336 9814 66434 9912 4 vdd
rlabel metal3 s 65831 9223 65929 9321 4 vdd
rlabel metal3 s 56352 9814 56450 9912 4 vdd
rlabel metal3 s 64464 9814 64562 9912 4 vdd
rlabel metal3 s 55104 9814 55202 9912 4 vdd
rlabel metal3 s 58343 9223 58441 9321 4 vdd
rlabel metal3 s 53737 9223 53835 9321 4 vdd
rlabel metal3 s 60096 9814 60194 9912 4 vdd
rlabel metal3 s 61968 9814 62066 9912 4 vdd
rlabel metal3 s 60839 9223 60937 9321 4 vdd
rlabel metal3 s 61225 9223 61323 9321 4 vdd
rlabel metal3 s 53856 9814 53954 9912 4 vdd
rlabel metal3 s 64969 9223 65067 9321 4 vdd
rlabel metal3 s 58224 9814 58322 9912 4 vdd
rlabel metal3 s 57481 9223 57579 9321 4 vdd
rlabel metal3 s 59591 9223 59689 9321 4 vdd
rlabel metal3 s 57095 9223 57193 9321 4 vdd
rlabel metal3 s 60720 9814 60818 9912 4 vdd
rlabel metal3 s 54599 9223 54697 9321 4 vdd
rlabel metal3 s 63840 9814 63938 9912 4 vdd
rlabel metal3 s 63216 9814 63314 9912 4 vdd
rlabel metal3 s 65712 9814 65810 9912 4 vdd
rlabel metal3 s 62473 9223 62571 9321 4 vdd
rlabel metal3 s 54480 9814 54578 9912 4 vdd
rlabel metal3 s 59472 9814 59570 9912 4 vdd
rlabel metal3 s 59977 9223 60075 9321 4 vdd
rlabel metal3 s 64583 9223 64681 9321 4 vdd
rlabel metal3 s 56233 9223 56331 9321 4 vdd
rlabel metal3 s 61344 9814 61442 9912 4 vdd
rlabel metal3 s 57600 9814 57698 9912 4 vdd
rlabel metal3 s 62087 9223 62185 9321 4 vdd
rlabel metal3 s 65088 9814 65186 9912 4 vdd
rlabel metal3 s 55728 9814 55826 9912 4 vdd
rlabel metal3 s 63335 9223 63433 9321 4 vdd
rlabel metal3 s 56976 9814 57074 9912 4 vdd
rlabel metal3 s 54985 9223 55083 9321 4 vdd
rlabel metal3 s 66217 9223 66315 9321 4 vdd
rlabel metal3 s 58848 9814 58946 9912 4 vdd
rlabel metal3 s 55847 9223 55945 9321 4 vdd
rlabel metal3 s 63721 9223 63819 9321 4 vdd
rlabel metal3 s 63795 2950 63893 3048 4 gnd
rlabel metal3 s 58917 3743 59015 3841 4 gnd
rlabel metal3 s 55416 7674 55514 7772 4 gnd
rlabel metal3 s 56302 1979 56400 2077 4 gnd
rlabel metal3 s 53921 2181 54019 2279 4 gnd
rlabel metal3 s 57912 7674 58010 7772 4 gnd
rlabel metal3 s 63790 1979 63888 2077 4 gnd
rlabel metal3 s 61656 7674 61754 7772 4 gnd
rlabel metal3 s 65400 7674 65498 7772 4 gnd
rlabel metal3 s 56316 1563 56414 1661 4 vdd
rlabel metal3 s 63979 5677 64077 5775 4 gnd
rlabel metal3 s 66280 2513 66378 2611 4 vdd
rlabel metal3 s 62904 7674 63002 7772 4 gnd
rlabel metal3 s 58812 1563 58910 1661 4 vdd
rlabel metal3 s 56409 4903 56507 5001 4 vdd
rlabel metal3 s 53925 4065 54023 4163 4 vdd
rlabel metal3 s 53925 3743 54023 3841 4 gnd
rlabel metal3 s 61288 2513 61386 2611 4 vdd
rlabel metal3 s 66291 2950 66389 3048 4 gnd
rlabel metal3 s 60408 7674 60506 7772 4 gnd
rlabel metal3 s 61413 4065 61511 4163 4 vdd
rlabel metal3 s 58913 2181 59011 2279 4 gnd
rlabel metal3 s 66401 2181 66499 2279 4 gnd
rlabel metal3 s 54168 7674 54266 7772 4 gnd
rlabel metal3 s 66286 1979 66384 2077 4 gnd
rlabel metal3 s 63909 3743 64007 3841 4 gnd
rlabel metal3 s 56296 2513 56394 2611 4 vdd
rlabel metal3 s 56491 5677 56589 5775 4 gnd
rlabel metal3 s 61483 5677 61581 5775 4 gnd
rlabel metal3 s 63784 2513 63882 2611 4 vdd
rlabel metal3 s 53820 1563 53918 1661 4 vdd
rlabel metal3 s 56664 7674 56762 7772 4 gnd
rlabel metal3 s 58792 2513 58890 2611 4 vdd
rlabel metal3 s 61409 2181 61507 2279 4 gnd
rlabel metal3 s 58798 1979 58896 2077 4 gnd
rlabel metal3 s 61308 1563 61406 1661 4 vdd
rlabel metal3 s 53995 5677 54093 5775 4 gnd
rlabel metal3 s 53806 1979 53904 2077 4 gnd
rlabel metal3 s 66475 5677 66573 5775 4 gnd
rlabel metal3 s 63909 4065 64007 4163 4 vdd
rlabel metal3 s 56417 2181 56515 2279 4 gnd
rlabel metal3 s 66300 1563 66398 1661 4 vdd
rlabel metal3 s 58803 2950 58901 3048 4 gnd
rlabel metal3 s 58905 4903 59003 5001 4 vdd
rlabel metal3 s 61413 3743 61511 3841 4 gnd
rlabel metal3 s 59160 7674 59258 7772 4 gnd
rlabel metal3 s 61294 1979 61392 2077 4 gnd
rlabel metal3 s 58987 5677 59085 5775 4 gnd
rlabel metal3 s 53913 4903 54011 5001 4 vdd
rlabel metal3 s 61299 2950 61397 3048 4 gnd
rlabel metal3 s 56421 3743 56519 3841 4 gnd
rlabel metal3 s 58917 4065 59015 4163 4 vdd
rlabel metal3 s 63804 1563 63902 1661 4 vdd
rlabel metal3 s 66405 3743 66503 3841 4 gnd
rlabel metal3 s 63905 2181 64003 2279 4 gnd
rlabel metal3 s 53800 2513 53898 2611 4 vdd
rlabel metal3 s 66393 4903 66491 5001 4 vdd
rlabel metal3 s 56307 2950 56405 3048 4 gnd
rlabel metal3 s 61401 4903 61499 5001 4 vdd
rlabel metal3 s 53811 2950 53909 3048 4 gnd
rlabel metal3 s 64152 7674 64250 7772 4 gnd
rlabel metal3 s 56421 4065 56519 4163 4 vdd
rlabel metal3 s 63897 4903 63995 5001 4 vdd
rlabel metal3 s 66405 4065 66503 4163 4 vdd
rlabel metal3 s 73779 2950 73877 3048 4 gnd
rlabel metal3 s 71397 4065 71495 4163 4 vdd
rlabel metal3 s 77880 7674 77978 7772 4 gnd
rlabel metal3 s 71385 4903 71483 5001 4 vdd
rlabel metal3 s 67896 7674 67994 7772 4 gnd
rlabel metal3 s 73788 1563 73886 1661 4 vdd
rlabel metal3 s 71397 3743 71495 3841 4 gnd
rlabel metal3 s 72888 7674 72986 7772 4 gnd
rlabel metal3 s 76377 4903 76475 5001 4 vdd
rlabel metal3 s 68782 1979 68880 2077 4 gnd
rlabel metal3 s 68901 4065 68999 4163 4 vdd
rlabel metal3 s 78771 2950 78869 3048 4 gnd
rlabel metal3 s 68889 4903 68987 5001 4 vdd
rlabel metal3 s 71292 1563 71390 1661 4 vdd
rlabel metal3 s 76270 1979 76368 2077 4 gnd
rlabel metal3 s 70392 7674 70490 7772 4 gnd
rlabel metal3 s 74136 7674 74234 7772 4 gnd
rlabel metal3 s 78780 1563 78878 1661 4 vdd
rlabel metal3 s 76389 4065 76487 4163 4 vdd
rlabel metal3 s 68971 5677 69069 5775 4 gnd
rlabel metal3 s 73889 2181 73987 2279 4 gnd
rlabel metal3 s 78955 5677 79053 5775 4 gnd
rlabel metal3 s 78885 4065 78983 4163 4 vdd
rlabel metal3 s 73768 2513 73866 2611 4 vdd
rlabel metal3 s 78873 4903 78971 5001 4 vdd
rlabel metal3 s 78885 3743 78983 3841 4 gnd
rlabel metal3 s 69144 7674 69242 7772 4 gnd
rlabel metal3 s 71467 5677 71565 5775 4 gnd
rlabel metal3 s 79128 7674 79226 7772 4 gnd
rlabel metal3 s 71272 2513 71370 2611 4 vdd
rlabel metal3 s 76389 3743 76487 3841 4 gnd
rlabel metal3 s 68796 1563 68894 1661 4 vdd
rlabel metal3 s 71393 2181 71491 2279 4 gnd
rlabel metal3 s 78881 2181 78979 2279 4 gnd
rlabel metal3 s 78760 2513 78858 2611 4 vdd
rlabel metal3 s 66648 7674 66746 7772 4 gnd
rlabel metal3 s 76275 2950 76373 3048 4 gnd
rlabel metal3 s 73774 1979 73872 2077 4 gnd
rlabel metal3 s 76284 1563 76382 1661 4 vdd
rlabel metal3 s 71640 7674 71738 7772 4 gnd
rlabel metal3 s 73881 4903 73979 5001 4 vdd
rlabel metal3 s 76264 2513 76362 2611 4 vdd
rlabel metal3 s 71278 1979 71376 2077 4 gnd
rlabel metal3 s 76385 2181 76483 2279 4 gnd
rlabel metal3 s 68897 2181 68995 2279 4 gnd
rlabel metal3 s 76632 7674 76730 7772 4 gnd
rlabel metal3 s 68776 2513 68874 2611 4 vdd
rlabel metal3 s 68787 2950 68885 3048 4 gnd
rlabel metal3 s 68901 3743 68999 3841 4 gnd
rlabel metal3 s 73893 4065 73991 4163 4 vdd
rlabel metal3 s 71283 2950 71381 3048 4 gnd
rlabel metal3 s 76459 5677 76557 5775 4 gnd
rlabel metal3 s 73893 3743 73991 3841 4 gnd
rlabel metal3 s 78766 1979 78864 2077 4 gnd
rlabel metal3 s 75384 7674 75482 7772 4 gnd
rlabel metal3 s 73963 5677 74061 5775 4 gnd
rlabel metal3 s 103620 15533 103718 15631 4 vdd
rlabel metal3 s 100638 13521 100736 13619 4 vdd
rlabel metal3 s 99824 14720 99922 14818 4 gnd
rlabel metal3 s 99428 15510 99526 15608 4 vdd
rlabel metal3 s 104940 13140 105038 13238 4 vdd
rlabel metal3 s 100206 15101 100304 15199 4 vdd
rlabel metal3 s 102842 16300 102940 16398 4 vdd
rlabel metal3 s 99428 16300 99526 16398 4 vdd
rlabel metal3 s 100206 15891 100304 15989 4 vdd
rlabel metal3 s 99428 14720 99526 14818 4 vdd
rlabel metal3 s 99824 17090 99922 17188 4 gnd
rlabel metal3 s 100206 14743 100304 14841 4 vdd
rlabel metal3 s 104052 16323 104150 16421 4 vdd
rlabel metal3 s 101063 17113 101161 17211 4 gnd
rlabel metal3 s 99824 13535 99922 13633 4 gnd
rlabel metal3 s 103238 16300 103336 16398 4 gnd
rlabel metal3 s 104042 13937 104140 14035 4 gnd
rlabel metal3 s 103238 13930 103336 14028 4 gnd
rlabel metal3 s 100206 13163 100304 13261 4 vdd
rlabel metal3 s 104477 17113 104575 17211 4 gnd
rlabel metal3 s 100206 13953 100304 14051 4 vdd
rlabel metal3 s 99824 13140 99922 13238 4 gnd
rlabel metal3 s 100638 13953 100736 14051 4 vdd
rlabel metal3 s 99428 17090 99526 17188 4 vdd
rlabel metal3 s 100206 16323 100304 16421 4 vdd
rlabel metal3 s 99428 13535 99526 13633 4 vdd
rlabel metal3 s 100638 14311 100736 14409 4 vdd
rlabel metal3 s 100206 14311 100304 14409 4 vdd
rlabel metal3 s 104477 16323 104575 16421 4 gnd
rlabel metal3 s 102842 13140 102940 13238 4 vdd
rlabel metal3 s 103617 13147 103715 13245 4 vdd
rlabel metal3 s 99824 16300 99922 16398 4 gnd
rlabel metal3 s 100206 17113 100304 17211 4 vdd
rlabel metal3 s 105536 15510 105634 15608 4 vdd
rlabel metal3 s 100638 16323 100736 16421 4 vdd
rlabel metal3 s 101063 14743 101161 14841 4 gnd
rlabel metal3 s 100638 16681 100736 16779 4 vdd
rlabel metal3 s 99428 15115 99526 15213 4 vdd
rlabel metal3 s 99824 13930 99922 14028 4 gnd
rlabel metal3 s 99824 16695 99922 16793 4 gnd
rlabel metal3 s 99428 13930 99526 14028 4 vdd
rlabel metal3 s 104052 17113 104150 17211 4 vdd
rlabel metal3 s 99824 15510 99922 15608 4 gnd
rlabel metal3 s 100638 15101 100736 15199 4 vdd
rlabel metal3 s 101063 13579 101161 13677 4 gnd
rlabel metal3 s 101063 15949 101161 16047 4 gnd
rlabel metal3 s 102842 17090 102940 17188 4 vdd
rlabel metal3 s 101063 14369 101161 14467 4 gnd
rlabel metal3 s 101063 16323 101161 16421 4 gnd
rlabel metal3 s 100206 13521 100304 13619 4 vdd
rlabel metal3 s 104052 15533 104150 15631 4 vdd
rlabel metal3 s 100638 13163 100736 13261 4 vdd
rlabel metal3 s 99824 15115 99922 15213 4 gnd
rlabel metal3 s 100638 15533 100736 15631 4 vdd
rlabel metal3 s 99428 13140 99526 13238 4 vdd
rlabel metal3 s 101063 13953 101161 14051 4 gnd
rlabel metal3 s 103617 13937 103715 14035 4 vdd
rlabel metal3 s 103238 15510 103336 15608 4 gnd
rlabel metal3 s 100638 15891 100736 15989 4 vdd
rlabel metal3 s 101063 15159 101161 15257 4 gnd
rlabel metal3 s 100206 16681 100304 16779 4 vdd
rlabel metal3 s 104042 13147 104140 13245 4 gnd
rlabel metal3 s 101063 15533 101161 15631 4 gnd
rlabel metal3 s 100638 14743 100736 14841 4 vdd
rlabel metal3 s 99428 14325 99526 14423 4 vdd
rlabel metal3 s 100206 15533 100304 15631 4 vdd
rlabel metal3 s 100638 17113 100736 17211 4 vdd
rlabel metal3 s 99428 16695 99526 16793 4 vdd
rlabel metal3 s 103620 16323 103718 16421 4 vdd
rlabel metal3 s 104477 15533 104575 15631 4 gnd
rlabel metal3 s 101063 13163 101161 13261 4 gnd
rlabel metal3 s 102842 13930 102940 14028 4 vdd
rlabel metal3 s 99428 15905 99526 16003 4 vdd
rlabel metal3 s 103238 17090 103336 17188 4 gnd
rlabel metal3 s 102842 15510 102940 15608 4 vdd
rlabel metal3 s 99824 15905 99922 16003 4 gnd
rlabel metal3 s 103620 17113 103718 17211 4 vdd
rlabel metal3 s 103238 13140 103336 13238 4 gnd
rlabel metal3 s 105336 13140 105434 13238 4 gnd
rlabel metal3 s 105932 15510 106030 15608 4 gnd
rlabel metal3 s 99824 14325 99922 14423 4 gnd
rlabel metal3 s 101063 16739 101161 16837 4 gnd
rlabel metal3 s 94488 15352 94586 15450 4 gnd
rlabel metal3 s 94488 16695 94586 16793 4 gnd
rlabel metal3 s 94488 16458 94586 16556 4 gnd
rlabel metal3 s 94488 16142 94586 16240 4 gnd
rlabel metal3 s 94488 15115 94586 15213 4 gnd
rlabel metal3 s 94488 14562 94586 14660 4 gnd
rlabel metal3 s 94488 14325 94586 14423 4 gnd
rlabel metal3 s 94488 14878 94586 14976 4 gnd
rlabel metal3 s 94488 13535 94586 13633 4 gnd
rlabel metal3 s 94488 15905 94586 16003 4 gnd
rlabel metal3 s 94488 14088 94586 14186 4 gnd
rlabel metal3 s 94488 15668 94586 15766 4 gnd
rlabel metal3 s 94488 12982 94586 13080 4 gnd
rlabel metal3 s 94488 13772 94586 13870 4 gnd
rlabel metal3 s 94488 13298 94586 13396 4 gnd
rlabel metal3 s 94488 16932 94586 17030 4 gnd
rlabel metal3 s 94488 17248 94586 17346 4 gnd
rlabel metal3 s 93287 9223 93385 9321 4 vdd
rlabel metal3 s 94488 10928 94586 11026 4 gnd
rlabel metal3 s 94488 12508 94586 12606 4 gnd
rlabel metal3 s 94488 10375 94586 10473 4 gnd
rlabel metal3 s 94488 11165 94586 11263 4 gnd
rlabel metal3 s 94488 11402 94586 11500 4 gnd
rlabel metal3 s 94488 11718 94586 11816 4 gnd
rlabel metal3 s 94488 12192 94586 12290 4 gnd
rlabel metal3 s 94488 10612 94586 10710 4 gnd
rlabel metal3 s 94488 11955 94586 12053 4 gnd
rlabel metal3 s 93168 9814 93266 9912 4 vdd
rlabel metal3 s 93792 9814 93890 9912 4 vdd
rlabel metal3 s 94488 12745 94586 12843 4 gnd
rlabel metal3 s 94854 10248 94952 10346 4 gnd
rlabel metal3 s 99824 10770 99922 10868 4 gnd
rlabel metal3 s 99824 12350 99922 12448 4 gnd
rlabel metal3 s 101063 10793 101161 10891 4 gnd
rlabel metal3 s 99824 11560 99922 11658 4 gnd
rlabel metal3 s 99824 12745 99922 12843 4 gnd
rlabel metal3 s 100206 10793 100304 10891 4 vdd
rlabel metal3 s 101063 11999 101161 12097 4 gnd
rlabel metal3 s 99428 12350 99526 12448 4 vdd
rlabel metal3 s 100638 12731 100736 12829 4 vdd
rlabel metal3 s 103617 11567 103715 11665 4 vdd
rlabel metal3 s 100638 11583 100736 11681 4 vdd
rlabel metal3 s 100638 11941 100736 12039 4 vdd
rlabel metal3 s 99428 11165 99526 11263 4 vdd
rlabel metal3 s 101063 12373 101161 12471 4 gnd
rlabel metal3 s 103238 10770 103336 10868 4 gnd
rlabel metal3 s 100206 12731 100304 12829 4 vdd
rlabel metal3 s 104042 11567 104140 11665 4 gnd
rlabel metal3 s 102842 10770 102940 10868 4 vdd
rlabel metal3 s 100206 11941 100304 12039 4 vdd
rlabel metal3 s 99824 11165 99922 11263 4 gnd
rlabel metal3 s 101063 12789 101161 12887 4 gnd
rlabel metal3 s 99428 11955 99526 12053 4 vdd
rlabel metal3 s 100638 11151 100736 11249 4 vdd
rlabel metal3 s 105336 10770 105434 10868 4 gnd
rlabel metal3 s 101063 11583 101161 11681 4 gnd
rlabel metal3 s 100206 11151 100304 11249 4 vdd
rlabel metal3 s 101063 11209 101161 11307 4 gnd
rlabel metal3 s 100638 12373 100736 12471 4 vdd
rlabel metal3 s 102842 11560 102940 11658 4 vdd
rlabel metal3 s 100206 11583 100304 11681 4 vdd
rlabel metal3 s 104940 10770 105038 10868 4 vdd
rlabel metal3 s 99428 10770 99526 10868 4 vdd
rlabel metal3 s 99428 12745 99526 12843 4 vdd
rlabel metal3 s 99428 11560 99526 11658 4 vdd
rlabel metal3 s 103238 11560 103336 11658 4 gnd
rlabel metal3 s 104042 10777 104140 10875 4 gnd
rlabel metal3 s 100206 12373 100304 12471 4 vdd
rlabel metal3 s 100638 10793 100736 10891 4 vdd
rlabel metal3 s 99824 11955 99922 12053 4 gnd
rlabel metal3 s 103617 10777 103715 10875 4 vdd
rlabel metal3 s 88681 9223 88779 9321 4 vdd
rlabel metal3 s 91920 9814 92018 9912 4 vdd
rlabel metal3 s 81936 9814 82034 9912 4 vdd
rlabel metal3 s 80064 9814 80162 9912 4 vdd
rlabel metal3 s 88295 9223 88393 9321 4 vdd
rlabel metal3 s 87433 9223 87531 9321 4 vdd
rlabel metal3 s 79945 9223 80043 9321 4 vdd
rlabel metal3 s 90791 9223 90889 9321 4 vdd
rlabel metal3 s 84551 9223 84649 9321 4 vdd
rlabel metal3 s 86304 9814 86402 9912 4 vdd
rlabel metal3 s 90672 9814 90770 9912 4 vdd
rlabel metal3 s 91296 9814 91394 9912 4 vdd
rlabel metal3 s 83303 9223 83401 9321 4 vdd
rlabel metal3 s 88800 9814 88898 9912 4 vdd
rlabel metal3 s 84432 9814 84530 9912 4 vdd
rlabel metal3 s 81312 9814 81410 9912 4 vdd
rlabel metal3 s 86185 9223 86283 9321 4 vdd
rlabel metal3 s 80688 9814 80786 9912 4 vdd
rlabel metal3 s 91177 9223 91275 9321 4 vdd
rlabel metal3 s 83689 9223 83787 9321 4 vdd
rlabel metal3 s 86928 9814 87026 9912 4 vdd
rlabel metal3 s 92425 9223 92523 9321 4 vdd
rlabel metal3 s 82560 9814 82658 9912 4 vdd
rlabel metal3 s 87047 9223 87145 9321 4 vdd
rlabel metal3 s 83184 9814 83282 9912 4 vdd
rlabel metal3 s 88176 9814 88274 9912 4 vdd
rlabel metal3 s 83808 9814 83906 9912 4 vdd
rlabel metal3 s 85056 9814 85154 9912 4 vdd
rlabel metal3 s 92039 9223 92137 9321 4 vdd
rlabel metal3 s 92544 9814 92642 9912 4 vdd
rlabel metal3 s 89543 9223 89641 9321 4 vdd
rlabel metal3 s 89424 9814 89522 9912 4 vdd
rlabel metal3 s 85799 9223 85897 9321 4 vdd
rlabel metal3 s 82441 9223 82539 9321 4 vdd
rlabel metal3 s 90048 9814 90146 9912 4 vdd
rlabel metal3 s 81193 9223 81291 9321 4 vdd
rlabel metal3 s 85680 9814 85778 9912 4 vdd
rlabel metal3 s 89929 9223 90027 9321 4 vdd
rlabel metal3 s 84937 9223 85035 9321 4 vdd
rlabel metal3 s 87552 9814 87650 9912 4 vdd
rlabel metal3 s 80807 9223 80905 9321 4 vdd
rlabel metal3 s 82055 9223 82153 9321 4 vdd
rlabel metal3 s 91365 3743 91463 3841 4 gnd
rlabel metal3 s 83865 4903 83963 5001 4 vdd
rlabel metal3 s 91435 5677 91533 5775 4 gnd
rlabel metal3 s 91365 4065 91463 4163 4 vdd
rlabel metal3 s 83758 1979 83856 2077 4 gnd
rlabel metal3 s 83752 2513 83850 2611 4 vdd
rlabel metal3 s 86373 3743 86471 3841 4 gnd
rlabel metal3 s 81377 2181 81475 2279 4 gnd
rlabel metal3 s 86248 2513 86346 2611 4 vdd
rlabel metal3 s 88764 1563 88862 1661 4 vdd
rlabel metal3 s 86373 4065 86471 4163 4 vdd
rlabel metal3 s 81262 1979 81360 2077 4 gnd
rlabel metal3 s 91251 2950 91349 3048 4 gnd
rlabel metal3 s 91353 4903 91451 5001 4 vdd
rlabel metal3 s 81276 1563 81374 1661 4 vdd
rlabel metal3 s 89112 7674 89210 7772 4 gnd
rlabel metal3 s 90360 7674 90458 7772 4 gnd
rlabel metal3 s 81256 2513 81354 2611 4 vdd
rlabel metal3 s 83877 4065 83975 4163 4 vdd
rlabel metal3 s 91246 1979 91344 2077 4 gnd
rlabel metal3 s 88744 2513 88842 2611 4 vdd
rlabel metal3 s 81267 2950 81365 3048 4 gnd
rlabel metal3 s 86616 7674 86714 7772 4 gnd
rlabel metal3 s 80376 7674 80474 7772 4 gnd
rlabel metal3 s 91608 7674 91706 7772 4 gnd
rlabel metal3 s 88755 2950 88853 3048 4 gnd
rlabel metal3 s 86443 5677 86541 5775 4 gnd
rlabel metal3 s 83877 3743 83975 3841 4 gnd
rlabel metal3 s 87864 7674 87962 7772 4 gnd
rlabel metal3 s 91240 2513 91338 2611 4 vdd
rlabel metal3 s 85368 7674 85466 7772 4 gnd
rlabel metal3 s 82872 7674 82970 7772 4 gnd
rlabel metal3 s 81381 3743 81479 3841 4 gnd
rlabel metal3 s 81369 4903 81467 5001 4 vdd
rlabel metal3 s 81624 7674 81722 7772 4 gnd
rlabel metal3 s 88869 3743 88967 3841 4 gnd
rlabel metal3 s 83772 1563 83870 1661 4 vdd
rlabel metal3 s 81451 5677 81549 5775 4 gnd
rlabel metal3 s 86361 4903 86459 5001 4 vdd
rlabel metal3 s 81381 4065 81479 4163 4 vdd
rlabel metal3 s 86268 1563 86366 1661 4 vdd
rlabel metal3 s 91361 2181 91459 2279 4 gnd
rlabel metal3 s 88939 5677 89037 5775 4 gnd
rlabel metal3 s 83873 2181 83971 2279 4 gnd
rlabel metal3 s 88865 2181 88963 2279 4 gnd
rlabel metal3 s 83763 2950 83861 3048 4 gnd
rlabel metal3 s 84120 7674 84218 7772 4 gnd
rlabel metal3 s 86259 2950 86357 3048 4 gnd
rlabel metal3 s 86254 1979 86352 2077 4 gnd
rlabel metal3 s 88857 4903 88955 5001 4 vdd
rlabel metal3 s 83947 5677 84045 5775 4 gnd
rlabel metal3 s 91260 1563 91358 1661 4 vdd
rlabel metal3 s 86369 2181 86467 2279 4 gnd
rlabel metal3 s 88869 4065 88967 4163 4 vdd
rlabel metal3 s 88750 1979 88848 2077 4 gnd
rlabel metal3 s 93480 0 93578 98 4 gnd
rlabel metal3 s 93480 1120 93578 1218 4 vdd
rlabel metal3 s 92856 7674 92954 7772 4 gnd
rlabel metal2 s 11663 49 11691 9634 4 p_en_bar0
rlabel metal2 s 11787 49 11815 9634 4 s_en0
rlabel metal2 s 11911 49 11939 9634 4 w_en0
rlabel metal2 s 7960 10111 7988 10139 4 wl_en0
rlabel metal2 s 95213 61774 95241 69282 4 s_en1
rlabel metal2 s 95337 61774 95365 69282 4 p_en_bar1
rlabel metal2 s 99198 61269 99226 61297 4 wl_en1
rlabel metal2 s 13643 305 13671 333 4 bank_wmask0_0
rlabel metal2 s 33611 305 33639 333 4 bank_wmask0_1
rlabel metal2 s 53579 305 53607 333 4 bank_wmask0_2
rlabel metal2 s 73547 305 73575 333 4 bank_wmask0_3
rlabel metal1 s 53697 67470 53743 67724 4 dout1_16
rlabel metal1 s 56193 67470 56239 67724 4 dout1_17
rlabel metal1 s 58689 67470 58735 67724 4 dout1_18
rlabel metal1 s 61185 67470 61231 67724 4 dout1_19
rlabel metal1 s 63681 67470 63727 67724 4 dout1_20
rlabel metal1 s 66177 67470 66223 67724 4 dout1_21
rlabel metal1 s 68673 67470 68719 67724 4 dout1_22
rlabel metal1 s 71169 67470 71215 67724 4 dout1_23
rlabel metal1 s 73665 67470 73711 67724 4 dout1_24
rlabel metal1 s 76161 67470 76207 67724 4 dout1_25
rlabel metal1 s 78657 67470 78703 67724 4 dout1_26
rlabel metal1 s 81153 67470 81199 67724 4 dout1_27
rlabel metal1 s 83649 67470 83695 67724 4 dout1_28
rlabel metal1 s 86145 67470 86191 67724 4 dout1_29
rlabel metal1 s 88641 67470 88687 67724 4 dout1_30
rlabel metal1 s 91137 67470 91183 67724 4 dout1_31
rlabel metal1 s 101898 68500 101944 68558 4 addr1_0
rlabel metal1 s 101774 67010 101820 67068 4 addr1_1
rlabel metal1 s 18753 67470 18799 67724 4 dout1_2
rlabel metal1 s 21249 67470 21295 67724 4 dout1_3
rlabel metal1 s 23745 67470 23791 67724 4 dout1_4
rlabel metal1 s 26241 67470 26287 67724 4 dout1_5
rlabel metal1 s 28737 67470 28783 67724 4 dout1_6
rlabel metal1 s 31233 67470 31279 67724 4 dout1_7
rlabel metal1 s 33729 67470 33775 67724 4 dout1_8
rlabel metal1 s 36225 67470 36271 67724 4 dout1_9
rlabel metal1 s 38721 67470 38767 67724 4 dout1_10
rlabel metal1 s 41217 67470 41263 67724 4 dout1_11
rlabel metal1 s 43713 67470 43759 67724 4 dout1_12
rlabel metal1 s 46209 67470 46255 67724 4 dout1_13
rlabel metal1 s 48705 67470 48751 67724 4 dout1_14
rlabel metal1 s 51201 67470 51247 67724 4 dout1_15
rlabel metal1 s 13761 67470 13807 67724 4 dout1_0
rlabel metal1 s 16257 67470 16303 67724 4 dout1_1
rlabel metal1 s 179 10424 207 18324 4 addr0_4
rlabel metal1 s 259 10424 287 18324 4 addr0_5
rlabel metal1 s 339 10424 367 18324 4 addr0_6
rlabel metal1 s 419 10424 447 18324 4 addr0_7
rlabel metal1 s 499 10424 527 18324 4 addr0_8
rlabel metal1 s 5118 2850 5164 2908 4 addr0_0
rlabel metal1 s 5242 4340 5288 4398 4 addr0_1
rlabel metal1 s 13912 1425 13972 1481 4 din0_0
rlabel metal1 s 16408 1425 16468 1481 4 din0_1
rlabel metal1 s 18904 1425 18964 1481 4 din0_2
rlabel metal1 s 21400 1425 21460 1481 4 din0_3
rlabel metal1 s 23896 1425 23956 1481 4 din0_4
rlabel metal1 s 26392 1425 26452 1481 4 din0_5
rlabel metal1 s 28888 1425 28948 1481 4 din0_6
rlabel metal1 s 31384 1425 31444 1481 4 din0_7
rlabel metal1 s 33880 1425 33940 1481 4 din0_8
rlabel metal1 s 36376 1425 36436 1481 4 din0_9
rlabel metal1 s 38872 1425 38932 1481 4 din0_10
rlabel metal1 s 41368 1425 41428 1481 4 din0_11
rlabel metal1 s 43864 1425 43924 1481 4 din0_12
rlabel metal1 s 46360 1425 46420 1481 4 din0_13
rlabel metal1 s 48856 1425 48916 1481 4 din0_14
rlabel metal1 s 51352 1425 51412 1481 4 din0_15
rlabel metal1 s 13761 3684 13807 3938 4 dout0_0
rlabel metal1 s 16257 3684 16303 3938 4 dout0_1
rlabel metal1 s 18753 3684 18799 3938 4 dout0_2
rlabel metal1 s 21249 3684 21295 3938 4 dout0_3
rlabel metal1 s 23745 3684 23791 3938 4 dout0_4
rlabel metal1 s 26241 3684 26287 3938 4 dout0_5
rlabel metal1 s 28737 3684 28783 3938 4 dout0_6
rlabel metal1 s 31233 3684 31279 3938 4 dout0_7
rlabel metal1 s 33729 3684 33775 3938 4 dout0_8
rlabel metal1 s 36225 3684 36271 3938 4 dout0_9
rlabel metal1 s 38721 3684 38767 3938 4 dout0_10
rlabel metal1 s 41217 3684 41263 3938 4 dout0_11
rlabel metal1 s 43713 3684 43759 3938 4 dout0_12
rlabel metal1 s 46209 3684 46255 3938 4 dout0_13
rlabel metal1 s 48705 3684 48751 3938 4 dout0_14
rlabel metal1 s 51201 3684 51247 3938 4 dout0_15
rlabel metal1 s 19 10424 47 18324 4 addr0_2
rlabel metal1 s 99 10424 127 18324 4 addr0_3
rlabel metal1 s 81304 1425 81364 1481 4 din0_27
rlabel metal1 s 83800 1425 83860 1481 4 din0_28
rlabel metal1 s 86296 1425 86356 1481 4 din0_29
rlabel metal1 s 88792 1425 88852 1481 4 din0_30
rlabel metal1 s 91288 1425 91348 1481 4 din0_31
rlabel metal1 s 53697 3684 53743 3938 4 dout0_16
rlabel metal1 s 56193 3684 56239 3938 4 dout0_17
rlabel metal1 s 58689 3684 58735 3938 4 dout0_18
rlabel metal1 s 61185 3684 61231 3938 4 dout0_19
rlabel metal1 s 63681 3684 63727 3938 4 dout0_20
rlabel metal1 s 66177 3684 66223 3938 4 dout0_21
rlabel metal1 s 68673 3684 68719 3938 4 dout0_22
rlabel metal1 s 71169 3684 71215 3938 4 dout0_23
rlabel metal1 s 73665 3684 73711 3938 4 dout0_24
rlabel metal1 s 76161 3684 76207 3938 4 dout0_25
rlabel metal1 s 78657 3684 78703 3938 4 dout0_26
rlabel metal1 s 81153 3684 81199 3938 4 dout0_27
rlabel metal1 s 83649 3684 83695 3938 4 dout0_28
rlabel metal1 s 86145 3684 86191 3938 4 dout0_29
rlabel metal1 s 88641 3684 88687 3938 4 dout0_30
rlabel metal1 s 91137 3684 91183 3938 4 dout0_31
rlabel metal1 s 53848 1425 53908 1481 4 din0_16
rlabel metal1 s 56344 1425 56404 1481 4 din0_17
rlabel metal1 s 58840 1425 58900 1481 4 din0_18
rlabel metal1 s 61336 1425 61396 1481 4 din0_19
rlabel metal1 s 63832 1425 63892 1481 4 din0_20
rlabel metal1 s 66328 1425 66388 1481 4 din0_21
rlabel metal1 s 68824 1425 68884 1481 4 din0_22
rlabel metal1 s 71320 1425 71380 1481 4 din0_23
rlabel metal1 s 73816 1425 73876 1481 4 din0_24
rlabel metal1 s 107139 10424 107167 18324 4 addr1_2
rlabel metal1 s 107059 10424 107087 18324 4 addr1_3
rlabel metal1 s 106979 10424 107007 18324 4 addr1_4
rlabel metal1 s 106899 10424 106927 18324 4 addr1_5
rlabel metal1 s 106819 10424 106847 18324 4 addr1_6
rlabel metal1 s 106739 10424 106767 18324 4 addr1_7
rlabel metal1 s 106659 10424 106687 18324 4 addr1_8
rlabel metal1 s 76312 1425 76372 1481 4 din0_25
rlabel metal1 s 78808 1425 78868 1481 4 din0_26
<< properties >>
string FIXED_BBOX 0 0 107270 69233
<< end >>
