magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -2410 -2360 2310 2360
<< metal3 >>
rect -1150 -1100 1050 1100
<< mimcap >>
rect -1050 952 950 1000
rect -1050 -952 -1002 952
rect 902 -952 950 952
rect -1050 -1000 950 -952
<< mimcapcontact >>
rect -1002 -952 902 952
<< metal4 >>
rect -1011 952 911 961
rect -1011 -952 -1002 952
rect 902 -952 911 952
rect -1011 -961 911 -952
<< properties >>
string FIXED_BBOX -1150 -1100 1050 1100
<< end >>
