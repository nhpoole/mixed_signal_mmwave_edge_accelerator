***** XSPICE digital controlled oscillator d_osc as vco *************** 
* 12.4 kHz to 117.9 kHz
* name: d_osc_vco
* aout analog out
* dout digital out 
* vctrl control voltage
* vdd supply voltage

.subckt d_osc_vco aout dout vctrl vdd=1.8

* Linear interpolation, input data from measured analog ring oscillator VCO.
a1 vctrl dout vco_clock
.model vco_clock d_osc(cntl_array = [0.7 0.75 0.8 0.85 0.9 0.95 1.0 1.05 1.1 1.15]
+ freq_array = [1.239e+004 1.999e+004 2.978e+004 4.085e+004 5.375e+004 6.742e+004 8.118e+004 9.464e+004 1.072e+005 1.179e+005]
+ duty_cycle = 0.5 init_phase = 180.0
+ rise_delay = 1e-7 fall_delay=1e-7)

*generate an analog output for plotting
abridge-fit [dout] [aout] dac1
.model dac1 dac_bridge(out_low=0 out_high='vdd' out_undef='vdd/2'
+ input_load=5.0e-12 t_rise=1e-7 t_fall=1e-7)

.ends d_osc_vco
