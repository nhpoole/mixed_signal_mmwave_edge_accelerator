magic
tech sky130A
magscale 1 2
timestamp 1623661481
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 30 -17 64 17
<< locali >>
rect 119 333 153 493
rect 287 333 321 493
rect 24 299 321 333
rect 24 161 68 299
rect 442 215 621 259
rect 667 215 806 265
rect 856 215 1015 265
rect 24 127 321 161
rect 119 51 153 127
rect 287 51 321 127
rect 1126 215 1356 325
rect 1406 259 1445 327
rect 1406 215 1542 259
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 19 383 85 527
rect 187 383 253 527
rect 355 383 421 527
rect 455 417 489 493
rect 523 451 589 527
rect 643 417 677 493
rect 711 451 777 527
rect 811 417 845 493
rect 879 451 945 527
rect 979 451 1545 485
rect 979 417 1013 451
rect 455 383 1013 417
rect 1227 415 1461 417
rect 1056 383 1461 415
rect 1056 381 1240 383
rect 1056 333 1090 381
rect 1495 351 1545 451
rect 360 299 1090 333
rect 360 265 394 299
rect 114 199 394 265
rect 19 17 85 93
rect 187 17 253 93
rect 455 131 777 165
rect 1056 161 1090 299
rect 355 17 421 93
rect 455 51 489 131
rect 879 127 1285 161
rect 1327 129 1529 163
rect 1327 93 1361 129
rect 523 17 589 93
rect 627 59 1029 93
rect 1134 59 1361 93
rect 1327 51 1361 59
rect 1395 17 1461 93
rect 1495 51 1529 129
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
rlabel locali s 856 215 1015 265 6 A1
port 1 nsew signal input
rlabel locali s 667 215 806 265 6 A2
port 2 nsew signal input
rlabel locali s 442 215 621 259 6 A3
port 3 nsew signal input
rlabel locali s 1126 215 1356 325 6 B1
port 4 nsew signal input
rlabel locali s 1406 259 1445 327 6 B2
port 5 nsew signal input
rlabel locali s 1406 215 1542 259 6 B2
port 5 nsew signal input
rlabel locali s 287 333 321 493 6 X
port 6 nsew signal output
rlabel locali s 287 51 321 127 6 X
port 6 nsew signal output
rlabel locali s 119 333 153 493 6 X
port 6 nsew signal output
rlabel locali s 119 51 153 127 6 X
port 6 nsew signal output
rlabel locali s 24 299 321 333 6 X
port 6 nsew signal output
rlabel locali s 24 161 68 299 6 X
port 6 nsew signal output
rlabel locali s 24 127 321 161 6 X
port 6 nsew signal output
rlabel metal1 s 0 -48 1564 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 17 8 VNB
port 8 nsew ground bidirectional
rlabel nwell s -38 261 1602 582 6 VPB
port 9 nsew power bidirectional
rlabel metal1 s 0 496 1564 592 6 VPWR
port 10 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1564 544
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
