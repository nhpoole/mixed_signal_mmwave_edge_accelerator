magic
tech sky130A
magscale 1 2
timestamp 1620703184
<< nmoslvt >>
rect -5570 1745 -4610 2345
rect -4552 1745 -3592 2345
rect -3534 1745 -2574 2345
rect -2516 1745 -1556 2345
rect -1498 1745 -538 2345
rect -480 1745 480 2345
rect 538 1745 1498 2345
rect 1556 1745 2516 2345
rect 2574 1745 3534 2345
rect 3592 1745 4552 2345
rect 4610 1745 5570 2345
rect -5570 927 -4610 1527
rect -4552 927 -3592 1527
rect -3534 927 -2574 1527
rect -2516 927 -1556 1527
rect -1498 927 -538 1527
rect -480 927 480 1527
rect 538 927 1498 1527
rect 1556 927 2516 1527
rect 2574 927 3534 1527
rect 3592 927 4552 1527
rect 4610 927 5570 1527
rect -5570 109 -4610 709
rect -4552 109 -3592 709
rect -3534 109 -2574 709
rect -2516 109 -1556 709
rect -1498 109 -538 709
rect -480 109 480 709
rect 538 109 1498 709
rect 1556 109 2516 709
rect 2574 109 3534 709
rect 3592 109 4552 709
rect 4610 109 5570 709
rect -5570 -709 -4610 -109
rect -4552 -709 -3592 -109
rect -3534 -709 -2574 -109
rect -2516 -709 -1556 -109
rect -1498 -709 -538 -109
rect -480 -709 480 -109
rect 538 -709 1498 -109
rect 1556 -709 2516 -109
rect 2574 -709 3534 -109
rect 3592 -709 4552 -109
rect 4610 -709 5570 -109
rect -5570 -1527 -4610 -927
rect -4552 -1527 -3592 -927
rect -3534 -1527 -2574 -927
rect -2516 -1527 -1556 -927
rect -1498 -1527 -538 -927
rect -480 -1527 480 -927
rect 538 -1527 1498 -927
rect 1556 -1527 2516 -927
rect 2574 -1527 3534 -927
rect 3592 -1527 4552 -927
rect 4610 -1527 5570 -927
rect -5570 -2345 -4610 -1745
rect -4552 -2345 -3592 -1745
rect -3534 -2345 -2574 -1745
rect -2516 -2345 -1556 -1745
rect -1498 -2345 -538 -1745
rect -480 -2345 480 -1745
rect 538 -2345 1498 -1745
rect 1556 -2345 2516 -1745
rect 2574 -2345 3534 -1745
rect 3592 -2345 4552 -1745
rect 4610 -2345 5570 -1745
<< ndiff >>
rect -5628 2333 -5570 2345
rect -5628 1757 -5616 2333
rect -5582 1757 -5570 2333
rect -5628 1745 -5570 1757
rect -4610 2333 -4552 2345
rect -4610 1757 -4598 2333
rect -4564 1757 -4552 2333
rect -4610 1745 -4552 1757
rect -3592 2333 -3534 2345
rect -3592 1757 -3580 2333
rect -3546 1757 -3534 2333
rect -3592 1745 -3534 1757
rect -2574 2333 -2516 2345
rect -2574 1757 -2562 2333
rect -2528 1757 -2516 2333
rect -2574 1745 -2516 1757
rect -1556 2333 -1498 2345
rect -1556 1757 -1544 2333
rect -1510 1757 -1498 2333
rect -1556 1745 -1498 1757
rect -538 2333 -480 2345
rect -538 1757 -526 2333
rect -492 1757 -480 2333
rect -538 1745 -480 1757
rect 480 2333 538 2345
rect 480 1757 492 2333
rect 526 1757 538 2333
rect 480 1745 538 1757
rect 1498 2333 1556 2345
rect 1498 1757 1510 2333
rect 1544 1757 1556 2333
rect 1498 1745 1556 1757
rect 2516 2333 2574 2345
rect 2516 1757 2528 2333
rect 2562 1757 2574 2333
rect 2516 1745 2574 1757
rect 3534 2333 3592 2345
rect 3534 1757 3546 2333
rect 3580 1757 3592 2333
rect 3534 1745 3592 1757
rect 4552 2333 4610 2345
rect 4552 1757 4564 2333
rect 4598 1757 4610 2333
rect 4552 1745 4610 1757
rect 5570 2333 5628 2345
rect 5570 1757 5582 2333
rect 5616 1757 5628 2333
rect 5570 1745 5628 1757
rect -5628 1515 -5570 1527
rect -5628 939 -5616 1515
rect -5582 939 -5570 1515
rect -5628 927 -5570 939
rect -4610 1515 -4552 1527
rect -4610 939 -4598 1515
rect -4564 939 -4552 1515
rect -4610 927 -4552 939
rect -3592 1515 -3534 1527
rect -3592 939 -3580 1515
rect -3546 939 -3534 1515
rect -3592 927 -3534 939
rect -2574 1515 -2516 1527
rect -2574 939 -2562 1515
rect -2528 939 -2516 1515
rect -2574 927 -2516 939
rect -1556 1515 -1498 1527
rect -1556 939 -1544 1515
rect -1510 939 -1498 1515
rect -1556 927 -1498 939
rect -538 1515 -480 1527
rect -538 939 -526 1515
rect -492 939 -480 1515
rect -538 927 -480 939
rect 480 1515 538 1527
rect 480 939 492 1515
rect 526 939 538 1515
rect 480 927 538 939
rect 1498 1515 1556 1527
rect 1498 939 1510 1515
rect 1544 939 1556 1515
rect 1498 927 1556 939
rect 2516 1515 2574 1527
rect 2516 939 2528 1515
rect 2562 939 2574 1515
rect 2516 927 2574 939
rect 3534 1515 3592 1527
rect 3534 939 3546 1515
rect 3580 939 3592 1515
rect 3534 927 3592 939
rect 4552 1515 4610 1527
rect 4552 939 4564 1515
rect 4598 939 4610 1515
rect 4552 927 4610 939
rect 5570 1515 5628 1527
rect 5570 939 5582 1515
rect 5616 939 5628 1515
rect 5570 927 5628 939
rect -5628 697 -5570 709
rect -5628 121 -5616 697
rect -5582 121 -5570 697
rect -5628 109 -5570 121
rect -4610 697 -4552 709
rect -4610 121 -4598 697
rect -4564 121 -4552 697
rect -4610 109 -4552 121
rect -3592 697 -3534 709
rect -3592 121 -3580 697
rect -3546 121 -3534 697
rect -3592 109 -3534 121
rect -2574 697 -2516 709
rect -2574 121 -2562 697
rect -2528 121 -2516 697
rect -2574 109 -2516 121
rect -1556 697 -1498 709
rect -1556 121 -1544 697
rect -1510 121 -1498 697
rect -1556 109 -1498 121
rect -538 697 -480 709
rect -538 121 -526 697
rect -492 121 -480 697
rect -538 109 -480 121
rect 480 697 538 709
rect 480 121 492 697
rect 526 121 538 697
rect 480 109 538 121
rect 1498 697 1556 709
rect 1498 121 1510 697
rect 1544 121 1556 697
rect 1498 109 1556 121
rect 2516 697 2574 709
rect 2516 121 2528 697
rect 2562 121 2574 697
rect 2516 109 2574 121
rect 3534 697 3592 709
rect 3534 121 3546 697
rect 3580 121 3592 697
rect 3534 109 3592 121
rect 4552 697 4610 709
rect 4552 121 4564 697
rect 4598 121 4610 697
rect 4552 109 4610 121
rect 5570 697 5628 709
rect 5570 121 5582 697
rect 5616 121 5628 697
rect 5570 109 5628 121
rect -5628 -121 -5570 -109
rect -5628 -697 -5616 -121
rect -5582 -697 -5570 -121
rect -5628 -709 -5570 -697
rect -4610 -121 -4552 -109
rect -4610 -697 -4598 -121
rect -4564 -697 -4552 -121
rect -4610 -709 -4552 -697
rect -3592 -121 -3534 -109
rect -3592 -697 -3580 -121
rect -3546 -697 -3534 -121
rect -3592 -709 -3534 -697
rect -2574 -121 -2516 -109
rect -2574 -697 -2562 -121
rect -2528 -697 -2516 -121
rect -2574 -709 -2516 -697
rect -1556 -121 -1498 -109
rect -1556 -697 -1544 -121
rect -1510 -697 -1498 -121
rect -1556 -709 -1498 -697
rect -538 -121 -480 -109
rect -538 -697 -526 -121
rect -492 -697 -480 -121
rect -538 -709 -480 -697
rect 480 -121 538 -109
rect 480 -697 492 -121
rect 526 -697 538 -121
rect 480 -709 538 -697
rect 1498 -121 1556 -109
rect 1498 -697 1510 -121
rect 1544 -697 1556 -121
rect 1498 -709 1556 -697
rect 2516 -121 2574 -109
rect 2516 -697 2528 -121
rect 2562 -697 2574 -121
rect 2516 -709 2574 -697
rect 3534 -121 3592 -109
rect 3534 -697 3546 -121
rect 3580 -697 3592 -121
rect 3534 -709 3592 -697
rect 4552 -121 4610 -109
rect 4552 -697 4564 -121
rect 4598 -697 4610 -121
rect 4552 -709 4610 -697
rect 5570 -121 5628 -109
rect 5570 -697 5582 -121
rect 5616 -697 5628 -121
rect 5570 -709 5628 -697
rect -5628 -939 -5570 -927
rect -5628 -1515 -5616 -939
rect -5582 -1515 -5570 -939
rect -5628 -1527 -5570 -1515
rect -4610 -939 -4552 -927
rect -4610 -1515 -4598 -939
rect -4564 -1515 -4552 -939
rect -4610 -1527 -4552 -1515
rect -3592 -939 -3534 -927
rect -3592 -1515 -3580 -939
rect -3546 -1515 -3534 -939
rect -3592 -1527 -3534 -1515
rect -2574 -939 -2516 -927
rect -2574 -1515 -2562 -939
rect -2528 -1515 -2516 -939
rect -2574 -1527 -2516 -1515
rect -1556 -939 -1498 -927
rect -1556 -1515 -1544 -939
rect -1510 -1515 -1498 -939
rect -1556 -1527 -1498 -1515
rect -538 -939 -480 -927
rect -538 -1515 -526 -939
rect -492 -1515 -480 -939
rect -538 -1527 -480 -1515
rect 480 -939 538 -927
rect 480 -1515 492 -939
rect 526 -1515 538 -939
rect 480 -1527 538 -1515
rect 1498 -939 1556 -927
rect 1498 -1515 1510 -939
rect 1544 -1515 1556 -939
rect 1498 -1527 1556 -1515
rect 2516 -939 2574 -927
rect 2516 -1515 2528 -939
rect 2562 -1515 2574 -939
rect 2516 -1527 2574 -1515
rect 3534 -939 3592 -927
rect 3534 -1515 3546 -939
rect 3580 -1515 3592 -939
rect 3534 -1527 3592 -1515
rect 4552 -939 4610 -927
rect 4552 -1515 4564 -939
rect 4598 -1515 4610 -939
rect 4552 -1527 4610 -1515
rect 5570 -939 5628 -927
rect 5570 -1515 5582 -939
rect 5616 -1515 5628 -939
rect 5570 -1527 5628 -1515
rect -5628 -1757 -5570 -1745
rect -5628 -2333 -5616 -1757
rect -5582 -2333 -5570 -1757
rect -5628 -2345 -5570 -2333
rect -4610 -1757 -4552 -1745
rect -4610 -2333 -4598 -1757
rect -4564 -2333 -4552 -1757
rect -4610 -2345 -4552 -2333
rect -3592 -1757 -3534 -1745
rect -3592 -2333 -3580 -1757
rect -3546 -2333 -3534 -1757
rect -3592 -2345 -3534 -2333
rect -2574 -1757 -2516 -1745
rect -2574 -2333 -2562 -1757
rect -2528 -2333 -2516 -1757
rect -2574 -2345 -2516 -2333
rect -1556 -1757 -1498 -1745
rect -1556 -2333 -1544 -1757
rect -1510 -2333 -1498 -1757
rect -1556 -2345 -1498 -2333
rect -538 -1757 -480 -1745
rect -538 -2333 -526 -1757
rect -492 -2333 -480 -1757
rect -538 -2345 -480 -2333
rect 480 -1757 538 -1745
rect 480 -2333 492 -1757
rect 526 -2333 538 -1757
rect 480 -2345 538 -2333
rect 1498 -1757 1556 -1745
rect 1498 -2333 1510 -1757
rect 1544 -2333 1556 -1757
rect 1498 -2345 1556 -2333
rect 2516 -1757 2574 -1745
rect 2516 -2333 2528 -1757
rect 2562 -2333 2574 -1757
rect 2516 -2345 2574 -2333
rect 3534 -1757 3592 -1745
rect 3534 -2333 3546 -1757
rect 3580 -2333 3592 -1757
rect 3534 -2345 3592 -2333
rect 4552 -1757 4610 -1745
rect 4552 -2333 4564 -1757
rect 4598 -2333 4610 -1757
rect 4552 -2345 4610 -2333
rect 5570 -1757 5628 -1745
rect 5570 -2333 5582 -1757
rect 5616 -2333 5628 -1757
rect 5570 -2345 5628 -2333
<< ndiffc >>
rect -5616 1757 -5582 2333
rect -4598 1757 -4564 2333
rect -3580 1757 -3546 2333
rect -2562 1757 -2528 2333
rect -1544 1757 -1510 2333
rect -526 1757 -492 2333
rect 492 1757 526 2333
rect 1510 1757 1544 2333
rect 2528 1757 2562 2333
rect 3546 1757 3580 2333
rect 4564 1757 4598 2333
rect 5582 1757 5616 2333
rect -5616 939 -5582 1515
rect -4598 939 -4564 1515
rect -3580 939 -3546 1515
rect -2562 939 -2528 1515
rect -1544 939 -1510 1515
rect -526 939 -492 1515
rect 492 939 526 1515
rect 1510 939 1544 1515
rect 2528 939 2562 1515
rect 3546 939 3580 1515
rect 4564 939 4598 1515
rect 5582 939 5616 1515
rect -5616 121 -5582 697
rect -4598 121 -4564 697
rect -3580 121 -3546 697
rect -2562 121 -2528 697
rect -1544 121 -1510 697
rect -526 121 -492 697
rect 492 121 526 697
rect 1510 121 1544 697
rect 2528 121 2562 697
rect 3546 121 3580 697
rect 4564 121 4598 697
rect 5582 121 5616 697
rect -5616 -697 -5582 -121
rect -4598 -697 -4564 -121
rect -3580 -697 -3546 -121
rect -2562 -697 -2528 -121
rect -1544 -697 -1510 -121
rect -526 -697 -492 -121
rect 492 -697 526 -121
rect 1510 -697 1544 -121
rect 2528 -697 2562 -121
rect 3546 -697 3580 -121
rect 4564 -697 4598 -121
rect 5582 -697 5616 -121
rect -5616 -1515 -5582 -939
rect -4598 -1515 -4564 -939
rect -3580 -1515 -3546 -939
rect -2562 -1515 -2528 -939
rect -1544 -1515 -1510 -939
rect -526 -1515 -492 -939
rect 492 -1515 526 -939
rect 1510 -1515 1544 -939
rect 2528 -1515 2562 -939
rect 3546 -1515 3580 -939
rect 4564 -1515 4598 -939
rect 5582 -1515 5616 -939
rect -5616 -2333 -5582 -1757
rect -4598 -2333 -4564 -1757
rect -3580 -2333 -3546 -1757
rect -2562 -2333 -2528 -1757
rect -1544 -2333 -1510 -1757
rect -526 -2333 -492 -1757
rect 492 -2333 526 -1757
rect 1510 -2333 1544 -1757
rect 2528 -2333 2562 -1757
rect 3546 -2333 3580 -1757
rect 4564 -2333 4598 -1757
rect 5582 -2333 5616 -1757
<< poly >>
rect -5384 2417 -4796 2433
rect -5384 2400 -5368 2417
rect -5570 2383 -5368 2400
rect -4812 2400 -4796 2417
rect -4366 2417 -3778 2433
rect -4366 2400 -4350 2417
rect -4812 2383 -4610 2400
rect -5570 2345 -4610 2383
rect -4552 2383 -4350 2400
rect -3794 2400 -3778 2417
rect -3348 2417 -2760 2433
rect -3348 2400 -3332 2417
rect -3794 2383 -3592 2400
rect -4552 2345 -3592 2383
rect -3534 2383 -3332 2400
rect -2776 2400 -2760 2417
rect -2330 2417 -1742 2433
rect -2330 2400 -2314 2417
rect -2776 2383 -2574 2400
rect -3534 2345 -2574 2383
rect -2516 2383 -2314 2400
rect -1758 2400 -1742 2417
rect -1312 2417 -724 2433
rect -1312 2400 -1296 2417
rect -1758 2383 -1556 2400
rect -2516 2345 -1556 2383
rect -1498 2383 -1296 2400
rect -740 2400 -724 2417
rect -294 2417 294 2433
rect -294 2400 -278 2417
rect -740 2383 -538 2400
rect -1498 2345 -538 2383
rect -480 2383 -278 2400
rect 278 2400 294 2417
rect 724 2417 1312 2433
rect 724 2400 740 2417
rect 278 2383 480 2400
rect -480 2345 480 2383
rect 538 2383 740 2400
rect 1296 2400 1312 2417
rect 1742 2417 2330 2433
rect 1742 2400 1758 2417
rect 1296 2383 1498 2400
rect 538 2345 1498 2383
rect 1556 2383 1758 2400
rect 2314 2400 2330 2417
rect 2760 2417 3348 2433
rect 2760 2400 2776 2417
rect 2314 2383 2516 2400
rect 1556 2345 2516 2383
rect 2574 2383 2776 2400
rect 3332 2400 3348 2417
rect 3778 2417 4366 2433
rect 3778 2400 3794 2417
rect 3332 2383 3534 2400
rect 2574 2345 3534 2383
rect 3592 2383 3794 2400
rect 4350 2400 4366 2417
rect 4796 2417 5384 2433
rect 4796 2400 4812 2417
rect 4350 2383 4552 2400
rect 3592 2345 4552 2383
rect 4610 2383 4812 2400
rect 5368 2400 5384 2417
rect 5368 2383 5570 2400
rect 4610 2345 5570 2383
rect -5570 1707 -4610 1745
rect -5570 1690 -5368 1707
rect -5384 1673 -5368 1690
rect -4812 1690 -4610 1707
rect -4552 1707 -3592 1745
rect -4552 1690 -4350 1707
rect -4812 1673 -4796 1690
rect -5384 1657 -4796 1673
rect -4366 1673 -4350 1690
rect -3794 1690 -3592 1707
rect -3534 1707 -2574 1745
rect -3534 1690 -3332 1707
rect -3794 1673 -3778 1690
rect -4366 1657 -3778 1673
rect -3348 1673 -3332 1690
rect -2776 1690 -2574 1707
rect -2516 1707 -1556 1745
rect -2516 1690 -2314 1707
rect -2776 1673 -2760 1690
rect -3348 1657 -2760 1673
rect -2330 1673 -2314 1690
rect -1758 1690 -1556 1707
rect -1498 1707 -538 1745
rect -1498 1690 -1296 1707
rect -1758 1673 -1742 1690
rect -2330 1657 -1742 1673
rect -1312 1673 -1296 1690
rect -740 1690 -538 1707
rect -480 1707 480 1745
rect -480 1690 -278 1707
rect -740 1673 -724 1690
rect -1312 1657 -724 1673
rect -294 1673 -278 1690
rect 278 1690 480 1707
rect 538 1707 1498 1745
rect 538 1690 740 1707
rect 278 1673 294 1690
rect -294 1657 294 1673
rect 724 1673 740 1690
rect 1296 1690 1498 1707
rect 1556 1707 2516 1745
rect 1556 1690 1758 1707
rect 1296 1673 1312 1690
rect 724 1657 1312 1673
rect 1742 1673 1758 1690
rect 2314 1690 2516 1707
rect 2574 1707 3534 1745
rect 2574 1690 2776 1707
rect 2314 1673 2330 1690
rect 1742 1657 2330 1673
rect 2760 1673 2776 1690
rect 3332 1690 3534 1707
rect 3592 1707 4552 1745
rect 3592 1690 3794 1707
rect 3332 1673 3348 1690
rect 2760 1657 3348 1673
rect 3778 1673 3794 1690
rect 4350 1690 4552 1707
rect 4610 1707 5570 1745
rect 4610 1690 4812 1707
rect 4350 1673 4366 1690
rect 3778 1657 4366 1673
rect 4796 1673 4812 1690
rect 5368 1690 5570 1707
rect 5368 1673 5384 1690
rect 4796 1657 5384 1673
rect -5384 1599 -4796 1615
rect -5384 1582 -5368 1599
rect -5570 1565 -5368 1582
rect -4812 1582 -4796 1599
rect -4366 1599 -3778 1615
rect -4366 1582 -4350 1599
rect -4812 1565 -4610 1582
rect -5570 1527 -4610 1565
rect -4552 1565 -4350 1582
rect -3794 1582 -3778 1599
rect -3348 1599 -2760 1615
rect -3348 1582 -3332 1599
rect -3794 1565 -3592 1582
rect -4552 1527 -3592 1565
rect -3534 1565 -3332 1582
rect -2776 1582 -2760 1599
rect -2330 1599 -1742 1615
rect -2330 1582 -2314 1599
rect -2776 1565 -2574 1582
rect -3534 1527 -2574 1565
rect -2516 1565 -2314 1582
rect -1758 1582 -1742 1599
rect -1312 1599 -724 1615
rect -1312 1582 -1296 1599
rect -1758 1565 -1556 1582
rect -2516 1527 -1556 1565
rect -1498 1565 -1296 1582
rect -740 1582 -724 1599
rect -294 1599 294 1615
rect -294 1582 -278 1599
rect -740 1565 -538 1582
rect -1498 1527 -538 1565
rect -480 1565 -278 1582
rect 278 1582 294 1599
rect 724 1599 1312 1615
rect 724 1582 740 1599
rect 278 1565 480 1582
rect -480 1527 480 1565
rect 538 1565 740 1582
rect 1296 1582 1312 1599
rect 1742 1599 2330 1615
rect 1742 1582 1758 1599
rect 1296 1565 1498 1582
rect 538 1527 1498 1565
rect 1556 1565 1758 1582
rect 2314 1582 2330 1599
rect 2760 1599 3348 1615
rect 2760 1582 2776 1599
rect 2314 1565 2516 1582
rect 1556 1527 2516 1565
rect 2574 1565 2776 1582
rect 3332 1582 3348 1599
rect 3778 1599 4366 1615
rect 3778 1582 3794 1599
rect 3332 1565 3534 1582
rect 2574 1527 3534 1565
rect 3592 1565 3794 1582
rect 4350 1582 4366 1599
rect 4796 1599 5384 1615
rect 4796 1582 4812 1599
rect 4350 1565 4552 1582
rect 3592 1527 4552 1565
rect 4610 1565 4812 1582
rect 5368 1582 5384 1599
rect 5368 1565 5570 1582
rect 4610 1527 5570 1565
rect -5570 889 -4610 927
rect -5570 872 -5368 889
rect -5384 855 -5368 872
rect -4812 872 -4610 889
rect -4552 889 -3592 927
rect -4552 872 -4350 889
rect -4812 855 -4796 872
rect -5384 839 -4796 855
rect -4366 855 -4350 872
rect -3794 872 -3592 889
rect -3534 889 -2574 927
rect -3534 872 -3332 889
rect -3794 855 -3778 872
rect -4366 839 -3778 855
rect -3348 855 -3332 872
rect -2776 872 -2574 889
rect -2516 889 -1556 927
rect -2516 872 -2314 889
rect -2776 855 -2760 872
rect -3348 839 -2760 855
rect -2330 855 -2314 872
rect -1758 872 -1556 889
rect -1498 889 -538 927
rect -1498 872 -1296 889
rect -1758 855 -1742 872
rect -2330 839 -1742 855
rect -1312 855 -1296 872
rect -740 872 -538 889
rect -480 889 480 927
rect -480 872 -278 889
rect -740 855 -724 872
rect -1312 839 -724 855
rect -294 855 -278 872
rect 278 872 480 889
rect 538 889 1498 927
rect 538 872 740 889
rect 278 855 294 872
rect -294 839 294 855
rect 724 855 740 872
rect 1296 872 1498 889
rect 1556 889 2516 927
rect 1556 872 1758 889
rect 1296 855 1312 872
rect 724 839 1312 855
rect 1742 855 1758 872
rect 2314 872 2516 889
rect 2574 889 3534 927
rect 2574 872 2776 889
rect 2314 855 2330 872
rect 1742 839 2330 855
rect 2760 855 2776 872
rect 3332 872 3534 889
rect 3592 889 4552 927
rect 3592 872 3794 889
rect 3332 855 3348 872
rect 2760 839 3348 855
rect 3778 855 3794 872
rect 4350 872 4552 889
rect 4610 889 5570 927
rect 4610 872 4812 889
rect 4350 855 4366 872
rect 3778 839 4366 855
rect 4796 855 4812 872
rect 5368 872 5570 889
rect 5368 855 5384 872
rect 4796 839 5384 855
rect -5384 781 -4796 797
rect -5384 764 -5368 781
rect -5570 747 -5368 764
rect -4812 764 -4796 781
rect -4366 781 -3778 797
rect -4366 764 -4350 781
rect -4812 747 -4610 764
rect -5570 709 -4610 747
rect -4552 747 -4350 764
rect -3794 764 -3778 781
rect -3348 781 -2760 797
rect -3348 764 -3332 781
rect -3794 747 -3592 764
rect -4552 709 -3592 747
rect -3534 747 -3332 764
rect -2776 764 -2760 781
rect -2330 781 -1742 797
rect -2330 764 -2314 781
rect -2776 747 -2574 764
rect -3534 709 -2574 747
rect -2516 747 -2314 764
rect -1758 764 -1742 781
rect -1312 781 -724 797
rect -1312 764 -1296 781
rect -1758 747 -1556 764
rect -2516 709 -1556 747
rect -1498 747 -1296 764
rect -740 764 -724 781
rect -294 781 294 797
rect -294 764 -278 781
rect -740 747 -538 764
rect -1498 709 -538 747
rect -480 747 -278 764
rect 278 764 294 781
rect 724 781 1312 797
rect 724 764 740 781
rect 278 747 480 764
rect -480 709 480 747
rect 538 747 740 764
rect 1296 764 1312 781
rect 1742 781 2330 797
rect 1742 764 1758 781
rect 1296 747 1498 764
rect 538 709 1498 747
rect 1556 747 1758 764
rect 2314 764 2330 781
rect 2760 781 3348 797
rect 2760 764 2776 781
rect 2314 747 2516 764
rect 1556 709 2516 747
rect 2574 747 2776 764
rect 3332 764 3348 781
rect 3778 781 4366 797
rect 3778 764 3794 781
rect 3332 747 3534 764
rect 2574 709 3534 747
rect 3592 747 3794 764
rect 4350 764 4366 781
rect 4796 781 5384 797
rect 4796 764 4812 781
rect 4350 747 4552 764
rect 3592 709 4552 747
rect 4610 747 4812 764
rect 5368 764 5384 781
rect 5368 747 5570 764
rect 4610 709 5570 747
rect -5570 71 -4610 109
rect -5570 54 -5368 71
rect -5384 37 -5368 54
rect -4812 54 -4610 71
rect -4552 71 -3592 109
rect -4552 54 -4350 71
rect -4812 37 -4796 54
rect -5384 21 -4796 37
rect -4366 37 -4350 54
rect -3794 54 -3592 71
rect -3534 71 -2574 109
rect -3534 54 -3332 71
rect -3794 37 -3778 54
rect -4366 21 -3778 37
rect -3348 37 -3332 54
rect -2776 54 -2574 71
rect -2516 71 -1556 109
rect -2516 54 -2314 71
rect -2776 37 -2760 54
rect -3348 21 -2760 37
rect -2330 37 -2314 54
rect -1758 54 -1556 71
rect -1498 71 -538 109
rect -1498 54 -1296 71
rect -1758 37 -1742 54
rect -2330 21 -1742 37
rect -1312 37 -1296 54
rect -740 54 -538 71
rect -480 71 480 109
rect -480 54 -278 71
rect -740 37 -724 54
rect -1312 21 -724 37
rect -294 37 -278 54
rect 278 54 480 71
rect 538 71 1498 109
rect 538 54 740 71
rect 278 37 294 54
rect -294 21 294 37
rect 724 37 740 54
rect 1296 54 1498 71
rect 1556 71 2516 109
rect 1556 54 1758 71
rect 1296 37 1312 54
rect 724 21 1312 37
rect 1742 37 1758 54
rect 2314 54 2516 71
rect 2574 71 3534 109
rect 2574 54 2776 71
rect 2314 37 2330 54
rect 1742 21 2330 37
rect 2760 37 2776 54
rect 3332 54 3534 71
rect 3592 71 4552 109
rect 3592 54 3794 71
rect 3332 37 3348 54
rect 2760 21 3348 37
rect 3778 37 3794 54
rect 4350 54 4552 71
rect 4610 71 5570 109
rect 4610 54 4812 71
rect 4350 37 4366 54
rect 3778 21 4366 37
rect 4796 37 4812 54
rect 5368 54 5570 71
rect 5368 37 5384 54
rect 4796 21 5384 37
rect -5384 -37 -4796 -21
rect -5384 -54 -5368 -37
rect -5570 -71 -5368 -54
rect -4812 -54 -4796 -37
rect -4366 -37 -3778 -21
rect -4366 -54 -4350 -37
rect -4812 -71 -4610 -54
rect -5570 -109 -4610 -71
rect -4552 -71 -4350 -54
rect -3794 -54 -3778 -37
rect -3348 -37 -2760 -21
rect -3348 -54 -3332 -37
rect -3794 -71 -3592 -54
rect -4552 -109 -3592 -71
rect -3534 -71 -3332 -54
rect -2776 -54 -2760 -37
rect -2330 -37 -1742 -21
rect -2330 -54 -2314 -37
rect -2776 -71 -2574 -54
rect -3534 -109 -2574 -71
rect -2516 -71 -2314 -54
rect -1758 -54 -1742 -37
rect -1312 -37 -724 -21
rect -1312 -54 -1296 -37
rect -1758 -71 -1556 -54
rect -2516 -109 -1556 -71
rect -1498 -71 -1296 -54
rect -740 -54 -724 -37
rect -294 -37 294 -21
rect -294 -54 -278 -37
rect -740 -71 -538 -54
rect -1498 -109 -538 -71
rect -480 -71 -278 -54
rect 278 -54 294 -37
rect 724 -37 1312 -21
rect 724 -54 740 -37
rect 278 -71 480 -54
rect -480 -109 480 -71
rect 538 -71 740 -54
rect 1296 -54 1312 -37
rect 1742 -37 2330 -21
rect 1742 -54 1758 -37
rect 1296 -71 1498 -54
rect 538 -109 1498 -71
rect 1556 -71 1758 -54
rect 2314 -54 2330 -37
rect 2760 -37 3348 -21
rect 2760 -54 2776 -37
rect 2314 -71 2516 -54
rect 1556 -109 2516 -71
rect 2574 -71 2776 -54
rect 3332 -54 3348 -37
rect 3778 -37 4366 -21
rect 3778 -54 3794 -37
rect 3332 -71 3534 -54
rect 2574 -109 3534 -71
rect 3592 -71 3794 -54
rect 4350 -54 4366 -37
rect 4796 -37 5384 -21
rect 4796 -54 4812 -37
rect 4350 -71 4552 -54
rect 3592 -109 4552 -71
rect 4610 -71 4812 -54
rect 5368 -54 5384 -37
rect 5368 -71 5570 -54
rect 4610 -109 5570 -71
rect -5570 -747 -4610 -709
rect -5570 -764 -5368 -747
rect -5384 -781 -5368 -764
rect -4812 -764 -4610 -747
rect -4552 -747 -3592 -709
rect -4552 -764 -4350 -747
rect -4812 -781 -4796 -764
rect -5384 -797 -4796 -781
rect -4366 -781 -4350 -764
rect -3794 -764 -3592 -747
rect -3534 -747 -2574 -709
rect -3534 -764 -3332 -747
rect -3794 -781 -3778 -764
rect -4366 -797 -3778 -781
rect -3348 -781 -3332 -764
rect -2776 -764 -2574 -747
rect -2516 -747 -1556 -709
rect -2516 -764 -2314 -747
rect -2776 -781 -2760 -764
rect -3348 -797 -2760 -781
rect -2330 -781 -2314 -764
rect -1758 -764 -1556 -747
rect -1498 -747 -538 -709
rect -1498 -764 -1296 -747
rect -1758 -781 -1742 -764
rect -2330 -797 -1742 -781
rect -1312 -781 -1296 -764
rect -740 -764 -538 -747
rect -480 -747 480 -709
rect -480 -764 -278 -747
rect -740 -781 -724 -764
rect -1312 -797 -724 -781
rect -294 -781 -278 -764
rect 278 -764 480 -747
rect 538 -747 1498 -709
rect 538 -764 740 -747
rect 278 -781 294 -764
rect -294 -797 294 -781
rect 724 -781 740 -764
rect 1296 -764 1498 -747
rect 1556 -747 2516 -709
rect 1556 -764 1758 -747
rect 1296 -781 1312 -764
rect 724 -797 1312 -781
rect 1742 -781 1758 -764
rect 2314 -764 2516 -747
rect 2574 -747 3534 -709
rect 2574 -764 2776 -747
rect 2314 -781 2330 -764
rect 1742 -797 2330 -781
rect 2760 -781 2776 -764
rect 3332 -764 3534 -747
rect 3592 -747 4552 -709
rect 3592 -764 3794 -747
rect 3332 -781 3348 -764
rect 2760 -797 3348 -781
rect 3778 -781 3794 -764
rect 4350 -764 4552 -747
rect 4610 -747 5570 -709
rect 4610 -764 4812 -747
rect 4350 -781 4366 -764
rect 3778 -797 4366 -781
rect 4796 -781 4812 -764
rect 5368 -764 5570 -747
rect 5368 -781 5384 -764
rect 4796 -797 5384 -781
rect -5384 -855 -4796 -839
rect -5384 -872 -5368 -855
rect -5570 -889 -5368 -872
rect -4812 -872 -4796 -855
rect -4366 -855 -3778 -839
rect -4366 -872 -4350 -855
rect -4812 -889 -4610 -872
rect -5570 -927 -4610 -889
rect -4552 -889 -4350 -872
rect -3794 -872 -3778 -855
rect -3348 -855 -2760 -839
rect -3348 -872 -3332 -855
rect -3794 -889 -3592 -872
rect -4552 -927 -3592 -889
rect -3534 -889 -3332 -872
rect -2776 -872 -2760 -855
rect -2330 -855 -1742 -839
rect -2330 -872 -2314 -855
rect -2776 -889 -2574 -872
rect -3534 -927 -2574 -889
rect -2516 -889 -2314 -872
rect -1758 -872 -1742 -855
rect -1312 -855 -724 -839
rect -1312 -872 -1296 -855
rect -1758 -889 -1556 -872
rect -2516 -927 -1556 -889
rect -1498 -889 -1296 -872
rect -740 -872 -724 -855
rect -294 -855 294 -839
rect -294 -872 -278 -855
rect -740 -889 -538 -872
rect -1498 -927 -538 -889
rect -480 -889 -278 -872
rect 278 -872 294 -855
rect 724 -855 1312 -839
rect 724 -872 740 -855
rect 278 -889 480 -872
rect -480 -927 480 -889
rect 538 -889 740 -872
rect 1296 -872 1312 -855
rect 1742 -855 2330 -839
rect 1742 -872 1758 -855
rect 1296 -889 1498 -872
rect 538 -927 1498 -889
rect 1556 -889 1758 -872
rect 2314 -872 2330 -855
rect 2760 -855 3348 -839
rect 2760 -872 2776 -855
rect 2314 -889 2516 -872
rect 1556 -927 2516 -889
rect 2574 -889 2776 -872
rect 3332 -872 3348 -855
rect 3778 -855 4366 -839
rect 3778 -872 3794 -855
rect 3332 -889 3534 -872
rect 2574 -927 3534 -889
rect 3592 -889 3794 -872
rect 4350 -872 4366 -855
rect 4796 -855 5384 -839
rect 4796 -872 4812 -855
rect 4350 -889 4552 -872
rect 3592 -927 4552 -889
rect 4610 -889 4812 -872
rect 5368 -872 5384 -855
rect 5368 -889 5570 -872
rect 4610 -927 5570 -889
rect -5570 -1565 -4610 -1527
rect -5570 -1582 -5368 -1565
rect -5384 -1599 -5368 -1582
rect -4812 -1582 -4610 -1565
rect -4552 -1565 -3592 -1527
rect -4552 -1582 -4350 -1565
rect -4812 -1599 -4796 -1582
rect -5384 -1615 -4796 -1599
rect -4366 -1599 -4350 -1582
rect -3794 -1582 -3592 -1565
rect -3534 -1565 -2574 -1527
rect -3534 -1582 -3332 -1565
rect -3794 -1599 -3778 -1582
rect -4366 -1615 -3778 -1599
rect -3348 -1599 -3332 -1582
rect -2776 -1582 -2574 -1565
rect -2516 -1565 -1556 -1527
rect -2516 -1582 -2314 -1565
rect -2776 -1599 -2760 -1582
rect -3348 -1615 -2760 -1599
rect -2330 -1599 -2314 -1582
rect -1758 -1582 -1556 -1565
rect -1498 -1565 -538 -1527
rect -1498 -1582 -1296 -1565
rect -1758 -1599 -1742 -1582
rect -2330 -1615 -1742 -1599
rect -1312 -1599 -1296 -1582
rect -740 -1582 -538 -1565
rect -480 -1565 480 -1527
rect -480 -1582 -278 -1565
rect -740 -1599 -724 -1582
rect -1312 -1615 -724 -1599
rect -294 -1599 -278 -1582
rect 278 -1582 480 -1565
rect 538 -1565 1498 -1527
rect 538 -1582 740 -1565
rect 278 -1599 294 -1582
rect -294 -1615 294 -1599
rect 724 -1599 740 -1582
rect 1296 -1582 1498 -1565
rect 1556 -1565 2516 -1527
rect 1556 -1582 1758 -1565
rect 1296 -1599 1312 -1582
rect 724 -1615 1312 -1599
rect 1742 -1599 1758 -1582
rect 2314 -1582 2516 -1565
rect 2574 -1565 3534 -1527
rect 2574 -1582 2776 -1565
rect 2314 -1599 2330 -1582
rect 1742 -1615 2330 -1599
rect 2760 -1599 2776 -1582
rect 3332 -1582 3534 -1565
rect 3592 -1565 4552 -1527
rect 3592 -1582 3794 -1565
rect 3332 -1599 3348 -1582
rect 2760 -1615 3348 -1599
rect 3778 -1599 3794 -1582
rect 4350 -1582 4552 -1565
rect 4610 -1565 5570 -1527
rect 4610 -1582 4812 -1565
rect 4350 -1599 4366 -1582
rect 3778 -1615 4366 -1599
rect 4796 -1599 4812 -1582
rect 5368 -1582 5570 -1565
rect 5368 -1599 5384 -1582
rect 4796 -1615 5384 -1599
rect -5384 -1673 -4796 -1657
rect -5384 -1690 -5368 -1673
rect -5570 -1707 -5368 -1690
rect -4812 -1690 -4796 -1673
rect -4366 -1673 -3778 -1657
rect -4366 -1690 -4350 -1673
rect -4812 -1707 -4610 -1690
rect -5570 -1745 -4610 -1707
rect -4552 -1707 -4350 -1690
rect -3794 -1690 -3778 -1673
rect -3348 -1673 -2760 -1657
rect -3348 -1690 -3332 -1673
rect -3794 -1707 -3592 -1690
rect -4552 -1745 -3592 -1707
rect -3534 -1707 -3332 -1690
rect -2776 -1690 -2760 -1673
rect -2330 -1673 -1742 -1657
rect -2330 -1690 -2314 -1673
rect -2776 -1707 -2574 -1690
rect -3534 -1745 -2574 -1707
rect -2516 -1707 -2314 -1690
rect -1758 -1690 -1742 -1673
rect -1312 -1673 -724 -1657
rect -1312 -1690 -1296 -1673
rect -1758 -1707 -1556 -1690
rect -2516 -1745 -1556 -1707
rect -1498 -1707 -1296 -1690
rect -740 -1690 -724 -1673
rect -294 -1673 294 -1657
rect -294 -1690 -278 -1673
rect -740 -1707 -538 -1690
rect -1498 -1745 -538 -1707
rect -480 -1707 -278 -1690
rect 278 -1690 294 -1673
rect 724 -1673 1312 -1657
rect 724 -1690 740 -1673
rect 278 -1707 480 -1690
rect -480 -1745 480 -1707
rect 538 -1707 740 -1690
rect 1296 -1690 1312 -1673
rect 1742 -1673 2330 -1657
rect 1742 -1690 1758 -1673
rect 1296 -1707 1498 -1690
rect 538 -1745 1498 -1707
rect 1556 -1707 1758 -1690
rect 2314 -1690 2330 -1673
rect 2760 -1673 3348 -1657
rect 2760 -1690 2776 -1673
rect 2314 -1707 2516 -1690
rect 1556 -1745 2516 -1707
rect 2574 -1707 2776 -1690
rect 3332 -1690 3348 -1673
rect 3778 -1673 4366 -1657
rect 3778 -1690 3794 -1673
rect 3332 -1707 3534 -1690
rect 2574 -1745 3534 -1707
rect 3592 -1707 3794 -1690
rect 4350 -1690 4366 -1673
rect 4796 -1673 5384 -1657
rect 4796 -1690 4812 -1673
rect 4350 -1707 4552 -1690
rect 3592 -1745 4552 -1707
rect 4610 -1707 4812 -1690
rect 5368 -1690 5384 -1673
rect 5368 -1707 5570 -1690
rect 4610 -1745 5570 -1707
rect -5570 -2383 -4610 -2345
rect -5570 -2400 -5368 -2383
rect -5384 -2417 -5368 -2400
rect -4812 -2400 -4610 -2383
rect -4552 -2383 -3592 -2345
rect -4552 -2400 -4350 -2383
rect -4812 -2417 -4796 -2400
rect -5384 -2433 -4796 -2417
rect -4366 -2417 -4350 -2400
rect -3794 -2400 -3592 -2383
rect -3534 -2383 -2574 -2345
rect -3534 -2400 -3332 -2383
rect -3794 -2417 -3778 -2400
rect -4366 -2433 -3778 -2417
rect -3348 -2417 -3332 -2400
rect -2776 -2400 -2574 -2383
rect -2516 -2383 -1556 -2345
rect -2516 -2400 -2314 -2383
rect -2776 -2417 -2760 -2400
rect -3348 -2433 -2760 -2417
rect -2330 -2417 -2314 -2400
rect -1758 -2400 -1556 -2383
rect -1498 -2383 -538 -2345
rect -1498 -2400 -1296 -2383
rect -1758 -2417 -1742 -2400
rect -2330 -2433 -1742 -2417
rect -1312 -2417 -1296 -2400
rect -740 -2400 -538 -2383
rect -480 -2383 480 -2345
rect -480 -2400 -278 -2383
rect -740 -2417 -724 -2400
rect -1312 -2433 -724 -2417
rect -294 -2417 -278 -2400
rect 278 -2400 480 -2383
rect 538 -2383 1498 -2345
rect 538 -2400 740 -2383
rect 278 -2417 294 -2400
rect -294 -2433 294 -2417
rect 724 -2417 740 -2400
rect 1296 -2400 1498 -2383
rect 1556 -2383 2516 -2345
rect 1556 -2400 1758 -2383
rect 1296 -2417 1312 -2400
rect 724 -2433 1312 -2417
rect 1742 -2417 1758 -2400
rect 2314 -2400 2516 -2383
rect 2574 -2383 3534 -2345
rect 2574 -2400 2776 -2383
rect 2314 -2417 2330 -2400
rect 1742 -2433 2330 -2417
rect 2760 -2417 2776 -2400
rect 3332 -2400 3534 -2383
rect 3592 -2383 4552 -2345
rect 3592 -2400 3794 -2383
rect 3332 -2417 3348 -2400
rect 2760 -2433 3348 -2417
rect 3778 -2417 3794 -2400
rect 4350 -2400 4552 -2383
rect 4610 -2383 5570 -2345
rect 4610 -2400 4812 -2383
rect 4350 -2417 4366 -2400
rect 3778 -2433 4366 -2417
rect 4796 -2417 4812 -2400
rect 5368 -2400 5570 -2383
rect 5368 -2417 5384 -2400
rect 4796 -2433 5384 -2417
<< polycont >>
rect -5368 2383 -4812 2417
rect -4350 2383 -3794 2417
rect -3332 2383 -2776 2417
rect -2314 2383 -1758 2417
rect -1296 2383 -740 2417
rect -278 2383 278 2417
rect 740 2383 1296 2417
rect 1758 2383 2314 2417
rect 2776 2383 3332 2417
rect 3794 2383 4350 2417
rect 4812 2383 5368 2417
rect -5368 1673 -4812 1707
rect -4350 1673 -3794 1707
rect -3332 1673 -2776 1707
rect -2314 1673 -1758 1707
rect -1296 1673 -740 1707
rect -278 1673 278 1707
rect 740 1673 1296 1707
rect 1758 1673 2314 1707
rect 2776 1673 3332 1707
rect 3794 1673 4350 1707
rect 4812 1673 5368 1707
rect -5368 1565 -4812 1599
rect -4350 1565 -3794 1599
rect -3332 1565 -2776 1599
rect -2314 1565 -1758 1599
rect -1296 1565 -740 1599
rect -278 1565 278 1599
rect 740 1565 1296 1599
rect 1758 1565 2314 1599
rect 2776 1565 3332 1599
rect 3794 1565 4350 1599
rect 4812 1565 5368 1599
rect -5368 855 -4812 889
rect -4350 855 -3794 889
rect -3332 855 -2776 889
rect -2314 855 -1758 889
rect -1296 855 -740 889
rect -278 855 278 889
rect 740 855 1296 889
rect 1758 855 2314 889
rect 2776 855 3332 889
rect 3794 855 4350 889
rect 4812 855 5368 889
rect -5368 747 -4812 781
rect -4350 747 -3794 781
rect -3332 747 -2776 781
rect -2314 747 -1758 781
rect -1296 747 -740 781
rect -278 747 278 781
rect 740 747 1296 781
rect 1758 747 2314 781
rect 2776 747 3332 781
rect 3794 747 4350 781
rect 4812 747 5368 781
rect -5368 37 -4812 71
rect -4350 37 -3794 71
rect -3332 37 -2776 71
rect -2314 37 -1758 71
rect -1296 37 -740 71
rect -278 37 278 71
rect 740 37 1296 71
rect 1758 37 2314 71
rect 2776 37 3332 71
rect 3794 37 4350 71
rect 4812 37 5368 71
rect -5368 -71 -4812 -37
rect -4350 -71 -3794 -37
rect -3332 -71 -2776 -37
rect -2314 -71 -1758 -37
rect -1296 -71 -740 -37
rect -278 -71 278 -37
rect 740 -71 1296 -37
rect 1758 -71 2314 -37
rect 2776 -71 3332 -37
rect 3794 -71 4350 -37
rect 4812 -71 5368 -37
rect -5368 -781 -4812 -747
rect -4350 -781 -3794 -747
rect -3332 -781 -2776 -747
rect -2314 -781 -1758 -747
rect -1296 -781 -740 -747
rect -278 -781 278 -747
rect 740 -781 1296 -747
rect 1758 -781 2314 -747
rect 2776 -781 3332 -747
rect 3794 -781 4350 -747
rect 4812 -781 5368 -747
rect -5368 -889 -4812 -855
rect -4350 -889 -3794 -855
rect -3332 -889 -2776 -855
rect -2314 -889 -1758 -855
rect -1296 -889 -740 -855
rect -278 -889 278 -855
rect 740 -889 1296 -855
rect 1758 -889 2314 -855
rect 2776 -889 3332 -855
rect 3794 -889 4350 -855
rect 4812 -889 5368 -855
rect -5368 -1599 -4812 -1565
rect -4350 -1599 -3794 -1565
rect -3332 -1599 -2776 -1565
rect -2314 -1599 -1758 -1565
rect -1296 -1599 -740 -1565
rect -278 -1599 278 -1565
rect 740 -1599 1296 -1565
rect 1758 -1599 2314 -1565
rect 2776 -1599 3332 -1565
rect 3794 -1599 4350 -1565
rect 4812 -1599 5368 -1565
rect -5368 -1707 -4812 -1673
rect -4350 -1707 -3794 -1673
rect -3332 -1707 -2776 -1673
rect -2314 -1707 -1758 -1673
rect -1296 -1707 -740 -1673
rect -278 -1707 278 -1673
rect 740 -1707 1296 -1673
rect 1758 -1707 2314 -1673
rect 2776 -1707 3332 -1673
rect 3794 -1707 4350 -1673
rect 4812 -1707 5368 -1673
rect -5368 -2417 -4812 -2383
rect -4350 -2417 -3794 -2383
rect -3332 -2417 -2776 -2383
rect -2314 -2417 -1758 -2383
rect -1296 -2417 -740 -2383
rect -278 -2417 278 -2383
rect 740 -2417 1296 -2383
rect 1758 -2417 2314 -2383
rect 2776 -2417 3332 -2383
rect 3794 -2417 4350 -2383
rect 4812 -2417 5368 -2383
<< locali >>
rect -5384 2383 -5368 2417
rect -4812 2383 -4796 2417
rect -4366 2383 -4350 2417
rect -3794 2383 -3778 2417
rect -3348 2383 -3332 2417
rect -2776 2383 -2760 2417
rect -2330 2383 -2314 2417
rect -1758 2383 -1742 2417
rect -1312 2383 -1296 2417
rect -740 2383 -724 2417
rect -294 2383 -278 2417
rect 278 2383 294 2417
rect 724 2383 740 2417
rect 1296 2383 1312 2417
rect 1742 2383 1758 2417
rect 2314 2383 2330 2417
rect 2760 2383 2776 2417
rect 3332 2383 3348 2417
rect 3778 2383 3794 2417
rect 4350 2383 4366 2417
rect 4796 2383 4812 2417
rect 5368 2383 5384 2417
rect -5616 2333 -5582 2349
rect -5616 1741 -5582 1757
rect -4598 2333 -4564 2349
rect -4598 1741 -4564 1757
rect -3580 2333 -3546 2349
rect -3580 1741 -3546 1757
rect -2562 2333 -2528 2349
rect -2562 1741 -2528 1757
rect -1544 2333 -1510 2349
rect -1544 1741 -1510 1757
rect -526 2333 -492 2349
rect -526 1741 -492 1757
rect 492 2333 526 2349
rect 492 1741 526 1757
rect 1510 2333 1544 2349
rect 1510 1741 1544 1757
rect 2528 2333 2562 2349
rect 2528 1741 2562 1757
rect 3546 2333 3580 2349
rect 3546 1741 3580 1757
rect 4564 2333 4598 2349
rect 4564 1741 4598 1757
rect 5582 2333 5616 2349
rect 5582 1741 5616 1757
rect -5384 1673 -5368 1707
rect -4812 1673 -4796 1707
rect -4366 1673 -4350 1707
rect -3794 1673 -3778 1707
rect -3348 1673 -3332 1707
rect -2776 1673 -2760 1707
rect -2330 1673 -2314 1707
rect -1758 1673 -1742 1707
rect -1312 1673 -1296 1707
rect -740 1673 -724 1707
rect -294 1673 -278 1707
rect 278 1673 294 1707
rect 724 1673 740 1707
rect 1296 1673 1312 1707
rect 1742 1673 1758 1707
rect 2314 1673 2330 1707
rect 2760 1673 2776 1707
rect 3332 1673 3348 1707
rect 3778 1673 3794 1707
rect 4350 1673 4366 1707
rect 4796 1673 4812 1707
rect 5368 1673 5384 1707
rect -5384 1565 -5368 1599
rect -4812 1565 -4796 1599
rect -4366 1565 -4350 1599
rect -3794 1565 -3778 1599
rect -3348 1565 -3332 1599
rect -2776 1565 -2760 1599
rect -2330 1565 -2314 1599
rect -1758 1565 -1742 1599
rect -1312 1565 -1296 1599
rect -740 1565 -724 1599
rect -294 1565 -278 1599
rect 278 1565 294 1599
rect 724 1565 740 1599
rect 1296 1565 1312 1599
rect 1742 1565 1758 1599
rect 2314 1565 2330 1599
rect 2760 1565 2776 1599
rect 3332 1565 3348 1599
rect 3778 1565 3794 1599
rect 4350 1565 4366 1599
rect 4796 1565 4812 1599
rect 5368 1565 5384 1599
rect -5616 1515 -5582 1531
rect -5616 923 -5582 939
rect -4598 1515 -4564 1531
rect -4598 923 -4564 939
rect -3580 1515 -3546 1531
rect -3580 923 -3546 939
rect -2562 1515 -2528 1531
rect -2562 923 -2528 939
rect -1544 1515 -1510 1531
rect -1544 923 -1510 939
rect -526 1515 -492 1531
rect -526 923 -492 939
rect 492 1515 526 1531
rect 492 923 526 939
rect 1510 1515 1544 1531
rect 1510 923 1544 939
rect 2528 1515 2562 1531
rect 2528 923 2562 939
rect 3546 1515 3580 1531
rect 3546 923 3580 939
rect 4564 1515 4598 1531
rect 4564 923 4598 939
rect 5582 1515 5616 1531
rect 5582 923 5616 939
rect -5384 855 -5368 889
rect -4812 855 -4796 889
rect -4366 855 -4350 889
rect -3794 855 -3778 889
rect -3348 855 -3332 889
rect -2776 855 -2760 889
rect -2330 855 -2314 889
rect -1758 855 -1742 889
rect -1312 855 -1296 889
rect -740 855 -724 889
rect -294 855 -278 889
rect 278 855 294 889
rect 724 855 740 889
rect 1296 855 1312 889
rect 1742 855 1758 889
rect 2314 855 2330 889
rect 2760 855 2776 889
rect 3332 855 3348 889
rect 3778 855 3794 889
rect 4350 855 4366 889
rect 4796 855 4812 889
rect 5368 855 5384 889
rect -5384 747 -5368 781
rect -4812 747 -4796 781
rect -4366 747 -4350 781
rect -3794 747 -3778 781
rect -3348 747 -3332 781
rect -2776 747 -2760 781
rect -2330 747 -2314 781
rect -1758 747 -1742 781
rect -1312 747 -1296 781
rect -740 747 -724 781
rect -294 747 -278 781
rect 278 747 294 781
rect 724 747 740 781
rect 1296 747 1312 781
rect 1742 747 1758 781
rect 2314 747 2330 781
rect 2760 747 2776 781
rect 3332 747 3348 781
rect 3778 747 3794 781
rect 4350 747 4366 781
rect 4796 747 4812 781
rect 5368 747 5384 781
rect -5616 697 -5582 713
rect -5616 105 -5582 121
rect -4598 697 -4564 713
rect -4598 105 -4564 121
rect -3580 697 -3546 713
rect -3580 105 -3546 121
rect -2562 697 -2528 713
rect -2562 105 -2528 121
rect -1544 697 -1510 713
rect -1544 105 -1510 121
rect -526 697 -492 713
rect -526 105 -492 121
rect 492 697 526 713
rect 492 105 526 121
rect 1510 697 1544 713
rect 1510 105 1544 121
rect 2528 697 2562 713
rect 2528 105 2562 121
rect 3546 697 3580 713
rect 3546 105 3580 121
rect 4564 697 4598 713
rect 4564 105 4598 121
rect 5582 697 5616 713
rect 5582 105 5616 121
rect -5384 37 -5368 71
rect -4812 37 -4796 71
rect -4366 37 -4350 71
rect -3794 37 -3778 71
rect -3348 37 -3332 71
rect -2776 37 -2760 71
rect -2330 37 -2314 71
rect -1758 37 -1742 71
rect -1312 37 -1296 71
rect -740 37 -724 71
rect -294 37 -278 71
rect 278 37 294 71
rect 724 37 740 71
rect 1296 37 1312 71
rect 1742 37 1758 71
rect 2314 37 2330 71
rect 2760 37 2776 71
rect 3332 37 3348 71
rect 3778 37 3794 71
rect 4350 37 4366 71
rect 4796 37 4812 71
rect 5368 37 5384 71
rect -5384 -71 -5368 -37
rect -4812 -71 -4796 -37
rect -4366 -71 -4350 -37
rect -3794 -71 -3778 -37
rect -3348 -71 -3332 -37
rect -2776 -71 -2760 -37
rect -2330 -71 -2314 -37
rect -1758 -71 -1742 -37
rect -1312 -71 -1296 -37
rect -740 -71 -724 -37
rect -294 -71 -278 -37
rect 278 -71 294 -37
rect 724 -71 740 -37
rect 1296 -71 1312 -37
rect 1742 -71 1758 -37
rect 2314 -71 2330 -37
rect 2760 -71 2776 -37
rect 3332 -71 3348 -37
rect 3778 -71 3794 -37
rect 4350 -71 4366 -37
rect 4796 -71 4812 -37
rect 5368 -71 5384 -37
rect -5616 -121 -5582 -105
rect -5616 -713 -5582 -697
rect -4598 -121 -4564 -105
rect -4598 -713 -4564 -697
rect -3580 -121 -3546 -105
rect -3580 -713 -3546 -697
rect -2562 -121 -2528 -105
rect -2562 -713 -2528 -697
rect -1544 -121 -1510 -105
rect -1544 -713 -1510 -697
rect -526 -121 -492 -105
rect -526 -713 -492 -697
rect 492 -121 526 -105
rect 492 -713 526 -697
rect 1510 -121 1544 -105
rect 1510 -713 1544 -697
rect 2528 -121 2562 -105
rect 2528 -713 2562 -697
rect 3546 -121 3580 -105
rect 3546 -713 3580 -697
rect 4564 -121 4598 -105
rect 4564 -713 4598 -697
rect 5582 -121 5616 -105
rect 5582 -713 5616 -697
rect -5384 -781 -5368 -747
rect -4812 -781 -4796 -747
rect -4366 -781 -4350 -747
rect -3794 -781 -3778 -747
rect -3348 -781 -3332 -747
rect -2776 -781 -2760 -747
rect -2330 -781 -2314 -747
rect -1758 -781 -1742 -747
rect -1312 -781 -1296 -747
rect -740 -781 -724 -747
rect -294 -781 -278 -747
rect 278 -781 294 -747
rect 724 -781 740 -747
rect 1296 -781 1312 -747
rect 1742 -781 1758 -747
rect 2314 -781 2330 -747
rect 2760 -781 2776 -747
rect 3332 -781 3348 -747
rect 3778 -781 3794 -747
rect 4350 -781 4366 -747
rect 4796 -781 4812 -747
rect 5368 -781 5384 -747
rect -5384 -889 -5368 -855
rect -4812 -889 -4796 -855
rect -4366 -889 -4350 -855
rect -3794 -889 -3778 -855
rect -3348 -889 -3332 -855
rect -2776 -889 -2760 -855
rect -2330 -889 -2314 -855
rect -1758 -889 -1742 -855
rect -1312 -889 -1296 -855
rect -740 -889 -724 -855
rect -294 -889 -278 -855
rect 278 -889 294 -855
rect 724 -889 740 -855
rect 1296 -889 1312 -855
rect 1742 -889 1758 -855
rect 2314 -889 2330 -855
rect 2760 -889 2776 -855
rect 3332 -889 3348 -855
rect 3778 -889 3794 -855
rect 4350 -889 4366 -855
rect 4796 -889 4812 -855
rect 5368 -889 5384 -855
rect -5616 -939 -5582 -923
rect -5616 -1531 -5582 -1515
rect -4598 -939 -4564 -923
rect -4598 -1531 -4564 -1515
rect -3580 -939 -3546 -923
rect -3580 -1531 -3546 -1515
rect -2562 -939 -2528 -923
rect -2562 -1531 -2528 -1515
rect -1544 -939 -1510 -923
rect -1544 -1531 -1510 -1515
rect -526 -939 -492 -923
rect -526 -1531 -492 -1515
rect 492 -939 526 -923
rect 492 -1531 526 -1515
rect 1510 -939 1544 -923
rect 1510 -1531 1544 -1515
rect 2528 -939 2562 -923
rect 2528 -1531 2562 -1515
rect 3546 -939 3580 -923
rect 3546 -1531 3580 -1515
rect 4564 -939 4598 -923
rect 4564 -1531 4598 -1515
rect 5582 -939 5616 -923
rect 5582 -1531 5616 -1515
rect -5384 -1599 -5368 -1565
rect -4812 -1599 -4796 -1565
rect -4366 -1599 -4350 -1565
rect -3794 -1599 -3778 -1565
rect -3348 -1599 -3332 -1565
rect -2776 -1599 -2760 -1565
rect -2330 -1599 -2314 -1565
rect -1758 -1599 -1742 -1565
rect -1312 -1599 -1296 -1565
rect -740 -1599 -724 -1565
rect -294 -1599 -278 -1565
rect 278 -1599 294 -1565
rect 724 -1599 740 -1565
rect 1296 -1599 1312 -1565
rect 1742 -1599 1758 -1565
rect 2314 -1599 2330 -1565
rect 2760 -1599 2776 -1565
rect 3332 -1599 3348 -1565
rect 3778 -1599 3794 -1565
rect 4350 -1599 4366 -1565
rect 4796 -1599 4812 -1565
rect 5368 -1599 5384 -1565
rect -5384 -1707 -5368 -1673
rect -4812 -1707 -4796 -1673
rect -4366 -1707 -4350 -1673
rect -3794 -1707 -3778 -1673
rect -3348 -1707 -3332 -1673
rect -2776 -1707 -2760 -1673
rect -2330 -1707 -2314 -1673
rect -1758 -1707 -1742 -1673
rect -1312 -1707 -1296 -1673
rect -740 -1707 -724 -1673
rect -294 -1707 -278 -1673
rect 278 -1707 294 -1673
rect 724 -1707 740 -1673
rect 1296 -1707 1312 -1673
rect 1742 -1707 1758 -1673
rect 2314 -1707 2330 -1673
rect 2760 -1707 2776 -1673
rect 3332 -1707 3348 -1673
rect 3778 -1707 3794 -1673
rect 4350 -1707 4366 -1673
rect 4796 -1707 4812 -1673
rect 5368 -1707 5384 -1673
rect -5616 -1757 -5582 -1741
rect -5616 -2349 -5582 -2333
rect -4598 -1757 -4564 -1741
rect -4598 -2349 -4564 -2333
rect -3580 -1757 -3546 -1741
rect -3580 -2349 -3546 -2333
rect -2562 -1757 -2528 -1741
rect -2562 -2349 -2528 -2333
rect -1544 -1757 -1510 -1741
rect -1544 -2349 -1510 -2333
rect -526 -1757 -492 -1741
rect -526 -2349 -492 -2333
rect 492 -1757 526 -1741
rect 492 -2349 526 -2333
rect 1510 -1757 1544 -1741
rect 1510 -2349 1544 -2333
rect 2528 -1757 2562 -1741
rect 2528 -2349 2562 -2333
rect 3546 -1757 3580 -1741
rect 3546 -2349 3580 -2333
rect 4564 -1757 4598 -1741
rect 4564 -2349 4598 -2333
rect 5582 -1757 5616 -1741
rect 5582 -2349 5616 -2333
rect -5384 -2417 -5368 -2383
rect -4812 -2417 -4796 -2383
rect -4366 -2417 -4350 -2383
rect -3794 -2417 -3778 -2383
rect -3348 -2417 -3332 -2383
rect -2776 -2417 -2760 -2383
rect -2330 -2417 -2314 -2383
rect -1758 -2417 -1742 -2383
rect -1312 -2417 -1296 -2383
rect -740 -2417 -724 -2383
rect -294 -2417 -278 -2383
rect 278 -2417 294 -2383
rect 724 -2417 740 -2383
rect 1296 -2417 1312 -2383
rect 1742 -2417 1758 -2383
rect 2314 -2417 2330 -2383
rect 2760 -2417 2776 -2383
rect 3332 -2417 3348 -2383
rect 3778 -2417 3794 -2383
rect 4350 -2417 4366 -2383
rect 4796 -2417 4812 -2383
rect 5368 -2417 5384 -2383
<< viali >>
rect -5322 2383 -4858 2417
rect -4304 2383 -3840 2417
rect -3286 2383 -2822 2417
rect -2268 2383 -1804 2417
rect -1250 2383 -786 2417
rect -232 2383 232 2417
rect 786 2383 1250 2417
rect 1804 2383 2268 2417
rect 2822 2383 3286 2417
rect 3840 2383 4304 2417
rect 4858 2383 5322 2417
rect -5616 1757 -5582 2333
rect -4598 1757 -4564 2333
rect -3580 1757 -3546 2333
rect -2562 1757 -2528 2333
rect -1544 1757 -1510 2333
rect -526 1757 -492 2333
rect 492 1757 526 2333
rect 1510 1757 1544 2333
rect 2528 1757 2562 2333
rect 3546 1757 3580 2333
rect 4564 1757 4598 2333
rect 5582 1757 5616 2333
rect -5322 1673 -4858 1707
rect -4304 1673 -3840 1707
rect -3286 1673 -2822 1707
rect -2268 1673 -1804 1707
rect -1250 1673 -786 1707
rect -232 1673 232 1707
rect 786 1673 1250 1707
rect 1804 1673 2268 1707
rect 2822 1673 3286 1707
rect 3840 1673 4304 1707
rect 4858 1673 5322 1707
rect -5322 1565 -4858 1599
rect -4304 1565 -3840 1599
rect -3286 1565 -2822 1599
rect -2268 1565 -1804 1599
rect -1250 1565 -786 1599
rect -232 1565 232 1599
rect 786 1565 1250 1599
rect 1804 1565 2268 1599
rect 2822 1565 3286 1599
rect 3840 1565 4304 1599
rect 4858 1565 5322 1599
rect -5616 939 -5582 1515
rect -4598 939 -4564 1515
rect -3580 939 -3546 1515
rect -2562 939 -2528 1515
rect -1544 939 -1510 1515
rect -526 939 -492 1515
rect 492 939 526 1515
rect 1510 939 1544 1515
rect 2528 939 2562 1515
rect 3546 939 3580 1515
rect 4564 939 4598 1515
rect 5582 939 5616 1515
rect -5322 855 -4858 889
rect -4304 855 -3840 889
rect -3286 855 -2822 889
rect -2268 855 -1804 889
rect -1250 855 -786 889
rect -232 855 232 889
rect 786 855 1250 889
rect 1804 855 2268 889
rect 2822 855 3286 889
rect 3840 855 4304 889
rect 4858 855 5322 889
rect -5322 747 -4858 781
rect -4304 747 -3840 781
rect -3286 747 -2822 781
rect -2268 747 -1804 781
rect -1250 747 -786 781
rect -232 747 232 781
rect 786 747 1250 781
rect 1804 747 2268 781
rect 2822 747 3286 781
rect 3840 747 4304 781
rect 4858 747 5322 781
rect -5616 121 -5582 697
rect -4598 121 -4564 697
rect -3580 121 -3546 697
rect -2562 121 -2528 697
rect -1544 121 -1510 697
rect -526 121 -492 697
rect 492 121 526 697
rect 1510 121 1544 697
rect 2528 121 2562 697
rect 3546 121 3580 697
rect 4564 121 4598 697
rect 5582 121 5616 697
rect -5322 37 -4858 71
rect -4304 37 -3840 71
rect -3286 37 -2822 71
rect -2268 37 -1804 71
rect -1250 37 -786 71
rect -232 37 232 71
rect 786 37 1250 71
rect 1804 37 2268 71
rect 2822 37 3286 71
rect 3840 37 4304 71
rect 4858 37 5322 71
rect -5322 -71 -4858 -37
rect -4304 -71 -3840 -37
rect -3286 -71 -2822 -37
rect -2268 -71 -1804 -37
rect -1250 -71 -786 -37
rect -232 -71 232 -37
rect 786 -71 1250 -37
rect 1804 -71 2268 -37
rect 2822 -71 3286 -37
rect 3840 -71 4304 -37
rect 4858 -71 5322 -37
rect -5616 -697 -5582 -121
rect -4598 -697 -4564 -121
rect -3580 -697 -3546 -121
rect -2562 -697 -2528 -121
rect -1544 -697 -1510 -121
rect -526 -697 -492 -121
rect 492 -697 526 -121
rect 1510 -697 1544 -121
rect 2528 -697 2562 -121
rect 3546 -697 3580 -121
rect 4564 -697 4598 -121
rect 5582 -697 5616 -121
rect -5322 -781 -4858 -747
rect -4304 -781 -3840 -747
rect -3286 -781 -2822 -747
rect -2268 -781 -1804 -747
rect -1250 -781 -786 -747
rect -232 -781 232 -747
rect 786 -781 1250 -747
rect 1804 -781 2268 -747
rect 2822 -781 3286 -747
rect 3840 -781 4304 -747
rect 4858 -781 5322 -747
rect -5322 -889 -4858 -855
rect -4304 -889 -3840 -855
rect -3286 -889 -2822 -855
rect -2268 -889 -1804 -855
rect -1250 -889 -786 -855
rect -232 -889 232 -855
rect 786 -889 1250 -855
rect 1804 -889 2268 -855
rect 2822 -889 3286 -855
rect 3840 -889 4304 -855
rect 4858 -889 5322 -855
rect -5616 -1515 -5582 -939
rect -4598 -1515 -4564 -939
rect -3580 -1515 -3546 -939
rect -2562 -1515 -2528 -939
rect -1544 -1515 -1510 -939
rect -526 -1515 -492 -939
rect 492 -1515 526 -939
rect 1510 -1515 1544 -939
rect 2528 -1515 2562 -939
rect 3546 -1515 3580 -939
rect 4564 -1515 4598 -939
rect 5582 -1515 5616 -939
rect -5322 -1599 -4858 -1565
rect -4304 -1599 -3840 -1565
rect -3286 -1599 -2822 -1565
rect -2268 -1599 -1804 -1565
rect -1250 -1599 -786 -1565
rect -232 -1599 232 -1565
rect 786 -1599 1250 -1565
rect 1804 -1599 2268 -1565
rect 2822 -1599 3286 -1565
rect 3840 -1599 4304 -1565
rect 4858 -1599 5322 -1565
rect -5322 -1707 -4858 -1673
rect -4304 -1707 -3840 -1673
rect -3286 -1707 -2822 -1673
rect -2268 -1707 -1804 -1673
rect -1250 -1707 -786 -1673
rect -232 -1707 232 -1673
rect 786 -1707 1250 -1673
rect 1804 -1707 2268 -1673
rect 2822 -1707 3286 -1673
rect 3840 -1707 4304 -1673
rect 4858 -1707 5322 -1673
rect -5616 -2333 -5582 -1757
rect -4598 -2333 -4564 -1757
rect -3580 -2333 -3546 -1757
rect -2562 -2333 -2528 -1757
rect -1544 -2333 -1510 -1757
rect -526 -2333 -492 -1757
rect 492 -2333 526 -1757
rect 1510 -2333 1544 -1757
rect 2528 -2333 2562 -1757
rect 3546 -2333 3580 -1757
rect 4564 -2333 4598 -1757
rect 5582 -2333 5616 -1757
rect -5322 -2417 -4858 -2383
rect -4304 -2417 -3840 -2383
rect -3286 -2417 -2822 -2383
rect -2268 -2417 -1804 -2383
rect -1250 -2417 -786 -2383
rect -232 -2417 232 -2383
rect 786 -2417 1250 -2383
rect 1804 -2417 2268 -2383
rect 2822 -2417 3286 -2383
rect 3840 -2417 4304 -2383
rect 4858 -2417 5322 -2383
<< metal1 >>
rect -5334 2417 -4846 2423
rect -5334 2383 -5322 2417
rect -4858 2383 -4846 2417
rect -5334 2377 -4846 2383
rect -4316 2417 -3828 2423
rect -4316 2383 -4304 2417
rect -3840 2383 -3828 2417
rect -4316 2377 -3828 2383
rect -3298 2417 -2810 2423
rect -3298 2383 -3286 2417
rect -2822 2383 -2810 2417
rect -3298 2377 -2810 2383
rect -2280 2417 -1792 2423
rect -2280 2383 -2268 2417
rect -1804 2383 -1792 2417
rect -2280 2377 -1792 2383
rect -1262 2417 -774 2423
rect -1262 2383 -1250 2417
rect -786 2383 -774 2417
rect -1262 2377 -774 2383
rect -244 2417 244 2423
rect -244 2383 -232 2417
rect 232 2383 244 2417
rect -244 2377 244 2383
rect 774 2417 1262 2423
rect 774 2383 786 2417
rect 1250 2383 1262 2417
rect 774 2377 1262 2383
rect 1792 2417 2280 2423
rect 1792 2383 1804 2417
rect 2268 2383 2280 2417
rect 1792 2377 2280 2383
rect 2810 2417 3298 2423
rect 2810 2383 2822 2417
rect 3286 2383 3298 2417
rect 2810 2377 3298 2383
rect 3828 2417 4316 2423
rect 3828 2383 3840 2417
rect 4304 2383 4316 2417
rect 3828 2377 4316 2383
rect 4846 2417 5334 2423
rect 4846 2383 4858 2417
rect 5322 2383 5334 2417
rect 4846 2377 5334 2383
rect -5622 2333 -5576 2345
rect -5622 1757 -5616 2333
rect -5582 1757 -5576 2333
rect -5622 1745 -5576 1757
rect -4604 2333 -4558 2345
rect -4604 1757 -4598 2333
rect -4564 1757 -4558 2333
rect -4604 1745 -4558 1757
rect -3586 2333 -3540 2345
rect -3586 1757 -3580 2333
rect -3546 1757 -3540 2333
rect -3586 1745 -3540 1757
rect -2568 2333 -2522 2345
rect -2568 1757 -2562 2333
rect -2528 1757 -2522 2333
rect -2568 1745 -2522 1757
rect -1550 2333 -1504 2345
rect -1550 1757 -1544 2333
rect -1510 1757 -1504 2333
rect -1550 1745 -1504 1757
rect -532 2333 -486 2345
rect -532 1757 -526 2333
rect -492 1757 -486 2333
rect -532 1745 -486 1757
rect 486 2333 532 2345
rect 486 1757 492 2333
rect 526 1757 532 2333
rect 486 1745 532 1757
rect 1504 2333 1550 2345
rect 1504 1757 1510 2333
rect 1544 1757 1550 2333
rect 1504 1745 1550 1757
rect 2522 2333 2568 2345
rect 2522 1757 2528 2333
rect 2562 1757 2568 2333
rect 2522 1745 2568 1757
rect 3540 2333 3586 2345
rect 3540 1757 3546 2333
rect 3580 1757 3586 2333
rect 3540 1745 3586 1757
rect 4558 2333 4604 2345
rect 4558 1757 4564 2333
rect 4598 1757 4604 2333
rect 4558 1745 4604 1757
rect 5576 2333 5622 2345
rect 5576 1757 5582 2333
rect 5616 1757 5622 2333
rect 5576 1745 5622 1757
rect -5334 1707 -4846 1713
rect -5334 1673 -5322 1707
rect -4858 1673 -4846 1707
rect -5334 1667 -4846 1673
rect -4316 1707 -3828 1713
rect -4316 1673 -4304 1707
rect -3840 1673 -3828 1707
rect -4316 1667 -3828 1673
rect -3298 1707 -2810 1713
rect -3298 1673 -3286 1707
rect -2822 1673 -2810 1707
rect -3298 1667 -2810 1673
rect -2280 1707 -1792 1713
rect -2280 1673 -2268 1707
rect -1804 1673 -1792 1707
rect -2280 1667 -1792 1673
rect -1262 1707 -774 1713
rect -1262 1673 -1250 1707
rect -786 1673 -774 1707
rect -1262 1667 -774 1673
rect -244 1707 244 1713
rect -244 1673 -232 1707
rect 232 1673 244 1707
rect -244 1667 244 1673
rect 774 1707 1262 1713
rect 774 1673 786 1707
rect 1250 1673 1262 1707
rect 774 1667 1262 1673
rect 1792 1707 2280 1713
rect 1792 1673 1804 1707
rect 2268 1673 2280 1707
rect 1792 1667 2280 1673
rect 2810 1707 3298 1713
rect 2810 1673 2822 1707
rect 3286 1673 3298 1707
rect 2810 1667 3298 1673
rect 3828 1707 4316 1713
rect 3828 1673 3840 1707
rect 4304 1673 4316 1707
rect 3828 1667 4316 1673
rect 4846 1707 5334 1713
rect 4846 1673 4858 1707
rect 5322 1673 5334 1707
rect 4846 1667 5334 1673
rect -5334 1599 -4846 1605
rect -5334 1565 -5322 1599
rect -4858 1565 -4846 1599
rect -5334 1559 -4846 1565
rect -4316 1599 -3828 1605
rect -4316 1565 -4304 1599
rect -3840 1565 -3828 1599
rect -4316 1559 -3828 1565
rect -3298 1599 -2810 1605
rect -3298 1565 -3286 1599
rect -2822 1565 -2810 1599
rect -3298 1559 -2810 1565
rect -2280 1599 -1792 1605
rect -2280 1565 -2268 1599
rect -1804 1565 -1792 1599
rect -2280 1559 -1792 1565
rect -1262 1599 -774 1605
rect -1262 1565 -1250 1599
rect -786 1565 -774 1599
rect -1262 1559 -774 1565
rect -244 1599 244 1605
rect -244 1565 -232 1599
rect 232 1565 244 1599
rect -244 1559 244 1565
rect 774 1599 1262 1605
rect 774 1565 786 1599
rect 1250 1565 1262 1599
rect 774 1559 1262 1565
rect 1792 1599 2280 1605
rect 1792 1565 1804 1599
rect 2268 1565 2280 1599
rect 1792 1559 2280 1565
rect 2810 1599 3298 1605
rect 2810 1565 2822 1599
rect 3286 1565 3298 1599
rect 2810 1559 3298 1565
rect 3828 1599 4316 1605
rect 3828 1565 3840 1599
rect 4304 1565 4316 1599
rect 3828 1559 4316 1565
rect 4846 1599 5334 1605
rect 4846 1565 4858 1599
rect 5322 1565 5334 1599
rect 4846 1559 5334 1565
rect -5622 1515 -5576 1527
rect -5622 939 -5616 1515
rect -5582 939 -5576 1515
rect -5622 927 -5576 939
rect -4604 1515 -4558 1527
rect -4604 939 -4598 1515
rect -4564 939 -4558 1515
rect -4604 927 -4558 939
rect -3586 1515 -3540 1527
rect -3586 939 -3580 1515
rect -3546 939 -3540 1515
rect -3586 927 -3540 939
rect -2568 1515 -2522 1527
rect -2568 939 -2562 1515
rect -2528 939 -2522 1515
rect -2568 927 -2522 939
rect -1550 1515 -1504 1527
rect -1550 939 -1544 1515
rect -1510 939 -1504 1515
rect -1550 927 -1504 939
rect -532 1515 -486 1527
rect -532 939 -526 1515
rect -492 939 -486 1515
rect -532 927 -486 939
rect 486 1515 532 1527
rect 486 939 492 1515
rect 526 939 532 1515
rect 486 927 532 939
rect 1504 1515 1550 1527
rect 1504 939 1510 1515
rect 1544 939 1550 1515
rect 1504 927 1550 939
rect 2522 1515 2568 1527
rect 2522 939 2528 1515
rect 2562 939 2568 1515
rect 2522 927 2568 939
rect 3540 1515 3586 1527
rect 3540 939 3546 1515
rect 3580 939 3586 1515
rect 3540 927 3586 939
rect 4558 1515 4604 1527
rect 4558 939 4564 1515
rect 4598 939 4604 1515
rect 4558 927 4604 939
rect 5576 1515 5622 1527
rect 5576 939 5582 1515
rect 5616 939 5622 1515
rect 5576 927 5622 939
rect -5334 889 -4846 895
rect -5334 855 -5322 889
rect -4858 855 -4846 889
rect -5334 849 -4846 855
rect -4316 889 -3828 895
rect -4316 855 -4304 889
rect -3840 855 -3828 889
rect -4316 849 -3828 855
rect -3298 889 -2810 895
rect -3298 855 -3286 889
rect -2822 855 -2810 889
rect -3298 849 -2810 855
rect -2280 889 -1792 895
rect -2280 855 -2268 889
rect -1804 855 -1792 889
rect -2280 849 -1792 855
rect -1262 889 -774 895
rect -1262 855 -1250 889
rect -786 855 -774 889
rect -1262 849 -774 855
rect -244 889 244 895
rect -244 855 -232 889
rect 232 855 244 889
rect -244 849 244 855
rect 774 889 1262 895
rect 774 855 786 889
rect 1250 855 1262 889
rect 774 849 1262 855
rect 1792 889 2280 895
rect 1792 855 1804 889
rect 2268 855 2280 889
rect 1792 849 2280 855
rect 2810 889 3298 895
rect 2810 855 2822 889
rect 3286 855 3298 889
rect 2810 849 3298 855
rect 3828 889 4316 895
rect 3828 855 3840 889
rect 4304 855 4316 889
rect 3828 849 4316 855
rect 4846 889 5334 895
rect 4846 855 4858 889
rect 5322 855 5334 889
rect 4846 849 5334 855
rect -5334 781 -4846 787
rect -5334 747 -5322 781
rect -4858 747 -4846 781
rect -5334 741 -4846 747
rect -4316 781 -3828 787
rect -4316 747 -4304 781
rect -3840 747 -3828 781
rect -4316 741 -3828 747
rect -3298 781 -2810 787
rect -3298 747 -3286 781
rect -2822 747 -2810 781
rect -3298 741 -2810 747
rect -2280 781 -1792 787
rect -2280 747 -2268 781
rect -1804 747 -1792 781
rect -2280 741 -1792 747
rect -1262 781 -774 787
rect -1262 747 -1250 781
rect -786 747 -774 781
rect -1262 741 -774 747
rect -244 781 244 787
rect -244 747 -232 781
rect 232 747 244 781
rect -244 741 244 747
rect 774 781 1262 787
rect 774 747 786 781
rect 1250 747 1262 781
rect 774 741 1262 747
rect 1792 781 2280 787
rect 1792 747 1804 781
rect 2268 747 2280 781
rect 1792 741 2280 747
rect 2810 781 3298 787
rect 2810 747 2822 781
rect 3286 747 3298 781
rect 2810 741 3298 747
rect 3828 781 4316 787
rect 3828 747 3840 781
rect 4304 747 4316 781
rect 3828 741 4316 747
rect 4846 781 5334 787
rect 4846 747 4858 781
rect 5322 747 5334 781
rect 4846 741 5334 747
rect -5622 697 -5576 709
rect -5622 121 -5616 697
rect -5582 121 -5576 697
rect -5622 109 -5576 121
rect -4604 697 -4558 709
rect -4604 121 -4598 697
rect -4564 121 -4558 697
rect -4604 109 -4558 121
rect -3586 697 -3540 709
rect -3586 121 -3580 697
rect -3546 121 -3540 697
rect -3586 109 -3540 121
rect -2568 697 -2522 709
rect -2568 121 -2562 697
rect -2528 121 -2522 697
rect -2568 109 -2522 121
rect -1550 697 -1504 709
rect -1550 121 -1544 697
rect -1510 121 -1504 697
rect -1550 109 -1504 121
rect -532 697 -486 709
rect -532 121 -526 697
rect -492 121 -486 697
rect -532 109 -486 121
rect 486 697 532 709
rect 486 121 492 697
rect 526 121 532 697
rect 486 109 532 121
rect 1504 697 1550 709
rect 1504 121 1510 697
rect 1544 121 1550 697
rect 1504 109 1550 121
rect 2522 697 2568 709
rect 2522 121 2528 697
rect 2562 121 2568 697
rect 2522 109 2568 121
rect 3540 697 3586 709
rect 3540 121 3546 697
rect 3580 121 3586 697
rect 3540 109 3586 121
rect 4558 697 4604 709
rect 4558 121 4564 697
rect 4598 121 4604 697
rect 4558 109 4604 121
rect 5576 697 5622 709
rect 5576 121 5582 697
rect 5616 121 5622 697
rect 5576 109 5622 121
rect -5334 71 -4846 77
rect -5334 37 -5322 71
rect -4858 37 -4846 71
rect -5334 31 -4846 37
rect -4316 71 -3828 77
rect -4316 37 -4304 71
rect -3840 37 -3828 71
rect -4316 31 -3828 37
rect -3298 71 -2810 77
rect -3298 37 -3286 71
rect -2822 37 -2810 71
rect -3298 31 -2810 37
rect -2280 71 -1792 77
rect -2280 37 -2268 71
rect -1804 37 -1792 71
rect -2280 31 -1792 37
rect -1262 71 -774 77
rect -1262 37 -1250 71
rect -786 37 -774 71
rect -1262 31 -774 37
rect -244 71 244 77
rect -244 37 -232 71
rect 232 37 244 71
rect -244 31 244 37
rect 774 71 1262 77
rect 774 37 786 71
rect 1250 37 1262 71
rect 774 31 1262 37
rect 1792 71 2280 77
rect 1792 37 1804 71
rect 2268 37 2280 71
rect 1792 31 2280 37
rect 2810 71 3298 77
rect 2810 37 2822 71
rect 3286 37 3298 71
rect 2810 31 3298 37
rect 3828 71 4316 77
rect 3828 37 3840 71
rect 4304 37 4316 71
rect 3828 31 4316 37
rect 4846 71 5334 77
rect 4846 37 4858 71
rect 5322 37 5334 71
rect 4846 31 5334 37
rect -5334 -37 -4846 -31
rect -5334 -71 -5322 -37
rect -4858 -71 -4846 -37
rect -5334 -77 -4846 -71
rect -4316 -37 -3828 -31
rect -4316 -71 -4304 -37
rect -3840 -71 -3828 -37
rect -4316 -77 -3828 -71
rect -3298 -37 -2810 -31
rect -3298 -71 -3286 -37
rect -2822 -71 -2810 -37
rect -3298 -77 -2810 -71
rect -2280 -37 -1792 -31
rect -2280 -71 -2268 -37
rect -1804 -71 -1792 -37
rect -2280 -77 -1792 -71
rect -1262 -37 -774 -31
rect -1262 -71 -1250 -37
rect -786 -71 -774 -37
rect -1262 -77 -774 -71
rect -244 -37 244 -31
rect -244 -71 -232 -37
rect 232 -71 244 -37
rect -244 -77 244 -71
rect 774 -37 1262 -31
rect 774 -71 786 -37
rect 1250 -71 1262 -37
rect 774 -77 1262 -71
rect 1792 -37 2280 -31
rect 1792 -71 1804 -37
rect 2268 -71 2280 -37
rect 1792 -77 2280 -71
rect 2810 -37 3298 -31
rect 2810 -71 2822 -37
rect 3286 -71 3298 -37
rect 2810 -77 3298 -71
rect 3828 -37 4316 -31
rect 3828 -71 3840 -37
rect 4304 -71 4316 -37
rect 3828 -77 4316 -71
rect 4846 -37 5334 -31
rect 4846 -71 4858 -37
rect 5322 -71 5334 -37
rect 4846 -77 5334 -71
rect -5622 -121 -5576 -109
rect -5622 -697 -5616 -121
rect -5582 -697 -5576 -121
rect -5622 -709 -5576 -697
rect -4604 -121 -4558 -109
rect -4604 -697 -4598 -121
rect -4564 -697 -4558 -121
rect -4604 -709 -4558 -697
rect -3586 -121 -3540 -109
rect -3586 -697 -3580 -121
rect -3546 -697 -3540 -121
rect -3586 -709 -3540 -697
rect -2568 -121 -2522 -109
rect -2568 -697 -2562 -121
rect -2528 -697 -2522 -121
rect -2568 -709 -2522 -697
rect -1550 -121 -1504 -109
rect -1550 -697 -1544 -121
rect -1510 -697 -1504 -121
rect -1550 -709 -1504 -697
rect -532 -121 -486 -109
rect -532 -697 -526 -121
rect -492 -697 -486 -121
rect -532 -709 -486 -697
rect 486 -121 532 -109
rect 486 -697 492 -121
rect 526 -697 532 -121
rect 486 -709 532 -697
rect 1504 -121 1550 -109
rect 1504 -697 1510 -121
rect 1544 -697 1550 -121
rect 1504 -709 1550 -697
rect 2522 -121 2568 -109
rect 2522 -697 2528 -121
rect 2562 -697 2568 -121
rect 2522 -709 2568 -697
rect 3540 -121 3586 -109
rect 3540 -697 3546 -121
rect 3580 -697 3586 -121
rect 3540 -709 3586 -697
rect 4558 -121 4604 -109
rect 4558 -697 4564 -121
rect 4598 -697 4604 -121
rect 4558 -709 4604 -697
rect 5576 -121 5622 -109
rect 5576 -697 5582 -121
rect 5616 -697 5622 -121
rect 5576 -709 5622 -697
rect -5334 -747 -4846 -741
rect -5334 -781 -5322 -747
rect -4858 -781 -4846 -747
rect -5334 -787 -4846 -781
rect -4316 -747 -3828 -741
rect -4316 -781 -4304 -747
rect -3840 -781 -3828 -747
rect -4316 -787 -3828 -781
rect -3298 -747 -2810 -741
rect -3298 -781 -3286 -747
rect -2822 -781 -2810 -747
rect -3298 -787 -2810 -781
rect -2280 -747 -1792 -741
rect -2280 -781 -2268 -747
rect -1804 -781 -1792 -747
rect -2280 -787 -1792 -781
rect -1262 -747 -774 -741
rect -1262 -781 -1250 -747
rect -786 -781 -774 -747
rect -1262 -787 -774 -781
rect -244 -747 244 -741
rect -244 -781 -232 -747
rect 232 -781 244 -747
rect -244 -787 244 -781
rect 774 -747 1262 -741
rect 774 -781 786 -747
rect 1250 -781 1262 -747
rect 774 -787 1262 -781
rect 1792 -747 2280 -741
rect 1792 -781 1804 -747
rect 2268 -781 2280 -747
rect 1792 -787 2280 -781
rect 2810 -747 3298 -741
rect 2810 -781 2822 -747
rect 3286 -781 3298 -747
rect 2810 -787 3298 -781
rect 3828 -747 4316 -741
rect 3828 -781 3840 -747
rect 4304 -781 4316 -747
rect 3828 -787 4316 -781
rect 4846 -747 5334 -741
rect 4846 -781 4858 -747
rect 5322 -781 5334 -747
rect 4846 -787 5334 -781
rect -5334 -855 -4846 -849
rect -5334 -889 -5322 -855
rect -4858 -889 -4846 -855
rect -5334 -895 -4846 -889
rect -4316 -855 -3828 -849
rect -4316 -889 -4304 -855
rect -3840 -889 -3828 -855
rect -4316 -895 -3828 -889
rect -3298 -855 -2810 -849
rect -3298 -889 -3286 -855
rect -2822 -889 -2810 -855
rect -3298 -895 -2810 -889
rect -2280 -855 -1792 -849
rect -2280 -889 -2268 -855
rect -1804 -889 -1792 -855
rect -2280 -895 -1792 -889
rect -1262 -855 -774 -849
rect -1262 -889 -1250 -855
rect -786 -889 -774 -855
rect -1262 -895 -774 -889
rect -244 -855 244 -849
rect -244 -889 -232 -855
rect 232 -889 244 -855
rect -244 -895 244 -889
rect 774 -855 1262 -849
rect 774 -889 786 -855
rect 1250 -889 1262 -855
rect 774 -895 1262 -889
rect 1792 -855 2280 -849
rect 1792 -889 1804 -855
rect 2268 -889 2280 -855
rect 1792 -895 2280 -889
rect 2810 -855 3298 -849
rect 2810 -889 2822 -855
rect 3286 -889 3298 -855
rect 2810 -895 3298 -889
rect 3828 -855 4316 -849
rect 3828 -889 3840 -855
rect 4304 -889 4316 -855
rect 3828 -895 4316 -889
rect 4846 -855 5334 -849
rect 4846 -889 4858 -855
rect 5322 -889 5334 -855
rect 4846 -895 5334 -889
rect -5622 -939 -5576 -927
rect -5622 -1515 -5616 -939
rect -5582 -1515 -5576 -939
rect -5622 -1527 -5576 -1515
rect -4604 -939 -4558 -927
rect -4604 -1515 -4598 -939
rect -4564 -1515 -4558 -939
rect -4604 -1527 -4558 -1515
rect -3586 -939 -3540 -927
rect -3586 -1515 -3580 -939
rect -3546 -1515 -3540 -939
rect -3586 -1527 -3540 -1515
rect -2568 -939 -2522 -927
rect -2568 -1515 -2562 -939
rect -2528 -1515 -2522 -939
rect -2568 -1527 -2522 -1515
rect -1550 -939 -1504 -927
rect -1550 -1515 -1544 -939
rect -1510 -1515 -1504 -939
rect -1550 -1527 -1504 -1515
rect -532 -939 -486 -927
rect -532 -1515 -526 -939
rect -492 -1515 -486 -939
rect -532 -1527 -486 -1515
rect 486 -939 532 -927
rect 486 -1515 492 -939
rect 526 -1515 532 -939
rect 486 -1527 532 -1515
rect 1504 -939 1550 -927
rect 1504 -1515 1510 -939
rect 1544 -1515 1550 -939
rect 1504 -1527 1550 -1515
rect 2522 -939 2568 -927
rect 2522 -1515 2528 -939
rect 2562 -1515 2568 -939
rect 2522 -1527 2568 -1515
rect 3540 -939 3586 -927
rect 3540 -1515 3546 -939
rect 3580 -1515 3586 -939
rect 3540 -1527 3586 -1515
rect 4558 -939 4604 -927
rect 4558 -1515 4564 -939
rect 4598 -1515 4604 -939
rect 4558 -1527 4604 -1515
rect 5576 -939 5622 -927
rect 5576 -1515 5582 -939
rect 5616 -1515 5622 -939
rect 5576 -1527 5622 -1515
rect -5334 -1565 -4846 -1559
rect -5334 -1599 -5322 -1565
rect -4858 -1599 -4846 -1565
rect -5334 -1605 -4846 -1599
rect -4316 -1565 -3828 -1559
rect -4316 -1599 -4304 -1565
rect -3840 -1599 -3828 -1565
rect -4316 -1605 -3828 -1599
rect -3298 -1565 -2810 -1559
rect -3298 -1599 -3286 -1565
rect -2822 -1599 -2810 -1565
rect -3298 -1605 -2810 -1599
rect -2280 -1565 -1792 -1559
rect -2280 -1599 -2268 -1565
rect -1804 -1599 -1792 -1565
rect -2280 -1605 -1792 -1599
rect -1262 -1565 -774 -1559
rect -1262 -1599 -1250 -1565
rect -786 -1599 -774 -1565
rect -1262 -1605 -774 -1599
rect -244 -1565 244 -1559
rect -244 -1599 -232 -1565
rect 232 -1599 244 -1565
rect -244 -1605 244 -1599
rect 774 -1565 1262 -1559
rect 774 -1599 786 -1565
rect 1250 -1599 1262 -1565
rect 774 -1605 1262 -1599
rect 1792 -1565 2280 -1559
rect 1792 -1599 1804 -1565
rect 2268 -1599 2280 -1565
rect 1792 -1605 2280 -1599
rect 2810 -1565 3298 -1559
rect 2810 -1599 2822 -1565
rect 3286 -1599 3298 -1565
rect 2810 -1605 3298 -1599
rect 3828 -1565 4316 -1559
rect 3828 -1599 3840 -1565
rect 4304 -1599 4316 -1565
rect 3828 -1605 4316 -1599
rect 4846 -1565 5334 -1559
rect 4846 -1599 4858 -1565
rect 5322 -1599 5334 -1565
rect 4846 -1605 5334 -1599
rect -5334 -1673 -4846 -1667
rect -5334 -1707 -5322 -1673
rect -4858 -1707 -4846 -1673
rect -5334 -1713 -4846 -1707
rect -4316 -1673 -3828 -1667
rect -4316 -1707 -4304 -1673
rect -3840 -1707 -3828 -1673
rect -4316 -1713 -3828 -1707
rect -3298 -1673 -2810 -1667
rect -3298 -1707 -3286 -1673
rect -2822 -1707 -2810 -1673
rect -3298 -1713 -2810 -1707
rect -2280 -1673 -1792 -1667
rect -2280 -1707 -2268 -1673
rect -1804 -1707 -1792 -1673
rect -2280 -1713 -1792 -1707
rect -1262 -1673 -774 -1667
rect -1262 -1707 -1250 -1673
rect -786 -1707 -774 -1673
rect -1262 -1713 -774 -1707
rect -244 -1673 244 -1667
rect -244 -1707 -232 -1673
rect 232 -1707 244 -1673
rect -244 -1713 244 -1707
rect 774 -1673 1262 -1667
rect 774 -1707 786 -1673
rect 1250 -1707 1262 -1673
rect 774 -1713 1262 -1707
rect 1792 -1673 2280 -1667
rect 1792 -1707 1804 -1673
rect 2268 -1707 2280 -1673
rect 1792 -1713 2280 -1707
rect 2810 -1673 3298 -1667
rect 2810 -1707 2822 -1673
rect 3286 -1707 3298 -1673
rect 2810 -1713 3298 -1707
rect 3828 -1673 4316 -1667
rect 3828 -1707 3840 -1673
rect 4304 -1707 4316 -1673
rect 3828 -1713 4316 -1707
rect 4846 -1673 5334 -1667
rect 4846 -1707 4858 -1673
rect 5322 -1707 5334 -1673
rect 4846 -1713 5334 -1707
rect -5622 -1757 -5576 -1745
rect -5622 -2333 -5616 -1757
rect -5582 -2333 -5576 -1757
rect -5622 -2345 -5576 -2333
rect -4604 -1757 -4558 -1745
rect -4604 -2333 -4598 -1757
rect -4564 -2333 -4558 -1757
rect -4604 -2345 -4558 -2333
rect -3586 -1757 -3540 -1745
rect -3586 -2333 -3580 -1757
rect -3546 -2333 -3540 -1757
rect -3586 -2345 -3540 -2333
rect -2568 -1757 -2522 -1745
rect -2568 -2333 -2562 -1757
rect -2528 -2333 -2522 -1757
rect -2568 -2345 -2522 -2333
rect -1550 -1757 -1504 -1745
rect -1550 -2333 -1544 -1757
rect -1510 -2333 -1504 -1757
rect -1550 -2345 -1504 -2333
rect -532 -1757 -486 -1745
rect -532 -2333 -526 -1757
rect -492 -2333 -486 -1757
rect -532 -2345 -486 -2333
rect 486 -1757 532 -1745
rect 486 -2333 492 -1757
rect 526 -2333 532 -1757
rect 486 -2345 532 -2333
rect 1504 -1757 1550 -1745
rect 1504 -2333 1510 -1757
rect 1544 -2333 1550 -1757
rect 1504 -2345 1550 -2333
rect 2522 -1757 2568 -1745
rect 2522 -2333 2528 -1757
rect 2562 -2333 2568 -1757
rect 2522 -2345 2568 -2333
rect 3540 -1757 3586 -1745
rect 3540 -2333 3546 -1757
rect 3580 -2333 3586 -1757
rect 3540 -2345 3586 -2333
rect 4558 -1757 4604 -1745
rect 4558 -2333 4564 -1757
rect 4598 -2333 4604 -1757
rect 4558 -2345 4604 -2333
rect 5576 -1757 5622 -1745
rect 5576 -2333 5582 -1757
rect 5616 -2333 5622 -1757
rect 5576 -2345 5622 -2333
rect -5334 -2383 -4846 -2377
rect -5334 -2417 -5322 -2383
rect -4858 -2417 -4846 -2383
rect -5334 -2423 -4846 -2417
rect -4316 -2383 -3828 -2377
rect -4316 -2417 -4304 -2383
rect -3840 -2417 -3828 -2383
rect -4316 -2423 -3828 -2417
rect -3298 -2383 -2810 -2377
rect -3298 -2417 -3286 -2383
rect -2822 -2417 -2810 -2383
rect -3298 -2423 -2810 -2417
rect -2280 -2383 -1792 -2377
rect -2280 -2417 -2268 -2383
rect -1804 -2417 -1792 -2383
rect -2280 -2423 -1792 -2417
rect -1262 -2383 -774 -2377
rect -1262 -2417 -1250 -2383
rect -786 -2417 -774 -2383
rect -1262 -2423 -774 -2417
rect -244 -2383 244 -2377
rect -244 -2417 -232 -2383
rect 232 -2417 244 -2383
rect -244 -2423 244 -2417
rect 774 -2383 1262 -2377
rect 774 -2417 786 -2383
rect 1250 -2417 1262 -2383
rect 774 -2423 1262 -2417
rect 1792 -2383 2280 -2377
rect 1792 -2417 1804 -2383
rect 2268 -2417 2280 -2383
rect 1792 -2423 2280 -2417
rect 2810 -2383 3298 -2377
rect 2810 -2417 2822 -2383
rect 3286 -2417 3298 -2383
rect 2810 -2423 3298 -2417
rect 3828 -2383 4316 -2377
rect 3828 -2417 3840 -2383
rect 4304 -2417 4316 -2383
rect 3828 -2423 4316 -2417
rect 4846 -2383 5334 -2377
rect 4846 -2417 4858 -2383
rect 5322 -2417 5334 -2383
rect 4846 -2423 5334 -2417
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string parameters w 3 l 4.8 m 6 nf 11 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
