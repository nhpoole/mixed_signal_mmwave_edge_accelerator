magic
tech sky130A
magscale 1 2
timestamp 1623661481
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 27 -17 61 17
<< locali >>
rect 885 325 935 493
rect 1053 325 1103 493
rect 1325 325 1375 425
rect 1493 325 1543 425
rect 885 291 1543 325
rect 85 215 365 257
rect 419 215 701 257
rect 1175 181 1231 291
rect 1293 215 1575 257
rect 1609 215 2001 257
rect 883 129 1231 181
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 31 359 81 527
rect 115 325 165 493
rect 199 359 249 527
rect 283 325 333 493
rect 367 359 417 527
rect 451 325 501 493
rect 535 359 585 527
rect 619 325 669 493
rect 703 359 851 527
rect 969 359 1019 527
rect 1137 359 1187 527
rect 1235 459 1627 493
rect 1235 359 1291 459
rect 1409 359 1459 459
rect 17 291 783 325
rect 1577 325 1627 459
rect 1661 359 1711 527
rect 1745 325 1795 493
rect 1829 359 1879 527
rect 1913 325 1975 493
rect 1577 291 1975 325
rect 17 181 51 291
rect 749 257 783 291
rect 749 215 1141 257
rect 17 129 341 181
rect 375 145 761 181
rect 375 95 425 145
rect 20 51 425 95
rect 459 17 493 111
rect 527 51 593 145
rect 627 17 661 111
rect 695 51 761 145
rect 812 95 849 167
rect 1265 147 1971 181
rect 1265 95 1299 147
rect 1401 145 1971 147
rect 812 51 1299 95
rect 1333 17 1367 111
rect 1401 51 1467 145
rect 1501 17 1535 111
rect 1569 51 1635 145
rect 1669 17 1703 111
rect 1737 51 1803 145
rect 1837 17 1871 111
rect 1905 51 1971 145
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< labels >>
rlabel locali s 419 215 701 257 6 A1_N
port 1 nsew signal input
rlabel locali s 85 215 365 257 6 A2_N
port 2 nsew signal input
rlabel locali s 1609 215 2001 257 6 B1
port 3 nsew signal input
rlabel locali s 1293 215 1575 257 6 B2
port 4 nsew signal input
rlabel locali s 1493 325 1543 425 6 Y
port 5 nsew signal output
rlabel locali s 1325 325 1375 425 6 Y
port 5 nsew signal output
rlabel locali s 1175 181 1231 291 6 Y
port 5 nsew signal output
rlabel locali s 1053 325 1103 493 6 Y
port 5 nsew signal output
rlabel locali s 885 325 935 493 6 Y
port 5 nsew signal output
rlabel locali s 885 291 1543 325 6 Y
port 5 nsew signal output
rlabel locali s 883 129 1231 181 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 2024 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 27 -17 61 17 8 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 2062 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 2024 592 6 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2024 544
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
