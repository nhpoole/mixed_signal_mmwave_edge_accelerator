magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< error_s >>
rect 1422 679 1458 1471
<< locali >>
rect 9430 7053 12418 7087
rect 3537 6790 3756 6824
rect 3722 6308 3756 6790
rect 5872 5639 12418 5673
rect 4584 4225 12418 4259
rect 4584 2811 12418 2845
rect 3519 2541 3704 2575
rect 3519 2176 3553 2541
rect 3386 2142 3553 2176
rect 4952 1397 12418 1431
rect 11878 -17 12418 17
<< metal1 >>
rect 12386 8458 12450 8510
rect 2700 7801 3271 7829
rect 9734 7751 9798 7803
rect 12386 7044 12450 7096
rect 7934 6337 7998 6389
rect 2616 6160 3419 6188
rect 2784 5912 3319 5940
rect 12386 5630 12450 5682
rect 2616 5372 3286 5400
rect 2700 5248 3419 5276
rect 3036 5124 3552 5152
rect 4700 4923 4764 4975
rect 1553 4308 2616 4336
rect 12386 4216 12450 4268
rect 383 4148 2868 4176
rect 4058 3493 4122 3545
rect 3036 3332 3419 3360
rect 2868 3084 3319 3112
rect 12386 2802 12450 2854
rect 3755 2284 3819 2336
rect 2868 2145 3271 2173
rect 4426 2111 4490 2163
rect 12386 1388 12450 1440
rect 3239 643 3303 695
rect 9410 681 9474 733
rect 12386 -26 12450 26
<< metal2 >>
rect -57 17699 -29 17727
rect 1539 4322 1567 6401
rect 369 1414 397 4162
rect 137 538 203 590
rect 2518 0 2546 8524
rect 2602 0 2630 8524
rect 2686 0 2714 8524
rect 2770 0 2798 8524
rect 2854 0 2882 8524
rect 2938 0 2966 8524
rect 3022 0 3050 8524
rect 12390 8460 12446 8508
rect 9766 7763 12502 7791
rect 12390 7046 12446 7094
rect 7966 6349 12502 6377
rect 12390 5632 12446 5680
rect 4732 4935 12502 4963
rect 12390 4218 12446 4266
rect 4062 3495 4118 3543
rect 12390 2804 12446 2852
rect 3759 2286 3815 2334
rect 4444 1571 4472 2137
rect 12390 1390 12446 1438
rect 9442 707 12502 721
rect 9428 693 12502 707
rect 3257 655 3285 683
rect 9428 141 9456 693
rect 12390 -24 12446 24
<< metal3 >>
rect 607 18333 705 18431
rect 1343 18333 1441 18431
rect 607 16919 705 17017
rect 1343 16919 1441 17017
rect 607 15505 705 15603
rect 1343 15505 1441 15603
rect 607 14091 705 14189
rect 1343 14091 1441 14189
rect 607 12677 705 12775
rect 1343 12677 1441 12775
rect 607 11263 705 11361
rect 1343 11263 1441 11361
rect 607 9849 705 9947
rect 1343 9849 1441 9947
rect 607 8435 705 8533
rect 1343 8435 1441 8533
rect 12369 8435 12467 8533
rect 607 7021 705 7119
rect 1343 7021 1441 7119
rect 12369 7021 12467 7119
rect 607 5607 705 5705
rect 1343 5607 1441 5705
rect 12369 5607 12467 5705
rect 12369 4193 12467 4291
rect 2784 3489 4090 3549
rect 12369 2779 12467 2877
rect 3036 2280 3787 2340
rect 2700 1541 4458 1601
rect -49 1365 49 1463
rect 12369 1365 12467 1463
rect 1836 855 3036 915
rect 2342 473 2952 533
rect 2868 111 9442 171
rect -49 -49 49 49
rect 12369 -49 12467 49
use dff_buf_array_0  dff_buf_array_0_0
timestamp 1624494425
transform 1 0 0 0 1 0
box -49 -49 2554 1471
use contact_9  contact_9_16
timestamp 1624494425
transform 1 0 1803 0 1 848
box 0 0 66 74
use contact_9  contact_9_15
timestamp 1624494425
transform 1 0 2309 0 1 466
box 0 0 66 74
use pand2_1  pand2_1_1
timestamp 1624494425
transform 1 0 3558 0 -1 2828
box -36 -17 1430 1471
use pinv_1  pinv_1_0
timestamp 1624494425
transform 1 0 3190 0 -1 2828
box -36 -17 404 1471
use contact_7  contact_7_22
timestamp 1624494425
transform 1 0 3242 0 1 636
box 0 0 58 66
use contact_8  contact_8_22
timestamp 1624494425
transform 1 0 3239 0 1 637
box 0 0 64 64
use contact_31  contact_31_7
timestamp 1624494425
transform 1 0 3003 0 1 848
box 0 0 66 74
use contact_31  contact_31_6
timestamp 1624494425
transform 1 0 2919 0 1 466
box 0 0 66 74
use contact_31  contact_31_4
timestamp 1624494425
transform 1 0 2835 0 1 104
box 0 0 66 74
use contact_7  contact_7_21
timestamp 1624494425
transform 1 0 9413 0 1 674
box 0 0 58 66
use contact_7  contact_7_20
timestamp 1624494425
transform 1 0 9413 0 1 674
box 0 0 58 66
use contact_8  contact_8_21
timestamp 1624494425
transform 1 0 9410 0 1 675
box 0 0 64 64
use contact_8  contact_8_20
timestamp 1624494425
transform 1 0 9410 0 1 675
box 0 0 64 64
use contact_31  contact_31_5
timestamp 1624494425
transform 1 0 9409 0 1 104
box 0 0 66 74
use contact_7  contact_7_11
timestamp 1624494425
transform 1 0 12389 0 1 1381
box 0 0 58 66
use contact_7  contact_7_10
timestamp 1624494425
transform 1 0 12389 0 1 -33
box 0 0 58 66
use contact_7  contact_7_9
timestamp 1624494425
transform 1 0 12389 0 1 1381
box 0 0 58 66
use contact_8  contact_8_11
timestamp 1624494425
transform 1 0 12386 0 1 1382
box 0 0 64 64
use contact_8  contact_8_10
timestamp 1624494425
transform 1 0 12386 0 1 -32
box 0 0 64 64
use contact_8  contact_8_9
timestamp 1624494425
transform 1 0 12386 0 1 1382
box 0 0 64 64
use contact_9  contact_9_11
timestamp 1624494425
transform 1 0 12385 0 1 1377
box 0 0 66 74
use contact_9  contact_9_10
timestamp 1624494425
transform 1 0 12385 0 1 -37
box 0 0 66 74
use contact_9  contact_9_9
timestamp 1624494425
transform 1 0 12385 0 1 1377
box 0 0 66 74
use pdriver_7  pdriver_7_0
timestamp 1624494425
transform 1 0 3190 0 1 0
box -36 -17 8724 1471
use contact_31  contact_31_1
timestamp 1624494425
transform 1 0 2667 0 1 1534
box 0 0 66 74
use contact_8  contact_8_19
timestamp 1624494425
transform 1 0 2836 0 1 2127
box 0 0 64 64
use contact_31  contact_31_3
timestamp 1624494425
transform 1 0 3003 0 1 2273
box 0 0 66 74
use contact_9  contact_9_13
timestamp 1624494425
transform 1 0 3754 0 1 2273
box 0 0 66 74
use contact_9  contact_9_14
timestamp 1624494425
transform 1 0 3754 0 1 2273
box 0 0 66 74
use contact_8  contact_8_17
timestamp 1624494425
transform 1 0 3755 0 1 2278
box 0 0 64 64
use contact_8  contact_8_18
timestamp 1624494425
transform 1 0 3755 0 1 2278
box 0 0 64 64
use contact_7  contact_7_17
timestamp 1624494425
transform 1 0 3758 0 1 2277
box 0 0 58 66
use contact_7  contact_7_18
timestamp 1624494425
transform 1 0 3758 0 1 2277
box 0 0 58 66
use contact_7  contact_7_19
timestamp 1624494425
transform 1 0 3242 0 1 2126
box 0 0 58 66
use pand2_1  pand2_1_0
timestamp 1624494425
transform 1 0 3190 0 1 2828
box -36 -17 1430 1471
use contact_31  contact_31_2
timestamp 1624494425
transform 1 0 4425 0 1 1534
box 0 0 66 74
use contact_8  contact_8_16
timestamp 1624494425
transform 1 0 4426 0 1 2105
box 0 0 64 64
use contact_7  contact_7_16
timestamp 1624494425
transform 1 0 4429 0 1 2104
box 0 0 58 66
use contact_9  contact_9_6
timestamp 1624494425
transform 1 0 12385 0 1 2791
box 0 0 66 74
use contact_9  contact_9_8
timestamp 1624494425
transform 1 0 12385 0 1 2791
box 0 0 66 74
use contact_8  contact_8_6
timestamp 1624494425
transform 1 0 12386 0 1 2796
box 0 0 64 64
use contact_8  contact_8_8
timestamp 1624494425
transform 1 0 12386 0 1 2796
box 0 0 64 64
use contact_7  contact_7_6
timestamp 1624494425
transform 1 0 12389 0 1 2795
box 0 0 58 66
use contact_7  contact_7_8
timestamp 1624494425
transform 1 0 12389 0 1 2795
box 0 0 58 66
use contact_8  contact_8_26
timestamp 1624494425
transform 1 0 2584 0 1 4290
box 0 0 64 64
use contact_8  contact_8_27
timestamp 1624494425
transform 1 0 1521 0 1 4290
box 0 0 64 64
use contact_8  contact_8_35
timestamp 1624494425
transform 1 0 351 0 1 4130
box 0 0 64 64
use contact_31  contact_31_0
timestamp 1624494425
transform 1 0 2751 0 1 3482
box 0 0 66 74
use contact_8  contact_8_15
timestamp 1624494425
transform 1 0 2836 0 1 3066
box 0 0 64 64
use contact_8  contact_8_14
timestamp 1624494425
transform 1 0 3004 0 1 3314
box 0 0 64 64
use contact_7  contact_7_14
timestamp 1624494425
transform 1 0 3390 0 1 3313
box 0 0 58 66
use contact_7  contact_7_15
timestamp 1624494425
transform 1 0 3290 0 1 3065
box 0 0 58 66
use contact_9  contact_9_12
timestamp 1624494425
transform 1 0 4057 0 1 3482
box 0 0 66 74
use contact_8  contact_8_12
timestamp 1624494425
transform 1 0 4058 0 1 3487
box 0 0 64 64
use contact_8  contact_8_13
timestamp 1624494425
transform 1 0 4058 0 1 3487
box 0 0 64 64
use contact_7  contact_7_12
timestamp 1624494425
transform 1 0 4061 0 1 3486
box 0 0 58 66
use contact_7  contact_7_13
timestamp 1624494425
transform 1 0 4061 0 1 3486
box 0 0 58 66
use contact_8  contact_8_34
timestamp 1624494425
transform 1 0 2836 0 1 4130
box 0 0 64 64
use pand3_0  pand3_0_0
timestamp 1624494425
transform 1 0 3190 0 -1 5656
box -36 -17 2718 1471
use contact_9  contact_9_5
timestamp 1624494425
transform 1 0 12385 0 1 4205
box 0 0 66 74
use contact_9  contact_9_7
timestamp 1624494425
transform 1 0 12385 0 1 4205
box 0 0 66 74
use contact_8  contact_8_5
timestamp 1624494425
transform 1 0 12386 0 1 4210
box 0 0 64 64
use contact_8  contact_8_7
timestamp 1624494425
transform 1 0 12386 0 1 4210
box 0 0 64 64
use contact_7  contact_7_5
timestamp 1624494425
transform 1 0 12389 0 1 4209
box 0 0 58 66
use contact_7  contact_7_7
timestamp 1624494425
transform 1 0 12389 0 1 4209
box 0 0 58 66
use contact_8  contact_8_31
timestamp 1624494425
transform 1 0 2584 0 1 5354
box 0 0 64 64
use contact_8  contact_8_30
timestamp 1624494425
transform 1 0 2668 0 1 5230
box 0 0 64 64
use contact_8  contact_8_25
timestamp 1624494425
transform 1 0 2752 0 1 5894
box 0 0 64 64
use pnand2_1  pnand2_1_0
timestamp 1624494425
transform 1 0 3190 0 1 5656
box -36 -17 504 1471
use contact_7  contact_7_29
timestamp 1624494425
transform 1 0 3257 0 1 5353
box 0 0 58 66
use contact_7  contact_7_28
timestamp 1624494425
transform 1 0 3390 0 1 5229
box 0 0 58 66
use contact_7  contact_7_27
timestamp 1624494425
transform 1 0 3523 0 1 5105
box 0 0 58 66
use contact_7  contact_7_26
timestamp 1624494425
transform 1 0 4703 0 1 4916
box 0 0 58 66
use contact_7  contact_7_25
timestamp 1624494425
transform 1 0 3290 0 1 5893
box 0 0 58 66
use contact_8  contact_8_29
timestamp 1624494425
transform 1 0 3004 0 1 5106
box 0 0 64 64
use contact_8  contact_8_28
timestamp 1624494425
transform 1 0 4700 0 1 4917
box 0 0 64 64
use pdriver_6  pdriver_6_0
timestamp 1624494425
transform 1 0 3658 0 1 5656
box -36 -17 5808 1471
use contact_9  contact_9_2
timestamp 1624494425
transform 1 0 12385 0 1 5619
box 0 0 66 74
use contact_9  contact_9_4
timestamp 1624494425
transform 1 0 12385 0 1 5619
box 0 0 66 74
use contact_8  contact_8_2
timestamp 1624494425
transform 1 0 12386 0 1 5624
box 0 0 64 64
use contact_8  contact_8_4
timestamp 1624494425
transform 1 0 12386 0 1 5624
box 0 0 64 64
use contact_7  contact_7_2
timestamp 1624494425
transform 1 0 12389 0 1 5623
box 0 0 58 66
use contact_7  contact_7_4
timestamp 1624494425
transform 1 0 12389 0 1 5623
box 0 0 58 66
use contact_8  contact_8_23
timestamp 1624494425
transform 1 0 7934 0 1 6331
box 0 0 64 64
use contact_8  contact_8_24
timestamp 1624494425
transform 1 0 2584 0 1 6142
box 0 0 64 64
use contact_7  contact_7_23
timestamp 1624494425
transform 1 0 7937 0 1 6330
box 0 0 58 66
use contact_7  contact_7_24
timestamp 1624494425
transform 1 0 3390 0 1 6141
box 0 0 58 66
use contact_9  contact_9_1
timestamp 1624494425
transform 1 0 12385 0 1 7033
box 0 0 66 74
use contact_9  contact_9_3
timestamp 1624494425
transform 1 0 12385 0 1 7033
box 0 0 66 74
use contact_8  contact_8_1
timestamp 1624494425
transform 1 0 12386 0 1 7038
box 0 0 64 64
use contact_8  contact_8_3
timestamp 1624494425
transform 1 0 12386 0 1 7038
box 0 0 64 64
use contact_7  contact_7_1
timestamp 1624494425
transform 1 0 12389 0 1 7037
box 0 0 58 66
use contact_7  contact_7_3
timestamp 1624494425
transform 1 0 12389 0 1 7037
box 0 0 58 66
use pdriver_3  pdriver_3_0
timestamp 1624494425
transform 1 0 3190 0 -1 8484
box -36 -17 9264 1471
use contact_7  contact_7_31
timestamp 1624494425
transform 1 0 3242 0 1 7782
box 0 0 58 66
use contact_7  contact_7_30
timestamp 1624494425
transform 1 0 9737 0 1 7744
box 0 0 58 66
use contact_7  contact_7_0
timestamp 1624494425
transform 1 0 12389 0 1 8451
box 0 0 58 66
use contact_8  contact_8_33
timestamp 1624494425
transform 1 0 2668 0 1 7783
box 0 0 64 64
use contact_8  contact_8_32
timestamp 1624494425
transform 1 0 9734 0 1 7745
box 0 0 64 64
use contact_8  contact_8_0
timestamp 1624494425
transform 1 0 12386 0 1 8452
box 0 0 64 64
use contact_9  contact_9_0
timestamp 1624494425
transform 1 0 12385 0 1 8447
box 0 0 66 74
use delay_chain  delay_chain_0
timestamp 1624494425
transform 1 0 0 0 -1 18382
box -75 -49 1876 12783
<< labels >>
rlabel metal2 s 137 538 203 590 4 csb
rlabel metal2 s 9766 7763 12502 7791 4 wl_en
rlabel metal2 s 4732 4935 12502 4963 4 s_en
rlabel metal2 s -57 17699 -29 17727 4 rbl_bl
rlabel metal2 s 7966 6349 12502 6377 4 p_en_bar
rlabel metal2 s 3257 655 3285 683 4 clk
rlabel metal2 s 9442 693 12502 721 4 clk_buf
rlabel metal3 s 1343 5607 1441 5705 4 vdd
rlabel metal3 s 607 8435 705 8533 4 vdd
rlabel metal3 s 607 16919 705 17017 4 vdd
rlabel metal3 s 1343 16919 1441 17017 4 vdd
rlabel metal3 s 607 11263 705 11361 4 vdd
rlabel metal3 s 12369 4193 12467 4291 4 vdd
rlabel metal3 s 607 14091 705 14189 4 vdd
rlabel metal3 s 1343 14091 1441 14189 4 vdd
rlabel metal3 s 1343 11263 1441 11361 4 vdd
rlabel metal3 s -49 1365 49 1463 4 vdd
rlabel metal3 s 607 5607 705 5705 4 vdd
rlabel metal3 s 1343 8435 1441 8533 4 vdd
rlabel metal3 s 12369 7021 12467 7119 4 vdd
rlabel metal3 s 12369 1365 12467 1463 4 vdd
rlabel metal3 s 1343 7021 1441 7119 4 gnd
rlabel metal3 s 1343 15505 1441 15603 4 gnd
rlabel metal3 s 12369 2779 12467 2877 4 gnd
rlabel metal3 s 607 9849 705 9947 4 gnd
rlabel metal3 s 1343 9849 1441 9947 4 gnd
rlabel metal3 s 12369 -49 12467 49 4 gnd
rlabel metal3 s 12369 8435 12467 8533 4 gnd
rlabel metal3 s 1343 18333 1441 18431 4 gnd
rlabel metal3 s 607 15505 705 15603 4 gnd
rlabel metal3 s 607 7021 705 7119 4 gnd
rlabel metal3 s 607 18333 705 18431 4 gnd
rlabel metal3 s 607 12677 705 12775 4 gnd
rlabel metal3 s 1343 12677 1441 12775 4 gnd
rlabel metal3 s -49 -49 49 49 4 gnd
rlabel metal3 s 12369 5607 12467 5705 4 gnd
<< properties >>
string FIXED_BBOX 0 0 12502 18542
<< end >>
