magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< error_s >>
rect 182 102305 224 102331
rect 544 102322 586 102331
rect 174 102293 182 102305
rect 186 102297 220 102305
rect 186 102290 190 102297
rect 216 102290 220 102297
rect 224 102293 232 102305
rect 170 102289 236 102290
rect 120 102275 170 102277
rect 76 102271 130 102275
rect 110 102266 130 102271
rect 60 102241 67 102251
rect 76 102241 77 102261
rect 96 102232 99 102266
rect 109 102241 110 102261
rect 119 102241 126 102251
rect 76 102225 92 102231
rect 94 102225 110 102231
rect 170 102225 172 102275
rect 213 102177 224 102215
rect 251 102177 287 102205
rect 288 102177 292 102305
rect 439 102288 444 102322
rect 468 102288 473 102322
rect 511 102305 586 102322
rect 476 102251 480 102305
rect 511 102288 582 102305
rect 586 102293 594 102305
rect 544 102281 548 102288
rect 12 102172 62 102174
rect 28 102163 59 102171
rect 62 102163 64 102172
rect 251 102171 263 102177
rect 28 102155 64 102163
rect 127 102163 161 102171
rect 127 102156 182 102163
rect 127 102155 161 102156
rect 59 102139 64 102155
rect 253 102143 263 102171
rect 273 102143 293 102177
rect 476 102171 480 102239
rect 544 102201 548 102251
rect 544 102161 553 102189
rect 612 102174 624 102175
rect 599 102172 649 102174
rect 612 102171 624 102172
rect 607 102163 632 102171
rect 28 102131 64 102139
rect 127 102138 161 102139
rect 127 102131 182 102138
rect 62 102122 64 102131
rect 120 102069 170 102071
rect 76 102063 92 102069
rect 94 102063 110 102069
rect 76 102053 99 102062
rect 60 102043 67 102053
rect 76 102033 77 102053
rect 96 102028 99 102053
rect 109 102033 110 102053
rect 119 102043 126 102053
rect 76 102019 110 102023
rect 170 102019 172 102069
rect 182 102013 224 102014
rect 186 101989 220 102006
rect 223 101989 257 102006
rect 182 101972 257 101989
rect 182 101971 224 101972
rect 160 101965 246 101971
rect 288 101965 292 102143
rect 476 102093 480 102161
rect 485 102117 495 102151
rect 505 102123 525 102151
rect 505 102117 519 102123
rect 544 102117 555 102161
rect 586 102156 641 102163
rect 607 102155 641 102156
rect 616 102139 641 102155
rect 607 102138 641 102139
rect 586 102131 641 102138
rect 612 102123 632 102131
rect 612 102119 624 102123
rect 649 102122 651 102172
rect 485 102093 492 102117
rect 476 102013 480 102081
rect 544 102043 548 102093
rect 544 102008 548 102013
rect 295 101972 300 102006
rect 324 101972 329 102006
rect 544 102004 582 102008
rect 544 101989 552 102004
rect 578 101989 582 102004
rect 544 101971 586 101989
rect 522 101965 608 101971
rect 182 101949 224 101965
rect 544 101949 586 101965
rect 17 101935 67 101937
rect 119 101935 169 101937
rect 186 101935 220 101949
rect 548 101935 582 101949
rect 599 101935 649 101937
rect 42 101893 59 101927
rect 67 101885 69 101935
rect 160 101927 246 101935
rect 522 101927 608 101935
rect 76 101893 110 101927
rect 127 101893 144 101927
rect 152 101893 161 101927
rect 162 101925 195 101927
rect 224 101925 244 101927
rect 162 101893 244 101925
rect 524 101925 548 101927
rect 573 101925 582 101927
rect 586 101925 606 101927
rect 160 101885 246 101893
rect 186 101869 220 101885
rect 182 101855 224 101856
rect 160 101849 182 101855
rect 224 101849 246 101855
rect 186 101814 220 101848
rect 223 101814 257 101848
rect 120 101801 170 101803
rect 76 101797 130 101801
rect 110 101792 130 101797
rect 60 101767 67 101777
rect 76 101767 77 101787
rect 96 101758 99 101792
rect 109 101767 110 101787
rect 119 101767 126 101777
rect 76 101751 92 101757
rect 94 101751 110 101757
rect 170 101751 172 101801
rect 186 101735 190 101769
rect 216 101735 220 101769
rect 288 101735 292 101923
rect 476 101855 480 101923
rect 524 101893 606 101925
rect 607 101893 616 101927
rect 522 101885 608 101893
rect 649 101885 651 101935
rect 548 101869 582 101885
rect 522 101850 548 101855
rect 522 101849 582 101850
rect 586 101849 608 101855
rect 295 101814 300 101848
rect 324 101814 329 101848
rect 544 101846 582 101849
rect 378 101809 450 101817
rect 428 101779 430 101795
rect 400 101771 430 101779
rect 476 101777 480 101845
rect 544 101816 552 101846
rect 578 101816 582 101846
rect 544 101807 548 101816
rect 400 101767 436 101771
rect 400 101737 408 101767
rect 420 101737 436 101767
rect 544 101769 548 101777
rect 12 101698 62 101700
rect 28 101689 59 101697
rect 62 101689 64 101698
rect 28 101681 64 101689
rect 127 101689 158 101697
rect 127 101682 182 101689
rect 215 101687 224 101715
rect 127 101681 161 101682
rect 59 101665 64 101681
rect 158 101665 161 101681
rect 28 101657 64 101665
rect 127 101664 161 101665
rect 127 101657 182 101664
rect 62 101648 64 101657
rect 213 101649 224 101687
rect 282 101677 292 101735
rect 296 101729 368 101737
rect 319 101699 346 101710
rect 318 101686 324 101699
rect 346 101686 348 101699
rect 428 101690 430 101737
rect 443 101727 450 101729
rect 476 101697 480 101765
rect 544 101735 552 101769
rect 578 101735 582 101769
rect 481 101703 517 101731
rect 481 101697 495 101703
rect 367 101686 380 101690
rect 251 101643 263 101677
rect 273 101643 293 101677
rect 295 101662 324 101686
rect 303 101652 316 101662
rect 318 101646 324 101662
rect 333 101662 380 101686
rect 333 101652 353 101662
rect 367 101656 380 101662
rect 396 101656 408 101690
rect 420 101656 436 101690
rect 120 101595 170 101597
rect 76 101589 92 101595
rect 94 101589 110 101595
rect 76 101579 99 101588
rect 60 101569 67 101579
rect 76 101559 77 101579
rect 96 101554 99 101579
rect 109 101559 110 101579
rect 119 101569 126 101579
rect 76 101545 110 101549
rect 170 101545 172 101595
rect 186 101577 190 101611
rect 216 101577 220 101611
rect 186 101500 220 101534
rect 282 101531 292 101643
rect 318 101636 335 101646
rect 318 101567 324 101636
rect 346 101567 348 101652
rect 428 101609 430 101656
rect 476 101619 480 101687
rect 485 101669 495 101697
rect 505 101697 519 101703
rect 544 101697 555 101735
rect 505 101669 525 101697
rect 544 101669 553 101697
rect 544 101649 548 101669
rect 579 101628 582 101718
rect 612 101700 624 101701
rect 599 101698 649 101700
rect 612 101697 624 101698
rect 610 101690 632 101697
rect 607 101689 632 101690
rect 586 101682 644 101689
rect 607 101681 644 101682
rect 607 101665 610 101681
rect 616 101665 644 101681
rect 607 101664 644 101665
rect 586 101657 644 101664
rect 607 101656 610 101657
rect 612 101649 632 101657
rect 612 101645 624 101649
rect 649 101648 651 101698
rect 544 101611 548 101619
rect 400 101579 408 101609
rect 420 101579 436 101609
rect 400 101575 436 101579
rect 400 101567 430 101575
rect 428 101551 430 101567
rect 476 101539 480 101607
rect 544 101577 552 101611
rect 578 101577 582 101611
rect 544 101569 548 101577
rect 544 101539 586 101540
rect 288 101499 292 101531
rect 296 101529 368 101537
rect 378 101529 450 101537
rect 544 101532 548 101539
rect 439 101501 444 101529
rect 120 101485 170 101487
rect 76 101481 130 101485
rect 110 101476 130 101481
rect 60 101451 67 101461
rect 76 101451 77 101471
rect 96 101442 99 101476
rect 109 101451 110 101471
rect 119 101451 126 101461
rect 76 101435 92 101441
rect 94 101435 110 101441
rect 170 101435 172 101485
rect 186 101419 190 101453
rect 216 101419 220 101453
rect 213 101387 224 101419
rect 282 101415 292 101499
rect 296 101493 368 101501
rect 378 101493 450 101501
rect 468 101498 473 101532
rect 428 101463 430 101479
rect 251 101387 292 101415
rect 318 101394 324 101463
rect 12 101382 62 101384
rect 28 101373 59 101381
rect 62 101373 64 101382
rect 251 101381 263 101387
rect 28 101365 64 101373
rect 127 101373 158 101381
rect 127 101366 182 101373
rect 127 101365 161 101366
rect 59 101349 64 101365
rect 158 101349 161 101365
rect 253 101353 263 101381
rect 273 101353 293 101387
rect 318 101384 335 101394
rect 303 101368 316 101378
rect 318 101368 324 101384
rect 346 101378 348 101463
rect 400 101455 430 101463
rect 476 101461 480 101529
rect 511 101498 582 101532
rect 544 101491 548 101498
rect 400 101451 436 101455
rect 400 101421 408 101451
rect 420 101421 436 101451
rect 544 101453 548 101461
rect 28 101341 64 101349
rect 127 101348 161 101349
rect 127 101341 182 101348
rect 62 101332 64 101341
rect 282 101295 292 101353
rect 295 101344 324 101368
rect 333 101368 353 101378
rect 428 101374 430 101421
rect 476 101381 480 101449
rect 544 101419 552 101453
rect 578 101419 582 101453
rect 544 101411 548 101419
rect 367 101368 380 101374
rect 333 101344 380 101368
rect 318 101331 324 101344
rect 346 101331 348 101344
rect 367 101340 380 101344
rect 396 101340 408 101374
rect 420 101340 436 101374
rect 544 101371 553 101399
rect 319 101320 346 101331
rect 120 101279 170 101281
rect 76 101273 92 101279
rect 94 101273 110 101279
rect 76 101263 99 101272
rect 60 101253 67 101263
rect 76 101243 77 101263
rect 96 101238 99 101263
rect 109 101243 110 101263
rect 119 101253 126 101263
rect 76 101229 110 101233
rect 170 101229 172 101279
rect 186 101261 190 101295
rect 216 101261 220 101295
rect 182 101223 224 101224
rect 186 101199 220 101216
rect 223 101199 257 101216
rect 182 101182 257 101199
rect 182 101181 224 101182
rect 160 101175 246 101181
rect 288 101175 292 101295
rect 296 101293 368 101301
rect 428 101293 430 101340
rect 476 101303 480 101371
rect 485 101327 495 101361
rect 505 101333 525 101361
rect 505 101327 519 101333
rect 544 101327 555 101371
rect 485 101303 492 101327
rect 579 101312 582 101402
rect 612 101384 624 101385
rect 599 101382 649 101384
rect 612 101381 624 101382
rect 610 101374 632 101381
rect 607 101373 632 101374
rect 586 101366 644 101373
rect 607 101365 644 101366
rect 607 101349 610 101365
rect 616 101349 644 101365
rect 607 101348 644 101349
rect 586 101341 644 101348
rect 607 101340 610 101341
rect 612 101333 632 101341
rect 612 101329 624 101333
rect 649 101332 651 101382
rect 544 101295 548 101303
rect 400 101263 408 101293
rect 420 101263 436 101293
rect 400 101259 436 101263
rect 400 101251 430 101259
rect 428 101235 430 101251
rect 476 101223 480 101291
rect 544 101261 552 101295
rect 578 101261 582 101295
rect 544 101253 548 101261
rect 295 101182 300 101216
rect 324 101182 329 101216
rect 378 101213 450 101221
rect 544 101218 548 101223
rect 544 101214 582 101218
rect 544 101199 552 101214
rect 578 101199 582 101214
rect 544 101181 586 101199
rect 522 101175 608 101181
rect 182 101159 224 101175
rect 544 101159 586 101175
rect 17 101145 67 101147
rect 119 101145 169 101147
rect 186 101145 220 101159
rect 548 101145 582 101159
rect 599 101145 649 101147
rect 42 101103 59 101137
rect 67 101095 69 101145
rect 160 101137 246 101145
rect 522 101137 608 101145
rect 76 101103 110 101137
rect 127 101103 144 101137
rect 152 101103 161 101137
rect 162 101135 195 101137
rect 224 101135 244 101137
rect 162 101103 244 101135
rect 524 101135 548 101137
rect 573 101135 582 101137
rect 586 101135 606 101137
rect 160 101095 246 101103
rect 186 101079 220 101095
rect 182 101065 224 101066
rect 160 101059 182 101065
rect 224 101059 246 101065
rect 186 101024 220 101058
rect 223 101024 257 101058
rect 120 101011 170 101013
rect 76 101007 130 101011
rect 110 101002 130 101007
rect 60 100977 67 100987
rect 76 100977 77 100997
rect 96 100968 99 101002
rect 109 100977 110 100997
rect 119 100977 126 100987
rect 76 100961 92 100967
rect 94 100961 110 100967
rect 170 100961 172 101011
rect 186 100945 190 100979
rect 216 100945 220 100979
rect 288 100945 292 101133
rect 476 101065 480 101133
rect 524 101103 606 101135
rect 607 101103 616 101137
rect 522 101095 608 101103
rect 649 101095 651 101145
rect 548 101079 582 101095
rect 522 101060 548 101065
rect 522 101059 582 101060
rect 586 101059 608 101065
rect 295 101024 300 101058
rect 324 101024 329 101058
rect 544 101056 582 101059
rect 378 101019 450 101027
rect 428 100989 430 101005
rect 400 100981 430 100989
rect 476 100987 480 101055
rect 544 101026 552 101056
rect 578 101026 582 101056
rect 544 101017 548 101026
rect 400 100977 436 100981
rect 400 100947 408 100977
rect 420 100947 436 100977
rect 544 100979 548 100987
rect 12 100908 62 100910
rect 28 100899 59 100907
rect 62 100899 64 100908
rect 28 100891 64 100899
rect 127 100899 158 100907
rect 127 100892 182 100899
rect 215 100897 224 100925
rect 127 100891 161 100892
rect 59 100875 64 100891
rect 158 100875 161 100891
rect 28 100867 64 100875
rect 127 100874 161 100875
rect 127 100867 182 100874
rect 62 100858 64 100867
rect 213 100859 224 100897
rect 282 100887 292 100945
rect 296 100939 368 100947
rect 319 100909 346 100920
rect 318 100896 324 100909
rect 346 100896 348 100909
rect 428 100900 430 100947
rect 443 100937 450 100939
rect 476 100907 480 100975
rect 544 100945 552 100979
rect 578 100945 582 100979
rect 481 100913 517 100941
rect 481 100907 495 100913
rect 367 100896 380 100900
rect 251 100853 263 100887
rect 273 100853 293 100887
rect 295 100872 324 100896
rect 303 100862 316 100872
rect 318 100856 324 100872
rect 333 100872 380 100896
rect 333 100862 353 100872
rect 367 100866 380 100872
rect 396 100866 408 100900
rect 420 100866 436 100900
rect 120 100805 170 100807
rect 76 100799 92 100805
rect 94 100799 110 100805
rect 76 100789 99 100798
rect 60 100779 67 100789
rect 76 100769 77 100789
rect 96 100764 99 100789
rect 109 100769 110 100789
rect 119 100779 126 100789
rect 76 100755 110 100759
rect 170 100755 172 100805
rect 186 100787 190 100821
rect 216 100787 220 100821
rect 186 100710 220 100744
rect 282 100741 292 100853
rect 318 100846 335 100856
rect 318 100777 324 100846
rect 346 100777 348 100862
rect 428 100819 430 100866
rect 476 100829 480 100897
rect 485 100879 495 100907
rect 505 100907 519 100913
rect 544 100907 555 100945
rect 505 100879 525 100907
rect 544 100879 553 100907
rect 544 100859 548 100879
rect 579 100838 582 100928
rect 612 100910 624 100911
rect 599 100908 649 100910
rect 612 100907 624 100908
rect 610 100900 632 100907
rect 607 100899 632 100900
rect 586 100892 644 100899
rect 607 100891 644 100892
rect 607 100875 610 100891
rect 616 100875 644 100891
rect 607 100874 644 100875
rect 586 100867 644 100874
rect 607 100866 610 100867
rect 612 100859 632 100867
rect 612 100855 624 100859
rect 649 100858 651 100908
rect 544 100821 548 100829
rect 400 100789 408 100819
rect 420 100789 436 100819
rect 400 100785 436 100789
rect 400 100777 430 100785
rect 428 100761 430 100777
rect 476 100749 480 100800
rect 544 100787 552 100821
rect 578 100787 582 100821
rect 544 100779 548 100787
rect 544 100749 586 100750
rect 288 100709 292 100741
rect 296 100739 368 100747
rect 378 100739 450 100747
rect 544 100742 548 100749
rect 439 100711 444 100739
rect 120 100695 170 100697
rect 76 100691 130 100695
rect 110 100686 130 100691
rect 60 100661 67 100671
rect 76 100661 77 100681
rect 96 100652 99 100686
rect 109 100661 110 100681
rect 119 100661 126 100671
rect 76 100645 92 100651
rect 94 100645 110 100651
rect 170 100645 172 100695
rect 186 100629 190 100663
rect 216 100629 220 100663
rect 213 100597 224 100629
rect 282 100625 292 100709
rect 296 100703 368 100711
rect 378 100703 450 100711
rect 468 100708 473 100742
rect 428 100673 430 100689
rect 251 100597 292 100625
rect 318 100604 324 100673
rect 12 100592 62 100594
rect 28 100583 59 100591
rect 62 100583 64 100592
rect 251 100591 263 100597
rect 28 100575 64 100583
rect 127 100583 158 100591
rect 127 100576 182 100583
rect 127 100575 161 100576
rect 59 100559 64 100575
rect 158 100559 161 100575
rect 253 100563 263 100591
rect 273 100563 293 100597
rect 318 100594 335 100604
rect 303 100578 316 100588
rect 318 100578 324 100594
rect 346 100588 348 100673
rect 400 100665 430 100673
rect 476 100671 480 100739
rect 511 100708 582 100742
rect 544 100701 548 100708
rect 400 100661 436 100665
rect 400 100631 408 100661
rect 420 100631 436 100661
rect 544 100663 548 100671
rect 28 100551 64 100559
rect 127 100558 161 100559
rect 127 100551 182 100558
rect 62 100542 64 100551
rect 282 100505 292 100563
rect 295 100554 324 100578
rect 333 100578 353 100588
rect 428 100584 430 100631
rect 476 100591 480 100659
rect 544 100629 552 100663
rect 578 100629 582 100663
rect 544 100621 548 100629
rect 367 100578 380 100584
rect 333 100554 380 100578
rect 318 100541 324 100554
rect 346 100541 348 100554
rect 367 100550 380 100554
rect 396 100550 408 100584
rect 420 100550 436 100584
rect 544 100581 553 100609
rect 319 100530 346 100541
rect 120 100489 170 100491
rect 76 100483 92 100489
rect 94 100483 110 100489
rect 76 100473 99 100482
rect 60 100463 67 100473
rect 76 100453 77 100473
rect 96 100448 99 100473
rect 109 100453 110 100473
rect 119 100463 126 100473
rect 76 100439 110 100443
rect 170 100439 172 100489
rect 186 100471 190 100505
rect 216 100471 220 100505
rect 182 100433 224 100434
rect 186 100409 220 100426
rect 223 100409 257 100426
rect 182 100392 257 100409
rect 182 100391 224 100392
rect 160 100385 246 100391
rect 288 100385 292 100505
rect 296 100503 368 100511
rect 428 100503 430 100550
rect 476 100513 480 100581
rect 485 100537 495 100571
rect 505 100543 525 100571
rect 505 100537 519 100543
rect 544 100537 555 100581
rect 485 100513 492 100537
rect 579 100522 582 100612
rect 612 100594 624 100595
rect 599 100592 649 100594
rect 612 100591 624 100592
rect 610 100584 632 100591
rect 607 100583 632 100584
rect 586 100576 644 100583
rect 607 100575 644 100576
rect 607 100559 610 100575
rect 616 100559 644 100575
rect 607 100558 644 100559
rect 586 100551 644 100558
rect 607 100550 610 100551
rect 612 100543 632 100551
rect 612 100539 624 100543
rect 649 100542 651 100592
rect 544 100505 548 100513
rect 400 100473 408 100503
rect 420 100473 436 100503
rect 400 100469 436 100473
rect 400 100461 430 100469
rect 428 100445 430 100461
rect 476 100433 480 100501
rect 544 100471 552 100505
rect 578 100471 582 100505
rect 544 100463 548 100471
rect 295 100392 300 100426
rect 324 100392 329 100426
rect 378 100423 450 100431
rect 544 100428 548 100433
rect 544 100424 582 100428
rect 544 100409 552 100424
rect 578 100409 582 100424
rect 544 100391 586 100409
rect 522 100385 608 100391
rect 182 100369 224 100385
rect 544 100369 586 100385
rect 17 100355 67 100357
rect 119 100355 169 100357
rect 186 100355 220 100369
rect 548 100355 582 100369
rect 599 100355 649 100357
rect 42 100313 59 100347
rect 67 100305 69 100355
rect 160 100347 246 100355
rect 522 100347 608 100355
rect 76 100313 110 100347
rect 127 100313 144 100347
rect 152 100313 161 100347
rect 162 100345 195 100347
rect 224 100345 244 100347
rect 162 100313 244 100345
rect 524 100345 548 100347
rect 573 100345 582 100347
rect 586 100345 606 100347
rect 160 100305 246 100313
rect 186 100289 220 100305
rect 182 100275 224 100276
rect 160 100269 182 100275
rect 224 100269 246 100275
rect 186 100234 220 100268
rect 223 100234 257 100268
rect 120 100221 170 100223
rect 76 100217 130 100221
rect 110 100212 130 100217
rect 60 100187 67 100197
rect 76 100187 77 100207
rect 96 100178 99 100212
rect 109 100187 110 100207
rect 119 100187 126 100197
rect 76 100171 92 100177
rect 94 100171 110 100177
rect 170 100171 172 100221
rect 186 100155 190 100189
rect 216 100155 220 100189
rect 288 100155 292 100343
rect 476 100275 480 100343
rect 524 100313 606 100345
rect 607 100313 616 100347
rect 522 100305 608 100313
rect 649 100305 651 100355
rect 548 100289 582 100305
rect 522 100270 548 100275
rect 522 100269 582 100270
rect 586 100269 608 100275
rect 295 100234 300 100268
rect 324 100234 329 100268
rect 544 100266 582 100269
rect 378 100229 450 100237
rect 428 100199 430 100215
rect 400 100191 430 100199
rect 476 100197 480 100265
rect 544 100236 552 100266
rect 578 100236 582 100266
rect 544 100227 548 100236
rect 400 100187 436 100191
rect 400 100157 408 100187
rect 420 100157 436 100187
rect 544 100189 548 100197
rect 12 100118 62 100120
rect 28 100109 59 100117
rect 62 100109 64 100118
rect 28 100101 64 100109
rect 127 100109 158 100117
rect 127 100102 182 100109
rect 215 100107 224 100135
rect 127 100101 161 100102
rect 59 100085 64 100101
rect 158 100085 161 100101
rect 28 100077 64 100085
rect 127 100084 161 100085
rect 127 100077 182 100084
rect 62 100068 64 100077
rect 213 100069 224 100107
rect 282 100097 292 100155
rect 296 100149 368 100157
rect 319 100119 346 100130
rect 318 100106 324 100119
rect 346 100106 348 100119
rect 428 100110 430 100157
rect 443 100147 450 100149
rect 476 100117 480 100185
rect 544 100155 552 100189
rect 578 100155 582 100189
rect 481 100123 517 100151
rect 481 100117 495 100123
rect 367 100106 380 100110
rect 251 100063 263 100097
rect 273 100063 293 100097
rect 295 100082 324 100106
rect 303 100072 316 100082
rect 318 100066 324 100082
rect 333 100082 380 100106
rect 333 100072 353 100082
rect 367 100076 380 100082
rect 396 100076 408 100110
rect 420 100076 436 100110
rect 120 100015 170 100017
rect 76 100009 92 100015
rect 94 100009 110 100015
rect 76 99999 99 100008
rect 60 99989 67 99999
rect 76 99979 77 99999
rect 96 99974 99 99999
rect 109 99979 110 99999
rect 119 99989 126 99999
rect 76 99965 110 99969
rect 170 99965 172 100015
rect 186 99997 190 100031
rect 216 99997 220 100031
rect 186 99920 220 99954
rect 282 99951 292 100063
rect 318 100056 335 100066
rect 318 99987 324 100056
rect 346 99987 348 100072
rect 428 100029 430 100076
rect 476 100039 480 100107
rect 485 100089 495 100117
rect 505 100117 519 100123
rect 544 100117 555 100155
rect 505 100089 525 100117
rect 544 100089 553 100117
rect 544 100069 548 100089
rect 579 100048 582 100138
rect 612 100120 624 100121
rect 599 100118 649 100120
rect 612 100117 624 100118
rect 610 100110 632 100117
rect 607 100109 632 100110
rect 586 100102 644 100109
rect 607 100101 644 100102
rect 607 100085 610 100101
rect 616 100085 644 100101
rect 607 100084 644 100085
rect 586 100077 644 100084
rect 607 100076 610 100077
rect 612 100069 632 100077
rect 612 100065 624 100069
rect 649 100068 651 100118
rect 544 100031 548 100039
rect 400 99999 408 100029
rect 420 99999 436 100029
rect 400 99995 436 99999
rect 400 99987 430 99995
rect 428 99971 430 99987
rect 476 99959 480 100027
rect 544 99997 552 100031
rect 578 99997 582 100031
rect 544 99989 548 99997
rect 544 99959 586 99960
rect 288 99919 292 99951
rect 296 99949 368 99957
rect 378 99949 450 99957
rect 544 99952 548 99959
rect 439 99921 444 99949
rect 120 99905 170 99907
rect 76 99901 130 99905
rect 110 99896 130 99901
rect 60 99871 67 99881
rect 76 99871 77 99891
rect 96 99862 99 99896
rect 109 99871 110 99891
rect 119 99871 126 99881
rect 76 99855 92 99861
rect 94 99855 110 99861
rect 170 99855 172 99905
rect 186 99839 190 99873
rect 216 99839 220 99873
rect 213 99807 224 99839
rect 282 99835 292 99919
rect 296 99913 368 99921
rect 378 99913 450 99921
rect 468 99918 473 99952
rect 428 99883 430 99899
rect 251 99807 292 99835
rect 318 99814 324 99883
rect 12 99802 62 99804
rect 28 99793 59 99801
rect 62 99793 64 99802
rect 251 99801 263 99807
rect 28 99785 64 99793
rect 127 99793 158 99801
rect 127 99786 182 99793
rect 127 99785 161 99786
rect 59 99769 64 99785
rect 158 99769 161 99785
rect 253 99773 263 99801
rect 273 99773 293 99807
rect 318 99804 335 99814
rect 303 99788 316 99798
rect 318 99788 324 99804
rect 346 99798 348 99883
rect 400 99875 430 99883
rect 476 99881 480 99949
rect 511 99918 582 99952
rect 544 99911 548 99918
rect 400 99871 436 99875
rect 400 99841 408 99871
rect 420 99841 436 99871
rect 544 99873 548 99881
rect 28 99761 64 99769
rect 127 99768 161 99769
rect 127 99761 182 99768
rect 62 99752 64 99761
rect 282 99715 292 99773
rect 295 99764 324 99788
rect 333 99788 353 99798
rect 428 99794 430 99841
rect 476 99801 480 99869
rect 544 99839 552 99873
rect 578 99839 582 99873
rect 544 99831 548 99839
rect 367 99788 380 99794
rect 333 99764 380 99788
rect 318 99751 324 99764
rect 346 99751 348 99764
rect 367 99760 380 99764
rect 396 99760 408 99794
rect 420 99760 436 99794
rect 544 99791 553 99819
rect 319 99740 346 99751
rect 120 99699 170 99701
rect 76 99693 92 99699
rect 94 99693 110 99699
rect 76 99683 99 99692
rect 60 99673 67 99683
rect 76 99663 77 99683
rect 96 99658 99 99683
rect 109 99663 110 99683
rect 119 99673 126 99683
rect 76 99649 110 99653
rect 170 99649 172 99699
rect 186 99681 190 99715
rect 216 99681 220 99715
rect 182 99643 224 99644
rect 186 99619 220 99636
rect 223 99619 257 99636
rect 182 99602 257 99619
rect 182 99601 224 99602
rect 160 99595 246 99601
rect 288 99595 292 99715
rect 296 99713 368 99721
rect 428 99713 430 99760
rect 476 99723 480 99791
rect 485 99747 495 99781
rect 505 99753 525 99781
rect 505 99747 519 99753
rect 544 99747 555 99791
rect 485 99723 492 99747
rect 579 99732 582 99822
rect 612 99804 624 99805
rect 599 99802 649 99804
rect 612 99801 624 99802
rect 610 99794 632 99801
rect 607 99793 632 99794
rect 586 99786 644 99793
rect 607 99785 644 99786
rect 607 99769 610 99785
rect 616 99769 644 99785
rect 607 99768 644 99769
rect 586 99761 644 99768
rect 607 99760 610 99761
rect 612 99753 632 99761
rect 612 99749 624 99753
rect 649 99752 651 99802
rect 544 99715 548 99723
rect 400 99683 408 99713
rect 420 99683 436 99713
rect 400 99679 436 99683
rect 400 99671 430 99679
rect 428 99655 430 99671
rect 476 99643 480 99711
rect 544 99681 552 99715
rect 578 99681 582 99715
rect 544 99673 548 99681
rect 295 99602 300 99636
rect 324 99602 329 99636
rect 378 99633 450 99641
rect 544 99638 548 99643
rect 544 99634 582 99638
rect 544 99619 552 99634
rect 578 99619 582 99634
rect 544 99601 586 99619
rect 522 99595 608 99601
rect 182 99579 224 99595
rect 544 99579 586 99595
rect 17 99565 67 99567
rect 119 99565 169 99567
rect 186 99565 220 99579
rect 548 99565 582 99579
rect 599 99565 649 99567
rect 42 99523 59 99557
rect 67 99515 69 99565
rect 160 99557 246 99565
rect 522 99557 608 99565
rect 76 99523 110 99557
rect 127 99523 144 99557
rect 152 99523 161 99557
rect 162 99555 195 99557
rect 224 99555 244 99557
rect 162 99523 244 99555
rect 524 99555 548 99557
rect 573 99555 582 99557
rect 586 99555 606 99557
rect 160 99515 246 99523
rect 186 99499 220 99515
rect 182 99485 224 99486
rect 160 99479 182 99485
rect 224 99479 246 99485
rect 186 99444 220 99478
rect 223 99444 257 99478
rect 120 99431 170 99433
rect 76 99427 130 99431
rect 110 99422 130 99427
rect 60 99397 67 99407
rect 76 99397 77 99417
rect 96 99388 99 99422
rect 109 99397 110 99417
rect 119 99397 126 99407
rect 76 99381 92 99387
rect 94 99381 110 99387
rect 170 99381 172 99431
rect 186 99365 190 99399
rect 216 99365 220 99399
rect 288 99365 292 99553
rect 476 99485 480 99553
rect 524 99523 606 99555
rect 607 99523 616 99557
rect 522 99515 608 99523
rect 649 99515 651 99565
rect 548 99499 582 99515
rect 522 99480 548 99485
rect 522 99479 582 99480
rect 586 99479 608 99485
rect 295 99444 300 99478
rect 324 99444 329 99478
rect 544 99476 582 99479
rect 378 99439 450 99447
rect 428 99409 430 99425
rect 400 99401 430 99409
rect 476 99407 480 99475
rect 544 99446 552 99476
rect 578 99446 582 99476
rect 544 99437 548 99446
rect 400 99397 436 99401
rect 400 99367 408 99397
rect 420 99367 436 99397
rect 544 99399 548 99407
rect 12 99328 62 99330
rect 28 99319 59 99327
rect 62 99319 64 99328
rect 28 99311 64 99319
rect 127 99319 158 99327
rect 127 99312 182 99319
rect 215 99317 224 99345
rect 127 99311 161 99312
rect 59 99295 64 99311
rect 158 99295 161 99311
rect 28 99287 64 99295
rect 127 99294 161 99295
rect 127 99287 182 99294
rect 62 99278 64 99287
rect 213 99279 224 99317
rect 282 99307 292 99365
rect 296 99359 368 99367
rect 319 99329 346 99340
rect 318 99316 324 99329
rect 346 99316 348 99329
rect 428 99320 430 99367
rect 443 99357 450 99359
rect 476 99327 480 99395
rect 544 99365 552 99399
rect 578 99365 582 99399
rect 481 99333 517 99361
rect 481 99327 495 99333
rect 367 99316 380 99320
rect 251 99273 263 99307
rect 273 99273 293 99307
rect 295 99292 324 99316
rect 303 99282 316 99292
rect 318 99276 324 99292
rect 333 99292 380 99316
rect 333 99282 353 99292
rect 367 99286 380 99292
rect 396 99286 408 99320
rect 420 99286 436 99320
rect 120 99225 170 99227
rect 76 99219 92 99225
rect 94 99219 110 99225
rect 76 99209 99 99218
rect 60 99199 67 99209
rect 76 99189 77 99209
rect 96 99184 99 99209
rect 109 99189 110 99209
rect 119 99199 126 99209
rect 76 99175 110 99179
rect 170 99175 172 99225
rect 186 99207 190 99241
rect 216 99207 220 99241
rect 186 99130 220 99164
rect 282 99161 292 99273
rect 318 99266 335 99276
rect 318 99197 324 99266
rect 346 99197 348 99282
rect 428 99239 430 99286
rect 476 99249 480 99317
rect 485 99299 495 99327
rect 505 99327 519 99333
rect 544 99327 555 99365
rect 505 99299 525 99327
rect 544 99299 553 99327
rect 544 99279 548 99299
rect 579 99258 582 99348
rect 612 99330 624 99331
rect 599 99328 649 99330
rect 612 99327 624 99328
rect 610 99320 632 99327
rect 607 99319 632 99320
rect 586 99312 644 99319
rect 607 99311 644 99312
rect 607 99295 610 99311
rect 616 99295 644 99311
rect 607 99294 644 99295
rect 586 99287 644 99294
rect 607 99286 610 99287
rect 612 99279 632 99287
rect 612 99275 624 99279
rect 649 99278 651 99328
rect 544 99241 548 99249
rect 400 99209 408 99239
rect 420 99209 436 99239
rect 400 99205 436 99209
rect 400 99197 430 99205
rect 428 99181 430 99197
rect 476 99169 480 99237
rect 544 99207 552 99241
rect 578 99207 582 99241
rect 544 99199 548 99207
rect 544 99169 586 99170
rect 288 99129 292 99161
rect 296 99159 368 99167
rect 378 99159 450 99167
rect 544 99162 548 99169
rect 439 99131 444 99159
rect 120 99115 170 99117
rect 76 99111 130 99115
rect 110 99106 130 99111
rect 60 99081 67 99091
rect 76 99081 77 99101
rect 96 99072 99 99106
rect 109 99081 110 99101
rect 119 99081 126 99091
rect 76 99065 92 99071
rect 94 99065 110 99071
rect 170 99065 172 99115
rect 186 99049 190 99083
rect 216 99049 220 99083
rect 213 99017 224 99049
rect 282 99045 292 99129
rect 296 99123 368 99131
rect 378 99123 450 99131
rect 468 99128 473 99162
rect 428 99093 430 99109
rect 251 99017 292 99045
rect 318 99024 324 99093
rect 12 99012 62 99014
rect 28 99003 59 99011
rect 62 99003 64 99012
rect 251 99011 263 99017
rect 28 98995 64 99003
rect 127 99003 158 99011
rect 127 98996 182 99003
rect 127 98995 161 98996
rect 59 98979 64 98995
rect 158 98979 161 98995
rect 253 98983 263 99011
rect 273 98983 293 99017
rect 318 99014 335 99024
rect 303 98998 316 99008
rect 318 98998 324 99014
rect 346 99008 348 99093
rect 400 99085 430 99093
rect 476 99091 480 99159
rect 511 99128 582 99162
rect 544 99121 548 99128
rect 400 99081 436 99085
rect 400 99051 408 99081
rect 420 99051 436 99081
rect 544 99083 548 99091
rect 28 98971 64 98979
rect 127 98978 161 98979
rect 127 98971 182 98978
rect 62 98962 64 98971
rect 282 98925 292 98983
rect 295 98974 324 98998
rect 333 98998 353 99008
rect 428 99004 430 99051
rect 476 99011 480 99079
rect 544 99049 552 99083
rect 578 99049 582 99083
rect 544 99041 548 99049
rect 367 98998 380 99004
rect 333 98974 380 98998
rect 318 98961 324 98974
rect 346 98961 348 98974
rect 367 98970 380 98974
rect 396 98970 408 99004
rect 420 98970 436 99004
rect 544 99001 553 99029
rect 319 98950 346 98961
rect 120 98909 170 98911
rect 76 98903 92 98909
rect 94 98903 110 98909
rect 76 98893 99 98902
rect 60 98883 67 98893
rect 76 98873 77 98893
rect 96 98868 99 98893
rect 109 98873 110 98893
rect 119 98883 126 98893
rect 76 98859 110 98863
rect 170 98859 172 98909
rect 186 98891 190 98925
rect 216 98891 220 98925
rect 182 98853 224 98854
rect 186 98829 220 98846
rect 223 98829 257 98846
rect 182 98812 257 98829
rect 182 98811 224 98812
rect 160 98805 246 98811
rect 288 98805 292 98925
rect 296 98923 368 98931
rect 428 98923 430 98970
rect 476 98933 480 99001
rect 485 98957 495 98991
rect 505 98963 525 98991
rect 505 98957 519 98963
rect 544 98957 555 99001
rect 485 98933 492 98957
rect 579 98942 582 99032
rect 612 99014 624 99015
rect 599 99012 649 99014
rect 612 99011 624 99012
rect 610 99004 632 99011
rect 607 99003 632 99004
rect 586 98996 644 99003
rect 607 98995 644 98996
rect 607 98979 610 98995
rect 616 98979 644 98995
rect 607 98978 644 98979
rect 586 98971 644 98978
rect 607 98970 610 98971
rect 612 98963 632 98971
rect 612 98959 624 98963
rect 649 98962 651 99012
rect 544 98925 548 98933
rect 400 98893 408 98923
rect 420 98893 436 98923
rect 400 98889 436 98893
rect 400 98881 430 98889
rect 428 98865 430 98881
rect 476 98853 480 98921
rect 544 98891 552 98925
rect 578 98891 582 98925
rect 544 98883 548 98891
rect 295 98812 300 98846
rect 324 98812 329 98846
rect 378 98843 450 98851
rect 544 98848 548 98853
rect 544 98844 582 98848
rect 544 98829 552 98844
rect 578 98829 582 98844
rect 544 98811 586 98829
rect 522 98805 608 98811
rect 182 98789 224 98805
rect 544 98789 586 98805
rect 17 98775 67 98777
rect 119 98775 169 98777
rect 186 98775 220 98789
rect 548 98775 582 98789
rect 599 98775 649 98777
rect 42 98733 59 98767
rect 67 98725 69 98775
rect 160 98767 246 98775
rect 522 98767 608 98775
rect 76 98733 110 98767
rect 127 98733 144 98767
rect 152 98733 161 98767
rect 162 98765 195 98767
rect 224 98765 244 98767
rect 162 98733 244 98765
rect 524 98765 548 98767
rect 573 98765 582 98767
rect 586 98765 606 98767
rect 160 98725 246 98733
rect 186 98709 220 98725
rect 182 98695 224 98696
rect 160 98689 182 98695
rect 224 98689 246 98695
rect 186 98654 220 98688
rect 223 98654 257 98688
rect 120 98641 170 98643
rect 76 98637 130 98641
rect 110 98632 130 98637
rect 60 98607 67 98617
rect 76 98607 77 98627
rect 96 98598 99 98632
rect 109 98607 110 98627
rect 119 98607 126 98617
rect 76 98591 92 98597
rect 94 98591 110 98597
rect 170 98591 172 98641
rect 186 98575 190 98609
rect 216 98575 220 98609
rect 288 98575 292 98763
rect 476 98695 480 98763
rect 524 98733 606 98765
rect 607 98733 616 98767
rect 522 98725 608 98733
rect 649 98725 651 98775
rect 548 98709 582 98725
rect 522 98690 548 98695
rect 522 98689 582 98690
rect 586 98689 608 98695
rect 295 98654 300 98688
rect 324 98654 329 98688
rect 544 98686 582 98689
rect 378 98649 450 98657
rect 428 98619 430 98635
rect 400 98611 430 98619
rect 476 98617 480 98685
rect 544 98656 552 98686
rect 578 98656 582 98686
rect 544 98647 548 98656
rect 400 98607 436 98611
rect 400 98577 408 98607
rect 420 98577 436 98607
rect 544 98609 548 98617
rect 12 98538 62 98540
rect 28 98529 59 98537
rect 62 98529 64 98538
rect 28 98521 64 98529
rect 127 98529 158 98537
rect 127 98522 182 98529
rect 215 98527 224 98555
rect 127 98521 161 98522
rect 59 98505 64 98521
rect 158 98505 161 98521
rect 28 98497 64 98505
rect 127 98504 161 98505
rect 127 98497 182 98504
rect 62 98488 64 98497
rect 213 98489 224 98527
rect 282 98517 292 98575
rect 296 98569 368 98577
rect 319 98539 346 98550
rect 318 98526 324 98539
rect 346 98526 348 98539
rect 428 98530 430 98577
rect 443 98567 450 98569
rect 476 98537 480 98605
rect 544 98575 552 98609
rect 578 98575 582 98609
rect 481 98543 517 98571
rect 481 98537 495 98543
rect 367 98526 380 98530
rect 251 98483 263 98517
rect 273 98483 293 98517
rect 295 98502 324 98526
rect 303 98492 316 98502
rect 318 98486 324 98502
rect 333 98502 380 98526
rect 333 98492 353 98502
rect 367 98496 380 98502
rect 396 98496 408 98530
rect 420 98496 436 98530
rect 120 98435 170 98437
rect 76 98429 92 98435
rect 94 98429 110 98435
rect 76 98419 99 98428
rect 60 98409 67 98419
rect 76 98399 77 98419
rect 96 98394 99 98419
rect 109 98399 110 98419
rect 119 98409 126 98419
rect 76 98385 110 98389
rect 170 98385 172 98435
rect 186 98417 190 98451
rect 216 98417 220 98451
rect 186 98340 220 98374
rect 282 98371 292 98483
rect 318 98476 335 98486
rect 318 98407 324 98476
rect 346 98407 348 98492
rect 428 98449 430 98496
rect 476 98459 480 98527
rect 485 98509 495 98537
rect 505 98537 519 98543
rect 544 98537 555 98575
rect 505 98509 525 98537
rect 544 98509 553 98537
rect 544 98489 548 98509
rect 579 98468 582 98558
rect 612 98540 624 98541
rect 599 98538 649 98540
rect 612 98537 624 98538
rect 610 98530 632 98537
rect 607 98529 632 98530
rect 586 98522 644 98529
rect 607 98521 644 98522
rect 607 98505 610 98521
rect 616 98505 644 98521
rect 607 98504 644 98505
rect 586 98497 644 98504
rect 607 98496 610 98497
rect 612 98489 632 98497
rect 612 98485 624 98489
rect 649 98488 651 98538
rect 544 98451 548 98459
rect 400 98419 408 98449
rect 420 98419 436 98449
rect 400 98415 436 98419
rect 400 98407 430 98415
rect 428 98391 430 98407
rect 476 98379 480 98447
rect 544 98417 552 98451
rect 578 98417 582 98451
rect 544 98409 548 98417
rect 544 98379 586 98380
rect 288 98339 292 98371
rect 296 98369 368 98377
rect 378 98369 450 98377
rect 544 98372 548 98379
rect 439 98341 444 98369
rect 120 98325 170 98327
rect 76 98321 130 98325
rect 110 98316 130 98321
rect 60 98291 67 98301
rect 76 98291 77 98311
rect 96 98282 99 98316
rect 109 98291 110 98311
rect 119 98291 126 98301
rect 76 98275 92 98281
rect 94 98275 110 98281
rect 170 98275 172 98325
rect 186 98259 190 98293
rect 216 98259 220 98293
rect 213 98227 224 98259
rect 282 98255 292 98339
rect 296 98333 368 98341
rect 378 98333 450 98341
rect 468 98338 473 98372
rect 428 98303 430 98319
rect 251 98227 292 98255
rect 318 98234 324 98303
rect 12 98222 62 98224
rect 28 98213 59 98221
rect 62 98213 64 98222
rect 251 98221 263 98227
rect 28 98205 64 98213
rect 127 98213 158 98221
rect 127 98206 182 98213
rect 127 98205 161 98206
rect 59 98189 64 98205
rect 158 98189 161 98205
rect 253 98193 263 98221
rect 273 98193 293 98227
rect 318 98224 335 98234
rect 303 98208 316 98218
rect 318 98208 324 98224
rect 346 98218 348 98303
rect 400 98295 430 98303
rect 476 98301 480 98369
rect 511 98338 582 98372
rect 544 98331 548 98338
rect 400 98291 436 98295
rect 400 98261 408 98291
rect 420 98261 436 98291
rect 544 98293 548 98301
rect 28 98181 64 98189
rect 127 98188 161 98189
rect 127 98181 182 98188
rect 62 98172 64 98181
rect 282 98135 292 98193
rect 295 98184 324 98208
rect 333 98208 353 98218
rect 428 98214 430 98261
rect 476 98221 480 98289
rect 544 98259 552 98293
rect 578 98259 582 98293
rect 544 98251 548 98259
rect 367 98208 380 98214
rect 333 98184 380 98208
rect 318 98171 324 98184
rect 346 98171 348 98184
rect 367 98180 380 98184
rect 396 98180 408 98214
rect 420 98180 436 98214
rect 544 98211 553 98239
rect 319 98160 346 98171
rect 120 98119 170 98121
rect 76 98113 92 98119
rect 94 98113 110 98119
rect 76 98103 99 98112
rect 60 98093 67 98103
rect 76 98083 77 98103
rect 96 98078 99 98103
rect 109 98083 110 98103
rect 119 98093 126 98103
rect 76 98069 110 98073
rect 170 98069 172 98119
rect 186 98101 190 98135
rect 216 98101 220 98135
rect 182 98063 224 98064
rect 186 98039 220 98056
rect 223 98039 257 98056
rect 182 98022 257 98039
rect 182 98021 224 98022
rect 160 98015 246 98021
rect 288 98015 292 98135
rect 296 98133 368 98141
rect 428 98133 430 98180
rect 476 98143 480 98211
rect 485 98167 495 98201
rect 505 98173 525 98201
rect 505 98167 519 98173
rect 544 98167 555 98211
rect 485 98143 492 98167
rect 579 98152 582 98242
rect 612 98224 624 98225
rect 599 98222 649 98224
rect 612 98221 624 98222
rect 610 98214 632 98221
rect 607 98213 632 98214
rect 586 98206 644 98213
rect 607 98205 644 98206
rect 607 98189 610 98205
rect 616 98189 644 98205
rect 607 98188 644 98189
rect 586 98181 644 98188
rect 607 98180 610 98181
rect 612 98173 632 98181
rect 612 98169 624 98173
rect 649 98172 651 98222
rect 544 98135 548 98143
rect 400 98103 408 98133
rect 420 98103 436 98133
rect 400 98099 436 98103
rect 400 98091 430 98099
rect 428 98075 430 98091
rect 476 98063 480 98131
rect 544 98101 552 98135
rect 578 98101 582 98135
rect 544 98093 548 98101
rect 295 98022 300 98056
rect 324 98022 329 98056
rect 378 98053 450 98061
rect 544 98058 548 98063
rect 544 98054 582 98058
rect 544 98039 552 98054
rect 578 98039 582 98054
rect 544 98021 586 98039
rect 522 98015 608 98021
rect 182 97999 224 98015
rect 544 97999 586 98015
rect 17 97985 67 97987
rect 119 97985 169 97987
rect 186 97985 220 97999
rect 548 97985 582 97999
rect 599 97985 649 97987
rect 42 97943 59 97977
rect 67 97935 69 97985
rect 160 97977 246 97985
rect 522 97977 608 97985
rect 76 97943 110 97977
rect 127 97943 144 97977
rect 152 97943 161 97977
rect 162 97975 195 97977
rect 224 97975 244 97977
rect 162 97943 244 97975
rect 524 97975 548 97977
rect 573 97975 582 97977
rect 586 97975 606 97977
rect 160 97935 246 97943
rect 186 97919 220 97935
rect 182 97905 224 97906
rect 160 97899 182 97905
rect 224 97899 246 97905
rect 186 97864 220 97898
rect 223 97864 257 97898
rect 120 97851 170 97853
rect 76 97847 130 97851
rect 110 97842 130 97847
rect 60 97817 67 97827
rect 76 97817 77 97837
rect 96 97808 99 97842
rect 109 97817 110 97837
rect 119 97817 126 97827
rect 76 97801 92 97807
rect 94 97801 110 97807
rect 170 97801 172 97851
rect 186 97785 190 97819
rect 216 97785 220 97819
rect 288 97785 292 97973
rect 476 97905 480 97973
rect 524 97943 606 97975
rect 607 97943 616 97977
rect 522 97935 608 97943
rect 649 97935 651 97985
rect 548 97919 582 97935
rect 522 97900 548 97905
rect 522 97899 582 97900
rect 586 97899 608 97905
rect 295 97864 300 97898
rect 324 97864 329 97898
rect 544 97896 582 97899
rect 378 97859 450 97867
rect 428 97829 430 97845
rect 400 97821 430 97829
rect 476 97827 480 97895
rect 544 97866 552 97896
rect 578 97866 582 97896
rect 544 97857 548 97866
rect 400 97817 436 97821
rect 400 97787 408 97817
rect 420 97787 436 97817
rect 544 97819 548 97827
rect 12 97748 62 97750
rect 28 97739 59 97747
rect 62 97739 64 97748
rect 28 97731 64 97739
rect 127 97739 158 97747
rect 127 97732 182 97739
rect 215 97737 224 97765
rect 127 97731 161 97732
rect 59 97715 64 97731
rect 158 97715 161 97731
rect 28 97707 64 97715
rect 127 97714 161 97715
rect 127 97707 182 97714
rect 62 97698 64 97707
rect 213 97699 224 97737
rect 282 97727 292 97785
rect 296 97779 368 97787
rect 319 97749 346 97760
rect 318 97736 324 97749
rect 346 97736 348 97749
rect 428 97740 430 97787
rect 443 97777 450 97779
rect 476 97747 480 97815
rect 544 97785 552 97819
rect 578 97785 582 97819
rect 481 97753 517 97781
rect 481 97747 495 97753
rect 367 97736 380 97740
rect 251 97693 263 97727
rect 273 97693 293 97727
rect 295 97712 324 97736
rect 303 97702 316 97712
rect 318 97696 324 97712
rect 333 97712 380 97736
rect 333 97702 353 97712
rect 367 97706 380 97712
rect 396 97706 408 97740
rect 420 97706 436 97740
rect 120 97645 170 97647
rect 76 97639 92 97645
rect 94 97639 110 97645
rect 76 97629 99 97638
rect 60 97619 67 97629
rect 76 97609 77 97629
rect 96 97604 99 97629
rect 109 97609 110 97629
rect 119 97619 126 97629
rect 76 97595 110 97599
rect 170 97595 172 97645
rect 186 97627 190 97661
rect 216 97627 220 97661
rect 186 97550 220 97584
rect 282 97581 292 97693
rect 318 97686 335 97696
rect 318 97617 324 97686
rect 346 97617 348 97702
rect 428 97659 430 97706
rect 476 97669 480 97737
rect 485 97719 495 97747
rect 505 97747 519 97753
rect 544 97747 555 97785
rect 505 97719 525 97747
rect 544 97719 553 97747
rect 544 97699 548 97719
rect 579 97678 582 97768
rect 612 97750 624 97751
rect 599 97748 649 97750
rect 612 97747 624 97748
rect 610 97740 632 97747
rect 607 97739 632 97740
rect 586 97732 644 97739
rect 607 97731 644 97732
rect 607 97715 610 97731
rect 616 97715 644 97731
rect 607 97714 644 97715
rect 586 97707 644 97714
rect 607 97706 610 97707
rect 612 97699 632 97707
rect 612 97695 624 97699
rect 649 97698 651 97748
rect 544 97661 548 97669
rect 400 97629 408 97659
rect 420 97629 436 97659
rect 400 97625 436 97629
rect 400 97617 430 97625
rect 428 97601 430 97617
rect 476 97589 480 97657
rect 544 97627 552 97661
rect 578 97627 582 97661
rect 544 97619 548 97627
rect 544 97589 586 97590
rect 288 97549 292 97581
rect 296 97579 368 97587
rect 378 97579 450 97587
rect 544 97582 548 97589
rect 439 97551 444 97579
rect 120 97535 170 97537
rect 76 97531 130 97535
rect 110 97526 130 97531
rect 60 97501 67 97511
rect 76 97501 77 97521
rect 96 97492 99 97526
rect 109 97501 110 97521
rect 119 97501 126 97511
rect 76 97485 92 97491
rect 94 97485 110 97491
rect 170 97485 172 97535
rect 186 97469 190 97503
rect 216 97469 220 97503
rect 213 97437 224 97469
rect 282 97465 292 97549
rect 296 97543 368 97551
rect 378 97543 450 97551
rect 468 97548 473 97582
rect 428 97513 430 97529
rect 251 97437 292 97465
rect 318 97444 324 97513
rect 12 97432 62 97434
rect 28 97423 59 97431
rect 62 97423 64 97432
rect 251 97431 263 97437
rect 28 97415 64 97423
rect 127 97423 158 97431
rect 127 97416 182 97423
rect 127 97415 161 97416
rect 59 97399 64 97415
rect 158 97399 161 97415
rect 253 97403 263 97431
rect 273 97403 293 97437
rect 318 97434 335 97444
rect 303 97418 316 97428
rect 318 97418 324 97434
rect 346 97428 348 97513
rect 400 97505 430 97513
rect 476 97511 480 97579
rect 511 97548 582 97582
rect 544 97541 548 97548
rect 400 97501 436 97505
rect 400 97471 408 97501
rect 420 97471 436 97501
rect 544 97503 548 97511
rect 28 97391 64 97399
rect 127 97398 161 97399
rect 127 97391 182 97398
rect 62 97382 64 97391
rect 282 97345 292 97403
rect 295 97394 324 97418
rect 333 97418 353 97428
rect 428 97424 430 97471
rect 476 97431 480 97499
rect 544 97469 552 97503
rect 578 97469 582 97503
rect 544 97461 548 97469
rect 367 97418 380 97424
rect 333 97394 380 97418
rect 318 97381 324 97394
rect 346 97381 348 97394
rect 367 97390 380 97394
rect 396 97390 408 97424
rect 420 97390 436 97424
rect 544 97421 553 97449
rect 319 97370 346 97381
rect 120 97329 170 97331
rect 76 97323 92 97329
rect 94 97323 110 97329
rect 76 97313 99 97322
rect 60 97303 67 97313
rect 76 97293 77 97313
rect 96 97288 99 97313
rect 109 97293 110 97313
rect 119 97303 126 97313
rect 76 97279 110 97283
rect 170 97279 172 97329
rect 186 97311 190 97345
rect 216 97311 220 97345
rect 182 97273 224 97274
rect 186 97249 220 97266
rect 223 97249 257 97266
rect 182 97232 257 97249
rect 182 97231 224 97232
rect 160 97225 246 97231
rect 288 97225 292 97345
rect 296 97343 368 97351
rect 428 97343 430 97390
rect 476 97353 480 97421
rect 485 97377 495 97411
rect 505 97383 525 97411
rect 505 97377 519 97383
rect 544 97377 555 97421
rect 485 97353 492 97377
rect 579 97362 582 97452
rect 612 97434 624 97435
rect 599 97432 649 97434
rect 612 97431 624 97432
rect 610 97424 632 97431
rect 607 97423 632 97424
rect 586 97416 644 97423
rect 607 97415 644 97416
rect 607 97399 610 97415
rect 616 97399 644 97415
rect 607 97398 644 97399
rect 586 97391 644 97398
rect 607 97390 610 97391
rect 612 97383 632 97391
rect 612 97379 624 97383
rect 649 97382 651 97432
rect 544 97345 548 97353
rect 400 97313 408 97343
rect 420 97313 436 97343
rect 400 97309 436 97313
rect 400 97301 430 97309
rect 428 97285 430 97301
rect 476 97273 480 97341
rect 544 97311 552 97345
rect 578 97311 582 97345
rect 544 97303 548 97311
rect 295 97232 300 97266
rect 324 97232 329 97266
rect 378 97263 450 97271
rect 544 97268 548 97273
rect 544 97264 582 97268
rect 544 97249 552 97264
rect 578 97249 582 97264
rect 544 97231 586 97249
rect 522 97225 608 97231
rect 182 97209 224 97225
rect 544 97209 586 97225
rect 17 97195 67 97197
rect 119 97195 169 97197
rect 186 97195 220 97209
rect 548 97195 582 97209
rect 599 97195 649 97197
rect 42 97153 59 97187
rect 67 97145 69 97195
rect 160 97187 246 97195
rect 522 97187 608 97195
rect 76 97153 110 97187
rect 127 97153 144 97187
rect 152 97153 161 97187
rect 162 97185 195 97187
rect 224 97185 244 97187
rect 162 97153 244 97185
rect 524 97185 548 97187
rect 573 97185 582 97187
rect 586 97185 606 97187
rect 160 97145 246 97153
rect 186 97129 220 97145
rect 182 97115 224 97116
rect 160 97109 182 97115
rect 224 97109 246 97115
rect 186 97074 220 97108
rect 223 97074 257 97108
rect 120 97061 170 97063
rect 76 97057 130 97061
rect 110 97052 130 97057
rect 60 97027 67 97037
rect 76 97027 77 97047
rect 96 97018 99 97052
rect 109 97027 110 97047
rect 119 97027 126 97037
rect 76 97011 92 97017
rect 94 97011 110 97017
rect 170 97011 172 97061
rect 186 96995 190 97029
rect 216 96995 220 97029
rect 288 96995 292 97183
rect 476 97115 480 97183
rect 524 97153 606 97185
rect 607 97153 616 97187
rect 522 97145 608 97153
rect 649 97145 651 97195
rect 548 97129 582 97145
rect 522 97110 548 97115
rect 522 97109 582 97110
rect 586 97109 608 97115
rect 295 97074 300 97108
rect 324 97074 329 97108
rect 544 97106 582 97109
rect 378 97069 450 97077
rect 428 97039 430 97055
rect 400 97031 430 97039
rect 476 97037 480 97105
rect 544 97076 552 97106
rect 578 97076 582 97106
rect 544 97067 548 97076
rect 400 97027 436 97031
rect 400 96997 408 97027
rect 420 96997 436 97027
rect 544 97029 548 97037
rect 12 96958 62 96960
rect 28 96949 59 96957
rect 62 96949 64 96958
rect 28 96941 64 96949
rect 127 96949 158 96957
rect 127 96942 182 96949
rect 215 96947 224 96975
rect 127 96941 161 96942
rect 59 96925 64 96941
rect 158 96925 161 96941
rect 28 96917 64 96925
rect 127 96924 161 96925
rect 127 96917 182 96924
rect 62 96908 64 96917
rect 213 96909 224 96947
rect 282 96937 292 96995
rect 296 96989 368 96997
rect 319 96959 346 96970
rect 318 96946 324 96959
rect 346 96946 348 96959
rect 428 96950 430 96997
rect 443 96987 450 96989
rect 476 96957 480 97025
rect 544 96995 552 97029
rect 578 96995 582 97029
rect 481 96963 517 96991
rect 481 96957 495 96963
rect 367 96946 380 96950
rect 251 96903 263 96937
rect 273 96903 293 96937
rect 295 96922 324 96946
rect 303 96912 316 96922
rect 318 96906 324 96922
rect 333 96922 380 96946
rect 333 96912 353 96922
rect 367 96916 380 96922
rect 396 96916 408 96950
rect 420 96916 436 96950
rect 120 96855 170 96857
rect 76 96849 92 96855
rect 94 96849 110 96855
rect 76 96839 99 96848
rect 60 96829 67 96839
rect 76 96819 77 96839
rect 96 96814 99 96839
rect 109 96819 110 96839
rect 119 96829 126 96839
rect 76 96805 110 96809
rect 170 96805 172 96855
rect 186 96837 190 96871
rect 216 96837 220 96871
rect 186 96760 220 96794
rect 282 96791 292 96903
rect 318 96896 335 96906
rect 318 96827 324 96896
rect 346 96827 348 96912
rect 428 96869 430 96916
rect 476 96879 480 96947
rect 485 96929 495 96957
rect 505 96957 519 96963
rect 544 96957 555 96995
rect 505 96929 525 96957
rect 544 96929 553 96957
rect 544 96909 548 96929
rect 579 96888 582 96978
rect 612 96960 624 96961
rect 599 96958 649 96960
rect 612 96957 624 96958
rect 610 96950 632 96957
rect 607 96949 632 96950
rect 586 96942 644 96949
rect 607 96941 644 96942
rect 607 96925 610 96941
rect 616 96925 644 96941
rect 607 96924 644 96925
rect 586 96917 644 96924
rect 607 96916 610 96917
rect 612 96909 632 96917
rect 612 96905 624 96909
rect 649 96908 651 96958
rect 544 96871 548 96879
rect 400 96839 408 96869
rect 420 96839 436 96869
rect 400 96835 436 96839
rect 400 96827 430 96835
rect 428 96811 430 96827
rect 476 96799 480 96867
rect 544 96837 552 96871
rect 578 96837 582 96871
rect 544 96829 548 96837
rect 544 96799 586 96800
rect 288 96759 292 96791
rect 296 96789 368 96797
rect 378 96789 450 96797
rect 544 96792 548 96799
rect 439 96761 444 96789
rect 120 96745 170 96747
rect 76 96741 130 96745
rect 110 96736 130 96741
rect 60 96711 67 96721
rect 76 96711 77 96731
rect 96 96702 99 96736
rect 109 96711 110 96731
rect 119 96711 126 96721
rect 76 96695 92 96701
rect 94 96695 110 96701
rect 170 96695 172 96745
rect 186 96679 190 96713
rect 216 96679 220 96713
rect 213 96647 224 96679
rect 282 96675 292 96759
rect 296 96753 368 96761
rect 378 96753 450 96761
rect 468 96758 473 96792
rect 428 96723 430 96739
rect 251 96647 292 96675
rect 318 96654 324 96723
rect 12 96642 62 96644
rect 28 96633 59 96641
rect 62 96633 64 96642
rect 251 96641 263 96647
rect 28 96625 64 96633
rect 127 96633 158 96641
rect 127 96626 182 96633
rect 127 96625 161 96626
rect 59 96609 64 96625
rect 158 96609 161 96625
rect 253 96613 263 96641
rect 273 96613 293 96647
rect 318 96644 335 96654
rect 303 96628 316 96638
rect 318 96628 324 96644
rect 346 96638 348 96723
rect 400 96715 430 96723
rect 476 96721 480 96789
rect 511 96758 582 96792
rect 544 96751 548 96758
rect 400 96711 436 96715
rect 400 96681 408 96711
rect 420 96681 436 96711
rect 544 96713 548 96721
rect 28 96601 64 96609
rect 127 96608 161 96609
rect 127 96601 182 96608
rect 62 96592 64 96601
rect 282 96555 292 96613
rect 295 96604 324 96628
rect 333 96628 353 96638
rect 428 96634 430 96681
rect 476 96641 480 96709
rect 544 96679 552 96713
rect 578 96679 582 96713
rect 544 96671 548 96679
rect 367 96628 380 96634
rect 333 96604 380 96628
rect 318 96591 324 96604
rect 346 96591 348 96604
rect 367 96600 380 96604
rect 396 96600 408 96634
rect 420 96600 436 96634
rect 544 96631 553 96659
rect 319 96580 346 96591
rect 120 96539 170 96541
rect 76 96533 92 96539
rect 94 96533 110 96539
rect 76 96523 99 96532
rect 60 96513 67 96523
rect 76 96503 77 96523
rect 96 96498 99 96523
rect 109 96503 110 96523
rect 119 96513 126 96523
rect 76 96489 110 96493
rect 170 96489 172 96539
rect 186 96521 190 96555
rect 216 96521 220 96555
rect 182 96483 224 96484
rect 186 96459 220 96476
rect 223 96459 257 96476
rect 182 96442 257 96459
rect 182 96441 224 96442
rect 160 96435 246 96441
rect 288 96435 292 96555
rect 296 96553 368 96561
rect 428 96553 430 96600
rect 476 96563 480 96631
rect 485 96587 495 96621
rect 505 96593 525 96621
rect 505 96587 519 96593
rect 544 96587 555 96631
rect 485 96563 492 96587
rect 579 96572 582 96662
rect 612 96644 624 96645
rect 599 96642 649 96644
rect 612 96641 624 96642
rect 610 96634 632 96641
rect 607 96633 632 96634
rect 586 96626 644 96633
rect 607 96625 644 96626
rect 607 96609 610 96625
rect 616 96609 644 96625
rect 607 96608 644 96609
rect 586 96601 644 96608
rect 607 96600 610 96601
rect 612 96593 632 96601
rect 612 96589 624 96593
rect 649 96592 651 96642
rect 544 96555 548 96563
rect 400 96523 408 96553
rect 420 96523 436 96553
rect 400 96519 436 96523
rect 400 96511 430 96519
rect 428 96495 430 96511
rect 476 96483 480 96551
rect 544 96521 552 96555
rect 578 96521 582 96555
rect 544 96513 548 96521
rect 295 96442 300 96476
rect 324 96442 329 96476
rect 378 96473 450 96481
rect 544 96478 548 96483
rect 544 96474 582 96478
rect 544 96459 552 96474
rect 578 96459 582 96474
rect 544 96441 586 96459
rect 522 96435 608 96441
rect 182 96419 224 96435
rect 544 96419 586 96435
rect 17 96405 67 96407
rect 119 96405 169 96407
rect 186 96405 220 96419
rect 548 96405 582 96419
rect 599 96405 649 96407
rect 42 96363 59 96397
rect 67 96355 69 96405
rect 160 96397 246 96405
rect 522 96397 608 96405
rect 76 96363 110 96397
rect 127 96363 144 96397
rect 152 96363 161 96397
rect 162 96395 195 96397
rect 224 96395 244 96397
rect 162 96363 244 96395
rect 524 96395 548 96397
rect 573 96395 582 96397
rect 586 96395 606 96397
rect 160 96355 246 96363
rect 186 96339 220 96355
rect 182 96325 224 96326
rect 160 96319 182 96325
rect 224 96319 246 96325
rect 186 96284 220 96318
rect 223 96284 257 96318
rect 120 96271 170 96273
rect 76 96267 130 96271
rect 110 96262 130 96267
rect 60 96237 67 96247
rect 76 96237 77 96257
rect 96 96228 99 96262
rect 109 96237 110 96257
rect 119 96237 126 96247
rect 76 96221 92 96227
rect 94 96221 110 96227
rect 170 96221 172 96271
rect 186 96205 190 96239
rect 216 96205 220 96239
rect 288 96205 292 96393
rect 476 96325 480 96393
rect 524 96363 606 96395
rect 607 96363 616 96397
rect 522 96355 608 96363
rect 649 96355 651 96405
rect 548 96339 582 96355
rect 522 96320 548 96325
rect 522 96319 582 96320
rect 586 96319 608 96325
rect 295 96284 300 96318
rect 324 96284 329 96318
rect 544 96316 582 96319
rect 378 96279 450 96287
rect 428 96249 430 96265
rect 400 96241 430 96249
rect 476 96247 480 96315
rect 544 96286 552 96316
rect 578 96286 582 96316
rect 544 96277 548 96286
rect 400 96237 436 96241
rect 400 96207 408 96237
rect 420 96207 436 96237
rect 544 96239 548 96247
rect 12 96168 62 96170
rect 28 96159 59 96167
rect 62 96159 64 96168
rect 28 96151 64 96159
rect 127 96159 158 96167
rect 127 96152 182 96159
rect 215 96157 224 96185
rect 127 96151 161 96152
rect 59 96135 64 96151
rect 158 96135 161 96151
rect 28 96127 64 96135
rect 127 96134 161 96135
rect 127 96127 182 96134
rect 62 96118 64 96127
rect 213 96119 224 96157
rect 282 96147 292 96205
rect 296 96199 368 96207
rect 319 96169 346 96180
rect 318 96156 324 96169
rect 346 96156 348 96169
rect 428 96160 430 96207
rect 443 96197 450 96199
rect 476 96167 480 96235
rect 544 96205 552 96239
rect 578 96205 582 96239
rect 481 96173 517 96201
rect 481 96167 495 96173
rect 367 96156 380 96160
rect 251 96113 263 96147
rect 273 96113 293 96147
rect 295 96132 324 96156
rect 303 96122 316 96132
rect 318 96116 324 96132
rect 333 96132 380 96156
rect 333 96122 353 96132
rect 367 96126 380 96132
rect 396 96126 408 96160
rect 420 96126 436 96160
rect 120 96065 170 96067
rect 76 96059 92 96065
rect 94 96059 110 96065
rect 76 96049 99 96058
rect 60 96039 67 96049
rect 76 96029 77 96049
rect 96 96024 99 96049
rect 109 96029 110 96049
rect 119 96039 126 96049
rect 76 96015 110 96019
rect 170 96015 172 96065
rect 186 96047 190 96081
rect 216 96047 220 96081
rect 186 95970 220 96004
rect 282 96001 292 96113
rect 318 96106 335 96116
rect 318 96037 324 96106
rect 346 96037 348 96122
rect 428 96079 430 96126
rect 476 96089 480 96157
rect 485 96139 495 96167
rect 505 96167 519 96173
rect 544 96167 555 96205
rect 505 96139 525 96167
rect 544 96139 553 96167
rect 544 96119 548 96139
rect 579 96098 582 96188
rect 612 96170 624 96171
rect 599 96168 649 96170
rect 612 96167 624 96168
rect 610 96160 632 96167
rect 607 96159 632 96160
rect 586 96152 644 96159
rect 607 96151 644 96152
rect 607 96135 610 96151
rect 616 96135 644 96151
rect 607 96134 644 96135
rect 586 96127 644 96134
rect 607 96126 610 96127
rect 612 96119 632 96127
rect 612 96115 624 96119
rect 649 96118 651 96168
rect 544 96081 548 96089
rect 400 96049 408 96079
rect 420 96049 436 96079
rect 400 96045 436 96049
rect 400 96037 430 96045
rect 428 96021 430 96037
rect 476 96009 480 96077
rect 544 96047 552 96081
rect 578 96047 582 96081
rect 544 96039 548 96047
rect 544 96009 586 96010
rect 288 95969 292 96001
rect 296 95999 368 96007
rect 378 95999 450 96007
rect 544 96002 548 96009
rect 439 95971 444 95999
rect 120 95955 170 95957
rect 76 95951 130 95955
rect 110 95946 130 95951
rect 60 95921 67 95931
rect 76 95921 77 95941
rect 96 95912 99 95946
rect 109 95921 110 95941
rect 119 95921 126 95931
rect 76 95905 92 95911
rect 94 95905 110 95911
rect 170 95905 172 95955
rect 186 95889 190 95923
rect 216 95889 220 95923
rect 213 95857 224 95889
rect 282 95885 292 95969
rect 296 95963 368 95971
rect 378 95963 450 95971
rect 468 95968 473 96002
rect 428 95933 430 95949
rect 251 95857 292 95885
rect 318 95864 324 95933
rect 12 95852 62 95854
rect 28 95843 59 95851
rect 62 95843 64 95852
rect 251 95851 263 95857
rect 28 95835 64 95843
rect 127 95843 158 95851
rect 127 95836 182 95843
rect 127 95835 161 95836
rect 59 95819 64 95835
rect 158 95819 161 95835
rect 253 95823 263 95851
rect 273 95823 293 95857
rect 318 95854 335 95864
rect 303 95838 316 95848
rect 318 95838 324 95854
rect 346 95848 348 95933
rect 400 95925 430 95933
rect 476 95931 480 95999
rect 511 95968 582 96002
rect 544 95961 548 95968
rect 400 95921 436 95925
rect 400 95891 408 95921
rect 420 95891 436 95921
rect 544 95923 548 95931
rect 28 95811 64 95819
rect 127 95818 161 95819
rect 127 95811 182 95818
rect 62 95802 64 95811
rect 282 95765 292 95823
rect 295 95814 324 95838
rect 333 95838 353 95848
rect 428 95844 430 95891
rect 476 95851 480 95919
rect 544 95889 552 95923
rect 578 95889 582 95923
rect 544 95881 548 95889
rect 367 95838 380 95844
rect 333 95814 380 95838
rect 318 95801 324 95814
rect 346 95801 348 95814
rect 367 95810 380 95814
rect 396 95810 408 95844
rect 420 95810 436 95844
rect 544 95841 553 95869
rect 319 95790 346 95801
rect 120 95749 170 95751
rect 76 95743 92 95749
rect 94 95743 110 95749
rect 76 95733 99 95742
rect 60 95723 67 95733
rect 76 95713 77 95733
rect 96 95708 99 95733
rect 109 95713 110 95733
rect 119 95723 126 95733
rect 76 95699 110 95703
rect 170 95699 172 95749
rect 186 95731 190 95765
rect 216 95731 220 95765
rect 182 95693 224 95694
rect 186 95669 220 95686
rect 223 95669 257 95686
rect 182 95652 257 95669
rect 182 95651 224 95652
rect 160 95645 246 95651
rect 288 95645 292 95765
rect 296 95763 368 95771
rect 428 95763 430 95810
rect 476 95773 480 95841
rect 485 95797 495 95831
rect 505 95803 525 95831
rect 505 95797 519 95803
rect 544 95797 555 95841
rect 485 95773 492 95797
rect 579 95782 582 95872
rect 612 95854 624 95855
rect 599 95852 649 95854
rect 612 95851 624 95852
rect 610 95844 632 95851
rect 607 95843 632 95844
rect 586 95836 644 95843
rect 607 95835 644 95836
rect 607 95819 610 95835
rect 616 95819 644 95835
rect 607 95818 644 95819
rect 586 95811 644 95818
rect 607 95810 610 95811
rect 612 95803 632 95811
rect 612 95799 624 95803
rect 649 95802 651 95852
rect 544 95765 548 95773
rect 400 95733 408 95763
rect 420 95733 436 95763
rect 400 95729 436 95733
rect 400 95721 430 95729
rect 428 95705 430 95721
rect 476 95693 480 95761
rect 544 95731 552 95765
rect 578 95731 582 95765
rect 544 95723 548 95731
rect 295 95652 300 95686
rect 324 95652 329 95686
rect 378 95683 450 95691
rect 544 95688 548 95693
rect 544 95684 582 95688
rect 544 95669 552 95684
rect 578 95669 582 95684
rect 544 95651 586 95669
rect 522 95645 608 95651
rect 182 95629 224 95645
rect 544 95629 586 95645
rect 17 95615 67 95617
rect 119 95615 169 95617
rect 186 95615 220 95629
rect 548 95615 582 95629
rect 599 95615 649 95617
rect 42 95573 59 95607
rect 67 95565 69 95615
rect 160 95607 246 95615
rect 522 95607 608 95615
rect 76 95573 110 95607
rect 127 95573 144 95607
rect 152 95573 161 95607
rect 162 95605 195 95607
rect 224 95605 244 95607
rect 162 95573 244 95605
rect 524 95605 548 95607
rect 573 95605 582 95607
rect 586 95605 606 95607
rect 160 95565 246 95573
rect 186 95549 220 95565
rect 182 95535 224 95536
rect 160 95529 182 95535
rect 224 95529 246 95535
rect 186 95494 220 95528
rect 223 95494 257 95528
rect 120 95481 170 95483
rect 76 95477 130 95481
rect 110 95472 130 95477
rect 60 95447 67 95457
rect 76 95447 77 95467
rect 96 95438 99 95472
rect 109 95447 110 95467
rect 119 95447 126 95457
rect 76 95431 92 95437
rect 94 95431 110 95437
rect 170 95431 172 95481
rect 186 95415 190 95449
rect 216 95415 220 95449
rect 288 95415 292 95603
rect 476 95535 480 95603
rect 524 95573 606 95605
rect 607 95573 616 95607
rect 522 95565 608 95573
rect 649 95565 651 95615
rect 548 95549 582 95565
rect 522 95530 548 95535
rect 522 95529 582 95530
rect 586 95529 608 95535
rect 295 95494 300 95528
rect 324 95494 329 95528
rect 544 95526 582 95529
rect 378 95489 450 95497
rect 428 95459 430 95475
rect 400 95451 430 95459
rect 476 95457 480 95525
rect 544 95496 552 95526
rect 578 95496 582 95526
rect 544 95487 548 95496
rect 400 95447 436 95451
rect 400 95417 408 95447
rect 420 95417 436 95447
rect 544 95449 548 95457
rect 12 95378 62 95380
rect 28 95369 59 95377
rect 62 95369 64 95378
rect 28 95361 64 95369
rect 127 95369 158 95377
rect 127 95362 182 95369
rect 215 95367 224 95395
rect 127 95361 161 95362
rect 59 95345 64 95361
rect 158 95345 161 95361
rect 28 95337 64 95345
rect 127 95344 161 95345
rect 127 95337 182 95344
rect 62 95328 64 95337
rect 213 95329 224 95367
rect 282 95357 292 95415
rect 296 95409 368 95417
rect 319 95379 346 95390
rect 318 95366 324 95379
rect 346 95366 348 95379
rect 428 95370 430 95417
rect 443 95407 450 95409
rect 476 95377 480 95445
rect 544 95415 552 95449
rect 578 95415 582 95449
rect 481 95383 517 95411
rect 481 95377 495 95383
rect 367 95366 380 95370
rect 251 95323 263 95357
rect 273 95323 293 95357
rect 295 95342 324 95366
rect 303 95332 316 95342
rect 318 95326 324 95342
rect 333 95342 380 95366
rect 333 95332 353 95342
rect 367 95336 380 95342
rect 396 95336 408 95370
rect 420 95336 436 95370
rect 120 95275 170 95277
rect 76 95269 92 95275
rect 94 95269 110 95275
rect 76 95259 99 95268
rect 60 95249 67 95259
rect 76 95239 77 95259
rect 96 95234 99 95259
rect 109 95239 110 95259
rect 119 95249 126 95259
rect 76 95225 110 95229
rect 170 95225 172 95275
rect 186 95257 190 95291
rect 216 95257 220 95291
rect 186 95180 220 95214
rect 282 95211 292 95323
rect 318 95316 335 95326
rect 318 95247 324 95316
rect 346 95247 348 95332
rect 428 95289 430 95336
rect 476 95299 480 95367
rect 485 95349 495 95377
rect 505 95377 519 95383
rect 544 95377 555 95415
rect 505 95349 525 95377
rect 544 95349 553 95377
rect 544 95329 548 95349
rect 579 95308 582 95398
rect 612 95380 624 95381
rect 599 95378 649 95380
rect 612 95377 624 95378
rect 610 95370 632 95377
rect 607 95369 632 95370
rect 586 95362 644 95369
rect 607 95361 644 95362
rect 607 95345 610 95361
rect 616 95345 644 95361
rect 607 95344 644 95345
rect 586 95337 644 95344
rect 607 95336 610 95337
rect 612 95329 632 95337
rect 612 95325 624 95329
rect 649 95328 651 95378
rect 544 95291 548 95299
rect 400 95259 408 95289
rect 420 95259 436 95289
rect 400 95255 436 95259
rect 400 95247 430 95255
rect 428 95231 430 95247
rect 476 95219 480 95287
rect 544 95257 552 95291
rect 578 95257 582 95291
rect 544 95249 548 95257
rect 544 95219 586 95220
rect 288 95179 292 95211
rect 296 95209 368 95217
rect 378 95209 450 95217
rect 544 95212 548 95219
rect 439 95181 444 95209
rect 120 95165 170 95167
rect 76 95161 130 95165
rect 110 95156 130 95161
rect 60 95131 67 95141
rect 76 95131 77 95151
rect 96 95122 99 95156
rect 109 95131 110 95151
rect 119 95131 126 95141
rect 76 95115 92 95121
rect 94 95115 110 95121
rect 170 95115 172 95165
rect 186 95099 190 95133
rect 216 95099 220 95133
rect 213 95067 224 95099
rect 282 95095 292 95179
rect 296 95173 368 95181
rect 378 95173 450 95181
rect 468 95178 473 95212
rect 428 95143 430 95159
rect 251 95067 292 95095
rect 318 95074 324 95143
rect 12 95062 62 95064
rect 28 95053 59 95061
rect 62 95053 64 95062
rect 251 95061 263 95067
rect 28 95045 64 95053
rect 127 95053 158 95061
rect 127 95046 182 95053
rect 127 95045 161 95046
rect 59 95029 64 95045
rect 158 95029 161 95045
rect 253 95033 263 95061
rect 273 95033 293 95067
rect 318 95064 335 95074
rect 303 95048 316 95058
rect 318 95048 324 95064
rect 346 95058 348 95143
rect 400 95135 430 95143
rect 476 95141 480 95209
rect 511 95178 582 95212
rect 544 95171 548 95178
rect 400 95131 436 95135
rect 400 95101 408 95131
rect 420 95101 436 95131
rect 544 95133 548 95141
rect 28 95021 64 95029
rect 127 95028 161 95029
rect 127 95021 182 95028
rect 62 95012 64 95021
rect 282 94975 292 95033
rect 295 95024 324 95048
rect 333 95048 353 95058
rect 428 95054 430 95101
rect 476 95061 480 95129
rect 544 95099 552 95133
rect 578 95099 582 95133
rect 544 95091 548 95099
rect 367 95048 380 95054
rect 333 95024 380 95048
rect 318 95011 324 95024
rect 346 95011 348 95024
rect 367 95020 380 95024
rect 396 95020 408 95054
rect 420 95020 436 95054
rect 544 95051 553 95079
rect 319 95000 346 95011
rect 120 94959 170 94961
rect 76 94953 92 94959
rect 94 94953 110 94959
rect 76 94943 99 94952
rect 60 94933 67 94943
rect 76 94923 77 94943
rect 96 94918 99 94943
rect 109 94923 110 94943
rect 119 94933 126 94943
rect 76 94909 110 94913
rect 170 94909 172 94959
rect 186 94941 190 94975
rect 216 94941 220 94975
rect 182 94903 224 94904
rect 186 94879 220 94896
rect 223 94879 257 94896
rect 182 94862 257 94879
rect 182 94861 224 94862
rect 160 94855 246 94861
rect 288 94855 292 94975
rect 296 94973 368 94981
rect 428 94973 430 95020
rect 476 94983 480 95051
rect 485 95007 495 95041
rect 505 95013 525 95041
rect 505 95007 519 95013
rect 544 95007 555 95051
rect 485 94983 492 95007
rect 579 94992 582 95082
rect 612 95064 624 95065
rect 599 95062 649 95064
rect 612 95061 624 95062
rect 610 95054 632 95061
rect 607 95053 632 95054
rect 586 95046 644 95053
rect 607 95045 644 95046
rect 607 95029 610 95045
rect 616 95029 644 95045
rect 607 95028 644 95029
rect 586 95021 644 95028
rect 607 95020 610 95021
rect 612 95013 632 95021
rect 612 95009 624 95013
rect 649 95012 651 95062
rect 544 94975 548 94983
rect 400 94943 408 94973
rect 420 94943 436 94973
rect 400 94939 436 94943
rect 400 94931 430 94939
rect 428 94915 430 94931
rect 476 94903 480 94971
rect 544 94941 552 94975
rect 578 94941 582 94975
rect 544 94933 548 94941
rect 295 94862 300 94896
rect 324 94862 329 94896
rect 378 94893 450 94901
rect 544 94898 548 94903
rect 544 94894 582 94898
rect 544 94879 552 94894
rect 578 94879 582 94894
rect 544 94861 586 94879
rect 522 94855 608 94861
rect 182 94839 224 94855
rect 544 94839 586 94855
rect 17 94825 67 94827
rect 119 94825 169 94827
rect 186 94825 220 94839
rect 548 94825 582 94839
rect 599 94825 649 94827
rect 42 94783 59 94817
rect 67 94775 69 94825
rect 160 94817 246 94825
rect 522 94817 608 94825
rect 76 94783 110 94817
rect 127 94783 144 94817
rect 152 94783 161 94817
rect 162 94815 195 94817
rect 224 94815 244 94817
rect 162 94783 244 94815
rect 524 94815 548 94817
rect 573 94815 582 94817
rect 586 94815 606 94817
rect 160 94775 246 94783
rect 186 94759 220 94775
rect 182 94745 224 94746
rect 160 94739 182 94745
rect 224 94739 246 94745
rect 186 94704 220 94738
rect 223 94704 257 94738
rect 120 94691 170 94693
rect 76 94687 130 94691
rect 110 94682 130 94687
rect 60 94657 67 94667
rect 76 94657 77 94677
rect 96 94648 99 94682
rect 109 94657 110 94677
rect 119 94657 126 94667
rect 76 94641 92 94647
rect 94 94641 110 94647
rect 170 94641 172 94691
rect 186 94625 190 94659
rect 216 94625 220 94659
rect 288 94625 292 94813
rect 476 94745 480 94813
rect 524 94783 606 94815
rect 607 94783 616 94817
rect 522 94775 608 94783
rect 649 94775 651 94825
rect 548 94759 582 94775
rect 522 94740 548 94745
rect 522 94739 582 94740
rect 586 94739 608 94745
rect 295 94704 300 94738
rect 324 94704 329 94738
rect 544 94736 582 94739
rect 378 94699 450 94707
rect 428 94669 430 94685
rect 400 94661 430 94669
rect 476 94667 480 94735
rect 544 94706 552 94736
rect 578 94706 582 94736
rect 544 94697 548 94706
rect 400 94657 436 94661
rect 400 94627 408 94657
rect 420 94627 436 94657
rect 544 94659 548 94667
rect 12 94588 62 94590
rect 28 94579 59 94587
rect 62 94579 64 94588
rect 28 94571 64 94579
rect 127 94579 158 94587
rect 127 94572 182 94579
rect 215 94577 224 94605
rect 127 94571 161 94572
rect 59 94555 64 94571
rect 158 94555 161 94571
rect 28 94547 64 94555
rect 127 94554 161 94555
rect 127 94547 182 94554
rect 62 94538 64 94547
rect 213 94539 224 94577
rect 282 94567 292 94625
rect 296 94619 368 94627
rect 319 94589 346 94600
rect 318 94576 324 94589
rect 346 94576 348 94589
rect 428 94580 430 94627
rect 443 94617 450 94619
rect 476 94587 480 94655
rect 544 94625 552 94659
rect 578 94625 582 94659
rect 481 94593 517 94621
rect 481 94587 495 94593
rect 367 94576 380 94580
rect 251 94533 263 94567
rect 273 94533 293 94567
rect 295 94552 324 94576
rect 303 94542 316 94552
rect 318 94536 324 94552
rect 333 94552 380 94576
rect 333 94542 353 94552
rect 367 94546 380 94552
rect 396 94546 408 94580
rect 420 94546 436 94580
rect 120 94485 170 94487
rect 76 94479 92 94485
rect 94 94479 110 94485
rect 76 94469 99 94478
rect 60 94459 67 94469
rect 76 94449 77 94469
rect 96 94444 99 94469
rect 109 94449 110 94469
rect 119 94459 126 94469
rect 76 94435 110 94439
rect 170 94435 172 94485
rect 186 94467 190 94501
rect 216 94467 220 94501
rect 186 94390 220 94424
rect 282 94421 292 94533
rect 318 94526 335 94536
rect 318 94457 324 94526
rect 346 94457 348 94542
rect 428 94499 430 94546
rect 476 94509 480 94577
rect 485 94559 495 94587
rect 505 94587 519 94593
rect 544 94587 555 94625
rect 505 94559 525 94587
rect 544 94559 553 94587
rect 544 94539 548 94559
rect 579 94518 582 94608
rect 612 94590 624 94591
rect 599 94588 649 94590
rect 612 94587 624 94588
rect 610 94580 632 94587
rect 607 94579 632 94580
rect 586 94572 644 94579
rect 607 94571 644 94572
rect 607 94555 610 94571
rect 616 94555 644 94571
rect 607 94554 644 94555
rect 586 94547 644 94554
rect 607 94546 610 94547
rect 612 94539 632 94547
rect 612 94535 624 94539
rect 649 94538 651 94588
rect 544 94501 548 94509
rect 400 94469 408 94499
rect 420 94469 436 94499
rect 400 94465 436 94469
rect 400 94457 430 94465
rect 428 94441 430 94457
rect 476 94429 480 94497
rect 544 94467 552 94501
rect 578 94467 582 94501
rect 544 94459 548 94467
rect 544 94429 586 94430
rect 288 94389 292 94421
rect 296 94419 368 94427
rect 378 94419 450 94427
rect 544 94422 548 94429
rect 439 94391 444 94419
rect 120 94375 170 94377
rect 76 94371 130 94375
rect 110 94366 130 94371
rect 60 94341 67 94351
rect 76 94341 77 94361
rect 96 94332 99 94366
rect 109 94341 110 94361
rect 119 94341 126 94351
rect 76 94325 92 94331
rect 94 94325 110 94331
rect 170 94325 172 94375
rect 186 94309 190 94343
rect 216 94309 220 94343
rect 213 94277 224 94309
rect 282 94305 292 94389
rect 296 94383 368 94391
rect 378 94383 450 94391
rect 468 94388 473 94422
rect 428 94353 430 94369
rect 251 94277 292 94305
rect 318 94284 324 94353
rect 12 94272 62 94274
rect 28 94263 59 94271
rect 62 94263 64 94272
rect 251 94271 263 94277
rect 28 94255 64 94263
rect 127 94263 158 94271
rect 127 94256 182 94263
rect 127 94255 161 94256
rect 59 94239 64 94255
rect 158 94239 161 94255
rect 253 94243 263 94271
rect 273 94243 293 94277
rect 318 94274 335 94284
rect 303 94258 316 94268
rect 318 94258 324 94274
rect 346 94268 348 94353
rect 400 94345 430 94353
rect 476 94351 480 94419
rect 511 94388 582 94422
rect 544 94381 548 94388
rect 400 94341 436 94345
rect 400 94311 408 94341
rect 420 94311 436 94341
rect 544 94343 548 94351
rect 28 94231 64 94239
rect 127 94238 161 94239
rect 127 94231 182 94238
rect 62 94222 64 94231
rect 282 94185 292 94243
rect 295 94234 324 94258
rect 333 94258 353 94268
rect 428 94264 430 94311
rect 476 94271 480 94339
rect 544 94309 552 94343
rect 578 94309 582 94343
rect 544 94301 548 94309
rect 367 94258 380 94264
rect 333 94234 380 94258
rect 318 94221 324 94234
rect 346 94221 348 94234
rect 367 94230 380 94234
rect 396 94230 408 94264
rect 420 94230 436 94264
rect 544 94261 553 94289
rect 319 94210 346 94221
rect 120 94169 170 94171
rect 76 94163 92 94169
rect 94 94163 110 94169
rect 76 94153 99 94162
rect 60 94143 67 94153
rect 76 94133 77 94153
rect 96 94128 99 94153
rect 109 94133 110 94153
rect 119 94143 126 94153
rect 76 94119 110 94123
rect 170 94119 172 94169
rect 186 94151 190 94185
rect 216 94151 220 94185
rect 182 94113 224 94114
rect 186 94089 220 94106
rect 223 94089 257 94106
rect 182 94072 257 94089
rect 182 94071 224 94072
rect 160 94065 246 94071
rect 288 94065 292 94185
rect 296 94183 368 94191
rect 428 94183 430 94230
rect 476 94193 480 94261
rect 485 94217 495 94251
rect 505 94223 525 94251
rect 505 94217 519 94223
rect 544 94217 555 94261
rect 485 94193 492 94217
rect 579 94202 582 94292
rect 612 94274 624 94275
rect 599 94272 649 94274
rect 612 94271 624 94272
rect 610 94264 632 94271
rect 607 94263 632 94264
rect 586 94256 644 94263
rect 607 94255 644 94256
rect 607 94239 610 94255
rect 616 94239 644 94255
rect 607 94238 644 94239
rect 586 94231 644 94238
rect 607 94230 610 94231
rect 612 94223 632 94231
rect 612 94219 624 94223
rect 649 94222 651 94272
rect 544 94185 548 94193
rect 400 94153 408 94183
rect 420 94153 436 94183
rect 400 94149 436 94153
rect 400 94141 430 94149
rect 428 94125 430 94141
rect 476 94113 480 94181
rect 544 94151 552 94185
rect 578 94151 582 94185
rect 544 94143 548 94151
rect 295 94072 300 94106
rect 324 94072 329 94106
rect 378 94103 450 94111
rect 544 94108 548 94113
rect 544 94104 582 94108
rect 544 94089 552 94104
rect 578 94089 582 94104
rect 544 94071 586 94089
rect 522 94065 608 94071
rect 182 94049 224 94065
rect 544 94049 586 94065
rect 17 94035 67 94037
rect 119 94035 169 94037
rect 186 94035 220 94049
rect 548 94035 582 94049
rect 599 94035 649 94037
rect 42 93993 59 94027
rect 67 93985 69 94035
rect 160 94027 246 94035
rect 522 94027 608 94035
rect 76 93993 110 94027
rect 127 93993 144 94027
rect 152 93993 161 94027
rect 162 94025 195 94027
rect 224 94025 244 94027
rect 162 93993 244 94025
rect 524 94025 548 94027
rect 573 94025 582 94027
rect 586 94025 606 94027
rect 160 93985 246 93993
rect 186 93969 220 93985
rect 182 93955 224 93956
rect 160 93949 182 93955
rect 224 93949 246 93955
rect 186 93914 220 93948
rect 223 93914 257 93948
rect 120 93901 170 93903
rect 76 93897 130 93901
rect 110 93892 130 93897
rect 60 93867 67 93877
rect 76 93867 77 93887
rect 96 93858 99 93892
rect 109 93867 110 93887
rect 119 93867 126 93877
rect 76 93851 92 93857
rect 94 93851 110 93857
rect 170 93851 172 93901
rect 186 93835 190 93869
rect 216 93835 220 93869
rect 288 93835 292 94023
rect 476 93955 480 94023
rect 524 93993 606 94025
rect 607 93993 616 94027
rect 522 93985 608 93993
rect 649 93985 651 94035
rect 548 93969 582 93985
rect 522 93950 548 93955
rect 522 93949 582 93950
rect 586 93949 608 93955
rect 295 93914 300 93948
rect 324 93914 329 93948
rect 544 93946 582 93949
rect 378 93909 450 93917
rect 428 93879 430 93895
rect 400 93871 430 93879
rect 476 93877 480 93945
rect 544 93916 552 93946
rect 578 93916 582 93946
rect 544 93907 548 93916
rect 400 93867 436 93871
rect 400 93837 408 93867
rect 420 93837 436 93867
rect 544 93869 548 93877
rect 12 93798 62 93800
rect 28 93789 59 93797
rect 62 93789 64 93798
rect 28 93781 64 93789
rect 127 93789 158 93797
rect 127 93782 182 93789
rect 215 93787 224 93815
rect 127 93781 161 93782
rect 59 93765 64 93781
rect 158 93765 161 93781
rect 28 93757 64 93765
rect 127 93764 161 93765
rect 127 93757 182 93764
rect 62 93748 64 93757
rect 213 93749 224 93787
rect 282 93777 292 93835
rect 296 93829 368 93837
rect 319 93799 346 93810
rect 318 93786 324 93799
rect 346 93786 348 93799
rect 428 93790 430 93837
rect 443 93827 450 93829
rect 476 93797 480 93865
rect 544 93835 552 93869
rect 578 93835 582 93869
rect 481 93803 517 93831
rect 481 93797 495 93803
rect 367 93786 380 93790
rect 251 93743 263 93777
rect 273 93743 293 93777
rect 295 93762 324 93786
rect 303 93752 316 93762
rect 318 93746 324 93762
rect 333 93762 380 93786
rect 333 93752 353 93762
rect 367 93756 380 93762
rect 396 93756 408 93790
rect 420 93756 436 93790
rect 120 93695 170 93697
rect 76 93689 92 93695
rect 94 93689 110 93695
rect 76 93679 99 93688
rect 60 93669 67 93679
rect 76 93659 77 93679
rect 96 93654 99 93679
rect 109 93659 110 93679
rect 119 93669 126 93679
rect 76 93645 110 93649
rect 170 93645 172 93695
rect 186 93677 190 93711
rect 216 93677 220 93711
rect 186 93600 220 93634
rect 282 93631 292 93743
rect 318 93736 335 93746
rect 318 93667 324 93736
rect 346 93667 348 93752
rect 428 93709 430 93756
rect 476 93719 480 93787
rect 485 93769 495 93797
rect 505 93797 519 93803
rect 544 93797 555 93835
rect 505 93769 525 93797
rect 544 93769 553 93797
rect 544 93749 548 93769
rect 579 93728 582 93818
rect 612 93800 624 93801
rect 599 93798 649 93800
rect 612 93797 624 93798
rect 610 93790 632 93797
rect 607 93789 632 93790
rect 586 93782 644 93789
rect 607 93781 644 93782
rect 607 93765 610 93781
rect 616 93765 644 93781
rect 607 93764 644 93765
rect 586 93757 644 93764
rect 607 93756 610 93757
rect 612 93749 632 93757
rect 612 93745 624 93749
rect 649 93748 651 93798
rect 544 93711 548 93719
rect 400 93679 408 93709
rect 420 93679 436 93709
rect 400 93675 436 93679
rect 400 93667 430 93675
rect 428 93651 430 93667
rect 476 93639 480 93707
rect 544 93677 552 93711
rect 578 93677 582 93711
rect 544 93669 548 93677
rect 544 93639 586 93640
rect 288 93599 292 93631
rect 296 93629 368 93637
rect 378 93629 450 93637
rect 544 93632 548 93639
rect 439 93601 444 93629
rect 120 93585 170 93587
rect 76 93581 130 93585
rect 110 93576 130 93581
rect 60 93551 67 93561
rect 76 93551 77 93571
rect 96 93542 99 93576
rect 109 93551 110 93571
rect 119 93551 126 93561
rect 76 93535 92 93541
rect 94 93535 110 93541
rect 170 93535 172 93585
rect 186 93519 190 93553
rect 216 93519 220 93553
rect 213 93487 224 93519
rect 282 93515 292 93599
rect 296 93593 368 93601
rect 378 93593 450 93601
rect 468 93598 473 93632
rect 428 93563 430 93579
rect 251 93487 292 93515
rect 318 93494 324 93563
rect 12 93482 62 93484
rect 28 93473 59 93481
rect 62 93473 64 93482
rect 251 93481 263 93487
rect 28 93465 64 93473
rect 127 93473 158 93481
rect 127 93466 182 93473
rect 127 93465 161 93466
rect 59 93449 64 93465
rect 158 93449 161 93465
rect 253 93453 263 93481
rect 273 93453 293 93487
rect 318 93484 335 93494
rect 303 93468 316 93478
rect 318 93468 324 93484
rect 346 93478 348 93563
rect 400 93555 430 93563
rect 476 93561 480 93629
rect 511 93598 582 93632
rect 544 93591 548 93598
rect 400 93551 436 93555
rect 400 93521 408 93551
rect 420 93521 436 93551
rect 544 93553 548 93561
rect 28 93441 64 93449
rect 127 93448 161 93449
rect 127 93441 182 93448
rect 62 93432 64 93441
rect 282 93395 292 93453
rect 295 93444 324 93468
rect 333 93468 353 93478
rect 428 93474 430 93521
rect 476 93481 480 93549
rect 544 93519 552 93553
rect 578 93519 582 93553
rect 544 93511 548 93519
rect 367 93468 380 93474
rect 333 93444 380 93468
rect 318 93431 324 93444
rect 346 93431 348 93444
rect 367 93440 380 93444
rect 396 93440 408 93474
rect 420 93440 436 93474
rect 544 93471 553 93499
rect 319 93420 346 93431
rect 120 93379 170 93381
rect 76 93373 92 93379
rect 94 93373 110 93379
rect 76 93363 99 93372
rect 60 93353 67 93363
rect 76 93343 77 93363
rect 96 93338 99 93363
rect 109 93343 110 93363
rect 119 93353 126 93363
rect 76 93329 110 93333
rect 170 93329 172 93379
rect 186 93361 190 93395
rect 216 93361 220 93395
rect 182 93323 224 93324
rect 186 93299 220 93316
rect 223 93299 257 93316
rect 182 93282 257 93299
rect 182 93281 224 93282
rect 160 93275 246 93281
rect 288 93275 292 93395
rect 296 93393 368 93401
rect 428 93393 430 93440
rect 476 93403 480 93471
rect 485 93427 495 93461
rect 505 93433 525 93461
rect 505 93427 519 93433
rect 544 93427 555 93471
rect 485 93403 492 93427
rect 579 93412 582 93502
rect 612 93484 624 93485
rect 599 93482 649 93484
rect 612 93481 624 93482
rect 610 93474 632 93481
rect 607 93473 632 93474
rect 586 93466 644 93473
rect 607 93465 644 93466
rect 607 93449 610 93465
rect 616 93449 644 93465
rect 607 93448 644 93449
rect 586 93441 644 93448
rect 607 93440 610 93441
rect 612 93433 632 93441
rect 612 93429 624 93433
rect 649 93432 651 93482
rect 544 93395 548 93403
rect 400 93363 408 93393
rect 420 93363 436 93393
rect 400 93359 436 93363
rect 400 93351 430 93359
rect 428 93335 430 93351
rect 476 93323 480 93391
rect 544 93361 552 93395
rect 578 93361 582 93395
rect 544 93353 548 93361
rect 295 93282 300 93316
rect 324 93282 329 93316
rect 378 93313 450 93321
rect 544 93318 548 93323
rect 544 93314 582 93318
rect 544 93299 552 93314
rect 578 93299 582 93314
rect 544 93281 586 93299
rect 522 93275 608 93281
rect 182 93259 224 93275
rect 544 93259 586 93275
rect 17 93245 67 93247
rect 119 93245 169 93247
rect 186 93245 220 93259
rect 548 93245 582 93259
rect 599 93245 649 93247
rect 42 93203 59 93237
rect 67 93195 69 93245
rect 160 93237 246 93245
rect 522 93237 608 93245
rect 76 93203 110 93237
rect 127 93203 144 93237
rect 152 93203 161 93237
rect 162 93235 195 93237
rect 224 93235 244 93237
rect 162 93203 244 93235
rect 524 93235 548 93237
rect 573 93235 582 93237
rect 586 93235 606 93237
rect 160 93195 246 93203
rect 186 93179 220 93195
rect 182 93165 224 93166
rect 160 93159 182 93165
rect 224 93159 246 93165
rect 186 93124 220 93158
rect 223 93124 257 93158
rect 120 93111 170 93113
rect 76 93107 130 93111
rect 110 93102 130 93107
rect 60 93077 67 93087
rect 76 93077 77 93097
rect 96 93068 99 93102
rect 109 93077 110 93097
rect 119 93077 126 93087
rect 76 93061 92 93067
rect 94 93061 110 93067
rect 170 93061 172 93111
rect 186 93045 190 93079
rect 216 93045 220 93079
rect 288 93045 292 93233
rect 476 93165 480 93233
rect 524 93203 606 93235
rect 607 93203 616 93237
rect 522 93195 608 93203
rect 649 93195 651 93245
rect 548 93179 582 93195
rect 522 93160 548 93165
rect 522 93159 582 93160
rect 586 93159 608 93165
rect 295 93124 300 93158
rect 324 93124 329 93158
rect 544 93156 582 93159
rect 378 93119 450 93127
rect 428 93089 430 93105
rect 400 93081 430 93089
rect 476 93087 480 93155
rect 544 93126 552 93156
rect 578 93126 582 93156
rect 544 93117 548 93126
rect 400 93077 436 93081
rect 400 93047 408 93077
rect 420 93047 436 93077
rect 544 93079 548 93087
rect 12 93008 62 93010
rect 28 92999 59 93007
rect 62 92999 64 93008
rect 28 92991 64 92999
rect 127 92999 158 93007
rect 127 92992 182 92999
rect 215 92997 224 93025
rect 127 92991 161 92992
rect 59 92975 64 92991
rect 158 92975 161 92991
rect 28 92967 64 92975
rect 127 92974 161 92975
rect 127 92967 182 92974
rect 62 92958 64 92967
rect 213 92959 224 92997
rect 282 92987 292 93045
rect 296 93039 368 93047
rect 319 93009 346 93020
rect 318 92996 324 93009
rect 346 92996 348 93009
rect 428 93000 430 93047
rect 443 93037 450 93039
rect 476 93007 480 93075
rect 544 93045 552 93079
rect 578 93045 582 93079
rect 481 93013 517 93041
rect 481 93007 495 93013
rect 367 92996 380 93000
rect 251 92953 263 92987
rect 273 92953 293 92987
rect 295 92972 324 92996
rect 303 92962 316 92972
rect 318 92956 324 92972
rect 333 92972 380 92996
rect 333 92962 353 92972
rect 367 92966 380 92972
rect 396 92966 408 93000
rect 420 92966 436 93000
rect 120 92905 170 92907
rect 76 92899 92 92905
rect 94 92899 110 92905
rect 76 92889 99 92898
rect 60 92879 67 92889
rect 76 92869 77 92889
rect 96 92864 99 92889
rect 109 92869 110 92889
rect 119 92879 126 92889
rect 76 92855 110 92859
rect 170 92855 172 92905
rect 186 92887 190 92921
rect 216 92887 220 92921
rect 186 92810 220 92844
rect 282 92841 292 92953
rect 318 92946 335 92956
rect 318 92877 324 92946
rect 346 92877 348 92962
rect 428 92919 430 92966
rect 476 92929 480 92997
rect 485 92979 495 93007
rect 505 93007 519 93013
rect 544 93007 555 93045
rect 505 92979 525 93007
rect 544 92979 553 93007
rect 544 92959 548 92979
rect 579 92938 582 93028
rect 612 93010 624 93011
rect 599 93008 649 93010
rect 612 93007 624 93008
rect 610 93000 632 93007
rect 607 92999 632 93000
rect 586 92992 644 92999
rect 607 92991 644 92992
rect 607 92975 610 92991
rect 616 92975 644 92991
rect 607 92974 644 92975
rect 586 92967 644 92974
rect 607 92966 610 92967
rect 612 92959 632 92967
rect 612 92955 624 92959
rect 649 92958 651 93008
rect 544 92921 548 92929
rect 400 92889 408 92919
rect 420 92889 436 92919
rect 400 92885 436 92889
rect 400 92877 430 92885
rect 428 92861 430 92877
rect 476 92849 480 92917
rect 544 92887 552 92921
rect 578 92887 582 92921
rect 544 92879 548 92887
rect 544 92849 586 92850
rect 288 92809 292 92841
rect 296 92839 368 92847
rect 378 92839 450 92847
rect 544 92842 548 92849
rect 439 92811 444 92839
rect 120 92795 170 92797
rect 76 92791 130 92795
rect 110 92786 130 92791
rect 60 92761 67 92771
rect 76 92761 77 92781
rect 96 92752 99 92786
rect 109 92761 110 92781
rect 119 92761 126 92771
rect 76 92745 92 92751
rect 94 92745 110 92751
rect 170 92745 172 92795
rect 186 92729 190 92763
rect 216 92729 220 92763
rect 213 92697 224 92729
rect 282 92725 292 92809
rect 296 92803 368 92811
rect 378 92803 450 92811
rect 468 92808 473 92842
rect 428 92773 430 92789
rect 251 92697 292 92725
rect 318 92704 324 92773
rect 12 92692 62 92694
rect 28 92683 59 92691
rect 62 92683 64 92692
rect 251 92691 263 92697
rect 28 92675 64 92683
rect 127 92683 158 92691
rect 127 92676 182 92683
rect 127 92675 161 92676
rect 59 92659 64 92675
rect 158 92659 161 92675
rect 253 92663 263 92691
rect 273 92663 293 92697
rect 318 92694 335 92704
rect 303 92678 316 92688
rect 318 92678 324 92694
rect 346 92688 348 92773
rect 400 92765 430 92773
rect 476 92771 480 92839
rect 511 92808 582 92842
rect 544 92801 548 92808
rect 400 92761 436 92765
rect 400 92731 408 92761
rect 420 92731 436 92761
rect 544 92763 548 92771
rect 28 92651 64 92659
rect 127 92658 161 92659
rect 127 92651 182 92658
rect 62 92642 64 92651
rect 282 92605 292 92663
rect 295 92654 324 92678
rect 333 92678 353 92688
rect 428 92684 430 92731
rect 476 92691 480 92759
rect 544 92729 552 92763
rect 578 92729 582 92763
rect 544 92721 548 92729
rect 367 92678 380 92684
rect 333 92654 380 92678
rect 318 92641 324 92654
rect 346 92641 348 92654
rect 367 92650 380 92654
rect 396 92650 408 92684
rect 420 92650 436 92684
rect 544 92681 553 92709
rect 319 92630 346 92641
rect 120 92589 170 92591
rect 76 92583 92 92589
rect 94 92583 110 92589
rect 76 92573 99 92582
rect 60 92563 67 92573
rect 76 92553 77 92573
rect 96 92548 99 92573
rect 109 92553 110 92573
rect 119 92563 126 92573
rect 76 92539 110 92543
rect 170 92539 172 92589
rect 186 92571 190 92605
rect 216 92571 220 92605
rect 182 92533 224 92534
rect 186 92509 220 92526
rect 223 92509 257 92526
rect 182 92492 257 92509
rect 182 92491 224 92492
rect 160 92485 246 92491
rect 288 92485 292 92605
rect 296 92603 368 92611
rect 428 92603 430 92650
rect 476 92613 480 92681
rect 485 92637 495 92671
rect 505 92643 525 92671
rect 505 92637 519 92643
rect 544 92637 555 92681
rect 485 92613 492 92637
rect 579 92622 582 92712
rect 612 92694 624 92695
rect 599 92692 649 92694
rect 612 92691 624 92692
rect 610 92684 632 92691
rect 607 92683 632 92684
rect 586 92676 644 92683
rect 607 92675 644 92676
rect 607 92659 610 92675
rect 616 92659 644 92675
rect 607 92658 644 92659
rect 586 92651 644 92658
rect 607 92650 610 92651
rect 612 92643 632 92651
rect 612 92639 624 92643
rect 649 92642 651 92692
rect 544 92605 548 92613
rect 400 92573 408 92603
rect 420 92573 436 92603
rect 400 92569 436 92573
rect 400 92561 430 92569
rect 428 92545 430 92561
rect 476 92533 480 92601
rect 544 92571 552 92605
rect 578 92571 582 92605
rect 544 92563 548 92571
rect 295 92492 300 92526
rect 324 92492 329 92526
rect 378 92523 450 92531
rect 544 92528 548 92533
rect 544 92524 582 92528
rect 544 92509 552 92524
rect 578 92509 582 92524
rect 544 92491 586 92509
rect 522 92485 608 92491
rect 182 92469 224 92485
rect 544 92469 586 92485
rect 17 92455 67 92457
rect 119 92455 169 92457
rect 186 92455 220 92469
rect 548 92455 582 92469
rect 599 92455 649 92457
rect 42 92413 59 92447
rect 67 92405 69 92455
rect 160 92447 246 92455
rect 522 92447 608 92455
rect 76 92413 110 92447
rect 127 92413 144 92447
rect 152 92413 161 92447
rect 162 92445 195 92447
rect 224 92445 244 92447
rect 162 92413 244 92445
rect 524 92445 548 92447
rect 573 92445 582 92447
rect 586 92445 606 92447
rect 160 92405 246 92413
rect 186 92389 220 92405
rect 182 92375 224 92376
rect 160 92369 182 92375
rect 224 92369 246 92375
rect 186 92334 220 92368
rect 223 92334 257 92368
rect 120 92321 170 92323
rect 76 92317 130 92321
rect 110 92312 130 92317
rect 60 92287 67 92297
rect 76 92287 77 92307
rect 96 92278 99 92312
rect 109 92287 110 92307
rect 119 92287 126 92297
rect 76 92271 92 92277
rect 94 92271 110 92277
rect 170 92271 172 92321
rect 186 92255 190 92289
rect 216 92255 220 92289
rect 288 92255 292 92443
rect 476 92375 480 92443
rect 524 92413 606 92445
rect 607 92413 616 92447
rect 522 92405 608 92413
rect 649 92405 651 92455
rect 548 92389 582 92405
rect 522 92370 548 92375
rect 522 92369 582 92370
rect 586 92369 608 92375
rect 295 92334 300 92368
rect 324 92334 329 92368
rect 544 92366 582 92369
rect 378 92329 450 92337
rect 428 92299 430 92315
rect 400 92291 430 92299
rect 476 92297 480 92365
rect 544 92336 552 92366
rect 578 92336 582 92366
rect 544 92327 548 92336
rect 400 92287 436 92291
rect 400 92257 408 92287
rect 420 92257 436 92287
rect 544 92289 548 92297
rect 12 92218 62 92220
rect 28 92209 59 92217
rect 62 92209 64 92218
rect 28 92201 64 92209
rect 127 92209 158 92217
rect 127 92202 182 92209
rect 215 92207 224 92235
rect 127 92201 161 92202
rect 59 92185 64 92201
rect 158 92185 161 92201
rect 28 92177 64 92185
rect 127 92184 161 92185
rect 127 92177 182 92184
rect 62 92168 64 92177
rect 213 92169 224 92207
rect 282 92197 292 92255
rect 296 92249 368 92257
rect 319 92219 346 92230
rect 318 92206 324 92219
rect 346 92206 348 92219
rect 428 92210 430 92257
rect 443 92247 450 92249
rect 476 92217 480 92285
rect 544 92255 552 92289
rect 578 92255 582 92289
rect 481 92223 517 92251
rect 481 92217 495 92223
rect 367 92206 380 92210
rect 251 92163 263 92197
rect 273 92163 293 92197
rect 295 92182 324 92206
rect 303 92172 316 92182
rect 318 92166 324 92182
rect 333 92182 380 92206
rect 333 92172 353 92182
rect 367 92176 380 92182
rect 396 92176 408 92210
rect 420 92176 436 92210
rect 120 92115 170 92117
rect 76 92109 92 92115
rect 94 92109 110 92115
rect 76 92099 99 92108
rect 60 92089 67 92099
rect 76 92079 77 92099
rect 96 92074 99 92099
rect 109 92079 110 92099
rect 119 92089 126 92099
rect 76 92065 110 92069
rect 170 92065 172 92115
rect 186 92097 190 92131
rect 216 92097 220 92131
rect 186 92020 220 92054
rect 282 92051 292 92163
rect 318 92156 335 92166
rect 318 92087 324 92156
rect 346 92087 348 92172
rect 428 92129 430 92176
rect 476 92139 480 92207
rect 485 92189 495 92217
rect 505 92217 519 92223
rect 544 92217 555 92255
rect 505 92189 525 92217
rect 544 92189 553 92217
rect 544 92169 548 92189
rect 579 92148 582 92238
rect 612 92220 624 92221
rect 599 92218 649 92220
rect 612 92217 624 92218
rect 610 92210 632 92217
rect 607 92209 632 92210
rect 586 92202 644 92209
rect 607 92201 644 92202
rect 607 92185 610 92201
rect 616 92185 644 92201
rect 607 92184 644 92185
rect 586 92177 644 92184
rect 607 92176 610 92177
rect 612 92169 632 92177
rect 612 92165 624 92169
rect 649 92168 651 92218
rect 544 92131 548 92139
rect 400 92099 408 92129
rect 420 92099 436 92129
rect 400 92095 436 92099
rect 400 92087 430 92095
rect 428 92071 430 92087
rect 476 92059 480 92127
rect 544 92097 552 92131
rect 578 92097 582 92131
rect 544 92089 548 92097
rect 544 92059 586 92060
rect 288 92019 292 92051
rect 296 92049 368 92057
rect 378 92049 450 92057
rect 544 92052 548 92059
rect 439 92021 444 92049
rect 120 92005 170 92007
rect 76 92001 130 92005
rect 110 91996 130 92001
rect 60 91971 67 91981
rect 76 91971 77 91991
rect 96 91962 99 91996
rect 109 91971 110 91991
rect 119 91971 126 91981
rect 76 91955 92 91961
rect 94 91955 110 91961
rect 170 91955 172 92005
rect 186 91939 190 91973
rect 216 91939 220 91973
rect 213 91907 224 91939
rect 282 91935 292 92019
rect 296 92013 368 92021
rect 378 92013 450 92021
rect 468 92018 473 92052
rect 428 91983 430 91999
rect 251 91907 292 91935
rect 318 91914 324 91983
rect 12 91902 62 91904
rect 28 91893 59 91901
rect 62 91893 64 91902
rect 251 91901 263 91907
rect 28 91885 64 91893
rect 127 91893 158 91901
rect 127 91886 182 91893
rect 127 91885 161 91886
rect 59 91869 64 91885
rect 158 91869 161 91885
rect 253 91873 263 91901
rect 273 91873 293 91907
rect 318 91904 335 91914
rect 303 91888 316 91898
rect 318 91888 324 91904
rect 346 91898 348 91983
rect 400 91975 430 91983
rect 476 91981 480 92049
rect 511 92018 582 92052
rect 544 92011 548 92018
rect 400 91971 436 91975
rect 400 91941 408 91971
rect 420 91941 436 91971
rect 544 91973 548 91981
rect 28 91861 64 91869
rect 127 91868 161 91869
rect 127 91861 182 91868
rect 62 91852 64 91861
rect 282 91815 292 91873
rect 295 91864 324 91888
rect 333 91888 353 91898
rect 428 91894 430 91941
rect 476 91901 480 91969
rect 544 91939 552 91973
rect 578 91939 582 91973
rect 544 91931 548 91939
rect 367 91888 380 91894
rect 333 91864 380 91888
rect 318 91851 324 91864
rect 346 91851 348 91864
rect 367 91860 380 91864
rect 396 91860 408 91894
rect 420 91860 436 91894
rect 544 91891 553 91919
rect 319 91840 346 91851
rect 120 91799 170 91801
rect 76 91793 92 91799
rect 94 91793 110 91799
rect 76 91783 99 91792
rect 60 91773 67 91783
rect 76 91763 77 91783
rect 96 91758 99 91783
rect 109 91763 110 91783
rect 119 91773 126 91783
rect 76 91749 110 91753
rect 170 91749 172 91799
rect 186 91781 190 91815
rect 216 91781 220 91815
rect 182 91743 224 91744
rect 186 91719 220 91736
rect 223 91719 257 91736
rect 182 91702 257 91719
rect 182 91701 224 91702
rect 160 91695 246 91701
rect 288 91695 292 91815
rect 296 91813 368 91821
rect 428 91813 430 91860
rect 476 91823 480 91891
rect 485 91847 495 91881
rect 505 91853 525 91881
rect 505 91847 519 91853
rect 544 91847 555 91891
rect 485 91823 492 91847
rect 579 91832 582 91922
rect 612 91904 624 91905
rect 599 91902 649 91904
rect 612 91901 624 91902
rect 610 91894 632 91901
rect 607 91893 632 91894
rect 586 91886 644 91893
rect 607 91885 644 91886
rect 607 91869 610 91885
rect 616 91869 644 91885
rect 607 91868 644 91869
rect 586 91861 644 91868
rect 607 91860 610 91861
rect 612 91853 632 91861
rect 612 91849 624 91853
rect 649 91852 651 91902
rect 544 91815 548 91823
rect 400 91783 408 91813
rect 420 91783 436 91813
rect 400 91779 436 91783
rect 400 91771 430 91779
rect 428 91755 430 91771
rect 476 91743 480 91811
rect 544 91781 552 91815
rect 578 91781 582 91815
rect 544 91773 548 91781
rect 295 91702 300 91736
rect 324 91702 329 91736
rect 378 91733 450 91741
rect 544 91738 548 91743
rect 544 91734 582 91738
rect 544 91719 552 91734
rect 578 91719 582 91734
rect 544 91701 586 91719
rect 522 91695 608 91701
rect 182 91679 224 91695
rect 544 91679 586 91695
rect 17 91665 67 91667
rect 119 91665 169 91667
rect 186 91665 220 91679
rect 548 91665 582 91679
rect 599 91665 649 91667
rect 42 91623 59 91657
rect 67 91615 69 91665
rect 160 91657 246 91665
rect 522 91657 608 91665
rect 76 91623 110 91657
rect 127 91623 144 91657
rect 152 91623 161 91657
rect 162 91655 195 91657
rect 224 91655 244 91657
rect 162 91623 244 91655
rect 524 91655 548 91657
rect 573 91655 582 91657
rect 586 91655 606 91657
rect 160 91615 246 91623
rect 186 91599 220 91615
rect 182 91585 224 91586
rect 160 91579 182 91585
rect 224 91579 246 91585
rect 186 91544 220 91578
rect 223 91544 257 91578
rect 120 91531 170 91533
rect 76 91527 130 91531
rect 110 91522 130 91527
rect 60 91497 67 91507
rect 76 91497 77 91517
rect 96 91488 99 91522
rect 109 91497 110 91517
rect 119 91497 126 91507
rect 76 91481 92 91487
rect 94 91481 110 91487
rect 170 91481 172 91531
rect 186 91465 190 91499
rect 216 91465 220 91499
rect 288 91465 292 91653
rect 476 91585 480 91653
rect 524 91623 606 91655
rect 607 91623 616 91657
rect 522 91615 608 91623
rect 649 91615 651 91665
rect 548 91599 582 91615
rect 522 91580 548 91585
rect 522 91579 582 91580
rect 586 91579 608 91585
rect 295 91544 300 91578
rect 324 91544 329 91578
rect 544 91576 582 91579
rect 378 91539 450 91547
rect 428 91509 430 91525
rect 400 91501 430 91509
rect 476 91507 480 91575
rect 544 91546 552 91576
rect 578 91546 582 91576
rect 544 91537 548 91546
rect 400 91497 436 91501
rect 400 91467 408 91497
rect 420 91467 436 91497
rect 544 91499 548 91507
rect 12 91428 62 91430
rect 28 91419 59 91427
rect 62 91419 64 91428
rect 28 91411 64 91419
rect 127 91419 158 91427
rect 127 91412 182 91419
rect 215 91417 224 91445
rect 127 91411 161 91412
rect 59 91395 64 91411
rect 158 91395 161 91411
rect 28 91387 64 91395
rect 127 91394 161 91395
rect 127 91387 182 91394
rect 62 91378 64 91387
rect 213 91379 224 91417
rect 282 91407 292 91465
rect 296 91459 368 91467
rect 319 91429 346 91440
rect 318 91416 324 91429
rect 346 91416 348 91429
rect 428 91420 430 91467
rect 443 91457 450 91459
rect 476 91427 480 91495
rect 544 91465 552 91499
rect 578 91465 582 91499
rect 481 91433 517 91461
rect 481 91427 495 91433
rect 367 91416 380 91420
rect 251 91373 263 91407
rect 273 91373 293 91407
rect 295 91392 324 91416
rect 303 91382 316 91392
rect 318 91376 324 91392
rect 333 91392 380 91416
rect 333 91382 353 91392
rect 367 91386 380 91392
rect 396 91386 408 91420
rect 420 91386 436 91420
rect 120 91325 170 91327
rect 76 91319 92 91325
rect 94 91319 110 91325
rect 76 91309 99 91318
rect 60 91299 67 91309
rect 76 91289 77 91309
rect 96 91284 99 91309
rect 109 91289 110 91309
rect 119 91299 126 91309
rect 76 91275 110 91279
rect 170 91275 172 91325
rect 186 91307 190 91341
rect 216 91307 220 91341
rect 186 91230 220 91264
rect 282 91261 292 91373
rect 318 91366 335 91376
rect 318 91297 324 91366
rect 346 91297 348 91382
rect 428 91339 430 91386
rect 476 91349 480 91417
rect 485 91399 495 91427
rect 505 91427 519 91433
rect 544 91427 555 91465
rect 505 91399 525 91427
rect 544 91399 553 91427
rect 544 91379 548 91399
rect 579 91358 582 91448
rect 612 91430 624 91431
rect 599 91428 649 91430
rect 612 91427 624 91428
rect 610 91420 632 91427
rect 607 91419 632 91420
rect 586 91412 644 91419
rect 607 91411 644 91412
rect 607 91395 610 91411
rect 616 91395 644 91411
rect 607 91394 644 91395
rect 586 91387 644 91394
rect 607 91386 610 91387
rect 612 91379 632 91387
rect 612 91375 624 91379
rect 649 91378 651 91428
rect 544 91341 548 91349
rect 400 91309 408 91339
rect 420 91309 436 91339
rect 400 91305 436 91309
rect 400 91297 430 91305
rect 428 91281 430 91297
rect 476 91269 480 91337
rect 544 91307 552 91341
rect 578 91307 582 91341
rect 544 91299 548 91307
rect 544 91269 586 91270
rect 288 91229 292 91261
rect 296 91259 368 91267
rect 378 91259 450 91267
rect 544 91262 548 91269
rect 439 91231 444 91259
rect 120 91215 170 91217
rect 76 91211 130 91215
rect 110 91206 130 91211
rect 60 91181 67 91191
rect 76 91181 77 91201
rect 96 91172 99 91206
rect 109 91181 110 91201
rect 119 91181 126 91191
rect 76 91165 92 91171
rect 94 91165 110 91171
rect 170 91165 172 91215
rect 186 91149 190 91183
rect 216 91149 220 91183
rect 213 91117 224 91149
rect 282 91145 292 91229
rect 296 91223 368 91231
rect 378 91223 450 91231
rect 468 91228 473 91262
rect 428 91193 430 91209
rect 251 91117 292 91145
rect 318 91124 324 91193
rect 12 91112 62 91114
rect 28 91103 59 91111
rect 62 91103 64 91112
rect 251 91111 263 91117
rect 28 91095 64 91103
rect 127 91103 158 91111
rect 127 91096 182 91103
rect 127 91095 161 91096
rect 59 91079 64 91095
rect 158 91079 161 91095
rect 253 91083 263 91111
rect 273 91083 293 91117
rect 318 91114 335 91124
rect 303 91098 316 91108
rect 318 91098 324 91114
rect 346 91108 348 91193
rect 400 91185 430 91193
rect 476 91191 480 91259
rect 511 91228 582 91262
rect 544 91221 548 91228
rect 400 91181 436 91185
rect 400 91151 408 91181
rect 420 91151 436 91181
rect 544 91183 548 91191
rect 28 91071 64 91079
rect 127 91078 161 91079
rect 127 91071 182 91078
rect 62 91062 64 91071
rect 282 91025 292 91083
rect 295 91074 324 91098
rect 333 91098 353 91108
rect 428 91104 430 91151
rect 476 91111 480 91179
rect 544 91149 552 91183
rect 578 91149 582 91183
rect 544 91141 548 91149
rect 367 91098 380 91104
rect 333 91074 380 91098
rect 318 91061 324 91074
rect 346 91061 348 91074
rect 367 91070 380 91074
rect 396 91070 408 91104
rect 420 91070 436 91104
rect 544 91101 553 91129
rect 319 91050 346 91061
rect 120 91009 170 91011
rect 76 91003 92 91009
rect 94 91003 110 91009
rect 76 90993 99 91002
rect 60 90983 67 90993
rect 76 90973 77 90993
rect 96 90968 99 90993
rect 109 90973 110 90993
rect 119 90983 126 90993
rect 76 90959 110 90963
rect 170 90959 172 91009
rect 186 90991 190 91025
rect 216 90991 220 91025
rect 182 90953 224 90954
rect 186 90929 220 90946
rect 223 90929 257 90946
rect 182 90912 257 90929
rect 182 90911 224 90912
rect 160 90905 246 90911
rect 288 90905 292 91025
rect 296 91023 368 91031
rect 428 91023 430 91070
rect 476 91033 480 91101
rect 485 91057 495 91091
rect 505 91063 525 91091
rect 505 91057 519 91063
rect 544 91057 555 91101
rect 485 91033 492 91057
rect 579 91042 582 91132
rect 612 91114 624 91115
rect 599 91112 649 91114
rect 612 91111 624 91112
rect 610 91104 632 91111
rect 607 91103 632 91104
rect 586 91096 644 91103
rect 607 91095 644 91096
rect 607 91079 610 91095
rect 616 91079 644 91095
rect 607 91078 644 91079
rect 586 91071 644 91078
rect 607 91070 610 91071
rect 612 91063 632 91071
rect 612 91059 624 91063
rect 649 91062 651 91112
rect 544 91025 548 91033
rect 400 90993 408 91023
rect 420 90993 436 91023
rect 400 90989 436 90993
rect 400 90981 430 90989
rect 428 90965 430 90981
rect 476 90953 480 91021
rect 544 90991 552 91025
rect 578 90991 582 91025
rect 544 90983 548 90991
rect 295 90912 300 90946
rect 324 90912 329 90946
rect 378 90943 450 90951
rect 544 90948 548 90953
rect 544 90944 582 90948
rect 544 90929 552 90944
rect 578 90929 582 90944
rect 544 90911 586 90929
rect 522 90905 608 90911
rect 182 90889 224 90905
rect 544 90889 586 90905
rect 17 90875 67 90877
rect 119 90875 169 90877
rect 186 90875 220 90889
rect 548 90875 582 90889
rect 599 90875 649 90877
rect 42 90833 59 90867
rect 67 90825 69 90875
rect 160 90867 246 90875
rect 522 90867 608 90875
rect 76 90833 110 90867
rect 127 90833 144 90867
rect 152 90833 161 90867
rect 162 90865 195 90867
rect 224 90865 244 90867
rect 162 90833 244 90865
rect 524 90865 548 90867
rect 573 90865 582 90867
rect 586 90865 606 90867
rect 160 90825 246 90833
rect 186 90809 220 90825
rect 182 90795 224 90796
rect 160 90789 182 90795
rect 224 90789 246 90795
rect 186 90754 220 90788
rect 223 90754 257 90788
rect 120 90741 170 90743
rect 76 90737 130 90741
rect 110 90732 130 90737
rect 60 90707 67 90717
rect 76 90707 77 90727
rect 96 90698 99 90732
rect 109 90707 110 90727
rect 119 90707 126 90717
rect 76 90691 92 90697
rect 94 90691 110 90697
rect 170 90691 172 90741
rect 186 90675 190 90709
rect 216 90675 220 90709
rect 288 90675 292 90863
rect 476 90795 480 90863
rect 524 90833 606 90865
rect 607 90833 616 90867
rect 522 90825 608 90833
rect 649 90825 651 90875
rect 548 90809 582 90825
rect 522 90790 548 90795
rect 522 90789 582 90790
rect 586 90789 608 90795
rect 295 90754 300 90788
rect 324 90754 329 90788
rect 544 90786 582 90789
rect 378 90749 450 90757
rect 428 90719 430 90735
rect 400 90711 430 90719
rect 476 90717 480 90785
rect 544 90756 552 90786
rect 578 90756 582 90786
rect 544 90747 548 90756
rect 400 90707 436 90711
rect 400 90677 408 90707
rect 420 90677 436 90707
rect 544 90709 548 90717
rect 12 90638 62 90640
rect 28 90629 59 90637
rect 62 90629 64 90638
rect 28 90621 64 90629
rect 127 90629 158 90637
rect 127 90622 182 90629
rect 215 90627 224 90655
rect 127 90621 161 90622
rect 59 90605 64 90621
rect 158 90605 161 90621
rect 28 90597 64 90605
rect 127 90604 161 90605
rect 127 90597 182 90604
rect 62 90588 64 90597
rect 213 90589 224 90627
rect 282 90617 292 90675
rect 296 90669 368 90677
rect 319 90639 346 90650
rect 318 90626 324 90639
rect 346 90626 348 90639
rect 428 90630 430 90677
rect 443 90667 450 90669
rect 476 90637 480 90705
rect 544 90675 552 90709
rect 578 90675 582 90709
rect 481 90643 517 90671
rect 481 90637 495 90643
rect 367 90626 380 90630
rect 251 90583 263 90617
rect 273 90583 293 90617
rect 295 90602 324 90626
rect 303 90592 316 90602
rect 318 90586 324 90602
rect 333 90602 380 90626
rect 333 90592 353 90602
rect 367 90596 380 90602
rect 396 90596 408 90630
rect 420 90596 436 90630
rect 120 90535 170 90537
rect 76 90529 92 90535
rect 94 90529 110 90535
rect 76 90519 99 90528
rect 60 90509 67 90519
rect 76 90499 77 90519
rect 96 90494 99 90519
rect 109 90499 110 90519
rect 119 90509 126 90519
rect 76 90485 110 90489
rect 170 90485 172 90535
rect 186 90517 190 90551
rect 216 90517 220 90551
rect 186 90440 220 90474
rect 282 90471 292 90583
rect 318 90576 335 90586
rect 318 90507 324 90576
rect 346 90507 348 90592
rect 428 90549 430 90596
rect 476 90559 480 90627
rect 485 90609 495 90637
rect 505 90637 519 90643
rect 544 90637 555 90675
rect 505 90609 525 90637
rect 544 90609 553 90637
rect 544 90589 548 90609
rect 579 90568 582 90658
rect 612 90640 624 90641
rect 599 90638 649 90640
rect 612 90637 624 90638
rect 610 90630 632 90637
rect 607 90629 632 90630
rect 586 90622 644 90629
rect 607 90621 644 90622
rect 607 90605 610 90621
rect 616 90605 644 90621
rect 607 90604 644 90605
rect 586 90597 644 90604
rect 607 90596 610 90597
rect 612 90589 632 90597
rect 612 90585 624 90589
rect 649 90588 651 90638
rect 544 90551 548 90559
rect 400 90519 408 90549
rect 420 90519 436 90549
rect 400 90515 436 90519
rect 400 90507 430 90515
rect 428 90491 430 90507
rect 476 90479 480 90547
rect 544 90517 552 90551
rect 578 90517 582 90551
rect 544 90509 548 90517
rect 544 90479 586 90480
rect 288 90439 292 90471
rect 296 90469 368 90477
rect 378 90469 450 90477
rect 544 90472 548 90479
rect 439 90441 444 90469
rect 120 90425 170 90427
rect 76 90421 130 90425
rect 110 90416 130 90421
rect 60 90391 67 90401
rect 76 90391 77 90411
rect 96 90382 99 90416
rect 109 90391 110 90411
rect 119 90391 126 90401
rect 76 90375 92 90381
rect 94 90375 110 90381
rect 170 90375 172 90425
rect 186 90359 190 90393
rect 216 90359 220 90393
rect 213 90327 224 90359
rect 282 90355 292 90439
rect 296 90433 368 90441
rect 378 90433 450 90441
rect 468 90438 473 90472
rect 428 90403 430 90419
rect 251 90327 292 90355
rect 318 90334 324 90403
rect 12 90322 62 90324
rect 28 90313 59 90321
rect 62 90313 64 90322
rect 251 90321 263 90327
rect 28 90305 64 90313
rect 127 90313 158 90321
rect 127 90306 182 90313
rect 127 90305 161 90306
rect 59 90289 64 90305
rect 158 90289 161 90305
rect 253 90293 263 90321
rect 273 90293 293 90327
rect 318 90324 335 90334
rect 303 90308 316 90318
rect 318 90308 324 90324
rect 346 90318 348 90403
rect 400 90395 430 90403
rect 476 90401 480 90469
rect 511 90438 582 90472
rect 544 90431 548 90438
rect 400 90391 436 90395
rect 400 90361 408 90391
rect 420 90361 436 90391
rect 544 90393 548 90401
rect 28 90281 64 90289
rect 127 90288 161 90289
rect 127 90281 182 90288
rect 62 90272 64 90281
rect 282 90235 292 90293
rect 295 90284 324 90308
rect 333 90308 353 90318
rect 428 90314 430 90361
rect 476 90321 480 90389
rect 544 90359 552 90393
rect 578 90359 582 90393
rect 544 90351 548 90359
rect 367 90308 380 90314
rect 333 90284 380 90308
rect 318 90271 324 90284
rect 346 90271 348 90284
rect 367 90280 380 90284
rect 396 90280 408 90314
rect 420 90280 436 90314
rect 544 90311 553 90339
rect 319 90260 346 90271
rect 120 90219 170 90221
rect 76 90213 92 90219
rect 94 90213 110 90219
rect 76 90203 99 90212
rect 60 90193 67 90203
rect 76 90183 77 90203
rect 96 90178 99 90203
rect 109 90183 110 90203
rect 119 90193 126 90203
rect 76 90169 110 90173
rect 170 90169 172 90219
rect 186 90201 190 90235
rect 216 90201 220 90235
rect 182 90163 224 90164
rect 186 90139 220 90156
rect 223 90139 257 90156
rect 182 90122 257 90139
rect 182 90121 224 90122
rect 160 90115 246 90121
rect 288 90115 292 90235
rect 296 90233 368 90241
rect 428 90233 430 90280
rect 476 90243 480 90311
rect 485 90267 495 90301
rect 505 90273 525 90301
rect 505 90267 519 90273
rect 544 90267 555 90311
rect 485 90243 492 90267
rect 579 90252 582 90342
rect 612 90324 624 90325
rect 599 90322 649 90324
rect 612 90321 624 90322
rect 610 90314 632 90321
rect 607 90313 632 90314
rect 586 90306 644 90313
rect 607 90305 644 90306
rect 607 90289 610 90305
rect 616 90289 644 90305
rect 607 90288 644 90289
rect 586 90281 644 90288
rect 607 90280 610 90281
rect 612 90273 632 90281
rect 612 90269 624 90273
rect 649 90272 651 90322
rect 544 90235 548 90243
rect 400 90203 408 90233
rect 420 90203 436 90233
rect 400 90199 436 90203
rect 400 90191 430 90199
rect 428 90175 430 90191
rect 476 90163 480 90231
rect 544 90201 552 90235
rect 578 90201 582 90235
rect 544 90193 548 90201
rect 295 90122 300 90156
rect 324 90122 329 90156
rect 378 90153 450 90161
rect 544 90158 548 90163
rect 544 90154 582 90158
rect 544 90139 552 90154
rect 578 90139 582 90154
rect 544 90121 586 90139
rect 522 90115 608 90121
rect 182 90099 224 90115
rect 544 90099 586 90115
rect 17 90085 67 90087
rect 119 90085 169 90087
rect 186 90085 220 90099
rect 548 90085 582 90099
rect 599 90085 649 90087
rect 42 90043 59 90077
rect 67 90035 69 90085
rect 160 90077 246 90085
rect 522 90077 608 90085
rect 76 90043 110 90077
rect 127 90043 144 90077
rect 152 90043 161 90077
rect 162 90075 195 90077
rect 224 90075 244 90077
rect 162 90043 244 90075
rect 524 90075 548 90077
rect 573 90075 582 90077
rect 586 90075 606 90077
rect 160 90035 246 90043
rect 186 90019 220 90035
rect 182 90005 224 90006
rect 160 89999 182 90005
rect 224 89999 246 90005
rect 186 89964 220 89998
rect 223 89964 257 89998
rect 120 89951 170 89953
rect 76 89947 130 89951
rect 110 89942 130 89947
rect 60 89917 67 89927
rect 76 89917 77 89937
rect 96 89908 99 89942
rect 109 89917 110 89937
rect 119 89917 126 89927
rect 76 89901 92 89907
rect 94 89901 110 89907
rect 170 89901 172 89951
rect 186 89885 190 89919
rect 216 89885 220 89919
rect 288 89885 292 90073
rect 476 90005 480 90073
rect 524 90043 606 90075
rect 607 90043 616 90077
rect 522 90035 608 90043
rect 649 90035 651 90085
rect 548 90019 582 90035
rect 522 90000 548 90005
rect 522 89999 582 90000
rect 586 89999 608 90005
rect 295 89964 300 89998
rect 324 89964 329 89998
rect 544 89996 582 89999
rect 378 89959 450 89967
rect 428 89929 430 89945
rect 400 89921 430 89929
rect 476 89927 480 89995
rect 544 89966 552 89996
rect 578 89966 582 89996
rect 544 89957 548 89966
rect 400 89917 436 89921
rect 400 89887 408 89917
rect 420 89887 436 89917
rect 544 89919 548 89927
rect 12 89848 62 89850
rect 28 89839 59 89847
rect 62 89839 64 89848
rect 28 89831 64 89839
rect 127 89839 158 89847
rect 127 89832 182 89839
rect 215 89837 224 89865
rect 127 89831 161 89832
rect 59 89815 64 89831
rect 158 89815 161 89831
rect 28 89807 64 89815
rect 127 89814 161 89815
rect 127 89807 182 89814
rect 62 89798 64 89807
rect 213 89799 224 89837
rect 282 89827 292 89885
rect 296 89879 368 89887
rect 319 89849 346 89860
rect 318 89836 324 89849
rect 346 89836 348 89849
rect 428 89840 430 89887
rect 443 89877 450 89879
rect 476 89847 480 89915
rect 544 89885 552 89919
rect 578 89885 582 89919
rect 481 89853 517 89881
rect 481 89847 495 89853
rect 367 89836 380 89840
rect 251 89793 263 89827
rect 273 89793 293 89827
rect 295 89812 324 89836
rect 303 89802 316 89812
rect 318 89796 324 89812
rect 333 89812 380 89836
rect 333 89802 353 89812
rect 367 89806 380 89812
rect 396 89806 408 89840
rect 420 89806 436 89840
rect 120 89745 170 89747
rect 76 89739 92 89745
rect 94 89739 110 89745
rect 76 89729 99 89738
rect 60 89719 67 89729
rect 76 89709 77 89729
rect 96 89704 99 89729
rect 109 89709 110 89729
rect 119 89719 126 89729
rect 76 89695 110 89699
rect 170 89695 172 89745
rect 186 89727 190 89761
rect 216 89727 220 89761
rect 186 89650 220 89684
rect 282 89681 292 89793
rect 318 89786 335 89796
rect 318 89717 324 89786
rect 346 89717 348 89802
rect 428 89759 430 89806
rect 476 89769 480 89837
rect 485 89819 495 89847
rect 505 89847 519 89853
rect 544 89847 555 89885
rect 505 89819 525 89847
rect 544 89819 553 89847
rect 544 89799 548 89819
rect 579 89778 582 89868
rect 612 89850 624 89851
rect 599 89848 649 89850
rect 612 89847 624 89848
rect 610 89840 632 89847
rect 607 89839 632 89840
rect 586 89832 644 89839
rect 607 89831 644 89832
rect 607 89815 610 89831
rect 616 89815 644 89831
rect 607 89814 644 89815
rect 586 89807 644 89814
rect 607 89806 610 89807
rect 612 89799 632 89807
rect 612 89795 624 89799
rect 649 89798 651 89848
rect 544 89761 548 89769
rect 400 89729 408 89759
rect 420 89729 436 89759
rect 400 89725 436 89729
rect 400 89717 430 89725
rect 428 89701 430 89717
rect 476 89689 480 89757
rect 544 89727 552 89761
rect 578 89727 582 89761
rect 544 89719 548 89727
rect 544 89689 586 89690
rect 288 89649 292 89681
rect 296 89679 368 89687
rect 378 89679 450 89687
rect 544 89682 548 89689
rect 439 89651 444 89679
rect 120 89635 170 89637
rect 76 89631 130 89635
rect 110 89626 130 89631
rect 60 89601 67 89611
rect 76 89601 77 89621
rect 96 89592 99 89626
rect 109 89601 110 89621
rect 119 89601 126 89611
rect 76 89585 92 89591
rect 94 89585 110 89591
rect 170 89585 172 89635
rect 186 89569 190 89603
rect 216 89569 220 89603
rect 213 89537 224 89569
rect 282 89565 292 89649
rect 296 89643 368 89651
rect 378 89643 450 89651
rect 468 89648 473 89682
rect 428 89613 430 89629
rect 251 89537 292 89565
rect 318 89544 324 89613
rect 12 89532 62 89534
rect 28 89523 59 89531
rect 62 89523 64 89532
rect 251 89531 263 89537
rect 28 89515 64 89523
rect 127 89523 158 89531
rect 127 89516 182 89523
rect 127 89515 161 89516
rect 59 89499 64 89515
rect 158 89499 161 89515
rect 253 89503 263 89531
rect 273 89503 293 89537
rect 318 89534 335 89544
rect 303 89518 316 89528
rect 318 89518 324 89534
rect 346 89528 348 89613
rect 400 89605 430 89613
rect 476 89611 480 89679
rect 511 89648 582 89682
rect 544 89641 548 89648
rect 400 89601 436 89605
rect 400 89571 408 89601
rect 420 89571 436 89601
rect 544 89603 548 89611
rect 28 89491 64 89499
rect 127 89498 161 89499
rect 127 89491 182 89498
rect 62 89482 64 89491
rect 282 89445 292 89503
rect 295 89494 324 89518
rect 333 89518 353 89528
rect 428 89524 430 89571
rect 476 89531 480 89599
rect 544 89569 552 89603
rect 578 89569 582 89603
rect 544 89561 548 89569
rect 367 89518 380 89524
rect 333 89494 380 89518
rect 318 89481 324 89494
rect 346 89481 348 89494
rect 367 89490 380 89494
rect 396 89490 408 89524
rect 420 89490 436 89524
rect 544 89521 553 89549
rect 319 89470 346 89481
rect 120 89429 170 89431
rect 76 89423 92 89429
rect 94 89423 110 89429
rect 76 89413 99 89422
rect 60 89403 67 89413
rect 76 89393 77 89413
rect 96 89388 99 89413
rect 109 89393 110 89413
rect 119 89403 126 89413
rect 76 89379 110 89383
rect 170 89379 172 89429
rect 186 89411 190 89445
rect 216 89411 220 89445
rect 182 89373 224 89374
rect 186 89349 220 89366
rect 223 89349 257 89366
rect 182 89332 257 89349
rect 182 89331 224 89332
rect 160 89325 246 89331
rect 288 89325 292 89445
rect 296 89443 368 89451
rect 428 89443 430 89490
rect 476 89453 480 89521
rect 485 89477 495 89511
rect 505 89483 525 89511
rect 505 89477 519 89483
rect 544 89477 555 89521
rect 485 89453 492 89477
rect 579 89462 582 89552
rect 612 89534 624 89535
rect 599 89532 649 89534
rect 612 89531 624 89532
rect 610 89524 632 89531
rect 607 89523 632 89524
rect 586 89516 644 89523
rect 607 89515 644 89516
rect 607 89499 610 89515
rect 616 89499 644 89515
rect 607 89498 644 89499
rect 586 89491 644 89498
rect 607 89490 610 89491
rect 612 89483 632 89491
rect 612 89479 624 89483
rect 649 89482 651 89532
rect 544 89445 548 89453
rect 400 89413 408 89443
rect 420 89413 436 89443
rect 400 89409 436 89413
rect 400 89401 430 89409
rect 428 89385 430 89401
rect 476 89373 480 89441
rect 544 89411 552 89445
rect 578 89411 582 89445
rect 544 89403 548 89411
rect 295 89332 300 89366
rect 324 89332 329 89366
rect 378 89363 450 89371
rect 544 89368 548 89373
rect 544 89364 582 89368
rect 544 89349 552 89364
rect 578 89349 582 89364
rect 544 89331 586 89349
rect 522 89325 608 89331
rect 182 89309 224 89325
rect 544 89309 586 89325
rect 17 89295 67 89297
rect 119 89295 169 89297
rect 186 89295 220 89309
rect 548 89295 582 89309
rect 599 89295 649 89297
rect 42 89253 59 89287
rect 67 89245 69 89295
rect 160 89287 246 89295
rect 522 89287 608 89295
rect 76 89253 110 89287
rect 127 89253 144 89287
rect 152 89253 161 89287
rect 162 89285 195 89287
rect 224 89285 244 89287
rect 162 89253 244 89285
rect 524 89285 548 89287
rect 573 89285 582 89287
rect 586 89285 606 89287
rect 160 89245 246 89253
rect 186 89229 220 89245
rect 182 89215 224 89216
rect 160 89209 182 89215
rect 224 89209 246 89215
rect 186 89174 220 89208
rect 223 89174 257 89208
rect 120 89161 170 89163
rect 76 89157 130 89161
rect 110 89152 130 89157
rect 60 89127 67 89137
rect 76 89127 77 89147
rect 96 89118 99 89152
rect 109 89127 110 89147
rect 119 89127 126 89137
rect 76 89111 92 89117
rect 94 89111 110 89117
rect 170 89111 172 89161
rect 186 89095 190 89129
rect 216 89095 220 89129
rect 288 89095 292 89283
rect 476 89215 480 89283
rect 524 89253 606 89285
rect 607 89253 616 89287
rect 522 89245 608 89253
rect 649 89245 651 89295
rect 548 89229 582 89245
rect 522 89210 548 89215
rect 522 89209 582 89210
rect 586 89209 608 89215
rect 295 89174 300 89208
rect 324 89174 329 89208
rect 544 89206 582 89209
rect 378 89169 450 89177
rect 428 89139 430 89155
rect 400 89131 430 89139
rect 476 89137 480 89205
rect 544 89176 552 89206
rect 578 89176 582 89206
rect 544 89167 548 89176
rect 400 89127 436 89131
rect 400 89097 408 89127
rect 420 89097 436 89127
rect 544 89129 548 89137
rect 12 89058 62 89060
rect 28 89049 59 89057
rect 62 89049 64 89058
rect 28 89041 64 89049
rect 127 89049 158 89057
rect 127 89042 182 89049
rect 215 89047 224 89075
rect 127 89041 161 89042
rect 59 89025 64 89041
rect 158 89025 161 89041
rect 28 89017 64 89025
rect 127 89024 161 89025
rect 127 89017 182 89024
rect 62 89008 64 89017
rect 213 89009 224 89047
rect 282 89037 292 89095
rect 296 89089 368 89097
rect 319 89059 346 89070
rect 318 89046 324 89059
rect 346 89046 348 89059
rect 428 89050 430 89097
rect 443 89087 450 89089
rect 476 89057 480 89125
rect 544 89095 552 89129
rect 578 89095 582 89129
rect 481 89063 517 89091
rect 481 89057 495 89063
rect 367 89046 380 89050
rect 251 89003 263 89037
rect 273 89003 293 89037
rect 295 89022 324 89046
rect 303 89012 316 89022
rect 318 89006 324 89022
rect 333 89022 380 89046
rect 333 89012 353 89022
rect 367 89016 380 89022
rect 396 89016 408 89050
rect 420 89016 436 89050
rect 120 88955 170 88957
rect 76 88949 92 88955
rect 94 88949 110 88955
rect 76 88939 99 88948
rect 60 88929 67 88939
rect 76 88919 77 88939
rect 96 88914 99 88939
rect 109 88919 110 88939
rect 119 88929 126 88939
rect 76 88905 110 88909
rect 170 88905 172 88955
rect 186 88937 190 88971
rect 216 88937 220 88971
rect 186 88860 220 88894
rect 282 88891 292 89003
rect 318 88996 335 89006
rect 318 88927 324 88996
rect 346 88927 348 89012
rect 428 88969 430 89016
rect 476 88979 480 89047
rect 485 89029 495 89057
rect 505 89057 519 89063
rect 544 89057 555 89095
rect 505 89029 525 89057
rect 544 89029 553 89057
rect 544 89009 548 89029
rect 579 88988 582 89078
rect 612 89060 624 89061
rect 599 89058 649 89060
rect 612 89057 624 89058
rect 610 89050 632 89057
rect 607 89049 632 89050
rect 586 89042 644 89049
rect 607 89041 644 89042
rect 607 89025 610 89041
rect 616 89025 644 89041
rect 607 89024 644 89025
rect 586 89017 644 89024
rect 607 89016 610 89017
rect 612 89009 632 89017
rect 612 89005 624 89009
rect 649 89008 651 89058
rect 544 88971 548 88979
rect 400 88939 408 88969
rect 420 88939 436 88969
rect 400 88935 436 88939
rect 400 88927 430 88935
rect 428 88911 430 88927
rect 476 88899 480 88967
rect 544 88937 552 88971
rect 578 88937 582 88971
rect 544 88929 548 88937
rect 544 88899 586 88900
rect 288 88859 292 88891
rect 296 88889 368 88897
rect 378 88889 450 88897
rect 544 88892 548 88899
rect 439 88861 444 88889
rect 120 88845 170 88847
rect 76 88841 130 88845
rect 110 88836 130 88841
rect 60 88811 67 88821
rect 76 88811 77 88831
rect 96 88802 99 88836
rect 109 88811 110 88831
rect 119 88811 126 88821
rect 76 88795 92 88801
rect 94 88795 110 88801
rect 170 88795 172 88845
rect 186 88779 190 88813
rect 216 88779 220 88813
rect 213 88747 224 88779
rect 282 88775 292 88859
rect 296 88853 368 88861
rect 378 88853 450 88861
rect 468 88858 473 88892
rect 428 88823 430 88839
rect 251 88747 292 88775
rect 318 88754 324 88823
rect 12 88742 62 88744
rect 28 88733 59 88741
rect 62 88733 64 88742
rect 251 88741 263 88747
rect 28 88725 64 88733
rect 127 88733 158 88741
rect 127 88726 182 88733
rect 127 88725 161 88726
rect 59 88709 64 88725
rect 158 88709 161 88725
rect 253 88713 263 88741
rect 273 88713 293 88747
rect 318 88744 335 88754
rect 303 88728 316 88738
rect 318 88728 324 88744
rect 346 88738 348 88823
rect 400 88815 430 88823
rect 476 88821 480 88889
rect 511 88858 582 88892
rect 544 88851 548 88858
rect 400 88811 436 88815
rect 400 88781 408 88811
rect 420 88781 436 88811
rect 544 88813 548 88821
rect 28 88701 64 88709
rect 127 88708 161 88709
rect 127 88701 182 88708
rect 62 88692 64 88701
rect 282 88655 292 88713
rect 295 88704 324 88728
rect 333 88728 353 88738
rect 428 88734 430 88781
rect 476 88741 480 88809
rect 544 88779 552 88813
rect 578 88779 582 88813
rect 544 88771 548 88779
rect 367 88728 380 88734
rect 333 88704 380 88728
rect 318 88691 324 88704
rect 346 88691 348 88704
rect 367 88700 380 88704
rect 396 88700 408 88734
rect 420 88700 436 88734
rect 544 88731 553 88759
rect 319 88680 346 88691
rect 120 88639 170 88641
rect 76 88633 92 88639
rect 94 88633 110 88639
rect 76 88623 99 88632
rect 60 88613 67 88623
rect 76 88603 77 88623
rect 96 88598 99 88623
rect 109 88603 110 88623
rect 119 88613 126 88623
rect 76 88589 110 88593
rect 170 88589 172 88639
rect 186 88621 190 88655
rect 216 88621 220 88655
rect 182 88583 224 88584
rect 186 88559 220 88576
rect 223 88559 257 88576
rect 182 88542 257 88559
rect 182 88541 224 88542
rect 160 88535 246 88541
rect 288 88535 292 88655
rect 296 88653 368 88661
rect 428 88653 430 88700
rect 476 88663 480 88731
rect 485 88687 495 88721
rect 505 88693 525 88721
rect 505 88687 519 88693
rect 544 88687 555 88731
rect 485 88663 492 88687
rect 579 88672 582 88762
rect 612 88744 624 88745
rect 599 88742 649 88744
rect 612 88741 624 88742
rect 610 88734 632 88741
rect 607 88733 632 88734
rect 586 88726 644 88733
rect 607 88725 644 88726
rect 607 88709 610 88725
rect 616 88709 644 88725
rect 607 88708 644 88709
rect 586 88701 644 88708
rect 607 88700 610 88701
rect 612 88693 632 88701
rect 612 88689 624 88693
rect 649 88692 651 88742
rect 544 88655 548 88663
rect 400 88623 408 88653
rect 420 88623 436 88653
rect 400 88619 436 88623
rect 400 88611 430 88619
rect 428 88595 430 88611
rect 476 88583 480 88651
rect 544 88621 552 88655
rect 578 88621 582 88655
rect 544 88613 548 88621
rect 295 88542 300 88576
rect 324 88542 329 88576
rect 378 88573 450 88581
rect 544 88578 548 88583
rect 544 88574 582 88578
rect 544 88559 552 88574
rect 578 88559 582 88574
rect 544 88541 586 88559
rect 522 88535 608 88541
rect 182 88519 224 88535
rect 544 88519 586 88535
rect 17 88505 67 88507
rect 119 88505 169 88507
rect 186 88505 220 88519
rect 548 88505 582 88519
rect 599 88505 649 88507
rect 42 88463 59 88497
rect 67 88455 69 88505
rect 160 88497 246 88505
rect 522 88497 608 88505
rect 76 88463 110 88497
rect 127 88463 144 88497
rect 152 88463 161 88497
rect 162 88495 195 88497
rect 224 88495 244 88497
rect 162 88463 244 88495
rect 524 88495 548 88497
rect 573 88495 582 88497
rect 586 88495 606 88497
rect 160 88455 246 88463
rect 186 88439 220 88455
rect 182 88425 224 88426
rect 160 88419 182 88425
rect 224 88419 246 88425
rect 186 88384 220 88418
rect 223 88384 257 88418
rect 120 88371 170 88373
rect 76 88367 130 88371
rect 110 88362 130 88367
rect 60 88337 67 88347
rect 76 88337 77 88357
rect 96 88328 99 88362
rect 109 88337 110 88357
rect 119 88337 126 88347
rect 76 88321 92 88327
rect 94 88321 110 88327
rect 170 88321 172 88371
rect 186 88305 190 88339
rect 216 88305 220 88339
rect 288 88305 292 88493
rect 476 88425 480 88493
rect 524 88463 606 88495
rect 607 88463 616 88497
rect 522 88455 608 88463
rect 649 88455 651 88505
rect 548 88439 582 88455
rect 522 88420 548 88425
rect 522 88419 582 88420
rect 586 88419 608 88425
rect 295 88384 300 88418
rect 324 88384 329 88418
rect 544 88416 582 88419
rect 378 88379 450 88387
rect 428 88349 430 88365
rect 400 88341 430 88349
rect 476 88347 480 88415
rect 544 88386 552 88416
rect 578 88386 582 88416
rect 544 88377 548 88386
rect 400 88337 436 88341
rect 400 88307 408 88337
rect 420 88307 436 88337
rect 544 88339 548 88347
rect 12 88268 62 88270
rect 28 88259 59 88267
rect 62 88259 64 88268
rect 28 88251 64 88259
rect 127 88259 158 88267
rect 127 88252 182 88259
rect 215 88257 224 88285
rect 127 88251 161 88252
rect 59 88235 64 88251
rect 158 88235 161 88251
rect 28 88227 64 88235
rect 127 88234 161 88235
rect 127 88227 182 88234
rect 62 88218 64 88227
rect 213 88219 224 88257
rect 282 88247 292 88305
rect 296 88299 368 88307
rect 319 88269 346 88280
rect 318 88256 324 88269
rect 346 88256 348 88269
rect 428 88260 430 88307
rect 443 88297 450 88299
rect 476 88267 480 88335
rect 544 88305 552 88339
rect 578 88305 582 88339
rect 481 88273 517 88301
rect 481 88267 495 88273
rect 367 88256 380 88260
rect 251 88213 263 88247
rect 273 88213 293 88247
rect 295 88232 324 88256
rect 303 88222 316 88232
rect 318 88216 324 88232
rect 333 88232 380 88256
rect 333 88222 353 88232
rect 367 88226 380 88232
rect 396 88226 408 88260
rect 420 88226 436 88260
rect 120 88165 170 88167
rect 76 88159 92 88165
rect 94 88159 110 88165
rect 76 88149 99 88158
rect 60 88139 67 88149
rect 76 88129 77 88149
rect 96 88124 99 88149
rect 109 88129 110 88149
rect 119 88139 126 88149
rect 76 88115 110 88119
rect 170 88115 172 88165
rect 186 88147 190 88181
rect 216 88147 220 88181
rect 186 88070 220 88104
rect 282 88101 292 88213
rect 318 88206 335 88216
rect 318 88137 324 88206
rect 346 88137 348 88222
rect 428 88179 430 88226
rect 476 88189 480 88257
rect 485 88239 495 88267
rect 505 88267 519 88273
rect 544 88267 555 88305
rect 505 88239 525 88267
rect 544 88239 553 88267
rect 544 88219 548 88239
rect 579 88198 582 88288
rect 612 88270 624 88271
rect 599 88268 649 88270
rect 612 88267 624 88268
rect 610 88260 632 88267
rect 607 88259 632 88260
rect 586 88252 644 88259
rect 607 88251 644 88252
rect 607 88235 610 88251
rect 616 88235 644 88251
rect 607 88234 644 88235
rect 586 88227 644 88234
rect 607 88226 610 88227
rect 612 88219 632 88227
rect 612 88215 624 88219
rect 649 88218 651 88268
rect 544 88181 548 88189
rect 400 88149 408 88179
rect 420 88149 436 88179
rect 400 88145 436 88149
rect 400 88137 430 88145
rect 428 88121 430 88137
rect 476 88109 480 88177
rect 544 88147 552 88181
rect 578 88147 582 88181
rect 544 88139 548 88147
rect 544 88109 586 88110
rect 288 88069 292 88101
rect 296 88099 368 88107
rect 378 88099 450 88107
rect 544 88102 548 88109
rect 439 88071 444 88099
rect 120 88055 170 88057
rect 76 88051 130 88055
rect 110 88046 130 88051
rect 60 88021 67 88031
rect 76 88021 77 88041
rect 96 88012 99 88046
rect 109 88021 110 88041
rect 119 88021 126 88031
rect 76 88005 92 88011
rect 94 88005 110 88011
rect 170 88005 172 88055
rect 186 87989 190 88023
rect 216 87989 220 88023
rect 213 87957 224 87989
rect 282 87985 292 88069
rect 296 88063 368 88071
rect 378 88063 450 88071
rect 468 88068 473 88102
rect 428 88033 430 88049
rect 251 87957 292 87985
rect 318 87964 324 88033
rect 12 87952 62 87954
rect 28 87943 59 87951
rect 62 87943 64 87952
rect 251 87951 263 87957
rect 28 87935 64 87943
rect 127 87943 158 87951
rect 127 87936 182 87943
rect 127 87935 161 87936
rect 59 87919 64 87935
rect 158 87919 161 87935
rect 253 87923 263 87951
rect 273 87923 293 87957
rect 318 87954 335 87964
rect 303 87938 316 87948
rect 318 87938 324 87954
rect 346 87948 348 88033
rect 400 88025 430 88033
rect 476 88031 480 88099
rect 511 88068 582 88102
rect 544 88061 548 88068
rect 400 88021 436 88025
rect 400 87991 408 88021
rect 420 87991 436 88021
rect 544 88023 548 88031
rect 28 87911 64 87919
rect 127 87918 161 87919
rect 127 87911 182 87918
rect 62 87902 64 87911
rect 282 87865 292 87923
rect 295 87914 324 87938
rect 333 87938 353 87948
rect 428 87944 430 87991
rect 476 87951 480 88019
rect 544 87989 552 88023
rect 578 87989 582 88023
rect 544 87981 548 87989
rect 367 87938 380 87944
rect 333 87914 380 87938
rect 318 87901 324 87914
rect 346 87901 348 87914
rect 367 87910 380 87914
rect 396 87910 408 87944
rect 420 87910 436 87944
rect 544 87941 553 87969
rect 319 87890 346 87901
rect 120 87849 170 87851
rect 76 87843 92 87849
rect 94 87843 110 87849
rect 76 87833 99 87842
rect 60 87823 67 87833
rect 76 87813 77 87833
rect 96 87808 99 87833
rect 109 87813 110 87833
rect 119 87823 126 87833
rect 76 87799 110 87803
rect 170 87799 172 87849
rect 186 87831 190 87865
rect 216 87831 220 87865
rect 182 87793 224 87794
rect 186 87769 220 87786
rect 223 87769 257 87786
rect 182 87752 257 87769
rect 182 87751 224 87752
rect 160 87745 246 87751
rect 288 87745 292 87865
rect 296 87863 368 87871
rect 428 87863 430 87910
rect 476 87873 480 87941
rect 485 87897 495 87931
rect 505 87903 525 87931
rect 505 87897 519 87903
rect 544 87897 555 87941
rect 485 87873 492 87897
rect 579 87882 582 87972
rect 612 87954 624 87955
rect 599 87952 649 87954
rect 612 87951 624 87952
rect 610 87944 632 87951
rect 607 87943 632 87944
rect 586 87936 644 87943
rect 607 87935 644 87936
rect 607 87919 610 87935
rect 616 87919 644 87935
rect 607 87918 644 87919
rect 586 87911 644 87918
rect 607 87910 610 87911
rect 612 87903 632 87911
rect 612 87899 624 87903
rect 649 87902 651 87952
rect 544 87865 548 87873
rect 400 87833 408 87863
rect 420 87833 436 87863
rect 400 87829 436 87833
rect 400 87821 430 87829
rect 428 87805 430 87821
rect 476 87793 480 87861
rect 544 87831 552 87865
rect 578 87831 582 87865
rect 544 87823 548 87831
rect 295 87752 300 87786
rect 324 87752 329 87786
rect 378 87783 450 87791
rect 544 87788 548 87793
rect 544 87784 582 87788
rect 544 87769 552 87784
rect 578 87769 582 87784
rect 544 87751 586 87769
rect 522 87745 608 87751
rect 182 87729 224 87745
rect 544 87729 586 87745
rect 17 87715 67 87717
rect 119 87715 169 87717
rect 186 87715 220 87729
rect 548 87715 582 87729
rect 599 87715 649 87717
rect 42 87673 59 87707
rect 67 87665 69 87715
rect 160 87707 246 87715
rect 522 87707 608 87715
rect 76 87673 110 87707
rect 127 87673 144 87707
rect 152 87673 161 87707
rect 162 87705 195 87707
rect 224 87705 244 87707
rect 162 87673 244 87705
rect 524 87705 548 87707
rect 573 87705 582 87707
rect 586 87705 606 87707
rect 160 87665 246 87673
rect 186 87649 220 87665
rect 182 87635 224 87636
rect 160 87629 182 87635
rect 224 87629 246 87635
rect 186 87594 220 87628
rect 223 87594 257 87628
rect 120 87581 170 87583
rect 76 87577 130 87581
rect 110 87572 130 87577
rect 60 87547 67 87557
rect 76 87547 77 87567
rect 96 87538 99 87572
rect 109 87547 110 87567
rect 119 87547 126 87557
rect 76 87531 92 87537
rect 94 87531 110 87537
rect 170 87531 172 87581
rect 186 87515 190 87549
rect 216 87515 220 87549
rect 288 87515 292 87703
rect 476 87635 480 87703
rect 524 87673 606 87705
rect 607 87673 616 87707
rect 522 87665 608 87673
rect 649 87665 651 87715
rect 548 87649 582 87665
rect 522 87630 548 87635
rect 522 87629 582 87630
rect 586 87629 608 87635
rect 295 87594 300 87628
rect 324 87594 329 87628
rect 544 87626 582 87629
rect 378 87589 450 87597
rect 428 87559 430 87575
rect 400 87551 430 87559
rect 476 87557 480 87625
rect 544 87596 552 87626
rect 578 87596 582 87626
rect 544 87587 548 87596
rect 400 87547 436 87551
rect 400 87517 408 87547
rect 420 87517 436 87547
rect 544 87549 548 87557
rect 12 87478 62 87480
rect 28 87469 59 87477
rect 62 87469 64 87478
rect 28 87461 64 87469
rect 127 87469 158 87477
rect 127 87462 182 87469
rect 215 87467 224 87495
rect 127 87461 161 87462
rect 59 87445 64 87461
rect 158 87445 161 87461
rect 28 87437 64 87445
rect 127 87444 161 87445
rect 127 87437 182 87444
rect 62 87428 64 87437
rect 213 87429 224 87467
rect 282 87457 292 87515
rect 296 87509 368 87517
rect 319 87479 346 87490
rect 318 87466 324 87479
rect 346 87466 348 87479
rect 428 87470 430 87517
rect 443 87507 450 87509
rect 476 87477 480 87545
rect 544 87515 552 87549
rect 578 87515 582 87549
rect 481 87483 517 87511
rect 481 87477 495 87483
rect 367 87466 380 87470
rect 251 87423 263 87457
rect 273 87423 293 87457
rect 295 87442 324 87466
rect 303 87432 316 87442
rect 318 87426 324 87442
rect 333 87442 380 87466
rect 333 87432 353 87442
rect 367 87436 380 87442
rect 396 87436 408 87470
rect 420 87436 436 87470
rect 120 87375 170 87377
rect 76 87369 92 87375
rect 94 87369 110 87375
rect 76 87359 99 87368
rect 60 87349 67 87359
rect 76 87339 77 87359
rect 96 87334 99 87359
rect 109 87339 110 87359
rect 119 87349 126 87359
rect 76 87325 110 87329
rect 170 87325 172 87375
rect 186 87357 190 87391
rect 216 87357 220 87391
rect 186 87280 220 87314
rect 282 87311 292 87423
rect 318 87416 335 87426
rect 318 87347 324 87416
rect 346 87347 348 87432
rect 428 87389 430 87436
rect 476 87399 480 87467
rect 485 87449 495 87477
rect 505 87477 519 87483
rect 544 87477 555 87515
rect 505 87449 525 87477
rect 544 87449 553 87477
rect 544 87429 548 87449
rect 579 87408 582 87498
rect 612 87480 624 87481
rect 599 87478 649 87480
rect 612 87477 624 87478
rect 610 87470 632 87477
rect 607 87469 632 87470
rect 586 87462 644 87469
rect 607 87461 644 87462
rect 607 87445 610 87461
rect 616 87445 644 87461
rect 607 87444 644 87445
rect 586 87437 644 87444
rect 607 87436 610 87437
rect 612 87429 632 87437
rect 612 87425 624 87429
rect 649 87428 651 87478
rect 544 87391 548 87399
rect 400 87359 408 87389
rect 420 87359 436 87389
rect 400 87355 436 87359
rect 400 87347 430 87355
rect 428 87331 430 87347
rect 476 87319 480 87387
rect 544 87357 552 87391
rect 578 87357 582 87391
rect 544 87349 548 87357
rect 544 87319 586 87320
rect 288 87279 292 87311
rect 296 87309 368 87317
rect 378 87309 450 87317
rect 544 87312 548 87319
rect 439 87281 444 87309
rect 120 87265 170 87267
rect 76 87261 130 87265
rect 110 87256 130 87261
rect 60 87231 67 87241
rect 76 87231 77 87251
rect 96 87222 99 87256
rect 109 87231 110 87251
rect 119 87231 126 87241
rect 76 87215 92 87221
rect 94 87215 110 87221
rect 170 87215 172 87265
rect 186 87199 190 87233
rect 216 87199 220 87233
rect 213 87167 224 87199
rect 282 87195 292 87279
rect 296 87273 368 87281
rect 378 87273 450 87281
rect 468 87278 473 87312
rect 428 87243 430 87259
rect 251 87167 292 87195
rect 318 87174 324 87243
rect 12 87162 62 87164
rect 28 87153 59 87161
rect 62 87153 64 87162
rect 251 87161 263 87167
rect 28 87145 64 87153
rect 127 87153 158 87161
rect 127 87146 182 87153
rect 127 87145 161 87146
rect 59 87129 64 87145
rect 158 87129 161 87145
rect 253 87133 263 87161
rect 273 87133 293 87167
rect 318 87164 335 87174
rect 303 87148 316 87158
rect 318 87148 324 87164
rect 346 87158 348 87243
rect 400 87235 430 87243
rect 476 87241 480 87309
rect 511 87278 582 87312
rect 544 87271 548 87278
rect 400 87231 436 87235
rect 400 87201 408 87231
rect 420 87201 436 87231
rect 544 87233 548 87241
rect 28 87121 64 87129
rect 127 87128 161 87129
rect 127 87121 182 87128
rect 62 87112 64 87121
rect 282 87075 292 87133
rect 295 87124 324 87148
rect 333 87148 353 87158
rect 428 87154 430 87201
rect 476 87161 480 87229
rect 544 87199 552 87233
rect 578 87199 582 87233
rect 544 87191 548 87199
rect 367 87148 380 87154
rect 333 87124 380 87148
rect 318 87111 324 87124
rect 346 87111 348 87124
rect 367 87120 380 87124
rect 396 87120 408 87154
rect 420 87120 436 87154
rect 544 87151 553 87179
rect 319 87100 346 87111
rect 120 87059 170 87061
rect 76 87053 92 87059
rect 94 87053 110 87059
rect 76 87043 99 87052
rect 60 87033 67 87043
rect 76 87023 77 87043
rect 96 87018 99 87043
rect 109 87023 110 87043
rect 119 87033 126 87043
rect 76 87009 110 87013
rect 170 87009 172 87059
rect 186 87041 190 87075
rect 216 87041 220 87075
rect 182 87003 224 87004
rect 186 86979 220 86996
rect 223 86979 257 86996
rect 182 86962 257 86979
rect 182 86961 224 86962
rect 160 86955 246 86961
rect 288 86955 292 87075
rect 296 87073 368 87081
rect 428 87073 430 87120
rect 476 87083 480 87151
rect 485 87107 495 87141
rect 505 87113 525 87141
rect 505 87107 519 87113
rect 544 87107 555 87151
rect 485 87083 492 87107
rect 579 87092 582 87182
rect 612 87164 624 87165
rect 599 87162 649 87164
rect 612 87161 624 87162
rect 610 87154 632 87161
rect 607 87153 632 87154
rect 586 87146 644 87153
rect 607 87145 644 87146
rect 607 87129 610 87145
rect 616 87129 644 87145
rect 607 87128 644 87129
rect 586 87121 644 87128
rect 607 87120 610 87121
rect 612 87113 632 87121
rect 612 87109 624 87113
rect 649 87112 651 87162
rect 544 87075 548 87083
rect 400 87043 408 87073
rect 420 87043 436 87073
rect 400 87039 436 87043
rect 400 87031 430 87039
rect 428 87015 430 87031
rect 476 87003 480 87071
rect 544 87041 552 87075
rect 578 87041 582 87075
rect 544 87033 548 87041
rect 295 86962 300 86996
rect 324 86962 329 86996
rect 378 86993 450 87001
rect 544 86998 548 87003
rect 544 86994 582 86998
rect 544 86979 552 86994
rect 578 86979 582 86994
rect 544 86961 586 86979
rect 522 86955 608 86961
rect 182 86939 224 86955
rect 544 86939 586 86955
rect 17 86925 67 86927
rect 119 86925 169 86927
rect 186 86925 220 86939
rect 548 86925 582 86939
rect 599 86925 649 86927
rect 42 86883 59 86917
rect 67 86875 69 86925
rect 160 86917 246 86925
rect 522 86917 608 86925
rect 76 86883 110 86917
rect 127 86883 144 86917
rect 152 86883 161 86917
rect 162 86915 195 86917
rect 224 86915 244 86917
rect 162 86883 244 86915
rect 524 86915 548 86917
rect 573 86915 582 86917
rect 586 86915 606 86917
rect 160 86875 246 86883
rect 186 86859 220 86875
rect 182 86845 224 86846
rect 160 86839 182 86845
rect 224 86839 246 86845
rect 186 86804 220 86838
rect 223 86804 257 86838
rect 120 86791 170 86793
rect 76 86787 130 86791
rect 110 86782 130 86787
rect 60 86757 67 86767
rect 76 86757 77 86777
rect 96 86748 99 86782
rect 109 86757 110 86777
rect 119 86757 126 86767
rect 76 86741 92 86747
rect 94 86741 110 86747
rect 170 86741 172 86791
rect 186 86725 190 86759
rect 216 86725 220 86759
rect 288 86725 292 86913
rect 476 86845 480 86913
rect 524 86883 606 86915
rect 607 86883 616 86917
rect 522 86875 608 86883
rect 649 86875 651 86925
rect 548 86859 582 86875
rect 522 86840 548 86845
rect 522 86839 582 86840
rect 586 86839 608 86845
rect 295 86804 300 86838
rect 324 86804 329 86838
rect 544 86836 582 86839
rect 378 86799 450 86807
rect 428 86769 430 86785
rect 400 86761 430 86769
rect 476 86767 480 86835
rect 544 86806 552 86836
rect 578 86806 582 86836
rect 544 86797 548 86806
rect 400 86757 436 86761
rect 400 86727 408 86757
rect 420 86727 436 86757
rect 544 86759 548 86767
rect 12 86688 62 86690
rect 28 86679 59 86687
rect 62 86679 64 86688
rect 28 86671 64 86679
rect 127 86679 158 86687
rect 127 86672 182 86679
rect 215 86677 224 86705
rect 127 86671 161 86672
rect 59 86655 64 86671
rect 158 86655 161 86671
rect 28 86647 64 86655
rect 127 86654 161 86655
rect 127 86647 182 86654
rect 62 86638 64 86647
rect 213 86639 224 86677
rect 282 86667 292 86725
rect 296 86719 368 86727
rect 319 86689 346 86700
rect 318 86676 324 86689
rect 346 86676 348 86689
rect 428 86680 430 86727
rect 443 86717 450 86719
rect 476 86687 480 86755
rect 544 86725 552 86759
rect 578 86725 582 86759
rect 481 86693 517 86721
rect 481 86687 495 86693
rect 367 86676 380 86680
rect 251 86633 263 86667
rect 273 86633 293 86667
rect 295 86652 324 86676
rect 303 86642 316 86652
rect 318 86636 324 86652
rect 333 86652 380 86676
rect 333 86642 353 86652
rect 367 86646 380 86652
rect 396 86646 408 86680
rect 420 86646 436 86680
rect 120 86585 170 86587
rect 76 86579 92 86585
rect 94 86579 110 86585
rect 76 86569 99 86578
rect 60 86559 67 86569
rect 76 86549 77 86569
rect 96 86544 99 86569
rect 109 86549 110 86569
rect 119 86559 126 86569
rect 76 86535 110 86539
rect 170 86535 172 86585
rect 186 86567 190 86601
rect 216 86567 220 86601
rect 186 86490 220 86524
rect 282 86521 292 86633
rect 318 86626 335 86636
rect 318 86557 324 86626
rect 346 86557 348 86642
rect 428 86599 430 86646
rect 476 86609 480 86677
rect 485 86659 495 86687
rect 505 86687 519 86693
rect 544 86687 555 86725
rect 505 86659 525 86687
rect 544 86659 553 86687
rect 544 86639 548 86659
rect 579 86618 582 86708
rect 612 86690 624 86691
rect 599 86688 649 86690
rect 612 86687 624 86688
rect 610 86680 632 86687
rect 607 86679 632 86680
rect 586 86672 644 86679
rect 607 86671 644 86672
rect 607 86655 610 86671
rect 616 86655 644 86671
rect 607 86654 644 86655
rect 586 86647 644 86654
rect 607 86646 610 86647
rect 612 86639 632 86647
rect 612 86635 624 86639
rect 649 86638 651 86688
rect 544 86601 548 86609
rect 400 86569 408 86599
rect 420 86569 436 86599
rect 400 86565 436 86569
rect 400 86557 430 86565
rect 428 86541 430 86557
rect 476 86529 480 86597
rect 544 86567 552 86601
rect 578 86567 582 86601
rect 544 86559 548 86567
rect 544 86529 586 86530
rect 288 86489 292 86521
rect 296 86519 368 86527
rect 378 86519 450 86527
rect 544 86522 548 86529
rect 439 86491 444 86519
rect 120 86475 170 86477
rect 76 86471 130 86475
rect 110 86466 130 86471
rect 60 86441 67 86451
rect 76 86441 77 86461
rect 96 86432 99 86466
rect 109 86441 110 86461
rect 119 86441 126 86451
rect 76 86425 92 86431
rect 94 86425 110 86431
rect 170 86425 172 86475
rect 186 86409 190 86443
rect 216 86409 220 86443
rect 213 86377 224 86409
rect 282 86405 292 86489
rect 296 86483 368 86491
rect 378 86483 450 86491
rect 468 86488 473 86522
rect 428 86453 430 86469
rect 251 86377 292 86405
rect 318 86384 324 86453
rect 12 86372 62 86374
rect 28 86363 59 86371
rect 62 86363 64 86372
rect 251 86371 263 86377
rect 28 86355 64 86363
rect 127 86363 158 86371
rect 127 86356 182 86363
rect 127 86355 161 86356
rect 59 86339 64 86355
rect 158 86339 161 86355
rect 253 86343 263 86371
rect 273 86343 293 86377
rect 318 86374 335 86384
rect 303 86358 316 86368
rect 318 86358 324 86374
rect 346 86368 348 86453
rect 400 86445 430 86453
rect 476 86451 480 86519
rect 511 86488 582 86522
rect 544 86481 548 86488
rect 400 86441 436 86445
rect 400 86411 408 86441
rect 420 86411 436 86441
rect 544 86443 548 86451
rect 28 86331 64 86339
rect 127 86338 161 86339
rect 127 86331 182 86338
rect 62 86322 64 86331
rect 282 86285 292 86343
rect 295 86334 324 86358
rect 333 86358 353 86368
rect 428 86364 430 86411
rect 476 86371 480 86439
rect 544 86409 552 86443
rect 578 86409 582 86443
rect 544 86401 548 86409
rect 367 86358 380 86364
rect 333 86334 380 86358
rect 318 86321 324 86334
rect 346 86321 348 86334
rect 367 86330 380 86334
rect 396 86330 408 86364
rect 420 86330 436 86364
rect 544 86361 553 86389
rect 319 86310 346 86321
rect 120 86269 170 86271
rect 76 86263 92 86269
rect 94 86263 110 86269
rect 76 86253 99 86262
rect 60 86243 67 86253
rect 76 86233 77 86253
rect 96 86228 99 86253
rect 109 86233 110 86253
rect 119 86243 126 86253
rect 76 86219 110 86223
rect 170 86219 172 86269
rect 186 86251 190 86285
rect 216 86251 220 86285
rect 182 86213 224 86214
rect 186 86189 220 86206
rect 223 86189 257 86206
rect 182 86172 257 86189
rect 182 86171 224 86172
rect 160 86165 246 86171
rect 288 86165 292 86285
rect 296 86283 368 86291
rect 428 86283 430 86330
rect 476 86293 480 86361
rect 485 86317 495 86351
rect 505 86323 525 86351
rect 505 86317 519 86323
rect 544 86317 555 86361
rect 485 86293 492 86317
rect 579 86302 582 86392
rect 612 86374 624 86375
rect 599 86372 649 86374
rect 612 86371 624 86372
rect 610 86364 632 86371
rect 607 86363 632 86364
rect 586 86356 644 86363
rect 607 86355 644 86356
rect 607 86339 610 86355
rect 616 86339 644 86355
rect 607 86338 644 86339
rect 586 86331 644 86338
rect 607 86330 610 86331
rect 612 86323 632 86331
rect 612 86319 624 86323
rect 649 86322 651 86372
rect 544 86285 548 86293
rect 400 86253 408 86283
rect 420 86253 436 86283
rect 400 86249 436 86253
rect 400 86241 430 86249
rect 428 86225 430 86241
rect 476 86213 480 86281
rect 544 86251 552 86285
rect 578 86251 582 86285
rect 544 86243 548 86251
rect 295 86172 300 86206
rect 324 86172 329 86206
rect 378 86203 450 86211
rect 544 86208 548 86213
rect 544 86204 582 86208
rect 544 86189 552 86204
rect 578 86189 582 86204
rect 544 86171 586 86189
rect 522 86165 608 86171
rect 182 86149 224 86165
rect 544 86149 586 86165
rect 17 86135 67 86137
rect 119 86135 169 86137
rect 186 86135 220 86149
rect 548 86135 582 86149
rect 599 86135 649 86137
rect 42 86093 59 86127
rect 67 86085 69 86135
rect 160 86127 246 86135
rect 522 86127 608 86135
rect 76 86093 110 86127
rect 127 86093 144 86127
rect 152 86093 161 86127
rect 162 86125 195 86127
rect 224 86125 244 86127
rect 162 86093 244 86125
rect 524 86125 548 86127
rect 573 86125 582 86127
rect 586 86125 606 86127
rect 160 86085 246 86093
rect 186 86069 220 86085
rect 182 86055 224 86056
rect 160 86049 182 86055
rect 224 86049 246 86055
rect 186 86014 220 86048
rect 223 86014 257 86048
rect 120 86001 170 86003
rect 76 85997 130 86001
rect 110 85992 130 85997
rect 60 85967 67 85977
rect 76 85967 77 85987
rect 96 85958 99 85992
rect 109 85967 110 85987
rect 119 85967 126 85977
rect 76 85951 92 85957
rect 94 85951 110 85957
rect 170 85951 172 86001
rect 186 85935 190 85969
rect 216 85935 220 85969
rect 288 85935 292 86123
rect 476 86055 480 86123
rect 524 86093 606 86125
rect 607 86093 616 86127
rect 522 86085 608 86093
rect 649 86085 651 86135
rect 548 86069 582 86085
rect 522 86050 548 86055
rect 522 86049 582 86050
rect 586 86049 608 86055
rect 295 86014 300 86048
rect 324 86014 329 86048
rect 544 86046 582 86049
rect 378 86009 450 86017
rect 428 85979 430 85995
rect 400 85971 430 85979
rect 476 85977 480 86045
rect 544 86016 552 86046
rect 578 86016 582 86046
rect 544 86007 548 86016
rect 400 85967 436 85971
rect 400 85937 408 85967
rect 420 85937 436 85967
rect 544 85969 548 85977
rect 12 85898 62 85900
rect 28 85889 59 85897
rect 62 85889 64 85898
rect 28 85881 64 85889
rect 127 85889 158 85897
rect 127 85882 182 85889
rect 215 85887 224 85915
rect 127 85881 161 85882
rect 59 85865 64 85881
rect 158 85865 161 85881
rect 28 85857 64 85865
rect 127 85864 161 85865
rect 127 85857 182 85864
rect 62 85848 64 85857
rect 213 85849 224 85887
rect 282 85877 292 85935
rect 296 85929 368 85937
rect 319 85899 346 85910
rect 318 85886 324 85899
rect 346 85886 348 85899
rect 428 85890 430 85937
rect 443 85927 450 85929
rect 476 85897 480 85965
rect 544 85935 552 85969
rect 578 85935 582 85969
rect 481 85903 517 85931
rect 481 85897 495 85903
rect 367 85886 380 85890
rect 251 85843 263 85877
rect 273 85843 293 85877
rect 295 85862 324 85886
rect 303 85852 316 85862
rect 318 85846 324 85862
rect 333 85862 380 85886
rect 333 85852 353 85862
rect 367 85856 380 85862
rect 396 85856 408 85890
rect 420 85856 436 85890
rect 120 85795 170 85797
rect 76 85789 92 85795
rect 94 85789 110 85795
rect 76 85779 99 85788
rect 60 85769 67 85779
rect 76 85759 77 85779
rect 96 85754 99 85779
rect 109 85759 110 85779
rect 119 85769 126 85779
rect 76 85745 110 85749
rect 170 85745 172 85795
rect 186 85777 190 85811
rect 216 85777 220 85811
rect 186 85700 220 85734
rect 282 85731 292 85843
rect 318 85836 335 85846
rect 318 85767 324 85836
rect 346 85767 348 85852
rect 428 85809 430 85856
rect 476 85819 480 85887
rect 485 85869 495 85897
rect 505 85897 519 85903
rect 544 85897 555 85935
rect 505 85869 525 85897
rect 544 85869 553 85897
rect 544 85849 548 85869
rect 579 85828 582 85918
rect 612 85900 624 85901
rect 599 85898 649 85900
rect 612 85897 624 85898
rect 610 85890 632 85897
rect 607 85889 632 85890
rect 586 85882 644 85889
rect 607 85881 644 85882
rect 607 85865 610 85881
rect 616 85865 644 85881
rect 607 85864 644 85865
rect 586 85857 644 85864
rect 607 85856 610 85857
rect 612 85849 632 85857
rect 612 85845 624 85849
rect 649 85848 651 85898
rect 544 85811 548 85819
rect 400 85779 408 85809
rect 420 85779 436 85809
rect 400 85775 436 85779
rect 400 85767 430 85775
rect 428 85751 430 85767
rect 476 85739 480 85807
rect 544 85777 552 85811
rect 578 85777 582 85811
rect 544 85769 548 85777
rect 544 85739 586 85740
rect 288 85699 292 85731
rect 296 85729 368 85737
rect 378 85729 450 85737
rect 544 85732 548 85739
rect 439 85701 444 85729
rect 120 85685 170 85687
rect 76 85681 130 85685
rect 110 85676 130 85681
rect 60 85651 67 85661
rect 76 85651 77 85671
rect 96 85642 99 85676
rect 109 85651 110 85671
rect 119 85651 126 85661
rect 76 85635 92 85641
rect 94 85635 110 85641
rect 170 85635 172 85685
rect 186 85619 190 85653
rect 216 85619 220 85653
rect 213 85587 224 85619
rect 282 85615 292 85699
rect 296 85693 368 85701
rect 378 85693 450 85701
rect 468 85698 473 85732
rect 428 85663 430 85679
rect 251 85587 292 85615
rect 318 85594 324 85663
rect 12 85582 62 85584
rect 28 85573 59 85581
rect 62 85573 64 85582
rect 251 85581 263 85587
rect 28 85565 64 85573
rect 127 85573 158 85581
rect 127 85566 182 85573
rect 127 85565 161 85566
rect 59 85549 64 85565
rect 158 85549 161 85565
rect 253 85553 263 85581
rect 273 85553 293 85587
rect 318 85584 335 85594
rect 303 85568 316 85578
rect 318 85568 324 85584
rect 346 85578 348 85663
rect 400 85655 430 85663
rect 476 85661 480 85729
rect 511 85698 582 85732
rect 544 85691 548 85698
rect 400 85651 436 85655
rect 400 85621 408 85651
rect 420 85621 436 85651
rect 544 85653 548 85661
rect 28 85541 64 85549
rect 127 85548 161 85549
rect 127 85541 182 85548
rect 62 85532 64 85541
rect 282 85495 292 85553
rect 295 85544 324 85568
rect 333 85568 353 85578
rect 428 85574 430 85621
rect 476 85581 480 85649
rect 544 85619 552 85653
rect 578 85619 582 85653
rect 544 85611 548 85619
rect 367 85568 380 85574
rect 333 85544 380 85568
rect 318 85531 324 85544
rect 346 85531 348 85544
rect 367 85540 380 85544
rect 396 85540 408 85574
rect 420 85540 436 85574
rect 544 85571 553 85599
rect 319 85520 346 85531
rect 120 85479 170 85481
rect 76 85473 92 85479
rect 94 85473 110 85479
rect 76 85463 99 85472
rect 60 85453 67 85463
rect 76 85443 77 85463
rect 96 85438 99 85463
rect 109 85443 110 85463
rect 119 85453 126 85463
rect 76 85429 110 85433
rect 170 85429 172 85479
rect 186 85461 190 85495
rect 216 85461 220 85495
rect 182 85423 224 85424
rect 186 85399 220 85416
rect 223 85399 257 85416
rect 182 85382 257 85399
rect 182 85381 224 85382
rect 160 85375 246 85381
rect 288 85375 292 85495
rect 296 85493 368 85501
rect 428 85493 430 85540
rect 476 85503 480 85571
rect 485 85527 495 85561
rect 505 85533 525 85561
rect 505 85527 519 85533
rect 544 85527 555 85571
rect 485 85503 492 85527
rect 579 85512 582 85602
rect 612 85584 624 85585
rect 599 85582 649 85584
rect 612 85581 624 85582
rect 610 85574 632 85581
rect 607 85573 632 85574
rect 586 85566 644 85573
rect 607 85565 644 85566
rect 607 85549 610 85565
rect 616 85549 644 85565
rect 607 85548 644 85549
rect 586 85541 644 85548
rect 607 85540 610 85541
rect 612 85533 632 85541
rect 612 85529 624 85533
rect 649 85532 651 85582
rect 544 85495 548 85503
rect 400 85463 408 85493
rect 420 85463 436 85493
rect 400 85459 436 85463
rect 400 85451 430 85459
rect 428 85435 430 85451
rect 476 85423 480 85491
rect 544 85461 552 85495
rect 578 85461 582 85495
rect 544 85453 548 85461
rect 295 85382 300 85416
rect 324 85382 329 85416
rect 378 85413 450 85421
rect 544 85418 548 85423
rect 544 85414 582 85418
rect 544 85399 552 85414
rect 578 85399 582 85414
rect 544 85381 586 85399
rect 522 85375 608 85381
rect 182 85359 224 85375
rect 544 85359 586 85375
rect 17 85345 67 85347
rect 119 85345 169 85347
rect 186 85345 220 85359
rect 548 85345 582 85359
rect 599 85345 649 85347
rect 42 85303 59 85337
rect 67 85295 69 85345
rect 160 85337 246 85345
rect 522 85337 608 85345
rect 76 85303 110 85337
rect 127 85303 144 85337
rect 152 85303 161 85337
rect 162 85335 195 85337
rect 224 85335 244 85337
rect 162 85303 244 85335
rect 524 85335 548 85337
rect 573 85335 582 85337
rect 586 85335 606 85337
rect 160 85295 246 85303
rect 186 85279 220 85295
rect 182 85265 224 85266
rect 160 85259 182 85265
rect 224 85259 246 85265
rect 186 85224 220 85258
rect 223 85224 257 85258
rect 120 85211 170 85213
rect 76 85207 130 85211
rect 110 85202 130 85207
rect 60 85177 67 85187
rect 76 85177 77 85197
rect 96 85168 99 85202
rect 109 85177 110 85197
rect 119 85177 126 85187
rect 76 85161 92 85167
rect 94 85161 110 85167
rect 170 85161 172 85211
rect 186 85145 190 85179
rect 216 85145 220 85179
rect 288 85145 292 85333
rect 476 85265 480 85333
rect 524 85303 606 85335
rect 607 85303 616 85337
rect 522 85295 608 85303
rect 649 85295 651 85345
rect 548 85279 582 85295
rect 522 85260 548 85265
rect 522 85259 582 85260
rect 586 85259 608 85265
rect 295 85224 300 85258
rect 324 85224 329 85258
rect 544 85256 582 85259
rect 378 85219 450 85227
rect 428 85189 430 85205
rect 400 85181 430 85189
rect 476 85187 480 85255
rect 544 85226 552 85256
rect 578 85226 582 85256
rect 544 85217 548 85226
rect 400 85177 436 85181
rect 400 85147 408 85177
rect 420 85147 436 85177
rect 544 85179 548 85187
rect 12 85108 62 85110
rect 28 85099 59 85107
rect 62 85099 64 85108
rect 28 85091 64 85099
rect 127 85099 158 85107
rect 127 85092 182 85099
rect 215 85097 224 85125
rect 127 85091 161 85092
rect 59 85075 64 85091
rect 158 85075 161 85091
rect 28 85067 64 85075
rect 127 85074 161 85075
rect 127 85067 182 85074
rect 62 85058 64 85067
rect 213 85059 224 85097
rect 282 85087 292 85145
rect 296 85139 368 85147
rect 319 85109 346 85120
rect 318 85096 324 85109
rect 346 85096 348 85109
rect 428 85100 430 85147
rect 443 85137 450 85139
rect 476 85107 480 85175
rect 544 85145 552 85179
rect 578 85145 582 85179
rect 481 85113 517 85141
rect 481 85107 495 85113
rect 367 85096 380 85100
rect 251 85053 263 85087
rect 273 85053 293 85087
rect 295 85072 324 85096
rect 303 85062 316 85072
rect 318 85056 324 85072
rect 333 85072 380 85096
rect 333 85062 353 85072
rect 367 85066 380 85072
rect 396 85066 408 85100
rect 420 85066 436 85100
rect 120 85005 170 85007
rect 76 84999 92 85005
rect 94 84999 110 85005
rect 76 84989 99 84998
rect 60 84979 67 84989
rect 76 84969 77 84989
rect 96 84964 99 84989
rect 109 84969 110 84989
rect 119 84979 126 84989
rect 76 84955 110 84959
rect 170 84955 172 85005
rect 186 84987 190 85021
rect 216 84987 220 85021
rect 186 84910 220 84944
rect 282 84941 292 85053
rect 318 85046 335 85056
rect 318 84977 324 85046
rect 346 84977 348 85062
rect 428 85019 430 85066
rect 476 85029 480 85097
rect 485 85079 495 85107
rect 505 85107 519 85113
rect 544 85107 555 85145
rect 505 85079 525 85107
rect 544 85079 553 85107
rect 544 85059 548 85079
rect 579 85038 582 85128
rect 612 85110 624 85111
rect 599 85108 649 85110
rect 612 85107 624 85108
rect 610 85100 632 85107
rect 607 85099 632 85100
rect 586 85092 644 85099
rect 607 85091 644 85092
rect 607 85075 610 85091
rect 616 85075 644 85091
rect 607 85074 644 85075
rect 586 85067 644 85074
rect 607 85066 610 85067
rect 612 85059 632 85067
rect 612 85055 624 85059
rect 649 85058 651 85108
rect 544 85021 548 85029
rect 400 84989 408 85019
rect 420 84989 436 85019
rect 400 84985 436 84989
rect 400 84977 430 84985
rect 428 84961 430 84977
rect 476 84949 480 85017
rect 544 84987 552 85021
rect 578 84987 582 85021
rect 544 84979 548 84987
rect 544 84949 586 84950
rect 288 84909 292 84941
rect 296 84939 368 84947
rect 378 84939 450 84947
rect 544 84942 548 84949
rect 439 84911 444 84939
rect 120 84895 170 84897
rect 76 84891 130 84895
rect 110 84886 130 84891
rect 60 84861 67 84871
rect 76 84861 77 84881
rect 96 84852 99 84886
rect 109 84861 110 84881
rect 119 84861 126 84871
rect 76 84845 92 84851
rect 94 84845 110 84851
rect 170 84845 172 84895
rect 186 84829 190 84863
rect 216 84829 220 84863
rect 213 84797 224 84829
rect 282 84825 292 84909
rect 296 84903 368 84911
rect 378 84903 450 84911
rect 468 84908 473 84942
rect 428 84873 430 84889
rect 251 84797 292 84825
rect 318 84804 324 84873
rect 12 84792 62 84794
rect 28 84783 59 84791
rect 62 84783 64 84792
rect 251 84791 263 84797
rect 28 84775 64 84783
rect 127 84783 158 84791
rect 127 84776 182 84783
rect 127 84775 161 84776
rect 59 84759 64 84775
rect 158 84759 161 84775
rect 253 84763 263 84791
rect 273 84763 293 84797
rect 318 84794 335 84804
rect 303 84778 316 84788
rect 318 84778 324 84794
rect 346 84788 348 84873
rect 400 84865 430 84873
rect 476 84871 480 84939
rect 511 84908 582 84942
rect 544 84901 548 84908
rect 400 84861 436 84865
rect 400 84831 408 84861
rect 420 84831 436 84861
rect 544 84863 548 84871
rect 28 84751 64 84759
rect 127 84758 161 84759
rect 127 84751 182 84758
rect 62 84742 64 84751
rect 282 84705 292 84763
rect 295 84754 324 84778
rect 333 84778 353 84788
rect 428 84784 430 84831
rect 476 84791 480 84859
rect 544 84829 552 84863
rect 578 84829 582 84863
rect 544 84821 548 84829
rect 367 84778 380 84784
rect 333 84754 380 84778
rect 318 84741 324 84754
rect 346 84741 348 84754
rect 367 84750 380 84754
rect 396 84750 408 84784
rect 420 84750 436 84784
rect 544 84781 553 84809
rect 319 84730 346 84741
rect 120 84689 170 84691
rect 76 84683 92 84689
rect 94 84683 110 84689
rect 76 84673 99 84682
rect 60 84663 67 84673
rect 76 84653 77 84673
rect 96 84648 99 84673
rect 109 84653 110 84673
rect 119 84663 126 84673
rect 76 84639 110 84643
rect 170 84639 172 84689
rect 186 84671 190 84705
rect 216 84671 220 84705
rect 182 84633 224 84634
rect 186 84609 220 84626
rect 223 84609 257 84626
rect 182 84592 257 84609
rect 182 84591 224 84592
rect 160 84585 246 84591
rect 288 84585 292 84705
rect 296 84703 368 84711
rect 428 84703 430 84750
rect 476 84713 480 84781
rect 485 84737 495 84771
rect 505 84743 525 84771
rect 505 84737 519 84743
rect 544 84737 555 84781
rect 485 84713 492 84737
rect 579 84722 582 84812
rect 612 84794 624 84795
rect 599 84792 649 84794
rect 612 84791 624 84792
rect 610 84784 632 84791
rect 607 84783 632 84784
rect 586 84776 644 84783
rect 607 84775 644 84776
rect 607 84759 610 84775
rect 616 84759 644 84775
rect 607 84758 644 84759
rect 586 84751 644 84758
rect 607 84750 610 84751
rect 612 84743 632 84751
rect 612 84739 624 84743
rect 649 84742 651 84792
rect 544 84705 548 84713
rect 400 84673 408 84703
rect 420 84673 436 84703
rect 400 84669 436 84673
rect 400 84661 430 84669
rect 428 84645 430 84661
rect 476 84633 480 84701
rect 544 84671 552 84705
rect 578 84671 582 84705
rect 544 84663 548 84671
rect 295 84592 300 84626
rect 324 84592 329 84626
rect 378 84623 450 84631
rect 544 84628 548 84633
rect 544 84624 582 84628
rect 544 84609 552 84624
rect 578 84609 582 84624
rect 544 84591 586 84609
rect 522 84585 608 84591
rect 182 84569 224 84585
rect 544 84569 586 84585
rect 17 84555 67 84557
rect 119 84555 169 84557
rect 186 84555 220 84569
rect 548 84555 582 84569
rect 599 84555 649 84557
rect 42 84513 59 84547
rect 67 84505 69 84555
rect 160 84547 246 84555
rect 522 84547 608 84555
rect 76 84513 110 84547
rect 127 84513 144 84547
rect 152 84513 161 84547
rect 162 84545 195 84547
rect 224 84545 244 84547
rect 162 84513 244 84545
rect 524 84545 548 84547
rect 573 84545 582 84547
rect 586 84545 606 84547
rect 160 84505 246 84513
rect 186 84489 220 84505
rect 182 84475 224 84476
rect 160 84469 182 84475
rect 224 84469 246 84475
rect 186 84434 220 84468
rect 223 84434 257 84468
rect 120 84421 170 84423
rect 76 84417 130 84421
rect 110 84412 130 84417
rect 60 84387 67 84397
rect 76 84387 77 84407
rect 96 84378 99 84412
rect 109 84387 110 84407
rect 119 84387 126 84397
rect 76 84371 92 84377
rect 94 84371 110 84377
rect 170 84371 172 84421
rect 186 84355 190 84389
rect 216 84355 220 84389
rect 288 84355 292 84543
rect 476 84475 480 84543
rect 524 84513 606 84545
rect 607 84513 616 84547
rect 522 84505 608 84513
rect 649 84505 651 84555
rect 548 84489 582 84505
rect 522 84470 548 84475
rect 522 84469 582 84470
rect 586 84469 608 84475
rect 295 84434 300 84468
rect 324 84434 329 84468
rect 544 84466 582 84469
rect 378 84429 450 84437
rect 428 84399 430 84415
rect 400 84391 430 84399
rect 476 84397 480 84465
rect 544 84436 552 84466
rect 578 84436 582 84466
rect 544 84427 548 84436
rect 400 84387 436 84391
rect 400 84357 408 84387
rect 420 84357 436 84387
rect 544 84389 548 84397
rect 12 84318 62 84320
rect 28 84309 59 84317
rect 62 84309 64 84318
rect 28 84301 64 84309
rect 127 84309 158 84317
rect 127 84302 182 84309
rect 215 84307 224 84335
rect 127 84301 161 84302
rect 59 84285 64 84301
rect 158 84285 161 84301
rect 28 84277 64 84285
rect 127 84284 161 84285
rect 127 84277 182 84284
rect 62 84268 64 84277
rect 213 84269 224 84307
rect 282 84297 292 84355
rect 296 84349 368 84357
rect 319 84319 346 84330
rect 318 84306 324 84319
rect 346 84306 348 84319
rect 428 84310 430 84357
rect 443 84347 450 84349
rect 476 84317 480 84385
rect 544 84355 552 84389
rect 578 84355 582 84389
rect 481 84323 517 84351
rect 481 84317 495 84323
rect 367 84306 380 84310
rect 251 84263 263 84297
rect 273 84263 293 84297
rect 295 84282 324 84306
rect 303 84272 316 84282
rect 318 84266 324 84282
rect 333 84282 380 84306
rect 333 84272 353 84282
rect 367 84276 380 84282
rect 396 84276 408 84310
rect 420 84276 436 84310
rect 120 84215 170 84217
rect 76 84209 92 84215
rect 94 84209 110 84215
rect 76 84199 99 84208
rect 60 84189 67 84199
rect 76 84179 77 84199
rect 96 84174 99 84199
rect 109 84179 110 84199
rect 119 84189 126 84199
rect 76 84165 110 84169
rect 170 84165 172 84215
rect 186 84197 190 84231
rect 216 84197 220 84231
rect 186 84120 220 84154
rect 282 84151 292 84263
rect 318 84256 335 84266
rect 318 84187 324 84256
rect 346 84187 348 84272
rect 428 84229 430 84276
rect 476 84239 480 84307
rect 485 84289 495 84317
rect 505 84317 519 84323
rect 544 84317 555 84355
rect 505 84289 525 84317
rect 544 84289 553 84317
rect 544 84269 548 84289
rect 579 84248 582 84338
rect 612 84320 624 84321
rect 599 84318 649 84320
rect 612 84317 624 84318
rect 610 84310 632 84317
rect 607 84309 632 84310
rect 586 84302 644 84309
rect 607 84301 644 84302
rect 607 84285 610 84301
rect 616 84285 644 84301
rect 607 84284 644 84285
rect 586 84277 644 84284
rect 607 84276 610 84277
rect 612 84269 632 84277
rect 612 84265 624 84269
rect 649 84268 651 84318
rect 544 84231 548 84239
rect 400 84199 408 84229
rect 420 84199 436 84229
rect 400 84195 436 84199
rect 400 84187 430 84195
rect 428 84171 430 84187
rect 476 84159 480 84227
rect 544 84197 552 84231
rect 578 84197 582 84231
rect 544 84189 548 84197
rect 544 84159 586 84160
rect 288 84119 292 84151
rect 296 84149 368 84157
rect 378 84149 450 84157
rect 544 84152 548 84159
rect 439 84121 444 84149
rect 120 84105 170 84107
rect 76 84101 130 84105
rect 110 84096 130 84101
rect 60 84071 67 84081
rect 76 84071 77 84091
rect 96 84062 99 84096
rect 109 84071 110 84091
rect 119 84071 126 84081
rect 76 84055 92 84061
rect 94 84055 110 84061
rect 170 84055 172 84105
rect 186 84039 190 84073
rect 216 84039 220 84073
rect 213 84007 224 84039
rect 282 84035 292 84119
rect 296 84113 368 84121
rect 378 84113 450 84121
rect 468 84118 473 84152
rect 428 84083 430 84099
rect 251 84007 292 84035
rect 318 84014 324 84083
rect 12 84002 62 84004
rect 28 83993 59 84001
rect 62 83993 64 84002
rect 251 84001 263 84007
rect 28 83985 64 83993
rect 127 83993 158 84001
rect 127 83986 182 83993
rect 127 83985 161 83986
rect 59 83969 64 83985
rect 158 83969 161 83985
rect 253 83973 263 84001
rect 273 83973 293 84007
rect 318 84004 335 84014
rect 303 83988 316 83998
rect 318 83988 324 84004
rect 346 83998 348 84083
rect 400 84075 430 84083
rect 476 84081 480 84149
rect 511 84118 582 84152
rect 544 84111 548 84118
rect 400 84071 436 84075
rect 400 84041 408 84071
rect 420 84041 436 84071
rect 544 84073 548 84081
rect 28 83961 64 83969
rect 127 83968 161 83969
rect 127 83961 182 83968
rect 62 83952 64 83961
rect 282 83915 292 83973
rect 295 83964 324 83988
rect 333 83988 353 83998
rect 428 83994 430 84041
rect 476 84001 480 84069
rect 544 84039 552 84073
rect 578 84039 582 84073
rect 544 84031 548 84039
rect 367 83988 380 83994
rect 333 83964 380 83988
rect 318 83951 324 83964
rect 346 83951 348 83964
rect 367 83960 380 83964
rect 396 83960 408 83994
rect 420 83960 436 83994
rect 544 83991 553 84019
rect 319 83940 346 83951
rect 120 83899 170 83901
rect 76 83893 92 83899
rect 94 83893 110 83899
rect 76 83883 99 83892
rect 60 83873 67 83883
rect 76 83863 77 83883
rect 96 83858 99 83883
rect 109 83863 110 83883
rect 119 83873 126 83883
rect 76 83849 110 83853
rect 170 83849 172 83899
rect 186 83881 190 83915
rect 216 83881 220 83915
rect 182 83843 224 83844
rect 186 83819 220 83836
rect 223 83819 257 83836
rect 182 83802 257 83819
rect 182 83801 224 83802
rect 160 83795 246 83801
rect 288 83795 292 83915
rect 296 83913 368 83921
rect 428 83913 430 83960
rect 476 83923 480 83991
rect 485 83947 495 83981
rect 505 83953 525 83981
rect 505 83947 519 83953
rect 544 83947 555 83991
rect 485 83923 492 83947
rect 579 83932 582 84022
rect 612 84004 624 84005
rect 599 84002 649 84004
rect 612 84001 624 84002
rect 610 83994 632 84001
rect 607 83993 632 83994
rect 586 83986 644 83993
rect 607 83985 644 83986
rect 607 83969 610 83985
rect 616 83969 644 83985
rect 607 83968 644 83969
rect 586 83961 644 83968
rect 607 83960 610 83961
rect 612 83953 632 83961
rect 612 83949 624 83953
rect 649 83952 651 84002
rect 544 83915 548 83923
rect 400 83883 408 83913
rect 420 83883 436 83913
rect 400 83879 436 83883
rect 400 83871 430 83879
rect 428 83855 430 83871
rect 476 83843 480 83911
rect 544 83881 552 83915
rect 578 83881 582 83915
rect 544 83873 548 83881
rect 295 83802 300 83836
rect 324 83802 329 83836
rect 378 83833 450 83841
rect 544 83838 548 83843
rect 544 83834 582 83838
rect 544 83819 552 83834
rect 578 83819 582 83834
rect 544 83801 586 83819
rect 522 83795 608 83801
rect 182 83779 224 83795
rect 544 83779 586 83795
rect 17 83765 67 83767
rect 119 83765 169 83767
rect 186 83765 220 83779
rect 548 83765 582 83779
rect 599 83765 649 83767
rect 42 83723 59 83757
rect 67 83715 69 83765
rect 160 83757 246 83765
rect 522 83757 608 83765
rect 76 83723 110 83757
rect 127 83723 144 83757
rect 152 83723 161 83757
rect 162 83755 195 83757
rect 224 83755 244 83757
rect 162 83723 244 83755
rect 524 83755 548 83757
rect 573 83755 582 83757
rect 586 83755 606 83757
rect 160 83715 246 83723
rect 186 83699 220 83715
rect 182 83685 224 83686
rect 160 83679 182 83685
rect 224 83679 246 83685
rect 186 83644 220 83678
rect 223 83644 257 83678
rect 120 83631 170 83633
rect 76 83627 130 83631
rect 110 83622 130 83627
rect 60 83597 67 83607
rect 76 83597 77 83617
rect 96 83588 99 83622
rect 109 83597 110 83617
rect 119 83597 126 83607
rect 76 83581 92 83587
rect 94 83581 110 83587
rect 170 83581 172 83631
rect 186 83565 190 83599
rect 216 83565 220 83599
rect 288 83565 292 83753
rect 476 83685 480 83753
rect 524 83723 606 83755
rect 607 83723 616 83757
rect 522 83715 608 83723
rect 649 83715 651 83765
rect 548 83699 582 83715
rect 522 83680 548 83685
rect 522 83679 582 83680
rect 586 83679 608 83685
rect 295 83644 300 83678
rect 324 83644 329 83678
rect 544 83676 582 83679
rect 378 83639 450 83647
rect 428 83609 430 83625
rect 400 83601 430 83609
rect 476 83607 480 83675
rect 544 83646 552 83676
rect 578 83646 582 83676
rect 544 83637 548 83646
rect 400 83597 436 83601
rect 400 83567 408 83597
rect 420 83567 436 83597
rect 544 83599 548 83607
rect 12 83528 62 83530
rect 28 83519 59 83527
rect 62 83519 64 83528
rect 28 83511 64 83519
rect 127 83519 158 83527
rect 127 83512 182 83519
rect 215 83517 224 83545
rect 127 83511 161 83512
rect 59 83495 64 83511
rect 158 83495 161 83511
rect 28 83487 64 83495
rect 127 83494 161 83495
rect 127 83487 182 83494
rect 62 83478 64 83487
rect 213 83479 224 83517
rect 282 83507 292 83565
rect 296 83559 368 83567
rect 319 83529 346 83540
rect 318 83516 324 83529
rect 346 83516 348 83529
rect 428 83520 430 83567
rect 443 83557 450 83559
rect 476 83527 480 83595
rect 544 83565 552 83599
rect 578 83565 582 83599
rect 481 83533 517 83561
rect 481 83527 495 83533
rect 367 83516 380 83520
rect 251 83473 263 83507
rect 273 83473 293 83507
rect 295 83492 324 83516
rect 303 83482 316 83492
rect 318 83476 324 83492
rect 333 83492 380 83516
rect 333 83482 353 83492
rect 367 83486 380 83492
rect 396 83486 408 83520
rect 420 83486 436 83520
rect 120 83425 170 83427
rect 76 83419 92 83425
rect 94 83419 110 83425
rect 76 83409 99 83418
rect 60 83399 67 83409
rect 76 83389 77 83409
rect 96 83384 99 83409
rect 109 83389 110 83409
rect 119 83399 126 83409
rect 76 83375 110 83379
rect 170 83375 172 83425
rect 186 83407 190 83441
rect 216 83407 220 83441
rect 186 83330 220 83364
rect 282 83361 292 83473
rect 318 83466 335 83476
rect 318 83397 324 83466
rect 346 83397 348 83482
rect 428 83439 430 83486
rect 476 83449 480 83517
rect 485 83499 495 83527
rect 505 83527 519 83533
rect 544 83527 555 83565
rect 505 83499 525 83527
rect 544 83499 553 83527
rect 544 83479 548 83499
rect 579 83458 582 83548
rect 612 83530 624 83531
rect 599 83528 649 83530
rect 612 83527 624 83528
rect 610 83520 632 83527
rect 607 83519 632 83520
rect 586 83512 644 83519
rect 607 83511 644 83512
rect 607 83495 610 83511
rect 616 83495 644 83511
rect 607 83494 644 83495
rect 586 83487 644 83494
rect 607 83486 610 83487
rect 612 83479 632 83487
rect 612 83475 624 83479
rect 649 83478 651 83528
rect 544 83441 548 83449
rect 400 83409 408 83439
rect 420 83409 436 83439
rect 400 83405 436 83409
rect 400 83397 430 83405
rect 428 83381 430 83397
rect 476 83369 480 83437
rect 544 83407 552 83441
rect 578 83407 582 83441
rect 544 83399 548 83407
rect 544 83369 586 83370
rect 288 83329 292 83361
rect 296 83359 368 83367
rect 378 83359 450 83367
rect 544 83362 548 83369
rect 439 83331 444 83359
rect 120 83315 170 83317
rect 76 83311 130 83315
rect 110 83306 130 83311
rect 60 83281 67 83291
rect 76 83281 77 83301
rect 96 83272 99 83306
rect 109 83281 110 83301
rect 119 83281 126 83291
rect 76 83265 92 83271
rect 94 83265 110 83271
rect 170 83265 172 83315
rect 186 83249 190 83283
rect 216 83249 220 83283
rect 213 83217 224 83249
rect 282 83245 292 83329
rect 296 83323 368 83331
rect 378 83323 450 83331
rect 468 83328 473 83362
rect 428 83293 430 83309
rect 251 83217 292 83245
rect 318 83224 324 83293
rect 12 83212 62 83214
rect 28 83203 59 83211
rect 62 83203 64 83212
rect 251 83211 263 83217
rect 28 83195 64 83203
rect 127 83203 158 83211
rect 127 83196 182 83203
rect 127 83195 161 83196
rect 59 83179 64 83195
rect 158 83179 161 83195
rect 253 83183 263 83211
rect 273 83183 293 83217
rect 318 83214 335 83224
rect 303 83198 316 83208
rect 318 83198 324 83214
rect 346 83208 348 83293
rect 400 83285 430 83293
rect 476 83291 480 83359
rect 511 83328 582 83362
rect 544 83321 548 83328
rect 400 83281 436 83285
rect 400 83251 408 83281
rect 420 83251 436 83281
rect 544 83283 548 83291
rect 28 83171 64 83179
rect 127 83178 161 83179
rect 127 83171 182 83178
rect 62 83162 64 83171
rect 282 83125 292 83183
rect 295 83174 324 83198
rect 333 83198 353 83208
rect 428 83204 430 83251
rect 476 83211 480 83279
rect 544 83249 552 83283
rect 578 83249 582 83283
rect 544 83241 548 83249
rect 367 83198 380 83204
rect 333 83174 380 83198
rect 318 83161 324 83174
rect 346 83161 348 83174
rect 367 83170 380 83174
rect 396 83170 408 83204
rect 420 83170 436 83204
rect 544 83201 553 83229
rect 319 83150 346 83161
rect 120 83109 170 83111
rect 76 83103 92 83109
rect 94 83103 110 83109
rect 76 83093 99 83102
rect 60 83083 67 83093
rect 76 83073 77 83093
rect 96 83068 99 83093
rect 109 83073 110 83093
rect 119 83083 126 83093
rect 76 83059 110 83063
rect 170 83059 172 83109
rect 186 83091 190 83125
rect 216 83091 220 83125
rect 182 83053 224 83054
rect 186 83029 220 83046
rect 223 83029 257 83046
rect 182 83012 257 83029
rect 182 83011 224 83012
rect 160 83005 246 83011
rect 288 83005 292 83125
rect 296 83123 368 83131
rect 428 83123 430 83170
rect 476 83133 480 83201
rect 485 83157 495 83191
rect 505 83163 525 83191
rect 505 83157 519 83163
rect 544 83157 555 83201
rect 485 83133 492 83157
rect 579 83142 582 83232
rect 612 83214 624 83215
rect 599 83212 649 83214
rect 612 83211 624 83212
rect 610 83204 632 83211
rect 607 83203 632 83204
rect 586 83196 644 83203
rect 607 83195 644 83196
rect 607 83179 610 83195
rect 616 83179 644 83195
rect 607 83178 644 83179
rect 586 83171 644 83178
rect 607 83170 610 83171
rect 612 83163 632 83171
rect 612 83159 624 83163
rect 649 83162 651 83212
rect 544 83125 548 83133
rect 400 83093 408 83123
rect 420 83093 436 83123
rect 400 83089 436 83093
rect 400 83081 430 83089
rect 428 83065 430 83081
rect 476 83053 480 83121
rect 544 83091 552 83125
rect 578 83091 582 83125
rect 544 83083 548 83091
rect 295 83012 300 83046
rect 324 83012 329 83046
rect 378 83043 450 83051
rect 544 83048 548 83053
rect 544 83044 582 83048
rect 544 83029 552 83044
rect 578 83029 582 83044
rect 544 83011 586 83029
rect 522 83005 608 83011
rect 182 82989 224 83005
rect 544 82989 586 83005
rect 17 82975 67 82977
rect 119 82975 169 82977
rect 186 82975 220 82989
rect 548 82975 582 82989
rect 599 82975 649 82977
rect 42 82933 59 82967
rect 67 82925 69 82975
rect 160 82967 246 82975
rect 522 82967 608 82975
rect 76 82933 110 82967
rect 127 82933 144 82967
rect 152 82933 161 82967
rect 162 82965 195 82967
rect 224 82965 244 82967
rect 162 82933 244 82965
rect 524 82965 548 82967
rect 573 82965 582 82967
rect 586 82965 606 82967
rect 160 82925 246 82933
rect 186 82909 220 82925
rect 182 82895 224 82896
rect 160 82889 182 82895
rect 224 82889 246 82895
rect 186 82854 220 82888
rect 223 82854 257 82888
rect 120 82841 170 82843
rect 76 82837 130 82841
rect 110 82832 130 82837
rect 60 82807 67 82817
rect 76 82807 77 82827
rect 96 82798 99 82832
rect 109 82807 110 82827
rect 119 82807 126 82817
rect 76 82791 92 82797
rect 94 82791 110 82797
rect 170 82791 172 82841
rect 186 82775 190 82809
rect 216 82775 220 82809
rect 288 82775 292 82963
rect 476 82895 480 82963
rect 524 82933 606 82965
rect 607 82933 616 82967
rect 522 82925 608 82933
rect 649 82925 651 82975
rect 548 82909 582 82925
rect 522 82890 548 82895
rect 522 82889 582 82890
rect 586 82889 608 82895
rect 295 82854 300 82888
rect 324 82854 329 82888
rect 544 82886 582 82889
rect 378 82849 450 82857
rect 428 82819 430 82835
rect 400 82811 430 82819
rect 476 82817 480 82885
rect 544 82856 552 82886
rect 578 82856 582 82886
rect 544 82847 548 82856
rect 400 82807 436 82811
rect 400 82777 408 82807
rect 420 82777 436 82807
rect 544 82809 548 82817
rect 12 82738 62 82740
rect 28 82729 59 82737
rect 62 82729 64 82738
rect 28 82721 64 82729
rect 127 82729 158 82737
rect 127 82722 182 82729
rect 215 82727 224 82755
rect 127 82721 161 82722
rect 59 82705 64 82721
rect 158 82705 161 82721
rect 28 82697 64 82705
rect 127 82704 161 82705
rect 127 82697 182 82704
rect 62 82688 64 82697
rect 213 82689 224 82727
rect 282 82717 292 82775
rect 296 82769 368 82777
rect 319 82739 346 82750
rect 318 82726 324 82739
rect 346 82726 348 82739
rect 428 82730 430 82777
rect 443 82767 450 82769
rect 476 82737 480 82805
rect 544 82775 552 82809
rect 578 82775 582 82809
rect 481 82743 517 82771
rect 481 82737 495 82743
rect 367 82726 380 82730
rect 251 82683 263 82717
rect 273 82683 293 82717
rect 295 82702 324 82726
rect 303 82692 316 82702
rect 318 82686 324 82702
rect 333 82702 380 82726
rect 333 82692 353 82702
rect 367 82696 380 82702
rect 396 82696 408 82730
rect 420 82696 436 82730
rect 120 82635 170 82637
rect 76 82629 92 82635
rect 94 82629 110 82635
rect 76 82619 99 82628
rect 60 82609 67 82619
rect 76 82599 77 82619
rect 96 82594 99 82619
rect 109 82599 110 82619
rect 119 82609 126 82619
rect 76 82585 110 82589
rect 170 82585 172 82635
rect 186 82617 190 82651
rect 216 82617 220 82651
rect 186 82540 220 82574
rect 282 82571 292 82683
rect 318 82676 335 82686
rect 318 82607 324 82676
rect 346 82607 348 82692
rect 428 82649 430 82696
rect 476 82659 480 82727
rect 485 82709 495 82737
rect 505 82737 519 82743
rect 544 82737 555 82775
rect 505 82709 525 82737
rect 544 82709 553 82737
rect 544 82689 548 82709
rect 579 82668 582 82758
rect 612 82740 624 82741
rect 599 82738 649 82740
rect 612 82737 624 82738
rect 610 82730 632 82737
rect 607 82729 632 82730
rect 586 82722 644 82729
rect 607 82721 644 82722
rect 607 82705 610 82721
rect 616 82705 644 82721
rect 607 82704 644 82705
rect 586 82697 644 82704
rect 607 82696 610 82697
rect 612 82689 632 82697
rect 612 82685 624 82689
rect 649 82688 651 82738
rect 544 82651 548 82659
rect 400 82619 408 82649
rect 420 82619 436 82649
rect 400 82615 436 82619
rect 400 82607 430 82615
rect 428 82591 430 82607
rect 476 82579 480 82647
rect 544 82617 552 82651
rect 578 82617 582 82651
rect 544 82609 548 82617
rect 544 82579 586 82580
rect 288 82539 292 82571
rect 296 82569 368 82577
rect 378 82569 450 82577
rect 544 82572 548 82579
rect 439 82541 444 82569
rect 120 82525 170 82527
rect 76 82521 130 82525
rect 110 82516 130 82521
rect 60 82491 67 82501
rect 76 82491 77 82511
rect 96 82482 99 82516
rect 109 82491 110 82511
rect 119 82491 126 82501
rect 76 82475 92 82481
rect 94 82475 110 82481
rect 170 82475 172 82525
rect 186 82459 190 82493
rect 216 82459 220 82493
rect 213 82427 224 82459
rect 282 82455 292 82539
rect 296 82533 368 82541
rect 378 82533 450 82541
rect 468 82538 473 82572
rect 428 82503 430 82519
rect 251 82427 292 82455
rect 318 82434 324 82503
rect 12 82422 62 82424
rect 28 82413 59 82421
rect 62 82413 64 82422
rect 251 82421 263 82427
rect 28 82405 64 82413
rect 127 82413 158 82421
rect 127 82406 182 82413
rect 127 82405 161 82406
rect 59 82389 64 82405
rect 158 82389 161 82405
rect 253 82393 263 82421
rect 273 82393 293 82427
rect 318 82424 335 82434
rect 303 82408 316 82418
rect 318 82408 324 82424
rect 346 82418 348 82503
rect 400 82495 430 82503
rect 476 82501 480 82569
rect 511 82538 582 82572
rect 544 82531 548 82538
rect 400 82491 436 82495
rect 400 82461 408 82491
rect 420 82461 436 82491
rect 544 82493 548 82501
rect 28 82381 64 82389
rect 127 82388 161 82389
rect 127 82381 182 82388
rect 62 82372 64 82381
rect 282 82335 292 82393
rect 295 82384 324 82408
rect 333 82408 353 82418
rect 428 82414 430 82461
rect 476 82421 480 82489
rect 544 82459 552 82493
rect 578 82459 582 82493
rect 544 82451 548 82459
rect 367 82408 380 82414
rect 333 82384 380 82408
rect 318 82371 324 82384
rect 346 82371 348 82384
rect 367 82380 380 82384
rect 396 82380 408 82414
rect 420 82380 436 82414
rect 544 82411 553 82439
rect 319 82360 346 82371
rect 120 82319 170 82321
rect 76 82313 92 82319
rect 94 82313 110 82319
rect 76 82303 99 82312
rect 60 82293 67 82303
rect 76 82283 77 82303
rect 96 82278 99 82303
rect 109 82283 110 82303
rect 119 82293 126 82303
rect 76 82269 110 82273
rect 170 82269 172 82319
rect 186 82301 190 82335
rect 216 82301 220 82335
rect 182 82263 224 82264
rect 186 82239 220 82256
rect 223 82239 257 82256
rect 182 82222 257 82239
rect 182 82221 224 82222
rect 160 82215 246 82221
rect 288 82215 292 82335
rect 296 82333 368 82341
rect 428 82333 430 82380
rect 476 82343 480 82411
rect 485 82367 495 82401
rect 505 82373 525 82401
rect 505 82367 519 82373
rect 544 82367 555 82411
rect 485 82343 492 82367
rect 579 82352 582 82442
rect 612 82424 624 82425
rect 599 82422 649 82424
rect 612 82421 624 82422
rect 610 82414 632 82421
rect 607 82413 632 82414
rect 586 82406 644 82413
rect 607 82405 644 82406
rect 607 82389 610 82405
rect 616 82389 644 82405
rect 607 82388 644 82389
rect 586 82381 644 82388
rect 607 82380 610 82381
rect 612 82373 632 82381
rect 612 82369 624 82373
rect 649 82372 651 82422
rect 544 82335 548 82343
rect 400 82303 408 82333
rect 420 82303 436 82333
rect 400 82299 436 82303
rect 400 82291 430 82299
rect 428 82275 430 82291
rect 476 82263 480 82331
rect 544 82301 552 82335
rect 578 82301 582 82335
rect 544 82293 548 82301
rect 295 82222 300 82256
rect 324 82222 329 82256
rect 378 82253 450 82261
rect 544 82258 548 82263
rect 544 82254 582 82258
rect 544 82239 552 82254
rect 578 82239 582 82254
rect 544 82221 586 82239
rect 522 82215 608 82221
rect 182 82199 224 82215
rect 544 82199 586 82215
rect 17 82185 67 82187
rect 119 82185 169 82187
rect 186 82185 220 82199
rect 548 82185 582 82199
rect 599 82185 649 82187
rect 42 82143 59 82177
rect 67 82135 69 82185
rect 160 82177 246 82185
rect 522 82177 608 82185
rect 76 82143 110 82177
rect 127 82143 144 82177
rect 152 82143 161 82177
rect 162 82175 195 82177
rect 224 82175 244 82177
rect 162 82143 244 82175
rect 524 82175 548 82177
rect 573 82175 582 82177
rect 586 82175 606 82177
rect 160 82135 246 82143
rect 186 82119 220 82135
rect 182 82105 224 82106
rect 160 82099 182 82105
rect 224 82099 246 82105
rect 186 82064 220 82098
rect 223 82064 257 82098
rect 120 82051 170 82053
rect 76 82047 130 82051
rect 110 82042 130 82047
rect 60 82017 67 82027
rect 76 82017 77 82037
rect 96 82008 99 82042
rect 109 82017 110 82037
rect 119 82017 126 82027
rect 76 82001 92 82007
rect 94 82001 110 82007
rect 170 82001 172 82051
rect 186 81985 190 82019
rect 216 81985 220 82019
rect 288 81985 292 82173
rect 476 82105 480 82173
rect 524 82143 606 82175
rect 607 82143 616 82177
rect 522 82135 608 82143
rect 649 82135 651 82185
rect 548 82119 582 82135
rect 522 82100 548 82105
rect 522 82099 582 82100
rect 586 82099 608 82105
rect 295 82064 300 82098
rect 324 82064 329 82098
rect 544 82096 582 82099
rect 378 82059 450 82067
rect 428 82029 430 82045
rect 400 82021 430 82029
rect 476 82027 480 82095
rect 544 82066 552 82096
rect 578 82066 582 82096
rect 544 82057 548 82066
rect 400 82017 436 82021
rect 400 81987 408 82017
rect 420 81987 436 82017
rect 544 82019 548 82027
rect 12 81948 62 81950
rect 28 81939 59 81947
rect 62 81939 64 81948
rect 28 81931 64 81939
rect 127 81939 158 81947
rect 127 81932 182 81939
rect 215 81937 224 81965
rect 127 81931 161 81932
rect 59 81915 64 81931
rect 158 81915 161 81931
rect 28 81907 64 81915
rect 127 81914 161 81915
rect 127 81907 182 81914
rect 62 81898 64 81907
rect 213 81899 224 81937
rect 282 81927 292 81985
rect 296 81979 368 81987
rect 319 81949 346 81960
rect 318 81936 324 81949
rect 346 81936 348 81949
rect 428 81940 430 81987
rect 443 81977 450 81979
rect 476 81947 480 82015
rect 544 81985 552 82019
rect 578 81985 582 82019
rect 481 81953 517 81981
rect 481 81947 495 81953
rect 367 81936 380 81940
rect 251 81893 263 81927
rect 273 81893 293 81927
rect 295 81912 324 81936
rect 303 81902 316 81912
rect 318 81896 324 81912
rect 333 81912 380 81936
rect 333 81902 353 81912
rect 367 81906 380 81912
rect 396 81906 408 81940
rect 420 81906 436 81940
rect 120 81845 170 81847
rect 76 81839 92 81845
rect 94 81839 110 81845
rect 76 81829 99 81838
rect 60 81819 67 81829
rect 76 81809 77 81829
rect 96 81804 99 81829
rect 109 81809 110 81829
rect 119 81819 126 81829
rect 76 81795 110 81799
rect 170 81795 172 81845
rect 186 81827 190 81861
rect 216 81827 220 81861
rect 186 81750 220 81784
rect 282 81781 292 81893
rect 318 81886 335 81896
rect 318 81817 324 81886
rect 346 81817 348 81902
rect 428 81859 430 81906
rect 476 81869 480 81937
rect 485 81919 495 81947
rect 505 81947 519 81953
rect 544 81947 555 81985
rect 505 81919 525 81947
rect 544 81919 553 81947
rect 544 81899 548 81919
rect 579 81878 582 81968
rect 612 81950 624 81951
rect 599 81948 649 81950
rect 612 81947 624 81948
rect 610 81940 632 81947
rect 607 81939 632 81940
rect 586 81932 644 81939
rect 607 81931 644 81932
rect 607 81915 610 81931
rect 616 81915 644 81931
rect 607 81914 644 81915
rect 586 81907 644 81914
rect 607 81906 610 81907
rect 612 81899 632 81907
rect 612 81895 624 81899
rect 649 81898 651 81948
rect 544 81861 548 81869
rect 400 81829 408 81859
rect 420 81829 436 81859
rect 400 81825 436 81829
rect 400 81817 430 81825
rect 428 81801 430 81817
rect 476 81789 480 81857
rect 544 81827 552 81861
rect 578 81827 582 81861
rect 544 81819 548 81827
rect 544 81789 586 81790
rect 288 81749 292 81781
rect 296 81779 368 81787
rect 378 81779 450 81787
rect 544 81782 548 81789
rect 439 81751 444 81779
rect 120 81735 170 81737
rect 76 81731 130 81735
rect 110 81726 130 81731
rect 60 81701 67 81711
rect 76 81701 77 81721
rect 96 81692 99 81726
rect 109 81701 110 81721
rect 119 81701 126 81711
rect 76 81685 92 81691
rect 94 81685 110 81691
rect 170 81685 172 81735
rect 186 81669 190 81703
rect 216 81669 220 81703
rect 213 81637 224 81669
rect 282 81665 292 81749
rect 296 81743 368 81751
rect 378 81743 450 81751
rect 468 81748 473 81782
rect 428 81713 430 81729
rect 251 81637 292 81665
rect 318 81644 324 81713
rect 12 81632 62 81634
rect 28 81623 59 81631
rect 62 81623 64 81632
rect 251 81631 263 81637
rect 28 81615 64 81623
rect 127 81623 158 81631
rect 127 81616 182 81623
rect 127 81615 161 81616
rect 59 81599 64 81615
rect 158 81599 161 81615
rect 253 81603 263 81631
rect 273 81603 293 81637
rect 318 81634 335 81644
rect 303 81618 316 81628
rect 318 81618 324 81634
rect 346 81628 348 81713
rect 400 81705 430 81713
rect 476 81711 480 81779
rect 511 81748 582 81782
rect 544 81741 548 81748
rect 400 81701 436 81705
rect 400 81671 408 81701
rect 420 81671 436 81701
rect 544 81703 548 81711
rect 28 81591 64 81599
rect 127 81598 161 81599
rect 127 81591 182 81598
rect 62 81582 64 81591
rect 282 81545 292 81603
rect 295 81594 324 81618
rect 333 81618 353 81628
rect 428 81624 430 81671
rect 476 81631 480 81699
rect 544 81669 552 81703
rect 578 81669 582 81703
rect 544 81661 548 81669
rect 367 81618 380 81624
rect 333 81594 380 81618
rect 318 81581 324 81594
rect 346 81581 348 81594
rect 367 81590 380 81594
rect 396 81590 408 81624
rect 420 81590 436 81624
rect 544 81621 553 81649
rect 319 81570 346 81581
rect 120 81529 170 81531
rect 76 81523 92 81529
rect 94 81523 110 81529
rect 76 81513 99 81522
rect 60 81503 67 81513
rect 76 81493 77 81513
rect 96 81488 99 81513
rect 109 81493 110 81513
rect 119 81503 126 81513
rect 76 81479 110 81483
rect 170 81479 172 81529
rect 186 81511 190 81545
rect 216 81511 220 81545
rect 182 81473 224 81474
rect 186 81449 220 81466
rect 223 81449 257 81466
rect 182 81432 257 81449
rect 182 81431 224 81432
rect 160 81425 246 81431
rect 288 81425 292 81545
rect 296 81543 368 81551
rect 428 81543 430 81590
rect 476 81553 480 81621
rect 485 81577 495 81611
rect 505 81583 525 81611
rect 505 81577 519 81583
rect 544 81577 555 81621
rect 485 81553 492 81577
rect 579 81562 582 81652
rect 612 81634 624 81635
rect 599 81632 649 81634
rect 612 81631 624 81632
rect 610 81624 632 81631
rect 607 81623 632 81624
rect 586 81616 644 81623
rect 607 81615 644 81616
rect 607 81599 610 81615
rect 616 81599 644 81615
rect 607 81598 644 81599
rect 586 81591 644 81598
rect 607 81590 610 81591
rect 612 81583 632 81591
rect 612 81579 624 81583
rect 649 81582 651 81632
rect 544 81545 548 81553
rect 400 81513 408 81543
rect 420 81513 436 81543
rect 400 81509 436 81513
rect 400 81501 430 81509
rect 428 81485 430 81501
rect 476 81473 480 81541
rect 544 81511 552 81545
rect 578 81511 582 81545
rect 544 81503 548 81511
rect 295 81432 300 81466
rect 324 81432 329 81466
rect 378 81463 450 81471
rect 544 81468 548 81473
rect 544 81464 582 81468
rect 544 81449 552 81464
rect 578 81449 582 81464
rect 544 81431 586 81449
rect 522 81425 608 81431
rect 182 81409 224 81425
rect 544 81409 586 81425
rect 17 81395 67 81397
rect 119 81395 169 81397
rect 186 81395 220 81409
rect 548 81395 582 81409
rect 599 81395 649 81397
rect 42 81353 59 81387
rect 67 81345 69 81395
rect 160 81387 246 81395
rect 522 81387 608 81395
rect 76 81353 110 81387
rect 127 81353 144 81387
rect 152 81353 161 81387
rect 162 81385 195 81387
rect 224 81385 244 81387
rect 162 81353 244 81385
rect 524 81385 548 81387
rect 573 81385 582 81387
rect 586 81385 606 81387
rect 160 81345 246 81353
rect 186 81329 220 81345
rect 182 81315 224 81316
rect 160 81309 182 81315
rect 224 81309 246 81315
rect 186 81274 220 81308
rect 223 81274 257 81308
rect 120 81261 170 81263
rect 76 81257 130 81261
rect 110 81252 130 81257
rect 60 81227 67 81237
rect 76 81227 77 81247
rect 96 81218 99 81252
rect 109 81227 110 81247
rect 119 81227 126 81237
rect 76 81211 92 81217
rect 94 81211 110 81217
rect 170 81211 172 81261
rect 186 81195 190 81229
rect 216 81195 220 81229
rect 288 81195 292 81383
rect 476 81315 480 81383
rect 524 81353 606 81385
rect 607 81353 616 81387
rect 522 81345 608 81353
rect 649 81345 651 81395
rect 548 81329 582 81345
rect 522 81310 548 81315
rect 522 81309 582 81310
rect 586 81309 608 81315
rect 295 81274 300 81308
rect 324 81274 329 81308
rect 544 81306 582 81309
rect 378 81269 450 81277
rect 428 81239 430 81255
rect 400 81231 430 81239
rect 476 81237 480 81305
rect 544 81276 552 81306
rect 578 81276 582 81306
rect 544 81267 548 81276
rect 400 81227 436 81231
rect 400 81197 408 81227
rect 420 81197 436 81227
rect 544 81229 548 81237
rect 12 81158 62 81160
rect 28 81149 59 81157
rect 62 81149 64 81158
rect 28 81141 64 81149
rect 127 81149 158 81157
rect 127 81142 182 81149
rect 215 81147 224 81175
rect 127 81141 161 81142
rect 59 81125 64 81141
rect 158 81125 161 81141
rect 28 81117 64 81125
rect 127 81124 161 81125
rect 127 81117 182 81124
rect 62 81108 64 81117
rect 213 81109 224 81147
rect 282 81137 292 81195
rect 296 81189 368 81197
rect 319 81159 346 81170
rect 318 81146 324 81159
rect 346 81146 348 81159
rect 428 81150 430 81197
rect 443 81187 450 81189
rect 476 81157 480 81225
rect 544 81195 552 81229
rect 578 81195 582 81229
rect 481 81163 517 81191
rect 481 81157 495 81163
rect 367 81146 380 81150
rect 251 81103 263 81137
rect 273 81103 293 81137
rect 295 81122 324 81146
rect 303 81112 316 81122
rect 318 81106 324 81122
rect 333 81122 380 81146
rect 333 81112 353 81122
rect 367 81116 380 81122
rect 396 81116 408 81150
rect 420 81116 436 81150
rect 120 81055 170 81057
rect 76 81049 92 81055
rect 94 81049 110 81055
rect 76 81039 99 81048
rect 60 81029 67 81039
rect 76 81019 77 81039
rect 96 81014 99 81039
rect 109 81019 110 81039
rect 119 81029 126 81039
rect 76 81005 110 81009
rect 170 81005 172 81055
rect 186 81037 190 81071
rect 216 81037 220 81071
rect 186 80960 220 80994
rect 282 80991 292 81103
rect 318 81096 335 81106
rect 318 81027 324 81096
rect 346 81027 348 81112
rect 428 81069 430 81116
rect 476 81079 480 81147
rect 485 81129 495 81157
rect 505 81157 519 81163
rect 544 81157 555 81195
rect 505 81129 525 81157
rect 544 81129 553 81157
rect 544 81109 548 81129
rect 579 81088 582 81178
rect 612 81160 624 81161
rect 599 81158 649 81160
rect 612 81157 624 81158
rect 610 81150 632 81157
rect 607 81149 632 81150
rect 586 81142 644 81149
rect 607 81141 644 81142
rect 607 81125 610 81141
rect 616 81125 644 81141
rect 607 81124 644 81125
rect 586 81117 644 81124
rect 607 81116 610 81117
rect 612 81109 632 81117
rect 612 81105 624 81109
rect 649 81108 651 81158
rect 544 81071 548 81079
rect 400 81039 408 81069
rect 420 81039 436 81069
rect 400 81035 436 81039
rect 400 81027 430 81035
rect 428 81011 430 81027
rect 476 80999 480 81067
rect 544 81037 552 81071
rect 578 81037 582 81071
rect 544 81029 548 81037
rect 544 80999 586 81000
rect 288 80959 292 80991
rect 296 80989 368 80997
rect 378 80989 450 80997
rect 544 80992 548 80999
rect 439 80961 444 80989
rect 120 80945 170 80947
rect 76 80941 130 80945
rect 110 80936 130 80941
rect 60 80911 67 80921
rect 76 80911 77 80931
rect 96 80902 99 80936
rect 109 80911 110 80931
rect 119 80911 126 80921
rect 76 80895 92 80901
rect 94 80895 110 80901
rect 170 80895 172 80945
rect 186 80879 190 80913
rect 216 80879 220 80913
rect 213 80847 224 80879
rect 282 80875 292 80959
rect 296 80953 368 80961
rect 378 80953 450 80961
rect 468 80958 473 80992
rect 428 80923 430 80939
rect 251 80847 292 80875
rect 318 80854 324 80923
rect 12 80842 62 80844
rect 28 80833 59 80841
rect 62 80833 64 80842
rect 251 80841 263 80847
rect 28 80825 64 80833
rect 127 80833 158 80841
rect 127 80826 182 80833
rect 127 80825 161 80826
rect 59 80809 64 80825
rect 158 80809 161 80825
rect 253 80813 263 80841
rect 273 80813 293 80847
rect 318 80844 335 80854
rect 303 80828 316 80838
rect 318 80828 324 80844
rect 346 80838 348 80923
rect 400 80915 430 80923
rect 476 80921 480 80989
rect 511 80958 582 80992
rect 544 80951 548 80958
rect 400 80911 436 80915
rect 400 80881 408 80911
rect 420 80881 436 80911
rect 544 80913 548 80921
rect 28 80801 64 80809
rect 127 80808 161 80809
rect 127 80801 182 80808
rect 62 80792 64 80801
rect 282 80755 292 80813
rect 295 80804 324 80828
rect 333 80828 353 80838
rect 428 80834 430 80881
rect 476 80841 480 80909
rect 544 80879 552 80913
rect 578 80879 582 80913
rect 544 80871 548 80879
rect 367 80828 380 80834
rect 333 80804 380 80828
rect 318 80791 324 80804
rect 346 80791 348 80804
rect 367 80800 380 80804
rect 396 80800 408 80834
rect 420 80800 436 80834
rect 544 80831 553 80859
rect 319 80780 346 80791
rect 120 80739 170 80741
rect 76 80733 92 80739
rect 94 80733 110 80739
rect 76 80723 99 80732
rect 60 80713 67 80723
rect 76 80703 77 80723
rect 96 80698 99 80723
rect 109 80703 110 80723
rect 119 80713 126 80723
rect 76 80689 110 80693
rect 170 80689 172 80739
rect 186 80721 190 80755
rect 216 80721 220 80755
rect 182 80683 224 80684
rect 186 80659 220 80676
rect 223 80659 257 80676
rect 182 80642 257 80659
rect 182 80641 224 80642
rect 160 80635 246 80641
rect 288 80635 292 80755
rect 296 80753 368 80761
rect 428 80753 430 80800
rect 476 80763 480 80831
rect 485 80787 495 80821
rect 505 80793 525 80821
rect 505 80787 519 80793
rect 544 80787 555 80831
rect 485 80763 492 80787
rect 579 80772 582 80862
rect 612 80844 624 80845
rect 599 80842 649 80844
rect 612 80841 624 80842
rect 610 80834 632 80841
rect 607 80833 632 80834
rect 586 80826 644 80833
rect 607 80825 644 80826
rect 607 80809 610 80825
rect 616 80809 644 80825
rect 607 80808 644 80809
rect 586 80801 644 80808
rect 607 80800 610 80801
rect 612 80793 632 80801
rect 612 80789 624 80793
rect 649 80792 651 80842
rect 544 80755 548 80763
rect 400 80723 408 80753
rect 420 80723 436 80753
rect 400 80719 436 80723
rect 400 80711 430 80719
rect 428 80695 430 80711
rect 476 80683 480 80751
rect 544 80721 552 80755
rect 578 80721 582 80755
rect 544 80713 548 80721
rect 295 80642 300 80676
rect 324 80642 329 80676
rect 378 80673 450 80681
rect 544 80678 548 80683
rect 544 80674 582 80678
rect 544 80659 552 80674
rect 578 80659 582 80674
rect 544 80641 586 80659
rect 522 80635 608 80641
rect 182 80619 224 80635
rect 544 80619 586 80635
rect 17 80605 67 80607
rect 119 80605 169 80607
rect 186 80605 220 80619
rect 548 80605 582 80619
rect 599 80605 649 80607
rect 42 80563 59 80597
rect 67 80555 69 80605
rect 160 80597 246 80605
rect 522 80597 608 80605
rect 76 80563 110 80597
rect 127 80563 144 80597
rect 152 80563 161 80597
rect 162 80595 195 80597
rect 224 80595 244 80597
rect 162 80563 244 80595
rect 524 80595 548 80597
rect 573 80595 582 80597
rect 586 80595 606 80597
rect 160 80555 246 80563
rect 186 80539 220 80555
rect 182 80525 224 80526
rect 160 80519 182 80525
rect 224 80519 246 80525
rect 186 80484 220 80518
rect 223 80484 257 80518
rect 120 80471 170 80473
rect 76 80467 130 80471
rect 110 80462 130 80467
rect 60 80437 67 80447
rect 76 80437 77 80457
rect 96 80428 99 80462
rect 109 80437 110 80457
rect 119 80437 126 80447
rect 76 80421 92 80427
rect 94 80421 110 80427
rect 170 80421 172 80471
rect 186 80405 190 80439
rect 216 80405 220 80439
rect 288 80405 292 80593
rect 476 80525 480 80593
rect 524 80563 606 80595
rect 607 80563 616 80597
rect 522 80555 608 80563
rect 649 80555 651 80605
rect 548 80539 582 80555
rect 522 80520 548 80525
rect 522 80519 582 80520
rect 586 80519 608 80525
rect 295 80484 300 80518
rect 324 80484 329 80518
rect 544 80516 582 80519
rect 378 80479 450 80487
rect 428 80449 430 80465
rect 400 80441 430 80449
rect 476 80447 480 80515
rect 544 80486 552 80516
rect 578 80486 582 80516
rect 544 80477 548 80486
rect 400 80437 436 80441
rect 400 80407 408 80437
rect 420 80407 436 80437
rect 544 80439 548 80447
rect 12 80368 62 80370
rect 28 80359 59 80367
rect 62 80359 64 80368
rect 28 80351 64 80359
rect 127 80359 158 80367
rect 127 80352 182 80359
rect 215 80357 224 80385
rect 127 80351 161 80352
rect 59 80335 64 80351
rect 158 80335 161 80351
rect 28 80327 64 80335
rect 127 80334 161 80335
rect 127 80327 182 80334
rect 62 80318 64 80327
rect 213 80319 224 80357
rect 282 80347 292 80405
rect 296 80399 368 80407
rect 319 80369 346 80380
rect 318 80356 324 80369
rect 346 80356 348 80369
rect 428 80360 430 80407
rect 443 80397 450 80399
rect 476 80367 480 80435
rect 544 80405 552 80439
rect 578 80405 582 80439
rect 481 80373 517 80401
rect 481 80367 495 80373
rect 367 80356 380 80360
rect 251 80313 263 80347
rect 273 80313 293 80347
rect 295 80332 324 80356
rect 303 80322 316 80332
rect 318 80316 324 80332
rect 333 80332 380 80356
rect 333 80322 353 80332
rect 367 80326 380 80332
rect 396 80326 408 80360
rect 420 80326 436 80360
rect 120 80265 170 80267
rect 76 80259 92 80265
rect 94 80259 110 80265
rect 76 80249 99 80258
rect 60 80239 67 80249
rect 76 80229 77 80249
rect 96 80224 99 80249
rect 109 80229 110 80249
rect 119 80239 126 80249
rect 76 80215 110 80219
rect 170 80215 172 80265
rect 186 80247 190 80281
rect 216 80247 220 80281
rect 186 80170 220 80204
rect 282 80201 292 80313
rect 318 80306 335 80316
rect 318 80237 324 80306
rect 346 80237 348 80322
rect 428 80279 430 80326
rect 476 80289 480 80357
rect 485 80339 495 80367
rect 505 80367 519 80373
rect 544 80367 555 80405
rect 505 80339 525 80367
rect 544 80339 553 80367
rect 544 80319 548 80339
rect 579 80298 582 80388
rect 612 80370 624 80371
rect 599 80368 649 80370
rect 612 80367 624 80368
rect 610 80360 632 80367
rect 607 80359 632 80360
rect 586 80352 644 80359
rect 607 80351 644 80352
rect 607 80335 610 80351
rect 616 80335 644 80351
rect 607 80334 644 80335
rect 586 80327 644 80334
rect 607 80326 610 80327
rect 612 80319 632 80327
rect 612 80315 624 80319
rect 649 80318 651 80368
rect 544 80281 548 80289
rect 400 80249 408 80279
rect 420 80249 436 80279
rect 400 80245 436 80249
rect 400 80237 430 80245
rect 428 80221 430 80237
rect 476 80209 480 80277
rect 544 80247 552 80281
rect 578 80247 582 80281
rect 544 80239 548 80247
rect 544 80209 586 80210
rect 288 80169 292 80201
rect 296 80199 368 80207
rect 378 80199 450 80207
rect 544 80202 548 80209
rect 439 80171 444 80199
rect 120 80155 170 80157
rect 76 80151 130 80155
rect 110 80146 130 80151
rect 60 80121 67 80131
rect 76 80121 77 80141
rect 96 80112 99 80146
rect 109 80121 110 80141
rect 119 80121 126 80131
rect 76 80105 92 80111
rect 94 80105 110 80111
rect 170 80105 172 80155
rect 186 80089 190 80123
rect 216 80089 220 80123
rect 213 80057 224 80089
rect 282 80085 292 80169
rect 296 80163 368 80171
rect 378 80163 450 80171
rect 468 80168 473 80202
rect 428 80133 430 80149
rect 251 80057 292 80085
rect 318 80064 324 80133
rect 12 80052 62 80054
rect 28 80043 59 80051
rect 62 80043 64 80052
rect 251 80051 263 80057
rect 28 80035 64 80043
rect 127 80043 158 80051
rect 127 80036 182 80043
rect 127 80035 161 80036
rect 59 80019 64 80035
rect 158 80019 161 80035
rect 253 80023 263 80051
rect 273 80023 293 80057
rect 318 80054 335 80064
rect 303 80038 316 80048
rect 318 80038 324 80054
rect 346 80048 348 80133
rect 400 80125 430 80133
rect 476 80131 480 80199
rect 511 80168 582 80202
rect 544 80161 548 80168
rect 400 80121 436 80125
rect 400 80091 408 80121
rect 420 80091 436 80121
rect 544 80123 548 80131
rect 28 80011 64 80019
rect 127 80018 161 80019
rect 127 80011 182 80018
rect 62 80002 64 80011
rect 282 79965 292 80023
rect 295 80014 324 80038
rect 333 80038 353 80048
rect 428 80044 430 80091
rect 476 80051 480 80119
rect 544 80089 552 80123
rect 578 80089 582 80123
rect 544 80081 548 80089
rect 367 80038 380 80044
rect 333 80014 380 80038
rect 318 80001 324 80014
rect 346 80001 348 80014
rect 367 80010 380 80014
rect 396 80010 408 80044
rect 420 80010 436 80044
rect 544 80041 553 80069
rect 319 79990 346 80001
rect 120 79949 170 79951
rect 76 79943 92 79949
rect 94 79943 110 79949
rect 76 79933 99 79942
rect 60 79923 67 79933
rect 76 79913 77 79933
rect 96 79908 99 79933
rect 109 79913 110 79933
rect 119 79923 126 79933
rect 76 79899 110 79903
rect 170 79899 172 79949
rect 186 79931 190 79965
rect 216 79931 220 79965
rect 182 79893 224 79894
rect 186 79869 220 79886
rect 223 79869 257 79886
rect 182 79852 257 79869
rect 182 79851 224 79852
rect 160 79845 246 79851
rect 288 79845 292 79965
rect 296 79963 368 79971
rect 428 79963 430 80010
rect 476 79973 480 80041
rect 485 79997 495 80031
rect 505 80003 525 80031
rect 505 79997 519 80003
rect 544 79997 555 80041
rect 485 79973 492 79997
rect 579 79982 582 80072
rect 612 80054 624 80055
rect 599 80052 649 80054
rect 612 80051 624 80052
rect 610 80044 632 80051
rect 607 80043 632 80044
rect 586 80036 644 80043
rect 607 80035 644 80036
rect 607 80019 610 80035
rect 616 80019 644 80035
rect 607 80018 644 80019
rect 586 80011 644 80018
rect 607 80010 610 80011
rect 612 80003 632 80011
rect 612 79999 624 80003
rect 649 80002 651 80052
rect 544 79965 548 79973
rect 400 79933 408 79963
rect 420 79933 436 79963
rect 400 79929 436 79933
rect 400 79921 430 79929
rect 428 79905 430 79921
rect 476 79893 480 79961
rect 544 79931 552 79965
rect 578 79931 582 79965
rect 544 79923 548 79931
rect 295 79852 300 79886
rect 324 79852 329 79886
rect 378 79883 450 79891
rect 544 79888 548 79893
rect 544 79884 582 79888
rect 544 79869 552 79884
rect 578 79869 582 79884
rect 544 79851 586 79869
rect 522 79845 608 79851
rect 182 79829 224 79845
rect 544 79829 586 79845
rect 17 79815 67 79817
rect 119 79815 169 79817
rect 186 79815 220 79829
rect 548 79815 582 79829
rect 599 79815 649 79817
rect 42 79773 59 79807
rect 67 79765 69 79815
rect 160 79807 246 79815
rect 522 79807 608 79815
rect 76 79773 110 79807
rect 127 79773 144 79807
rect 152 79773 161 79807
rect 162 79805 195 79807
rect 224 79805 244 79807
rect 162 79773 244 79805
rect 524 79805 548 79807
rect 573 79805 582 79807
rect 586 79805 606 79807
rect 160 79765 246 79773
rect 186 79749 220 79765
rect 182 79735 224 79736
rect 160 79729 182 79735
rect 224 79729 246 79735
rect 186 79694 220 79728
rect 223 79694 257 79728
rect 120 79681 170 79683
rect 76 79677 130 79681
rect 110 79672 130 79677
rect 60 79647 67 79657
rect 76 79647 77 79667
rect 96 79638 99 79672
rect 109 79647 110 79667
rect 119 79647 126 79657
rect 76 79631 92 79637
rect 94 79631 110 79637
rect 170 79631 172 79681
rect 186 79615 190 79649
rect 216 79615 220 79649
rect 288 79615 292 79803
rect 476 79735 480 79803
rect 524 79773 606 79805
rect 607 79773 616 79807
rect 522 79765 608 79773
rect 649 79765 651 79815
rect 548 79749 582 79765
rect 522 79730 548 79735
rect 522 79729 582 79730
rect 586 79729 608 79735
rect 295 79694 300 79728
rect 324 79694 329 79728
rect 544 79726 582 79729
rect 378 79689 450 79697
rect 428 79659 430 79675
rect 400 79651 430 79659
rect 476 79657 480 79725
rect 544 79696 552 79726
rect 578 79696 582 79726
rect 544 79687 548 79696
rect 400 79647 436 79651
rect 400 79617 408 79647
rect 420 79617 436 79647
rect 544 79649 548 79657
rect 12 79578 62 79580
rect 28 79569 59 79577
rect 62 79569 64 79578
rect 28 79561 64 79569
rect 127 79569 158 79577
rect 127 79562 182 79569
rect 215 79567 224 79595
rect 127 79561 161 79562
rect 59 79545 64 79561
rect 158 79545 161 79561
rect 28 79537 64 79545
rect 127 79544 161 79545
rect 127 79537 182 79544
rect 62 79528 64 79537
rect 213 79529 224 79567
rect 282 79557 292 79615
rect 296 79609 368 79617
rect 319 79579 346 79590
rect 318 79566 324 79579
rect 346 79566 348 79579
rect 428 79570 430 79617
rect 443 79607 450 79609
rect 476 79577 480 79645
rect 544 79615 552 79649
rect 578 79615 582 79649
rect 481 79583 517 79611
rect 481 79577 495 79583
rect 367 79566 380 79570
rect 251 79523 263 79557
rect 273 79523 293 79557
rect 295 79542 324 79566
rect 303 79532 316 79542
rect 318 79526 324 79542
rect 333 79542 380 79566
rect 333 79532 353 79542
rect 367 79536 380 79542
rect 396 79536 408 79570
rect 420 79536 436 79570
rect 120 79475 170 79477
rect 76 79469 92 79475
rect 94 79469 110 79475
rect 76 79459 99 79468
rect 60 79449 67 79459
rect 76 79439 77 79459
rect 96 79434 99 79459
rect 109 79439 110 79459
rect 119 79449 126 79459
rect 76 79425 110 79429
rect 170 79425 172 79475
rect 186 79457 190 79491
rect 216 79457 220 79491
rect 186 79380 220 79414
rect 282 79411 292 79523
rect 318 79516 335 79526
rect 318 79447 324 79516
rect 346 79447 348 79532
rect 428 79489 430 79536
rect 476 79499 480 79567
rect 485 79549 495 79577
rect 505 79577 519 79583
rect 544 79577 555 79615
rect 505 79549 525 79577
rect 544 79549 553 79577
rect 544 79529 548 79549
rect 579 79508 582 79598
rect 612 79580 624 79581
rect 599 79578 649 79580
rect 612 79577 624 79578
rect 610 79570 632 79577
rect 607 79569 632 79570
rect 586 79562 644 79569
rect 607 79561 644 79562
rect 607 79545 610 79561
rect 616 79545 644 79561
rect 607 79544 644 79545
rect 586 79537 644 79544
rect 607 79536 610 79537
rect 612 79529 632 79537
rect 612 79525 624 79529
rect 649 79528 651 79578
rect 544 79491 548 79499
rect 400 79459 408 79489
rect 420 79459 436 79489
rect 400 79455 436 79459
rect 400 79447 430 79455
rect 428 79431 430 79447
rect 476 79419 480 79487
rect 544 79457 552 79491
rect 578 79457 582 79491
rect 544 79449 548 79457
rect 544 79419 586 79420
rect 288 79379 292 79411
rect 296 79409 368 79417
rect 378 79409 450 79417
rect 544 79412 548 79419
rect 439 79381 444 79409
rect 120 79365 170 79367
rect 76 79361 130 79365
rect 110 79356 130 79361
rect 60 79331 67 79341
rect 76 79331 77 79351
rect 96 79322 99 79356
rect 109 79331 110 79351
rect 119 79331 126 79341
rect 76 79315 92 79321
rect 94 79315 110 79321
rect 170 79315 172 79365
rect 186 79299 190 79333
rect 216 79299 220 79333
rect 213 79267 224 79299
rect 282 79295 292 79379
rect 296 79373 368 79381
rect 378 79373 450 79381
rect 468 79378 473 79412
rect 428 79343 430 79359
rect 251 79267 292 79295
rect 318 79274 324 79343
rect 12 79262 62 79264
rect 28 79253 59 79261
rect 62 79253 64 79262
rect 251 79261 263 79267
rect 28 79245 64 79253
rect 127 79253 158 79261
rect 127 79246 182 79253
rect 127 79245 161 79246
rect 59 79229 64 79245
rect 158 79229 161 79245
rect 253 79233 263 79261
rect 273 79233 293 79267
rect 318 79264 335 79274
rect 303 79248 316 79258
rect 318 79248 324 79264
rect 346 79258 348 79343
rect 400 79335 430 79343
rect 476 79341 480 79409
rect 511 79378 582 79412
rect 544 79371 548 79378
rect 400 79331 436 79335
rect 400 79301 408 79331
rect 420 79301 436 79331
rect 544 79333 548 79341
rect 28 79221 64 79229
rect 127 79228 161 79229
rect 127 79221 182 79228
rect 62 79212 64 79221
rect 282 79175 292 79233
rect 295 79224 324 79248
rect 333 79248 353 79258
rect 428 79254 430 79301
rect 476 79261 480 79329
rect 544 79299 552 79333
rect 578 79299 582 79333
rect 544 79291 548 79299
rect 367 79248 380 79254
rect 333 79224 380 79248
rect 318 79211 324 79224
rect 346 79211 348 79224
rect 367 79220 380 79224
rect 396 79220 408 79254
rect 420 79220 436 79254
rect 544 79251 553 79279
rect 319 79200 346 79211
rect 120 79159 170 79161
rect 76 79153 92 79159
rect 94 79153 110 79159
rect 76 79143 99 79152
rect 60 79133 67 79143
rect 76 79123 77 79143
rect 96 79118 99 79143
rect 109 79123 110 79143
rect 119 79133 126 79143
rect 76 79109 110 79113
rect 170 79109 172 79159
rect 186 79141 190 79175
rect 216 79141 220 79175
rect 182 79103 224 79104
rect 186 79079 220 79096
rect 223 79079 257 79096
rect 182 79062 257 79079
rect 182 79061 224 79062
rect 160 79055 246 79061
rect 288 79055 292 79175
rect 296 79173 368 79181
rect 428 79173 430 79220
rect 476 79183 480 79251
rect 485 79207 495 79241
rect 505 79213 525 79241
rect 505 79207 519 79213
rect 544 79207 555 79251
rect 485 79183 492 79207
rect 579 79192 582 79282
rect 612 79264 624 79265
rect 599 79262 649 79264
rect 612 79261 624 79262
rect 610 79254 632 79261
rect 607 79253 632 79254
rect 586 79246 644 79253
rect 607 79245 644 79246
rect 607 79229 610 79245
rect 616 79229 644 79245
rect 607 79228 644 79229
rect 586 79221 644 79228
rect 607 79220 610 79221
rect 612 79213 632 79221
rect 612 79209 624 79213
rect 649 79212 651 79262
rect 544 79175 548 79183
rect 400 79143 408 79173
rect 420 79143 436 79173
rect 400 79139 436 79143
rect 400 79131 430 79139
rect 428 79115 430 79131
rect 476 79103 480 79171
rect 544 79141 552 79175
rect 578 79141 582 79175
rect 544 79133 548 79141
rect 295 79062 300 79096
rect 324 79062 329 79096
rect 378 79093 450 79101
rect 544 79098 548 79103
rect 544 79094 582 79098
rect 544 79079 552 79094
rect 578 79079 582 79094
rect 544 79061 586 79079
rect 522 79055 608 79061
rect 182 79039 224 79055
rect 544 79039 586 79055
rect 17 79025 67 79027
rect 119 79025 169 79027
rect 186 79025 220 79039
rect 548 79025 582 79039
rect 599 79025 649 79027
rect 42 78983 59 79017
rect 67 78975 69 79025
rect 160 79017 246 79025
rect 522 79017 608 79025
rect 76 78983 110 79017
rect 127 78983 144 79017
rect 152 78983 161 79017
rect 162 79015 195 79017
rect 224 79015 244 79017
rect 162 78983 244 79015
rect 524 79015 548 79017
rect 573 79015 582 79017
rect 586 79015 606 79017
rect 160 78975 246 78983
rect 186 78959 220 78975
rect 182 78945 224 78946
rect 160 78939 182 78945
rect 224 78939 246 78945
rect 186 78904 220 78938
rect 223 78904 257 78938
rect 120 78891 170 78893
rect 76 78887 130 78891
rect 110 78882 130 78887
rect 60 78857 67 78867
rect 76 78857 77 78877
rect 96 78848 99 78882
rect 109 78857 110 78877
rect 119 78857 126 78867
rect 76 78841 92 78847
rect 94 78841 110 78847
rect 170 78841 172 78891
rect 186 78825 190 78859
rect 216 78825 220 78859
rect 288 78825 292 79013
rect 476 78945 480 79013
rect 524 78983 606 79015
rect 607 78983 616 79017
rect 522 78975 608 78983
rect 649 78975 651 79025
rect 548 78959 582 78975
rect 522 78940 548 78945
rect 522 78939 582 78940
rect 586 78939 608 78945
rect 295 78904 300 78938
rect 324 78904 329 78938
rect 544 78936 582 78939
rect 378 78899 450 78907
rect 428 78869 430 78885
rect 400 78861 430 78869
rect 476 78867 480 78935
rect 544 78906 552 78936
rect 578 78906 582 78936
rect 544 78897 548 78906
rect 400 78857 436 78861
rect 400 78827 408 78857
rect 420 78827 436 78857
rect 544 78859 548 78867
rect 12 78788 62 78790
rect 28 78779 59 78787
rect 62 78779 64 78788
rect 28 78771 64 78779
rect 127 78779 158 78787
rect 127 78772 182 78779
rect 215 78777 224 78805
rect 127 78771 161 78772
rect 59 78755 64 78771
rect 158 78755 161 78771
rect 28 78747 64 78755
rect 127 78754 161 78755
rect 127 78747 182 78754
rect 62 78738 64 78747
rect 213 78739 224 78777
rect 282 78767 292 78825
rect 296 78819 368 78827
rect 319 78789 346 78800
rect 318 78776 324 78789
rect 346 78776 348 78789
rect 428 78780 430 78827
rect 443 78817 450 78819
rect 476 78787 480 78855
rect 544 78825 552 78859
rect 578 78825 582 78859
rect 481 78793 517 78821
rect 481 78787 495 78793
rect 367 78776 380 78780
rect 251 78733 263 78767
rect 273 78733 293 78767
rect 295 78752 324 78776
rect 303 78742 316 78752
rect 318 78736 324 78752
rect 333 78752 380 78776
rect 333 78742 353 78752
rect 367 78746 380 78752
rect 396 78746 408 78780
rect 420 78746 436 78780
rect 120 78685 170 78687
rect 76 78679 92 78685
rect 94 78679 110 78685
rect 76 78669 99 78678
rect 60 78659 67 78669
rect 76 78649 77 78669
rect 96 78644 99 78669
rect 109 78649 110 78669
rect 119 78659 126 78669
rect 76 78635 110 78639
rect 170 78635 172 78685
rect 186 78667 190 78701
rect 216 78667 220 78701
rect 186 78590 220 78624
rect 282 78621 292 78733
rect 318 78726 335 78736
rect 318 78657 324 78726
rect 346 78657 348 78742
rect 428 78699 430 78746
rect 476 78709 480 78777
rect 485 78759 495 78787
rect 505 78787 519 78793
rect 544 78787 555 78825
rect 505 78759 525 78787
rect 544 78759 553 78787
rect 544 78739 548 78759
rect 579 78718 582 78808
rect 612 78790 624 78791
rect 599 78788 649 78790
rect 612 78787 624 78788
rect 610 78780 632 78787
rect 607 78779 632 78780
rect 586 78772 644 78779
rect 607 78771 644 78772
rect 607 78755 610 78771
rect 616 78755 644 78771
rect 607 78754 644 78755
rect 586 78747 644 78754
rect 607 78746 610 78747
rect 612 78739 632 78747
rect 612 78735 624 78739
rect 649 78738 651 78788
rect 544 78701 548 78709
rect 400 78669 408 78699
rect 420 78669 436 78699
rect 400 78665 436 78669
rect 400 78657 430 78665
rect 428 78641 430 78657
rect 476 78629 480 78697
rect 544 78667 552 78701
rect 578 78667 582 78701
rect 544 78659 548 78667
rect 544 78629 586 78630
rect 288 78589 292 78621
rect 296 78619 368 78627
rect 378 78619 450 78627
rect 544 78622 548 78629
rect 439 78591 444 78619
rect 120 78575 170 78577
rect 76 78571 130 78575
rect 110 78566 130 78571
rect 60 78541 67 78551
rect 76 78541 77 78561
rect 96 78532 99 78566
rect 109 78541 110 78561
rect 119 78541 126 78551
rect 76 78525 92 78531
rect 94 78525 110 78531
rect 170 78525 172 78575
rect 186 78509 190 78543
rect 216 78509 220 78543
rect 213 78477 224 78509
rect 282 78505 292 78589
rect 296 78583 368 78591
rect 378 78583 450 78591
rect 468 78588 473 78622
rect 428 78553 430 78569
rect 251 78477 292 78505
rect 318 78484 324 78553
rect 12 78472 62 78474
rect 28 78463 59 78471
rect 62 78463 64 78472
rect 251 78471 263 78477
rect 28 78455 64 78463
rect 127 78463 158 78471
rect 127 78456 182 78463
rect 127 78455 161 78456
rect 59 78439 64 78455
rect 158 78439 161 78455
rect 253 78443 263 78471
rect 273 78443 293 78477
rect 318 78474 335 78484
rect 303 78458 316 78468
rect 318 78458 324 78474
rect 346 78468 348 78553
rect 400 78545 430 78553
rect 476 78551 480 78619
rect 511 78588 582 78622
rect 544 78581 548 78588
rect 400 78541 436 78545
rect 400 78511 408 78541
rect 420 78511 436 78541
rect 544 78543 548 78551
rect 28 78431 64 78439
rect 127 78438 161 78439
rect 127 78431 182 78438
rect 62 78422 64 78431
rect 282 78385 292 78443
rect 295 78434 324 78458
rect 333 78458 353 78468
rect 428 78464 430 78511
rect 476 78471 480 78539
rect 544 78509 552 78543
rect 578 78509 582 78543
rect 544 78501 548 78509
rect 367 78458 380 78464
rect 333 78434 380 78458
rect 318 78421 324 78434
rect 346 78421 348 78434
rect 367 78430 380 78434
rect 396 78430 408 78464
rect 420 78430 436 78464
rect 544 78461 553 78489
rect 319 78410 346 78421
rect 120 78369 170 78371
rect 76 78363 92 78369
rect 94 78363 110 78369
rect 76 78353 99 78362
rect 60 78343 67 78353
rect 76 78333 77 78353
rect 96 78328 99 78353
rect 109 78333 110 78353
rect 119 78343 126 78353
rect 76 78319 110 78323
rect 170 78319 172 78369
rect 186 78351 190 78385
rect 216 78351 220 78385
rect 182 78313 224 78314
rect 186 78289 220 78306
rect 223 78289 257 78306
rect 182 78272 257 78289
rect 182 78271 224 78272
rect 160 78265 246 78271
rect 288 78265 292 78385
rect 296 78383 368 78391
rect 428 78383 430 78430
rect 476 78393 480 78461
rect 485 78417 495 78451
rect 505 78423 525 78451
rect 505 78417 519 78423
rect 544 78417 555 78461
rect 485 78393 492 78417
rect 579 78402 582 78492
rect 612 78474 624 78475
rect 599 78472 649 78474
rect 612 78471 624 78472
rect 610 78464 632 78471
rect 607 78463 632 78464
rect 586 78456 644 78463
rect 607 78455 644 78456
rect 607 78439 610 78455
rect 616 78439 644 78455
rect 607 78438 644 78439
rect 586 78431 644 78438
rect 607 78430 610 78431
rect 612 78423 632 78431
rect 612 78419 624 78423
rect 649 78422 651 78472
rect 544 78385 548 78393
rect 400 78353 408 78383
rect 420 78353 436 78383
rect 400 78349 436 78353
rect 400 78341 430 78349
rect 428 78325 430 78341
rect 476 78313 480 78381
rect 544 78351 552 78385
rect 578 78351 582 78385
rect 544 78343 548 78351
rect 295 78272 300 78306
rect 324 78272 329 78306
rect 378 78303 450 78311
rect 544 78308 548 78313
rect 544 78304 582 78308
rect 544 78289 552 78304
rect 578 78289 582 78304
rect 544 78271 586 78289
rect 522 78265 608 78271
rect 182 78249 224 78265
rect 544 78249 586 78265
rect 17 78235 67 78237
rect 119 78235 169 78237
rect 186 78235 220 78249
rect 548 78235 582 78249
rect 599 78235 649 78237
rect 42 78193 59 78227
rect 67 78185 69 78235
rect 160 78227 246 78235
rect 522 78227 608 78235
rect 76 78193 110 78227
rect 127 78193 144 78227
rect 152 78193 161 78227
rect 162 78225 195 78227
rect 224 78225 244 78227
rect 162 78193 244 78225
rect 524 78225 548 78227
rect 573 78225 582 78227
rect 586 78225 606 78227
rect 160 78185 246 78193
rect 186 78169 220 78185
rect 182 78155 224 78156
rect 160 78149 182 78155
rect 224 78149 246 78155
rect 186 78114 220 78148
rect 223 78114 257 78148
rect 120 78101 170 78103
rect 76 78097 130 78101
rect 110 78092 130 78097
rect 60 78067 67 78077
rect 76 78067 77 78087
rect 96 78058 99 78092
rect 109 78067 110 78087
rect 119 78067 126 78077
rect 76 78051 92 78057
rect 94 78051 110 78057
rect 170 78051 172 78101
rect 186 78035 190 78069
rect 216 78035 220 78069
rect 288 78035 292 78223
rect 476 78155 480 78223
rect 524 78193 606 78225
rect 607 78193 616 78227
rect 522 78185 608 78193
rect 649 78185 651 78235
rect 548 78169 582 78185
rect 522 78150 548 78155
rect 522 78149 582 78150
rect 586 78149 608 78155
rect 295 78114 300 78148
rect 324 78114 329 78148
rect 544 78146 582 78149
rect 378 78109 450 78117
rect 428 78079 430 78095
rect 400 78071 430 78079
rect 476 78077 480 78145
rect 544 78116 552 78146
rect 578 78116 582 78146
rect 544 78107 548 78116
rect 400 78067 436 78071
rect 400 78037 408 78067
rect 420 78037 436 78067
rect 544 78069 548 78077
rect 12 77998 62 78000
rect 28 77989 59 77997
rect 62 77989 64 77998
rect 28 77981 64 77989
rect 127 77989 158 77997
rect 127 77982 182 77989
rect 215 77987 224 78015
rect 127 77981 161 77982
rect 59 77965 64 77981
rect 158 77965 161 77981
rect 28 77957 64 77965
rect 127 77964 161 77965
rect 127 77957 182 77964
rect 62 77948 64 77957
rect 213 77949 224 77987
rect 282 77977 292 78035
rect 296 78029 368 78037
rect 319 77999 346 78010
rect 318 77986 324 77999
rect 346 77986 348 77999
rect 428 77990 430 78037
rect 443 78027 450 78029
rect 476 77997 480 78065
rect 544 78035 552 78069
rect 578 78035 582 78069
rect 481 78003 517 78031
rect 481 77997 495 78003
rect 367 77986 380 77990
rect 251 77943 263 77977
rect 273 77943 293 77977
rect 295 77962 324 77986
rect 303 77952 316 77962
rect 318 77946 324 77962
rect 333 77962 380 77986
rect 333 77952 353 77962
rect 367 77956 380 77962
rect 396 77956 408 77990
rect 420 77956 436 77990
rect 120 77895 170 77897
rect 76 77889 92 77895
rect 94 77889 110 77895
rect 76 77879 99 77888
rect 60 77869 67 77879
rect 76 77859 77 77879
rect 96 77854 99 77879
rect 109 77859 110 77879
rect 119 77869 126 77879
rect 76 77845 110 77849
rect 170 77845 172 77895
rect 186 77877 190 77911
rect 216 77877 220 77911
rect 186 77800 220 77834
rect 282 77831 292 77943
rect 318 77936 335 77946
rect 318 77867 324 77936
rect 346 77867 348 77952
rect 428 77909 430 77956
rect 476 77919 480 77987
rect 485 77969 495 77997
rect 505 77997 519 78003
rect 544 77997 555 78035
rect 505 77969 525 77997
rect 544 77969 553 77997
rect 544 77949 548 77969
rect 579 77928 582 78018
rect 612 78000 624 78001
rect 599 77998 649 78000
rect 612 77997 624 77998
rect 610 77990 632 77997
rect 607 77989 632 77990
rect 586 77982 644 77989
rect 607 77981 644 77982
rect 607 77965 610 77981
rect 616 77965 644 77981
rect 607 77964 644 77965
rect 586 77957 644 77964
rect 607 77956 610 77957
rect 612 77949 632 77957
rect 612 77945 624 77949
rect 649 77948 651 77998
rect 544 77911 548 77919
rect 400 77879 408 77909
rect 420 77879 436 77909
rect 400 77875 436 77879
rect 400 77867 430 77875
rect 428 77851 430 77867
rect 476 77839 480 77907
rect 544 77877 552 77911
rect 578 77877 582 77911
rect 544 77869 548 77877
rect 544 77839 586 77840
rect 288 77799 292 77831
rect 296 77829 368 77837
rect 378 77829 450 77837
rect 544 77832 548 77839
rect 439 77801 444 77829
rect 120 77785 170 77787
rect 76 77781 130 77785
rect 110 77776 130 77781
rect 60 77751 67 77761
rect 76 77751 77 77771
rect 96 77742 99 77776
rect 109 77751 110 77771
rect 119 77751 126 77761
rect 76 77735 92 77741
rect 94 77735 110 77741
rect 170 77735 172 77785
rect 186 77719 190 77753
rect 216 77719 220 77753
rect 213 77687 224 77719
rect 282 77715 292 77799
rect 296 77793 368 77801
rect 378 77793 450 77801
rect 468 77798 473 77832
rect 428 77763 430 77779
rect 251 77687 292 77715
rect 318 77694 324 77763
rect 12 77682 62 77684
rect 28 77673 59 77681
rect 62 77673 64 77682
rect 251 77681 263 77687
rect 28 77665 64 77673
rect 127 77673 158 77681
rect 127 77666 182 77673
rect 127 77665 161 77666
rect 59 77649 64 77665
rect 158 77649 161 77665
rect 253 77653 263 77681
rect 273 77653 293 77687
rect 318 77684 335 77694
rect 303 77668 316 77678
rect 318 77668 324 77684
rect 346 77678 348 77763
rect 400 77755 430 77763
rect 476 77761 480 77829
rect 511 77798 582 77832
rect 544 77791 548 77798
rect 400 77751 436 77755
rect 400 77721 408 77751
rect 420 77721 436 77751
rect 544 77753 548 77761
rect 28 77641 64 77649
rect 127 77648 161 77649
rect 127 77641 182 77648
rect 62 77632 64 77641
rect 282 77595 292 77653
rect 295 77644 324 77668
rect 333 77668 353 77678
rect 428 77674 430 77721
rect 476 77681 480 77749
rect 544 77719 552 77753
rect 578 77719 582 77753
rect 544 77711 548 77719
rect 367 77668 380 77674
rect 333 77644 380 77668
rect 318 77631 324 77644
rect 346 77631 348 77644
rect 367 77640 380 77644
rect 396 77640 408 77674
rect 420 77640 436 77674
rect 544 77671 553 77699
rect 319 77620 346 77631
rect 120 77579 170 77581
rect 76 77573 92 77579
rect 94 77573 110 77579
rect 76 77563 99 77572
rect 60 77553 67 77563
rect 76 77543 77 77563
rect 96 77538 99 77563
rect 109 77543 110 77563
rect 119 77553 126 77563
rect 76 77529 110 77533
rect 170 77529 172 77579
rect 186 77561 190 77595
rect 216 77561 220 77595
rect 182 77523 224 77524
rect 186 77499 220 77516
rect 223 77499 257 77516
rect 182 77482 257 77499
rect 182 77481 224 77482
rect 160 77475 246 77481
rect 288 77475 292 77595
rect 296 77593 368 77601
rect 428 77593 430 77640
rect 476 77603 480 77671
rect 485 77627 495 77661
rect 505 77633 525 77661
rect 505 77627 519 77633
rect 544 77627 555 77671
rect 485 77603 492 77627
rect 579 77612 582 77702
rect 612 77684 624 77685
rect 599 77682 649 77684
rect 612 77681 624 77682
rect 610 77674 632 77681
rect 607 77673 632 77674
rect 586 77666 644 77673
rect 607 77665 644 77666
rect 607 77649 610 77665
rect 616 77649 644 77665
rect 607 77648 644 77649
rect 586 77641 644 77648
rect 607 77640 610 77641
rect 612 77633 632 77641
rect 612 77629 624 77633
rect 649 77632 651 77682
rect 544 77595 548 77603
rect 400 77563 408 77593
rect 420 77563 436 77593
rect 400 77559 436 77563
rect 400 77551 430 77559
rect 428 77535 430 77551
rect 476 77523 480 77591
rect 544 77561 552 77595
rect 578 77561 582 77595
rect 544 77553 548 77561
rect 295 77482 300 77516
rect 324 77482 329 77516
rect 378 77513 450 77521
rect 544 77518 548 77523
rect 544 77514 582 77518
rect 544 77499 552 77514
rect 578 77499 582 77514
rect 544 77481 586 77499
rect 522 77475 608 77481
rect 182 77459 224 77475
rect 544 77459 586 77475
rect 17 77445 67 77447
rect 119 77445 169 77447
rect 186 77445 220 77459
rect 548 77445 582 77459
rect 599 77445 649 77447
rect 42 77403 59 77437
rect 67 77395 69 77445
rect 160 77437 246 77445
rect 522 77437 608 77445
rect 76 77403 110 77437
rect 127 77403 144 77437
rect 152 77403 161 77437
rect 162 77435 195 77437
rect 224 77435 244 77437
rect 162 77403 244 77435
rect 524 77435 548 77437
rect 573 77435 582 77437
rect 586 77435 606 77437
rect 160 77395 246 77403
rect 186 77379 220 77395
rect 182 77365 224 77366
rect 160 77359 182 77365
rect 224 77359 246 77365
rect 186 77324 220 77358
rect 223 77324 257 77358
rect 120 77311 170 77313
rect 76 77307 130 77311
rect 110 77302 130 77307
rect 60 77277 67 77287
rect 76 77277 77 77297
rect 96 77268 99 77302
rect 109 77277 110 77297
rect 119 77277 126 77287
rect 76 77261 92 77267
rect 94 77261 110 77267
rect 170 77261 172 77311
rect 186 77245 190 77279
rect 216 77245 220 77279
rect 288 77245 292 77433
rect 476 77365 480 77433
rect 524 77403 606 77435
rect 607 77403 616 77437
rect 522 77395 608 77403
rect 649 77395 651 77445
rect 548 77379 582 77395
rect 522 77360 548 77365
rect 522 77359 582 77360
rect 586 77359 608 77365
rect 295 77324 300 77358
rect 324 77324 329 77358
rect 544 77356 582 77359
rect 378 77319 450 77327
rect 428 77289 430 77305
rect 400 77281 430 77289
rect 476 77287 480 77355
rect 544 77326 552 77356
rect 578 77326 582 77356
rect 544 77317 548 77326
rect 400 77277 436 77281
rect 400 77247 408 77277
rect 420 77247 436 77277
rect 544 77279 548 77287
rect 12 77208 62 77210
rect 28 77199 59 77207
rect 62 77199 64 77208
rect 28 77191 64 77199
rect 127 77199 158 77207
rect 127 77192 182 77199
rect 215 77197 224 77225
rect 127 77191 161 77192
rect 59 77175 64 77191
rect 158 77175 161 77191
rect 28 77167 64 77175
rect 127 77174 161 77175
rect 127 77167 182 77174
rect 62 77158 64 77167
rect 213 77159 224 77197
rect 282 77187 292 77245
rect 296 77239 368 77247
rect 319 77209 346 77220
rect 318 77196 324 77209
rect 346 77196 348 77209
rect 428 77200 430 77247
rect 443 77237 450 77239
rect 476 77207 480 77275
rect 544 77245 552 77279
rect 578 77245 582 77279
rect 481 77213 517 77241
rect 481 77207 495 77213
rect 367 77196 380 77200
rect 251 77153 263 77187
rect 273 77153 293 77187
rect 295 77172 324 77196
rect 303 77162 316 77172
rect 318 77156 324 77172
rect 333 77172 380 77196
rect 333 77162 353 77172
rect 367 77166 380 77172
rect 396 77166 408 77200
rect 420 77166 436 77200
rect 120 77105 170 77107
rect 76 77099 92 77105
rect 94 77099 110 77105
rect 76 77089 99 77098
rect 60 77079 67 77089
rect 76 77069 77 77089
rect 96 77064 99 77089
rect 109 77069 110 77089
rect 119 77079 126 77089
rect 76 77055 110 77059
rect 170 77055 172 77105
rect 186 77087 190 77121
rect 216 77087 220 77121
rect 186 77010 220 77044
rect 282 77041 292 77153
rect 318 77146 335 77156
rect 318 77077 324 77146
rect 346 77077 348 77162
rect 428 77119 430 77166
rect 476 77129 480 77197
rect 485 77179 495 77207
rect 505 77207 519 77213
rect 544 77207 555 77245
rect 505 77179 525 77207
rect 544 77179 553 77207
rect 544 77159 548 77179
rect 579 77138 582 77228
rect 612 77210 624 77211
rect 599 77208 649 77210
rect 612 77207 624 77208
rect 610 77200 632 77207
rect 607 77199 632 77200
rect 586 77192 644 77199
rect 607 77191 644 77192
rect 607 77175 610 77191
rect 616 77175 644 77191
rect 607 77174 644 77175
rect 586 77167 644 77174
rect 607 77166 610 77167
rect 612 77159 632 77167
rect 612 77155 624 77159
rect 649 77158 651 77208
rect 544 77121 548 77129
rect 400 77089 408 77119
rect 420 77089 436 77119
rect 400 77085 436 77089
rect 400 77077 430 77085
rect 428 77061 430 77077
rect 476 77049 480 77117
rect 544 77087 552 77121
rect 578 77087 582 77121
rect 544 77079 548 77087
rect 544 77049 586 77050
rect 288 77009 292 77041
rect 296 77039 368 77047
rect 378 77039 450 77047
rect 544 77042 548 77049
rect 439 77011 444 77039
rect 120 76995 170 76997
rect 76 76991 130 76995
rect 110 76986 130 76991
rect 60 76961 67 76971
rect 76 76961 77 76981
rect 96 76952 99 76986
rect 109 76961 110 76981
rect 119 76961 126 76971
rect 76 76945 92 76951
rect 94 76945 110 76951
rect 170 76945 172 76995
rect 186 76929 190 76963
rect 216 76929 220 76963
rect 213 76897 224 76929
rect 282 76925 292 77009
rect 296 77003 368 77011
rect 378 77003 450 77011
rect 468 77008 473 77042
rect 428 76973 430 76989
rect 251 76897 292 76925
rect 318 76904 324 76973
rect 12 76892 62 76894
rect 28 76883 59 76891
rect 62 76883 64 76892
rect 251 76891 263 76897
rect 28 76875 64 76883
rect 127 76883 158 76891
rect 127 76876 182 76883
rect 127 76875 161 76876
rect 59 76859 64 76875
rect 158 76859 161 76875
rect 253 76863 263 76891
rect 273 76863 293 76897
rect 318 76894 335 76904
rect 303 76878 316 76888
rect 318 76878 324 76894
rect 346 76888 348 76973
rect 400 76965 430 76973
rect 476 76971 480 77039
rect 511 77008 582 77042
rect 544 77001 548 77008
rect 400 76961 436 76965
rect 400 76931 408 76961
rect 420 76931 436 76961
rect 544 76963 548 76971
rect 28 76851 64 76859
rect 127 76858 161 76859
rect 127 76851 182 76858
rect 62 76842 64 76851
rect 282 76805 292 76863
rect 295 76854 324 76878
rect 333 76878 353 76888
rect 428 76884 430 76931
rect 476 76891 480 76959
rect 544 76929 552 76963
rect 578 76929 582 76963
rect 544 76921 548 76929
rect 367 76878 380 76884
rect 333 76854 380 76878
rect 318 76841 324 76854
rect 346 76841 348 76854
rect 367 76850 380 76854
rect 396 76850 408 76884
rect 420 76850 436 76884
rect 544 76881 553 76909
rect 319 76830 346 76841
rect 120 76789 170 76791
rect 76 76783 92 76789
rect 94 76783 110 76789
rect 76 76773 99 76782
rect 60 76763 67 76773
rect 76 76753 77 76773
rect 96 76748 99 76773
rect 109 76753 110 76773
rect 119 76763 126 76773
rect 76 76739 110 76743
rect 170 76739 172 76789
rect 186 76771 190 76805
rect 216 76771 220 76805
rect 182 76733 224 76734
rect 186 76709 220 76726
rect 223 76709 257 76726
rect 182 76692 257 76709
rect 182 76691 224 76692
rect 160 76685 246 76691
rect 288 76685 292 76805
rect 296 76803 368 76811
rect 428 76803 430 76850
rect 476 76813 480 76881
rect 485 76837 495 76871
rect 505 76843 525 76871
rect 505 76837 519 76843
rect 544 76837 555 76881
rect 485 76813 492 76837
rect 579 76822 582 76912
rect 612 76894 624 76895
rect 599 76892 649 76894
rect 612 76891 624 76892
rect 610 76884 632 76891
rect 607 76883 632 76884
rect 586 76876 644 76883
rect 607 76875 644 76876
rect 607 76859 610 76875
rect 616 76859 644 76875
rect 607 76858 644 76859
rect 586 76851 644 76858
rect 607 76850 610 76851
rect 612 76843 632 76851
rect 612 76839 624 76843
rect 649 76842 651 76892
rect 544 76805 548 76813
rect 400 76773 408 76803
rect 420 76773 436 76803
rect 400 76769 436 76773
rect 400 76761 430 76769
rect 428 76745 430 76761
rect 476 76733 480 76801
rect 544 76771 552 76805
rect 578 76771 582 76805
rect 544 76763 548 76771
rect 295 76692 300 76726
rect 324 76692 329 76726
rect 378 76723 450 76731
rect 544 76728 548 76733
rect 544 76724 582 76728
rect 544 76709 552 76724
rect 578 76709 582 76724
rect 544 76691 586 76709
rect 522 76685 608 76691
rect 182 76669 224 76685
rect 544 76669 586 76685
rect 17 76655 67 76657
rect 119 76655 169 76657
rect 186 76655 220 76669
rect 548 76655 582 76669
rect 599 76655 649 76657
rect 42 76613 59 76647
rect 67 76605 69 76655
rect 160 76647 246 76655
rect 522 76647 608 76655
rect 76 76613 110 76647
rect 127 76613 144 76647
rect 152 76613 161 76647
rect 162 76645 195 76647
rect 224 76645 244 76647
rect 162 76613 244 76645
rect 524 76645 548 76647
rect 573 76645 582 76647
rect 586 76645 606 76647
rect 160 76605 246 76613
rect 186 76589 220 76605
rect 182 76575 224 76576
rect 160 76569 182 76575
rect 224 76569 246 76575
rect 186 76534 220 76568
rect 223 76534 257 76568
rect 120 76521 170 76523
rect 76 76517 130 76521
rect 110 76512 130 76517
rect 60 76487 67 76497
rect 76 76487 77 76507
rect 96 76478 99 76512
rect 109 76487 110 76507
rect 119 76487 126 76497
rect 76 76471 92 76477
rect 94 76471 110 76477
rect 170 76471 172 76521
rect 186 76455 190 76489
rect 216 76455 220 76489
rect 288 76455 292 76643
rect 476 76575 480 76643
rect 524 76613 606 76645
rect 607 76613 616 76647
rect 522 76605 608 76613
rect 649 76605 651 76655
rect 548 76589 582 76605
rect 522 76570 548 76575
rect 522 76569 582 76570
rect 586 76569 608 76575
rect 295 76534 300 76568
rect 324 76534 329 76568
rect 544 76566 582 76569
rect 378 76529 450 76537
rect 428 76499 430 76515
rect 400 76491 430 76499
rect 476 76497 480 76565
rect 544 76536 552 76566
rect 578 76536 582 76566
rect 544 76527 548 76536
rect 400 76487 436 76491
rect 400 76457 408 76487
rect 420 76457 436 76487
rect 544 76489 548 76497
rect 12 76418 62 76420
rect 28 76409 59 76417
rect 62 76409 64 76418
rect 28 76401 64 76409
rect 127 76409 158 76417
rect 127 76402 182 76409
rect 215 76407 224 76435
rect 127 76401 161 76402
rect 59 76385 64 76401
rect 158 76385 161 76401
rect 28 76377 64 76385
rect 127 76384 161 76385
rect 127 76377 182 76384
rect 62 76368 64 76377
rect 213 76369 224 76407
rect 282 76397 292 76455
rect 296 76449 368 76457
rect 319 76419 346 76430
rect 318 76406 324 76419
rect 346 76406 348 76419
rect 428 76410 430 76457
rect 443 76447 450 76449
rect 476 76417 480 76485
rect 544 76455 552 76489
rect 578 76455 582 76489
rect 481 76423 517 76451
rect 481 76417 495 76423
rect 367 76406 380 76410
rect 251 76363 263 76397
rect 273 76363 293 76397
rect 295 76382 324 76406
rect 303 76372 316 76382
rect 318 76366 324 76382
rect 333 76382 380 76406
rect 333 76372 353 76382
rect 367 76376 380 76382
rect 396 76376 408 76410
rect 420 76376 436 76410
rect 120 76315 170 76317
rect 76 76309 92 76315
rect 94 76309 110 76315
rect 76 76299 99 76308
rect 60 76289 67 76299
rect 76 76279 77 76299
rect 96 76274 99 76299
rect 109 76279 110 76299
rect 119 76289 126 76299
rect 76 76265 110 76269
rect 170 76265 172 76315
rect 186 76297 190 76331
rect 216 76297 220 76331
rect 186 76220 220 76254
rect 282 76251 292 76363
rect 318 76356 335 76366
rect 318 76287 324 76356
rect 346 76287 348 76372
rect 428 76329 430 76376
rect 476 76339 480 76407
rect 485 76389 495 76417
rect 505 76417 519 76423
rect 544 76417 555 76455
rect 505 76389 525 76417
rect 544 76389 553 76417
rect 544 76369 548 76389
rect 579 76348 582 76438
rect 612 76420 624 76421
rect 599 76418 649 76420
rect 612 76417 624 76418
rect 610 76410 632 76417
rect 607 76409 632 76410
rect 586 76402 644 76409
rect 607 76401 644 76402
rect 607 76385 610 76401
rect 616 76385 644 76401
rect 607 76384 644 76385
rect 586 76377 644 76384
rect 607 76376 610 76377
rect 612 76369 632 76377
rect 612 76365 624 76369
rect 649 76368 651 76418
rect 544 76331 548 76339
rect 400 76299 408 76329
rect 420 76299 436 76329
rect 400 76295 436 76299
rect 400 76287 430 76295
rect 428 76271 430 76287
rect 476 76259 480 76327
rect 544 76297 552 76331
rect 578 76297 582 76331
rect 544 76289 548 76297
rect 544 76259 586 76260
rect 288 76219 292 76251
rect 296 76249 368 76257
rect 378 76249 450 76257
rect 544 76252 548 76259
rect 439 76221 444 76249
rect 120 76205 170 76207
rect 76 76201 130 76205
rect 110 76196 130 76201
rect 60 76171 67 76181
rect 76 76171 77 76191
rect 96 76162 99 76196
rect 109 76171 110 76191
rect 119 76171 126 76181
rect 76 76155 92 76161
rect 94 76155 110 76161
rect 170 76155 172 76205
rect 186 76139 190 76173
rect 216 76139 220 76173
rect 213 76107 224 76139
rect 282 76135 292 76219
rect 296 76213 368 76221
rect 378 76213 450 76221
rect 468 76218 473 76252
rect 428 76183 430 76199
rect 251 76107 292 76135
rect 318 76114 324 76183
rect 12 76102 62 76104
rect 28 76093 59 76101
rect 62 76093 64 76102
rect 251 76101 263 76107
rect 28 76085 64 76093
rect 127 76093 158 76101
rect 127 76086 182 76093
rect 127 76085 161 76086
rect 59 76069 64 76085
rect 158 76069 161 76085
rect 253 76073 263 76101
rect 273 76073 293 76107
rect 318 76104 335 76114
rect 303 76088 316 76098
rect 318 76088 324 76104
rect 346 76098 348 76183
rect 400 76175 430 76183
rect 476 76181 480 76249
rect 511 76218 582 76252
rect 544 76211 548 76218
rect 400 76171 436 76175
rect 400 76141 408 76171
rect 420 76141 436 76171
rect 544 76173 548 76181
rect 28 76061 64 76069
rect 127 76068 161 76069
rect 127 76061 182 76068
rect 62 76052 64 76061
rect 282 76015 292 76073
rect 295 76064 324 76088
rect 333 76088 353 76098
rect 428 76094 430 76141
rect 476 76101 480 76169
rect 544 76139 552 76173
rect 578 76139 582 76173
rect 544 76131 548 76139
rect 367 76088 380 76094
rect 333 76064 380 76088
rect 318 76051 324 76064
rect 346 76051 348 76064
rect 367 76060 380 76064
rect 396 76060 408 76094
rect 420 76060 436 76094
rect 544 76091 553 76119
rect 319 76040 346 76051
rect 120 75999 170 76001
rect 76 75993 92 75999
rect 94 75993 110 75999
rect 76 75983 99 75992
rect 60 75973 67 75983
rect 76 75963 77 75983
rect 96 75958 99 75983
rect 109 75963 110 75983
rect 119 75973 126 75983
rect 76 75949 110 75953
rect 170 75949 172 75999
rect 186 75981 190 76015
rect 216 75981 220 76015
rect 182 75943 224 75944
rect 186 75919 220 75936
rect 223 75919 257 75936
rect 182 75902 257 75919
rect 182 75901 224 75902
rect 160 75895 246 75901
rect 288 75895 292 76015
rect 296 76013 368 76021
rect 428 76013 430 76060
rect 476 76023 480 76091
rect 485 76047 495 76081
rect 505 76053 525 76081
rect 505 76047 519 76053
rect 544 76047 555 76091
rect 485 76023 492 76047
rect 579 76032 582 76122
rect 612 76104 624 76105
rect 599 76102 649 76104
rect 612 76101 624 76102
rect 610 76094 632 76101
rect 607 76093 632 76094
rect 586 76086 644 76093
rect 607 76085 644 76086
rect 607 76069 610 76085
rect 616 76069 644 76085
rect 607 76068 644 76069
rect 586 76061 644 76068
rect 607 76060 610 76061
rect 612 76053 632 76061
rect 612 76049 624 76053
rect 649 76052 651 76102
rect 544 76015 548 76023
rect 400 75983 408 76013
rect 420 75983 436 76013
rect 400 75979 436 75983
rect 400 75971 430 75979
rect 428 75955 430 75971
rect 476 75943 480 76011
rect 544 75981 552 76015
rect 578 75981 582 76015
rect 544 75973 548 75981
rect 295 75902 300 75936
rect 324 75902 329 75936
rect 378 75933 450 75941
rect 544 75938 548 75943
rect 544 75934 582 75938
rect 544 75919 552 75934
rect 578 75919 582 75934
rect 544 75901 586 75919
rect 522 75895 608 75901
rect 182 75879 224 75895
rect 544 75879 586 75895
rect 17 75865 67 75867
rect 119 75865 169 75867
rect 186 75865 220 75879
rect 548 75865 582 75879
rect 599 75865 649 75867
rect 42 75823 59 75857
rect 67 75815 69 75865
rect 160 75857 246 75865
rect 522 75857 608 75865
rect 76 75823 110 75857
rect 127 75823 144 75857
rect 152 75823 161 75857
rect 162 75855 195 75857
rect 224 75855 244 75857
rect 162 75823 244 75855
rect 524 75855 548 75857
rect 573 75855 582 75857
rect 586 75855 606 75857
rect 160 75815 246 75823
rect 186 75799 220 75815
rect 182 75785 224 75786
rect 160 75779 182 75785
rect 224 75779 246 75785
rect 186 75744 220 75778
rect 223 75744 257 75778
rect 120 75731 170 75733
rect 76 75727 130 75731
rect 110 75722 130 75727
rect 60 75697 67 75707
rect 76 75697 77 75717
rect 96 75688 99 75722
rect 109 75697 110 75717
rect 119 75697 126 75707
rect 76 75681 92 75687
rect 94 75681 110 75687
rect 170 75681 172 75731
rect 186 75665 190 75699
rect 216 75665 220 75699
rect 288 75665 292 75853
rect 476 75785 480 75853
rect 524 75823 606 75855
rect 607 75823 616 75857
rect 522 75815 608 75823
rect 649 75815 651 75865
rect 548 75799 582 75815
rect 522 75780 548 75785
rect 522 75779 582 75780
rect 586 75779 608 75785
rect 295 75744 300 75778
rect 324 75744 329 75778
rect 544 75776 582 75779
rect 378 75739 450 75747
rect 428 75709 430 75725
rect 400 75701 430 75709
rect 476 75707 480 75775
rect 544 75746 552 75776
rect 578 75746 582 75776
rect 544 75737 548 75746
rect 400 75697 436 75701
rect 400 75667 408 75697
rect 420 75667 436 75697
rect 544 75699 548 75707
rect 12 75628 62 75630
rect 28 75619 59 75627
rect 62 75619 64 75628
rect 28 75611 64 75619
rect 127 75619 158 75627
rect 127 75612 182 75619
rect 215 75617 224 75645
rect 127 75611 161 75612
rect 59 75595 64 75611
rect 158 75595 161 75611
rect 28 75587 64 75595
rect 127 75594 161 75595
rect 127 75587 182 75594
rect 62 75578 64 75587
rect 213 75579 224 75617
rect 282 75607 292 75665
rect 296 75659 368 75667
rect 319 75629 346 75640
rect 318 75616 324 75629
rect 346 75616 348 75629
rect 428 75620 430 75667
rect 443 75657 450 75659
rect 476 75627 480 75695
rect 544 75665 552 75699
rect 578 75665 582 75699
rect 481 75633 517 75661
rect 481 75627 495 75633
rect 367 75616 380 75620
rect 251 75573 263 75607
rect 273 75573 293 75607
rect 295 75592 324 75616
rect 303 75582 316 75592
rect 318 75576 324 75592
rect 333 75592 380 75616
rect 333 75582 353 75592
rect 367 75586 380 75592
rect 396 75586 408 75620
rect 420 75586 436 75620
rect 120 75525 170 75527
rect 76 75519 92 75525
rect 94 75519 110 75525
rect 76 75509 99 75518
rect 60 75499 67 75509
rect 76 75489 77 75509
rect 96 75484 99 75509
rect 109 75489 110 75509
rect 119 75499 126 75509
rect 76 75475 110 75479
rect 170 75475 172 75525
rect 186 75507 190 75541
rect 216 75507 220 75541
rect 186 75430 220 75464
rect 282 75461 292 75573
rect 318 75566 335 75576
rect 318 75497 324 75566
rect 346 75497 348 75582
rect 428 75539 430 75586
rect 476 75549 480 75617
rect 485 75599 495 75627
rect 505 75627 519 75633
rect 544 75627 555 75665
rect 505 75599 525 75627
rect 544 75599 553 75627
rect 544 75579 548 75599
rect 579 75558 582 75648
rect 612 75630 624 75631
rect 599 75628 649 75630
rect 612 75627 624 75628
rect 610 75620 632 75627
rect 607 75619 632 75620
rect 586 75612 644 75619
rect 607 75611 644 75612
rect 607 75595 610 75611
rect 616 75595 644 75611
rect 607 75594 644 75595
rect 586 75587 644 75594
rect 607 75586 610 75587
rect 612 75579 632 75587
rect 612 75575 624 75579
rect 649 75578 651 75628
rect 544 75541 548 75549
rect 400 75509 408 75539
rect 420 75509 436 75539
rect 400 75505 436 75509
rect 400 75497 430 75505
rect 428 75481 430 75497
rect 476 75469 480 75537
rect 544 75507 552 75541
rect 578 75507 582 75541
rect 544 75499 548 75507
rect 544 75469 586 75470
rect 288 75429 292 75461
rect 296 75459 368 75467
rect 378 75459 450 75467
rect 544 75462 548 75469
rect 439 75431 444 75459
rect 120 75415 170 75417
rect 76 75411 130 75415
rect 110 75406 130 75411
rect 60 75381 67 75391
rect 76 75381 77 75401
rect 96 75372 99 75406
rect 109 75381 110 75401
rect 119 75381 126 75391
rect 76 75365 92 75371
rect 94 75365 110 75371
rect 170 75365 172 75415
rect 186 75349 190 75383
rect 216 75349 220 75383
rect 213 75317 224 75349
rect 282 75345 292 75429
rect 296 75423 368 75431
rect 378 75423 450 75431
rect 468 75428 473 75462
rect 428 75393 430 75409
rect 251 75317 292 75345
rect 318 75324 324 75393
rect 12 75312 62 75314
rect 28 75303 59 75311
rect 62 75303 64 75312
rect 251 75311 263 75317
rect 28 75295 64 75303
rect 127 75303 158 75311
rect 127 75296 182 75303
rect 127 75295 161 75296
rect 59 75279 64 75295
rect 158 75279 161 75295
rect 253 75283 263 75311
rect 273 75283 293 75317
rect 318 75314 335 75324
rect 303 75298 316 75308
rect 318 75298 324 75314
rect 346 75308 348 75393
rect 400 75385 430 75393
rect 476 75391 480 75459
rect 511 75428 582 75462
rect 544 75421 548 75428
rect 400 75381 436 75385
rect 400 75351 408 75381
rect 420 75351 436 75381
rect 544 75383 548 75391
rect 28 75271 64 75279
rect 127 75278 161 75279
rect 127 75271 182 75278
rect 62 75262 64 75271
rect 282 75225 292 75283
rect 295 75274 324 75298
rect 333 75298 353 75308
rect 428 75304 430 75351
rect 476 75311 480 75379
rect 544 75349 552 75383
rect 578 75349 582 75383
rect 544 75341 548 75349
rect 367 75298 380 75304
rect 333 75274 380 75298
rect 318 75261 324 75274
rect 346 75261 348 75274
rect 367 75270 380 75274
rect 396 75270 408 75304
rect 420 75270 436 75304
rect 544 75301 553 75329
rect 319 75250 346 75261
rect 120 75209 170 75211
rect 76 75203 92 75209
rect 94 75203 110 75209
rect 76 75193 99 75202
rect 60 75183 67 75193
rect 76 75173 77 75193
rect 96 75168 99 75193
rect 109 75173 110 75193
rect 119 75183 126 75193
rect 76 75159 110 75163
rect 170 75159 172 75209
rect 186 75191 190 75225
rect 216 75191 220 75225
rect 182 75153 224 75154
rect 186 75129 220 75146
rect 223 75129 257 75146
rect 182 75112 257 75129
rect 182 75111 224 75112
rect 160 75105 246 75111
rect 288 75105 292 75225
rect 296 75223 368 75231
rect 428 75223 430 75270
rect 476 75233 480 75301
rect 485 75257 495 75291
rect 505 75263 525 75291
rect 505 75257 519 75263
rect 544 75257 555 75301
rect 485 75233 492 75257
rect 579 75242 582 75332
rect 612 75314 624 75315
rect 599 75312 649 75314
rect 612 75311 624 75312
rect 610 75304 632 75311
rect 607 75303 632 75304
rect 586 75296 644 75303
rect 607 75295 644 75296
rect 607 75279 610 75295
rect 616 75279 644 75295
rect 607 75278 644 75279
rect 586 75271 644 75278
rect 607 75270 610 75271
rect 612 75263 632 75271
rect 612 75259 624 75263
rect 649 75262 651 75312
rect 544 75225 548 75233
rect 400 75193 408 75223
rect 420 75193 436 75223
rect 400 75189 436 75193
rect 400 75181 430 75189
rect 428 75165 430 75181
rect 476 75153 480 75221
rect 544 75191 552 75225
rect 578 75191 582 75225
rect 544 75183 548 75191
rect 295 75112 300 75146
rect 324 75112 329 75146
rect 378 75143 450 75151
rect 544 75148 548 75153
rect 544 75144 582 75148
rect 544 75129 552 75144
rect 578 75129 582 75144
rect 544 75111 586 75129
rect 522 75105 608 75111
rect 182 75089 224 75105
rect 544 75089 586 75105
rect 17 75075 67 75077
rect 119 75075 169 75077
rect 186 75075 220 75089
rect 548 75075 582 75089
rect 599 75075 649 75077
rect 42 75033 59 75067
rect 67 75025 69 75075
rect 160 75067 246 75075
rect 522 75067 608 75075
rect 76 75033 110 75067
rect 127 75033 144 75067
rect 152 75033 161 75067
rect 162 75065 195 75067
rect 224 75065 244 75067
rect 162 75033 244 75065
rect 524 75065 548 75067
rect 573 75065 582 75067
rect 586 75065 606 75067
rect 160 75025 246 75033
rect 186 75009 220 75025
rect 182 74995 224 74996
rect 160 74989 182 74995
rect 224 74989 246 74995
rect 186 74954 220 74988
rect 223 74954 257 74988
rect 120 74941 170 74943
rect 76 74937 130 74941
rect 110 74932 130 74937
rect 60 74907 67 74917
rect 76 74907 77 74927
rect 96 74898 99 74932
rect 109 74907 110 74927
rect 119 74907 126 74917
rect 76 74891 92 74897
rect 94 74891 110 74897
rect 170 74891 172 74941
rect 186 74875 190 74909
rect 216 74875 220 74909
rect 288 74875 292 75063
rect 476 74995 480 75063
rect 524 75033 606 75065
rect 607 75033 616 75067
rect 522 75025 608 75033
rect 649 75025 651 75075
rect 548 75009 582 75025
rect 522 74990 548 74995
rect 522 74989 582 74990
rect 586 74989 608 74995
rect 295 74954 300 74988
rect 324 74954 329 74988
rect 544 74986 582 74989
rect 378 74949 450 74957
rect 428 74919 430 74935
rect 400 74911 430 74919
rect 476 74917 480 74985
rect 544 74956 552 74986
rect 578 74956 582 74986
rect 544 74947 548 74956
rect 400 74907 436 74911
rect 400 74877 408 74907
rect 420 74877 436 74907
rect 544 74909 548 74917
rect 12 74838 62 74840
rect 28 74829 59 74837
rect 62 74829 64 74838
rect 28 74821 64 74829
rect 127 74829 158 74837
rect 127 74822 182 74829
rect 215 74827 224 74855
rect 127 74821 161 74822
rect 59 74805 64 74821
rect 158 74805 161 74821
rect 28 74797 64 74805
rect 127 74804 161 74805
rect 127 74797 182 74804
rect 62 74788 64 74797
rect 213 74789 224 74827
rect 282 74817 292 74875
rect 296 74869 368 74877
rect 319 74839 346 74850
rect 318 74826 324 74839
rect 346 74826 348 74839
rect 428 74830 430 74877
rect 443 74867 450 74869
rect 476 74837 480 74905
rect 544 74875 552 74909
rect 578 74875 582 74909
rect 481 74843 517 74871
rect 481 74837 495 74843
rect 367 74826 380 74830
rect 251 74783 263 74817
rect 273 74783 293 74817
rect 295 74802 324 74826
rect 303 74792 316 74802
rect 318 74786 324 74802
rect 333 74802 380 74826
rect 333 74792 353 74802
rect 367 74796 380 74802
rect 396 74796 408 74830
rect 420 74796 436 74830
rect 120 74735 170 74737
rect 76 74729 92 74735
rect 94 74729 110 74735
rect 76 74719 99 74728
rect 60 74709 67 74719
rect 76 74699 77 74719
rect 96 74694 99 74719
rect 109 74699 110 74719
rect 119 74709 126 74719
rect 76 74685 110 74689
rect 170 74685 172 74735
rect 186 74717 190 74751
rect 216 74717 220 74751
rect 186 74640 220 74674
rect 282 74671 292 74783
rect 318 74776 335 74786
rect 318 74707 324 74776
rect 346 74707 348 74792
rect 428 74749 430 74796
rect 476 74759 480 74827
rect 485 74809 495 74837
rect 505 74837 519 74843
rect 544 74837 555 74875
rect 505 74809 525 74837
rect 544 74809 553 74837
rect 544 74789 548 74809
rect 579 74768 582 74858
rect 612 74840 624 74841
rect 599 74838 649 74840
rect 612 74837 624 74838
rect 610 74830 632 74837
rect 607 74829 632 74830
rect 586 74822 644 74829
rect 607 74821 644 74822
rect 607 74805 610 74821
rect 616 74805 644 74821
rect 607 74804 644 74805
rect 586 74797 644 74804
rect 607 74796 610 74797
rect 612 74789 632 74797
rect 612 74785 624 74789
rect 649 74788 651 74838
rect 544 74751 548 74759
rect 400 74719 408 74749
rect 420 74719 436 74749
rect 400 74715 436 74719
rect 400 74707 430 74715
rect 428 74691 430 74707
rect 476 74679 480 74747
rect 544 74717 552 74751
rect 578 74717 582 74751
rect 544 74709 548 74717
rect 544 74679 586 74680
rect 288 74639 292 74671
rect 296 74669 368 74677
rect 378 74669 450 74677
rect 544 74672 548 74679
rect 439 74641 444 74669
rect 120 74625 170 74627
rect 76 74621 130 74625
rect 110 74616 130 74621
rect 60 74591 67 74601
rect 76 74591 77 74611
rect 96 74582 99 74616
rect 109 74591 110 74611
rect 119 74591 126 74601
rect 76 74575 92 74581
rect 94 74575 110 74581
rect 170 74575 172 74625
rect 186 74559 190 74593
rect 216 74559 220 74593
rect 213 74527 224 74559
rect 282 74555 292 74639
rect 296 74633 368 74641
rect 378 74633 450 74641
rect 468 74638 473 74672
rect 428 74603 430 74619
rect 251 74527 292 74555
rect 318 74534 324 74603
rect 12 74522 62 74524
rect 28 74513 59 74521
rect 62 74513 64 74522
rect 251 74521 263 74527
rect 28 74505 64 74513
rect 127 74513 158 74521
rect 127 74506 182 74513
rect 127 74505 161 74506
rect 59 74489 64 74505
rect 158 74489 161 74505
rect 253 74493 263 74521
rect 273 74493 293 74527
rect 318 74524 335 74534
rect 303 74508 316 74518
rect 318 74508 324 74524
rect 346 74518 348 74603
rect 400 74595 430 74603
rect 476 74601 480 74669
rect 511 74638 582 74672
rect 544 74631 548 74638
rect 400 74591 436 74595
rect 400 74561 408 74591
rect 420 74561 436 74591
rect 544 74593 548 74601
rect 28 74481 64 74489
rect 127 74488 161 74489
rect 127 74481 182 74488
rect 62 74472 64 74481
rect 282 74435 292 74493
rect 295 74484 324 74508
rect 333 74508 353 74518
rect 428 74514 430 74561
rect 476 74521 480 74589
rect 544 74559 552 74593
rect 578 74559 582 74593
rect 544 74551 548 74559
rect 367 74508 380 74514
rect 333 74484 380 74508
rect 318 74471 324 74484
rect 346 74471 348 74484
rect 367 74480 380 74484
rect 396 74480 408 74514
rect 420 74480 436 74514
rect 544 74511 553 74539
rect 319 74460 346 74471
rect 120 74419 170 74421
rect 76 74413 92 74419
rect 94 74413 110 74419
rect 76 74403 99 74412
rect 60 74393 67 74403
rect 76 74383 77 74403
rect 96 74378 99 74403
rect 109 74383 110 74403
rect 119 74393 126 74403
rect 76 74369 110 74373
rect 170 74369 172 74419
rect 186 74401 190 74435
rect 216 74401 220 74435
rect 182 74363 224 74364
rect 186 74339 220 74356
rect 223 74339 257 74356
rect 182 74322 257 74339
rect 182 74321 224 74322
rect 160 74315 246 74321
rect 288 74315 292 74435
rect 296 74433 368 74441
rect 428 74433 430 74480
rect 476 74443 480 74511
rect 485 74467 495 74501
rect 505 74473 525 74501
rect 505 74467 519 74473
rect 544 74467 555 74511
rect 485 74443 492 74467
rect 579 74452 582 74542
rect 612 74524 624 74525
rect 599 74522 649 74524
rect 612 74521 624 74522
rect 610 74514 632 74521
rect 607 74513 632 74514
rect 586 74506 644 74513
rect 607 74505 644 74506
rect 607 74489 610 74505
rect 616 74489 644 74505
rect 607 74488 644 74489
rect 586 74481 644 74488
rect 607 74480 610 74481
rect 612 74473 632 74481
rect 612 74469 624 74473
rect 649 74472 651 74522
rect 544 74435 548 74443
rect 400 74403 408 74433
rect 420 74403 436 74433
rect 400 74399 436 74403
rect 400 74391 430 74399
rect 428 74375 430 74391
rect 476 74363 480 74431
rect 544 74401 552 74435
rect 578 74401 582 74435
rect 544 74393 548 74401
rect 295 74322 300 74356
rect 324 74322 329 74356
rect 378 74353 450 74361
rect 544 74358 548 74363
rect 544 74354 582 74358
rect 544 74339 552 74354
rect 578 74339 582 74354
rect 544 74321 586 74339
rect 522 74315 608 74321
rect 182 74299 224 74315
rect 544 74299 586 74315
rect 17 74285 67 74287
rect 119 74285 169 74287
rect 186 74285 220 74299
rect 548 74285 582 74299
rect 599 74285 649 74287
rect 42 74243 59 74277
rect 67 74235 69 74285
rect 160 74277 246 74285
rect 522 74277 608 74285
rect 76 74243 110 74277
rect 127 74243 144 74277
rect 152 74243 161 74277
rect 162 74275 195 74277
rect 224 74275 244 74277
rect 162 74243 244 74275
rect 524 74275 548 74277
rect 573 74275 582 74277
rect 586 74275 606 74277
rect 160 74235 246 74243
rect 186 74219 220 74235
rect 182 74205 224 74206
rect 160 74199 182 74205
rect 224 74199 246 74205
rect 186 74164 220 74198
rect 223 74164 257 74198
rect 120 74151 170 74153
rect 76 74147 130 74151
rect 110 74142 130 74147
rect 60 74117 67 74127
rect 76 74117 77 74137
rect 96 74108 99 74142
rect 109 74117 110 74137
rect 119 74117 126 74127
rect 76 74101 92 74107
rect 94 74101 110 74107
rect 170 74101 172 74151
rect 186 74085 190 74119
rect 216 74085 220 74119
rect 288 74085 292 74273
rect 476 74205 480 74273
rect 524 74243 606 74275
rect 607 74243 616 74277
rect 522 74235 608 74243
rect 649 74235 651 74285
rect 548 74219 582 74235
rect 522 74200 548 74205
rect 522 74199 582 74200
rect 586 74199 608 74205
rect 295 74164 300 74198
rect 324 74164 329 74198
rect 544 74196 582 74199
rect 378 74159 450 74167
rect 428 74129 430 74145
rect 400 74121 430 74129
rect 476 74127 480 74195
rect 544 74166 552 74196
rect 578 74166 582 74196
rect 544 74157 548 74166
rect 400 74117 436 74121
rect 400 74087 408 74117
rect 420 74087 436 74117
rect 544 74119 548 74127
rect 12 74048 62 74050
rect 28 74039 59 74047
rect 62 74039 64 74048
rect 28 74031 64 74039
rect 127 74039 158 74047
rect 127 74032 182 74039
rect 215 74037 224 74065
rect 127 74031 161 74032
rect 59 74015 64 74031
rect 158 74015 161 74031
rect 28 74007 64 74015
rect 127 74014 161 74015
rect 127 74007 182 74014
rect 62 73998 64 74007
rect 213 73999 224 74037
rect 282 74027 292 74085
rect 296 74079 368 74087
rect 319 74049 346 74060
rect 318 74036 324 74049
rect 346 74036 348 74049
rect 428 74040 430 74087
rect 443 74077 450 74079
rect 476 74047 480 74115
rect 544 74085 552 74119
rect 578 74085 582 74119
rect 481 74053 517 74081
rect 481 74047 495 74053
rect 367 74036 380 74040
rect 251 73993 263 74027
rect 273 73993 293 74027
rect 295 74012 324 74036
rect 303 74002 316 74012
rect 318 73996 324 74012
rect 333 74012 380 74036
rect 333 74002 353 74012
rect 367 74006 380 74012
rect 396 74006 408 74040
rect 420 74006 436 74040
rect 120 73945 170 73947
rect 76 73939 92 73945
rect 94 73939 110 73945
rect 76 73929 99 73938
rect 60 73919 67 73929
rect 76 73909 77 73929
rect 96 73904 99 73929
rect 109 73909 110 73929
rect 119 73919 126 73929
rect 76 73895 110 73899
rect 170 73895 172 73945
rect 186 73927 190 73961
rect 216 73927 220 73961
rect 186 73850 220 73884
rect 282 73881 292 73993
rect 318 73986 335 73996
rect 318 73917 324 73986
rect 346 73917 348 74002
rect 428 73959 430 74006
rect 476 73969 480 74037
rect 485 74019 495 74047
rect 505 74047 519 74053
rect 544 74047 555 74085
rect 505 74019 525 74047
rect 544 74019 553 74047
rect 544 73999 548 74019
rect 579 73978 582 74068
rect 612 74050 624 74051
rect 599 74048 649 74050
rect 612 74047 624 74048
rect 610 74040 632 74047
rect 607 74039 632 74040
rect 586 74032 644 74039
rect 607 74031 644 74032
rect 607 74015 610 74031
rect 616 74015 644 74031
rect 607 74014 644 74015
rect 586 74007 644 74014
rect 607 74006 610 74007
rect 612 73999 632 74007
rect 612 73995 624 73999
rect 649 73998 651 74048
rect 544 73961 548 73969
rect 400 73929 408 73959
rect 420 73929 436 73959
rect 400 73925 436 73929
rect 400 73917 430 73925
rect 428 73901 430 73917
rect 476 73889 480 73957
rect 544 73927 552 73961
rect 578 73927 582 73961
rect 544 73919 548 73927
rect 544 73889 586 73890
rect 288 73849 292 73881
rect 296 73879 368 73887
rect 378 73879 450 73887
rect 544 73882 548 73889
rect 439 73851 444 73879
rect 120 73835 170 73837
rect 76 73831 130 73835
rect 110 73826 130 73831
rect 60 73801 67 73811
rect 76 73801 77 73821
rect 96 73792 99 73826
rect 109 73801 110 73821
rect 119 73801 126 73811
rect 76 73785 92 73791
rect 94 73785 110 73791
rect 170 73785 172 73835
rect 186 73769 190 73803
rect 216 73769 220 73803
rect 213 73737 224 73769
rect 282 73765 292 73849
rect 296 73843 368 73851
rect 378 73843 450 73851
rect 468 73848 473 73882
rect 428 73813 430 73829
rect 251 73737 292 73765
rect 318 73744 324 73813
rect 12 73732 62 73734
rect 28 73723 59 73731
rect 62 73723 64 73732
rect 251 73731 263 73737
rect 28 73715 64 73723
rect 127 73723 158 73731
rect 127 73716 182 73723
rect 127 73715 161 73716
rect 59 73699 64 73715
rect 158 73699 161 73715
rect 253 73703 263 73731
rect 273 73703 293 73737
rect 318 73734 335 73744
rect 303 73718 316 73728
rect 318 73718 324 73734
rect 346 73728 348 73813
rect 400 73805 430 73813
rect 476 73811 480 73879
rect 511 73848 582 73882
rect 544 73841 548 73848
rect 400 73801 436 73805
rect 400 73771 408 73801
rect 420 73771 436 73801
rect 544 73803 548 73811
rect 28 73691 64 73699
rect 127 73698 161 73699
rect 127 73691 182 73698
rect 62 73682 64 73691
rect 282 73645 292 73703
rect 295 73694 324 73718
rect 333 73718 353 73728
rect 428 73724 430 73771
rect 476 73731 480 73799
rect 544 73769 552 73803
rect 578 73769 582 73803
rect 544 73761 548 73769
rect 367 73718 380 73724
rect 333 73694 380 73718
rect 318 73681 324 73694
rect 346 73681 348 73694
rect 367 73690 380 73694
rect 396 73690 408 73724
rect 420 73690 436 73724
rect 544 73721 553 73749
rect 319 73670 346 73681
rect 120 73629 170 73631
rect 76 73623 92 73629
rect 94 73623 110 73629
rect 76 73613 99 73622
rect 60 73603 67 73613
rect 76 73593 77 73613
rect 96 73588 99 73613
rect 109 73593 110 73613
rect 119 73603 126 73613
rect 76 73579 110 73583
rect 170 73579 172 73629
rect 186 73611 190 73645
rect 216 73611 220 73645
rect 182 73573 224 73574
rect 186 73549 220 73566
rect 223 73549 257 73566
rect 182 73532 257 73549
rect 182 73531 224 73532
rect 160 73525 246 73531
rect 288 73525 292 73645
rect 296 73643 368 73651
rect 428 73643 430 73690
rect 476 73653 480 73721
rect 485 73677 495 73711
rect 505 73683 525 73711
rect 505 73677 519 73683
rect 544 73677 555 73721
rect 485 73653 492 73677
rect 579 73662 582 73752
rect 612 73734 624 73735
rect 599 73732 649 73734
rect 612 73731 624 73732
rect 610 73724 632 73731
rect 607 73723 632 73724
rect 586 73716 644 73723
rect 607 73715 644 73716
rect 607 73699 610 73715
rect 616 73699 644 73715
rect 607 73698 644 73699
rect 586 73691 644 73698
rect 607 73690 610 73691
rect 612 73683 632 73691
rect 612 73679 624 73683
rect 649 73682 651 73732
rect 544 73645 548 73653
rect 400 73613 408 73643
rect 420 73613 436 73643
rect 400 73609 436 73613
rect 400 73601 430 73609
rect 428 73585 430 73601
rect 476 73573 480 73641
rect 544 73611 552 73645
rect 578 73611 582 73645
rect 544 73603 548 73611
rect 295 73532 300 73566
rect 324 73532 329 73566
rect 378 73563 450 73571
rect 544 73568 548 73573
rect 544 73564 582 73568
rect 544 73549 552 73564
rect 578 73549 582 73564
rect 544 73531 586 73549
rect 522 73525 608 73531
rect 182 73509 224 73525
rect 544 73509 586 73525
rect 17 73495 67 73497
rect 119 73495 169 73497
rect 186 73495 220 73509
rect 548 73495 582 73509
rect 599 73495 649 73497
rect 42 73453 59 73487
rect 67 73445 69 73495
rect 160 73487 246 73495
rect 522 73487 608 73495
rect 76 73453 110 73487
rect 127 73453 144 73487
rect 152 73453 161 73487
rect 162 73485 195 73487
rect 224 73485 244 73487
rect 162 73453 244 73485
rect 524 73485 548 73487
rect 573 73485 582 73487
rect 586 73485 606 73487
rect 160 73445 246 73453
rect 186 73429 220 73445
rect 182 73415 224 73416
rect 160 73409 182 73415
rect 224 73409 246 73415
rect 186 73374 220 73408
rect 223 73374 257 73408
rect 120 73361 170 73363
rect 76 73357 130 73361
rect 110 73352 130 73357
rect 60 73327 67 73337
rect 76 73327 77 73347
rect 96 73318 99 73352
rect 109 73327 110 73347
rect 119 73327 126 73337
rect 76 73311 92 73317
rect 94 73311 110 73317
rect 170 73311 172 73361
rect 186 73295 190 73329
rect 216 73295 220 73329
rect 288 73295 292 73483
rect 476 73415 480 73483
rect 524 73453 606 73485
rect 607 73453 616 73487
rect 522 73445 608 73453
rect 649 73445 651 73495
rect 548 73429 582 73445
rect 522 73410 548 73415
rect 522 73409 582 73410
rect 586 73409 608 73415
rect 295 73374 300 73408
rect 324 73374 329 73408
rect 544 73406 582 73409
rect 378 73369 450 73377
rect 428 73339 430 73355
rect 400 73331 430 73339
rect 476 73337 480 73405
rect 544 73376 552 73406
rect 578 73376 582 73406
rect 544 73367 548 73376
rect 400 73327 436 73331
rect 400 73297 408 73327
rect 420 73297 436 73327
rect 544 73329 548 73337
rect 12 73258 62 73260
rect 28 73249 59 73257
rect 62 73249 64 73258
rect 28 73241 64 73249
rect 127 73249 158 73257
rect 127 73242 182 73249
rect 215 73247 224 73275
rect 127 73241 161 73242
rect 59 73225 64 73241
rect 158 73225 161 73241
rect 28 73217 64 73225
rect 127 73224 161 73225
rect 127 73217 182 73224
rect 62 73208 64 73217
rect 213 73209 224 73247
rect 282 73237 292 73295
rect 296 73289 368 73297
rect 319 73259 346 73270
rect 318 73246 324 73259
rect 346 73246 348 73259
rect 428 73250 430 73297
rect 443 73287 450 73289
rect 476 73257 480 73325
rect 544 73295 552 73329
rect 578 73295 582 73329
rect 481 73263 517 73291
rect 481 73257 495 73263
rect 367 73246 380 73250
rect 251 73203 263 73237
rect 273 73203 293 73237
rect 295 73222 324 73246
rect 303 73212 316 73222
rect 318 73206 324 73222
rect 333 73222 380 73246
rect 333 73212 353 73222
rect 367 73216 380 73222
rect 396 73216 408 73250
rect 420 73216 436 73250
rect 120 73155 170 73157
rect 76 73149 92 73155
rect 94 73149 110 73155
rect 76 73139 99 73148
rect 60 73129 67 73139
rect 76 73119 77 73139
rect 96 73114 99 73139
rect 109 73119 110 73139
rect 119 73129 126 73139
rect 76 73105 110 73109
rect 170 73105 172 73155
rect 186 73137 190 73171
rect 216 73137 220 73171
rect 186 73060 220 73094
rect 282 73091 292 73203
rect 318 73196 335 73206
rect 318 73127 324 73196
rect 346 73127 348 73212
rect 428 73169 430 73216
rect 476 73179 480 73247
rect 485 73229 495 73257
rect 505 73257 519 73263
rect 544 73257 555 73295
rect 505 73229 525 73257
rect 544 73229 553 73257
rect 544 73209 548 73229
rect 579 73188 582 73278
rect 612 73260 624 73261
rect 599 73258 649 73260
rect 612 73257 624 73258
rect 610 73250 632 73257
rect 607 73249 632 73250
rect 586 73242 644 73249
rect 607 73241 644 73242
rect 607 73225 610 73241
rect 616 73225 644 73241
rect 607 73224 644 73225
rect 586 73217 644 73224
rect 607 73216 610 73217
rect 612 73209 632 73217
rect 612 73205 624 73209
rect 649 73208 651 73258
rect 544 73171 548 73179
rect 400 73139 408 73169
rect 420 73139 436 73169
rect 400 73135 436 73139
rect 400 73127 430 73135
rect 428 73111 430 73127
rect 476 73099 480 73167
rect 544 73137 552 73171
rect 578 73137 582 73171
rect 544 73129 548 73137
rect 544 73099 586 73100
rect 288 73059 292 73091
rect 296 73089 368 73097
rect 378 73089 450 73097
rect 544 73092 548 73099
rect 439 73061 444 73089
rect 120 73045 170 73047
rect 76 73041 130 73045
rect 110 73036 130 73041
rect 60 73011 67 73021
rect 76 73011 77 73031
rect 96 73002 99 73036
rect 109 73011 110 73031
rect 119 73011 126 73021
rect 76 72995 92 73001
rect 94 72995 110 73001
rect 170 72995 172 73045
rect 186 72979 190 73013
rect 216 72979 220 73013
rect 213 72947 224 72979
rect 282 72975 292 73059
rect 296 73053 368 73061
rect 378 73053 450 73061
rect 468 73058 473 73092
rect 428 73023 430 73039
rect 251 72947 292 72975
rect 318 72954 324 73023
rect 12 72942 62 72944
rect 28 72933 59 72941
rect 62 72933 64 72942
rect 251 72941 263 72947
rect 28 72925 64 72933
rect 127 72933 158 72941
rect 127 72926 182 72933
rect 127 72925 161 72926
rect 59 72909 64 72925
rect 158 72909 161 72925
rect 253 72913 263 72941
rect 273 72913 293 72947
rect 318 72944 335 72954
rect 303 72928 316 72938
rect 318 72928 324 72944
rect 346 72938 348 73023
rect 400 73015 430 73023
rect 476 73021 480 73089
rect 511 73058 582 73092
rect 544 73051 548 73058
rect 400 73011 436 73015
rect 400 72981 408 73011
rect 420 72981 436 73011
rect 544 73013 548 73021
rect 28 72901 64 72909
rect 127 72908 161 72909
rect 127 72901 182 72908
rect 62 72892 64 72901
rect 282 72855 292 72913
rect 295 72904 324 72928
rect 333 72928 353 72938
rect 428 72934 430 72981
rect 476 72941 480 73009
rect 544 72979 552 73013
rect 578 72979 582 73013
rect 544 72971 548 72979
rect 367 72928 380 72934
rect 333 72904 380 72928
rect 318 72891 324 72904
rect 346 72891 348 72904
rect 367 72900 380 72904
rect 396 72900 408 72934
rect 420 72900 436 72934
rect 544 72931 553 72959
rect 319 72880 346 72891
rect 120 72839 170 72841
rect 76 72833 92 72839
rect 94 72833 110 72839
rect 76 72823 99 72832
rect 60 72813 67 72823
rect 76 72803 77 72823
rect 96 72798 99 72823
rect 109 72803 110 72823
rect 119 72813 126 72823
rect 76 72789 110 72793
rect 170 72789 172 72839
rect 186 72821 190 72855
rect 216 72821 220 72855
rect 182 72783 224 72784
rect 186 72759 220 72776
rect 223 72759 257 72776
rect 182 72742 257 72759
rect 182 72741 224 72742
rect 160 72735 246 72741
rect 288 72735 292 72855
rect 296 72853 368 72861
rect 428 72853 430 72900
rect 476 72863 480 72931
rect 485 72887 495 72921
rect 505 72893 525 72921
rect 505 72887 519 72893
rect 544 72887 555 72931
rect 485 72863 492 72887
rect 579 72872 582 72962
rect 612 72944 624 72945
rect 599 72942 649 72944
rect 612 72941 624 72942
rect 610 72934 632 72941
rect 607 72933 632 72934
rect 586 72926 644 72933
rect 607 72925 644 72926
rect 607 72909 610 72925
rect 616 72909 644 72925
rect 607 72908 644 72909
rect 586 72901 644 72908
rect 607 72900 610 72901
rect 612 72893 632 72901
rect 612 72889 624 72893
rect 649 72892 651 72942
rect 544 72855 548 72863
rect 400 72823 408 72853
rect 420 72823 436 72853
rect 400 72819 436 72823
rect 400 72811 430 72819
rect 428 72795 430 72811
rect 476 72783 480 72851
rect 544 72821 552 72855
rect 578 72821 582 72855
rect 544 72813 548 72821
rect 295 72742 300 72776
rect 324 72742 329 72776
rect 378 72773 450 72781
rect 544 72778 548 72783
rect 544 72774 582 72778
rect 544 72759 552 72774
rect 578 72759 582 72774
rect 544 72741 586 72759
rect 522 72735 608 72741
rect 182 72719 224 72735
rect 544 72719 586 72735
rect 17 72705 67 72707
rect 119 72705 169 72707
rect 186 72705 220 72719
rect 548 72705 582 72719
rect 599 72705 649 72707
rect 42 72663 59 72697
rect 67 72655 69 72705
rect 160 72697 246 72705
rect 522 72697 608 72705
rect 76 72663 110 72697
rect 127 72663 144 72697
rect 152 72663 161 72697
rect 162 72695 195 72697
rect 224 72695 244 72697
rect 162 72663 244 72695
rect 524 72695 548 72697
rect 573 72695 582 72697
rect 586 72695 606 72697
rect 160 72655 246 72663
rect 186 72639 220 72655
rect 182 72625 224 72626
rect 160 72619 182 72625
rect 224 72619 246 72625
rect 186 72584 220 72618
rect 223 72584 257 72618
rect 120 72571 170 72573
rect 76 72567 130 72571
rect 110 72562 130 72567
rect 60 72537 67 72547
rect 76 72537 77 72557
rect 96 72528 99 72562
rect 109 72537 110 72557
rect 119 72537 126 72547
rect 76 72521 92 72527
rect 94 72521 110 72527
rect 170 72521 172 72571
rect 186 72505 190 72539
rect 216 72505 220 72539
rect 288 72505 292 72693
rect 476 72625 480 72693
rect 524 72663 606 72695
rect 607 72663 616 72697
rect 522 72655 608 72663
rect 649 72655 651 72705
rect 548 72639 582 72655
rect 522 72620 548 72625
rect 522 72619 582 72620
rect 586 72619 608 72625
rect 295 72584 300 72618
rect 324 72584 329 72618
rect 544 72616 582 72619
rect 378 72579 450 72587
rect 428 72549 430 72565
rect 400 72541 430 72549
rect 476 72547 480 72615
rect 544 72586 552 72616
rect 578 72586 582 72616
rect 544 72577 548 72586
rect 400 72537 436 72541
rect 400 72507 408 72537
rect 420 72507 436 72537
rect 544 72539 548 72547
rect 12 72468 62 72470
rect 28 72459 59 72467
rect 62 72459 64 72468
rect 28 72451 64 72459
rect 127 72459 158 72467
rect 127 72452 182 72459
rect 215 72457 224 72485
rect 127 72451 161 72452
rect 59 72435 64 72451
rect 158 72435 161 72451
rect 28 72427 64 72435
rect 127 72434 161 72435
rect 127 72427 182 72434
rect 62 72418 64 72427
rect 213 72419 224 72457
rect 282 72447 292 72505
rect 296 72499 368 72507
rect 319 72469 346 72480
rect 318 72456 324 72469
rect 346 72456 348 72469
rect 428 72460 430 72507
rect 443 72497 450 72499
rect 476 72467 480 72535
rect 544 72505 552 72539
rect 578 72505 582 72539
rect 481 72473 517 72501
rect 481 72467 495 72473
rect 367 72456 380 72460
rect 251 72413 263 72447
rect 273 72413 293 72447
rect 295 72432 324 72456
rect 303 72422 316 72432
rect 318 72416 324 72432
rect 333 72432 380 72456
rect 333 72422 353 72432
rect 367 72426 380 72432
rect 396 72426 408 72460
rect 420 72426 436 72460
rect 120 72365 170 72367
rect 76 72359 92 72365
rect 94 72359 110 72365
rect 76 72349 99 72358
rect 60 72339 67 72349
rect 76 72329 77 72349
rect 96 72324 99 72349
rect 109 72329 110 72349
rect 119 72339 126 72349
rect 76 72315 110 72319
rect 170 72315 172 72365
rect 186 72347 190 72381
rect 216 72347 220 72381
rect 186 72270 220 72304
rect 282 72301 292 72413
rect 318 72406 335 72416
rect 318 72337 324 72406
rect 346 72337 348 72422
rect 428 72379 430 72426
rect 476 72389 480 72457
rect 485 72439 495 72467
rect 505 72467 519 72473
rect 544 72467 555 72505
rect 505 72439 525 72467
rect 544 72439 553 72467
rect 544 72419 548 72439
rect 579 72398 582 72488
rect 612 72470 624 72471
rect 599 72468 649 72470
rect 612 72467 624 72468
rect 610 72460 632 72467
rect 607 72459 632 72460
rect 586 72452 644 72459
rect 607 72451 644 72452
rect 607 72435 610 72451
rect 616 72435 644 72451
rect 607 72434 644 72435
rect 586 72427 644 72434
rect 607 72426 610 72427
rect 612 72419 632 72427
rect 612 72415 624 72419
rect 649 72418 651 72468
rect 544 72381 548 72389
rect 400 72349 408 72379
rect 420 72349 436 72379
rect 400 72345 436 72349
rect 400 72337 430 72345
rect 428 72321 430 72337
rect 476 72309 480 72377
rect 544 72347 552 72381
rect 578 72347 582 72381
rect 544 72339 548 72347
rect 544 72309 586 72310
rect 288 72269 292 72301
rect 296 72299 368 72307
rect 378 72299 450 72307
rect 544 72302 548 72309
rect 439 72271 444 72299
rect 120 72255 170 72257
rect 76 72251 130 72255
rect 110 72246 130 72251
rect 60 72221 67 72231
rect 76 72221 77 72241
rect 96 72212 99 72246
rect 109 72221 110 72241
rect 119 72221 126 72231
rect 76 72205 92 72211
rect 94 72205 110 72211
rect 170 72205 172 72255
rect 186 72189 190 72223
rect 216 72189 220 72223
rect 213 72157 224 72189
rect 282 72185 292 72269
rect 296 72263 368 72271
rect 378 72263 450 72271
rect 468 72268 473 72302
rect 428 72233 430 72249
rect 251 72157 292 72185
rect 318 72164 324 72233
rect 12 72152 62 72154
rect 28 72143 59 72151
rect 62 72143 64 72152
rect 251 72151 263 72157
rect 28 72135 64 72143
rect 127 72143 158 72151
rect 127 72136 182 72143
rect 127 72135 161 72136
rect 59 72119 64 72135
rect 158 72119 161 72135
rect 253 72123 263 72151
rect 273 72123 293 72157
rect 318 72154 335 72164
rect 303 72138 316 72148
rect 318 72138 324 72154
rect 346 72148 348 72233
rect 400 72225 430 72233
rect 476 72231 480 72299
rect 511 72268 582 72302
rect 544 72261 548 72268
rect 400 72221 436 72225
rect 400 72191 408 72221
rect 420 72191 436 72221
rect 544 72223 548 72231
rect 28 72111 64 72119
rect 127 72118 161 72119
rect 127 72111 182 72118
rect 62 72102 64 72111
rect 282 72065 292 72123
rect 295 72114 324 72138
rect 333 72138 353 72148
rect 428 72144 430 72191
rect 476 72151 480 72219
rect 544 72189 552 72223
rect 578 72189 582 72223
rect 544 72181 548 72189
rect 367 72138 380 72144
rect 333 72114 380 72138
rect 318 72101 324 72114
rect 346 72101 348 72114
rect 367 72110 380 72114
rect 396 72110 408 72144
rect 420 72110 436 72144
rect 544 72141 553 72169
rect 319 72090 346 72101
rect 120 72049 170 72051
rect 76 72043 92 72049
rect 94 72043 110 72049
rect 76 72033 99 72042
rect 60 72023 67 72033
rect 76 72013 77 72033
rect 96 72008 99 72033
rect 109 72013 110 72033
rect 119 72023 126 72033
rect 76 71999 110 72003
rect 170 71999 172 72049
rect 186 72031 190 72065
rect 216 72031 220 72065
rect 182 71993 224 71994
rect 186 71969 220 71986
rect 223 71969 257 71986
rect 182 71952 257 71969
rect 182 71951 224 71952
rect 160 71945 246 71951
rect 288 71945 292 72065
rect 296 72063 368 72071
rect 428 72063 430 72110
rect 476 72073 480 72141
rect 485 72097 495 72131
rect 505 72103 525 72131
rect 505 72097 519 72103
rect 544 72097 555 72141
rect 485 72073 492 72097
rect 579 72082 582 72172
rect 612 72154 624 72155
rect 599 72152 649 72154
rect 612 72151 624 72152
rect 610 72144 632 72151
rect 607 72143 632 72144
rect 586 72136 644 72143
rect 607 72135 644 72136
rect 607 72119 610 72135
rect 616 72119 644 72135
rect 607 72118 644 72119
rect 586 72111 644 72118
rect 607 72110 610 72111
rect 612 72103 632 72111
rect 612 72099 624 72103
rect 649 72102 651 72152
rect 544 72065 548 72073
rect 400 72033 408 72063
rect 420 72033 436 72063
rect 400 72029 436 72033
rect 400 72021 430 72029
rect 428 72005 430 72021
rect 476 71993 480 72061
rect 544 72031 552 72065
rect 578 72031 582 72065
rect 544 72023 548 72031
rect 295 71952 300 71986
rect 324 71952 329 71986
rect 378 71983 450 71991
rect 544 71988 548 71993
rect 544 71984 582 71988
rect 544 71969 552 71984
rect 578 71969 582 71984
rect 544 71951 586 71969
rect 522 71945 608 71951
rect 182 71929 224 71945
rect 544 71929 586 71945
rect 17 71915 67 71917
rect 119 71915 169 71917
rect 186 71915 220 71929
rect 548 71915 582 71929
rect 599 71915 649 71917
rect 42 71873 59 71907
rect 67 71865 69 71915
rect 160 71907 246 71915
rect 522 71907 608 71915
rect 76 71873 110 71907
rect 127 71873 144 71907
rect 152 71873 161 71907
rect 162 71905 195 71907
rect 224 71905 244 71907
rect 162 71873 244 71905
rect 524 71905 548 71907
rect 573 71905 582 71907
rect 586 71905 606 71907
rect 160 71865 246 71873
rect 186 71849 220 71865
rect 182 71835 224 71836
rect 160 71829 182 71835
rect 224 71829 246 71835
rect 186 71794 220 71828
rect 223 71794 257 71828
rect 120 71781 170 71783
rect 76 71777 130 71781
rect 110 71772 130 71777
rect 60 71747 67 71757
rect 76 71747 77 71767
rect 96 71738 99 71772
rect 109 71747 110 71767
rect 119 71747 126 71757
rect 76 71731 92 71737
rect 94 71731 110 71737
rect 170 71731 172 71781
rect 186 71715 190 71749
rect 216 71715 220 71749
rect 288 71715 292 71903
rect 476 71835 480 71903
rect 524 71873 606 71905
rect 607 71873 616 71907
rect 522 71865 608 71873
rect 649 71865 651 71915
rect 548 71849 582 71865
rect 522 71830 548 71835
rect 522 71829 582 71830
rect 586 71829 608 71835
rect 295 71794 300 71828
rect 324 71794 329 71828
rect 544 71826 582 71829
rect 378 71789 450 71797
rect 428 71759 430 71775
rect 400 71751 430 71759
rect 476 71757 480 71825
rect 544 71796 552 71826
rect 578 71796 582 71826
rect 544 71787 548 71796
rect 400 71747 436 71751
rect 400 71717 408 71747
rect 420 71717 436 71747
rect 544 71749 548 71757
rect 12 71678 62 71680
rect 28 71669 59 71677
rect 62 71669 64 71678
rect 28 71661 64 71669
rect 127 71669 158 71677
rect 127 71662 182 71669
rect 215 71667 224 71695
rect 127 71661 161 71662
rect 59 71645 64 71661
rect 158 71645 161 71661
rect 28 71637 64 71645
rect 127 71644 161 71645
rect 127 71637 182 71644
rect 62 71628 64 71637
rect 213 71629 224 71667
rect 282 71657 292 71715
rect 296 71709 368 71717
rect 319 71679 346 71690
rect 318 71666 324 71679
rect 346 71666 348 71679
rect 428 71670 430 71717
rect 443 71707 450 71709
rect 476 71677 480 71745
rect 544 71715 552 71749
rect 578 71715 582 71749
rect 481 71683 517 71711
rect 481 71677 495 71683
rect 367 71666 380 71670
rect 251 71623 263 71657
rect 273 71623 293 71657
rect 295 71642 324 71666
rect 303 71632 316 71642
rect 318 71626 324 71642
rect 333 71642 380 71666
rect 333 71632 353 71642
rect 367 71636 380 71642
rect 396 71636 408 71670
rect 420 71636 436 71670
rect 120 71575 170 71577
rect 76 71569 92 71575
rect 94 71569 110 71575
rect 76 71559 99 71568
rect 60 71549 67 71559
rect 76 71539 77 71559
rect 96 71534 99 71559
rect 109 71539 110 71559
rect 119 71549 126 71559
rect 76 71525 110 71529
rect 170 71525 172 71575
rect 186 71557 190 71591
rect 216 71557 220 71591
rect 186 71480 220 71514
rect 282 71511 292 71623
rect 318 71616 335 71626
rect 318 71547 324 71616
rect 346 71547 348 71632
rect 428 71589 430 71636
rect 476 71599 480 71667
rect 485 71649 495 71677
rect 505 71677 519 71683
rect 544 71677 555 71715
rect 505 71649 525 71677
rect 544 71649 553 71677
rect 544 71629 548 71649
rect 579 71608 582 71698
rect 612 71680 624 71681
rect 599 71678 649 71680
rect 612 71677 624 71678
rect 610 71670 632 71677
rect 607 71669 632 71670
rect 586 71662 644 71669
rect 607 71661 644 71662
rect 607 71645 610 71661
rect 616 71645 644 71661
rect 607 71644 644 71645
rect 586 71637 644 71644
rect 607 71636 610 71637
rect 612 71629 632 71637
rect 612 71625 624 71629
rect 649 71628 651 71678
rect 544 71591 548 71599
rect 400 71559 408 71589
rect 420 71559 436 71589
rect 400 71555 436 71559
rect 400 71547 430 71555
rect 428 71531 430 71547
rect 476 71519 480 71587
rect 544 71557 552 71591
rect 578 71557 582 71591
rect 544 71549 548 71557
rect 544 71519 586 71520
rect 288 71479 292 71511
rect 296 71509 368 71517
rect 378 71509 450 71517
rect 544 71512 548 71519
rect 439 71481 444 71509
rect 120 71465 170 71467
rect 76 71461 130 71465
rect 110 71456 130 71461
rect 60 71431 67 71441
rect 76 71431 77 71451
rect 96 71422 99 71456
rect 109 71431 110 71451
rect 119 71431 126 71441
rect 76 71415 92 71421
rect 94 71415 110 71421
rect 170 71415 172 71465
rect 186 71399 190 71433
rect 216 71399 220 71433
rect 213 71367 224 71399
rect 282 71395 292 71479
rect 296 71473 368 71481
rect 378 71473 450 71481
rect 468 71478 473 71512
rect 428 71443 430 71459
rect 251 71367 292 71395
rect 318 71374 324 71443
rect 12 71362 62 71364
rect 28 71353 59 71361
rect 62 71353 64 71362
rect 251 71361 263 71367
rect 28 71345 64 71353
rect 127 71353 158 71361
rect 127 71346 182 71353
rect 127 71345 161 71346
rect 59 71329 64 71345
rect 158 71329 161 71345
rect 253 71333 263 71361
rect 273 71333 293 71367
rect 318 71364 335 71374
rect 303 71348 316 71358
rect 318 71348 324 71364
rect 346 71358 348 71443
rect 400 71435 430 71443
rect 476 71441 480 71509
rect 511 71478 582 71512
rect 544 71471 548 71478
rect 400 71431 436 71435
rect 400 71401 408 71431
rect 420 71401 436 71431
rect 544 71433 548 71441
rect 28 71321 64 71329
rect 127 71328 161 71329
rect 127 71321 182 71328
rect 62 71312 64 71321
rect 282 71275 292 71333
rect 295 71324 324 71348
rect 333 71348 353 71358
rect 428 71354 430 71401
rect 476 71361 480 71429
rect 544 71399 552 71433
rect 578 71399 582 71433
rect 544 71391 548 71399
rect 367 71348 380 71354
rect 333 71324 380 71348
rect 318 71311 324 71324
rect 346 71311 348 71324
rect 367 71320 380 71324
rect 396 71320 408 71354
rect 420 71320 436 71354
rect 544 71351 553 71379
rect 319 71300 346 71311
rect 120 71259 170 71261
rect 76 71253 92 71259
rect 94 71253 110 71259
rect 76 71243 99 71252
rect 60 71233 67 71243
rect 76 71223 77 71243
rect 96 71218 99 71243
rect 109 71223 110 71243
rect 119 71233 126 71243
rect 76 71209 110 71213
rect 170 71209 172 71259
rect 186 71241 190 71275
rect 216 71241 220 71275
rect 182 71203 224 71204
rect 186 71179 220 71196
rect 223 71179 257 71196
rect 182 71162 257 71179
rect 182 71161 224 71162
rect 160 71155 246 71161
rect 288 71155 292 71275
rect 296 71273 368 71281
rect 428 71273 430 71320
rect 476 71283 480 71351
rect 485 71307 495 71341
rect 505 71313 525 71341
rect 505 71307 519 71313
rect 544 71307 555 71351
rect 485 71283 492 71307
rect 579 71292 582 71382
rect 612 71364 624 71365
rect 599 71362 649 71364
rect 612 71361 624 71362
rect 610 71354 632 71361
rect 607 71353 632 71354
rect 586 71346 644 71353
rect 607 71345 644 71346
rect 607 71329 610 71345
rect 616 71329 644 71345
rect 607 71328 644 71329
rect 586 71321 644 71328
rect 607 71320 610 71321
rect 612 71313 632 71321
rect 612 71309 624 71313
rect 649 71312 651 71362
rect 544 71275 548 71283
rect 400 71243 408 71273
rect 420 71243 436 71273
rect 400 71239 436 71243
rect 400 71231 430 71239
rect 428 71215 430 71231
rect 476 71203 480 71271
rect 544 71241 552 71275
rect 578 71241 582 71275
rect 544 71233 548 71241
rect 295 71162 300 71196
rect 324 71162 329 71196
rect 378 71193 450 71201
rect 544 71198 548 71203
rect 544 71194 582 71198
rect 544 71179 552 71194
rect 578 71179 582 71194
rect 544 71161 586 71179
rect 522 71155 608 71161
rect 182 71139 224 71155
rect 544 71139 586 71155
rect 17 71125 67 71127
rect 119 71125 169 71127
rect 186 71125 220 71139
rect 548 71125 582 71139
rect 599 71125 649 71127
rect 42 71083 59 71117
rect 67 71075 69 71125
rect 160 71117 246 71125
rect 522 71117 608 71125
rect 76 71083 110 71117
rect 127 71083 144 71117
rect 152 71083 161 71117
rect 162 71115 195 71117
rect 224 71115 244 71117
rect 162 71083 244 71115
rect 524 71115 548 71117
rect 573 71115 582 71117
rect 586 71115 606 71117
rect 160 71075 246 71083
rect 186 71059 220 71075
rect 182 71045 224 71046
rect 160 71039 182 71045
rect 224 71039 246 71045
rect 186 71004 220 71038
rect 223 71004 257 71038
rect 120 70991 170 70993
rect 76 70987 130 70991
rect 110 70982 130 70987
rect 60 70957 67 70967
rect 76 70957 77 70977
rect 96 70948 99 70982
rect 109 70957 110 70977
rect 119 70957 126 70967
rect 76 70941 92 70947
rect 94 70941 110 70947
rect 170 70941 172 70991
rect 186 70925 190 70959
rect 216 70925 220 70959
rect 288 70925 292 71113
rect 476 71045 480 71113
rect 524 71083 606 71115
rect 607 71083 616 71117
rect 522 71075 608 71083
rect 649 71075 651 71125
rect 548 71059 582 71075
rect 522 71040 548 71045
rect 522 71039 582 71040
rect 586 71039 608 71045
rect 295 71004 300 71038
rect 324 71004 329 71038
rect 544 71036 582 71039
rect 378 70999 450 71007
rect 428 70969 430 70985
rect 400 70961 430 70969
rect 476 70967 480 71035
rect 544 71006 552 71036
rect 578 71006 582 71036
rect 544 70997 548 71006
rect 400 70957 436 70961
rect 400 70927 408 70957
rect 420 70927 436 70957
rect 544 70959 548 70967
rect 12 70888 62 70890
rect 28 70879 59 70887
rect 62 70879 64 70888
rect 28 70871 64 70879
rect 127 70879 158 70887
rect 127 70872 182 70879
rect 215 70877 224 70905
rect 127 70871 161 70872
rect 59 70855 64 70871
rect 158 70855 161 70871
rect 28 70847 64 70855
rect 127 70854 161 70855
rect 127 70847 182 70854
rect 62 70838 64 70847
rect 213 70839 224 70877
rect 282 70867 292 70925
rect 296 70919 368 70927
rect 319 70889 346 70900
rect 318 70876 324 70889
rect 346 70876 348 70889
rect 428 70880 430 70927
rect 443 70917 450 70919
rect 476 70887 480 70955
rect 544 70925 552 70959
rect 578 70925 582 70959
rect 481 70893 517 70921
rect 481 70887 495 70893
rect 367 70876 380 70880
rect 251 70833 263 70867
rect 273 70833 293 70867
rect 295 70852 324 70876
rect 303 70842 316 70852
rect 318 70836 324 70852
rect 333 70852 380 70876
rect 333 70842 353 70852
rect 367 70846 380 70852
rect 396 70846 408 70880
rect 420 70846 436 70880
rect 120 70785 170 70787
rect 76 70779 92 70785
rect 94 70779 110 70785
rect 76 70769 99 70778
rect 60 70759 67 70769
rect 76 70749 77 70769
rect 96 70744 99 70769
rect 109 70749 110 70769
rect 119 70759 126 70769
rect 76 70735 110 70739
rect 170 70735 172 70785
rect 186 70767 190 70801
rect 216 70767 220 70801
rect 186 70690 220 70724
rect 282 70721 292 70833
rect 318 70826 335 70836
rect 318 70757 324 70826
rect 346 70757 348 70842
rect 428 70799 430 70846
rect 476 70809 480 70877
rect 485 70859 495 70887
rect 505 70887 519 70893
rect 544 70887 555 70925
rect 505 70859 525 70887
rect 544 70859 553 70887
rect 544 70839 548 70859
rect 579 70818 582 70908
rect 612 70890 624 70891
rect 599 70888 649 70890
rect 612 70887 624 70888
rect 610 70880 632 70887
rect 607 70879 632 70880
rect 586 70872 644 70879
rect 607 70871 644 70872
rect 607 70855 610 70871
rect 616 70855 644 70871
rect 607 70854 644 70855
rect 586 70847 644 70854
rect 607 70846 610 70847
rect 612 70839 632 70847
rect 612 70835 624 70839
rect 649 70838 651 70888
rect 544 70801 548 70809
rect 400 70769 408 70799
rect 420 70769 436 70799
rect 400 70765 436 70769
rect 400 70757 430 70765
rect 428 70741 430 70757
rect 476 70729 480 70797
rect 544 70767 552 70801
rect 578 70767 582 70801
rect 544 70759 548 70767
rect 544 70729 586 70730
rect 288 70689 292 70721
rect 296 70719 368 70727
rect 378 70719 450 70727
rect 544 70722 548 70729
rect 439 70691 444 70719
rect 120 70675 170 70677
rect 76 70671 130 70675
rect 110 70666 130 70671
rect 60 70641 67 70651
rect 76 70641 77 70661
rect 96 70632 99 70666
rect 109 70641 110 70661
rect 119 70641 126 70651
rect 76 70625 92 70631
rect 94 70625 110 70631
rect 170 70625 172 70675
rect 186 70609 190 70643
rect 216 70609 220 70643
rect 213 70577 224 70609
rect 282 70605 292 70689
rect 296 70683 368 70691
rect 378 70683 450 70691
rect 468 70688 473 70722
rect 428 70653 430 70669
rect 251 70577 292 70605
rect 318 70584 324 70653
rect 12 70572 62 70574
rect 28 70563 59 70571
rect 62 70563 64 70572
rect 251 70571 263 70577
rect 28 70555 64 70563
rect 127 70563 158 70571
rect 127 70556 182 70563
rect 127 70555 161 70556
rect 59 70539 64 70555
rect 158 70539 161 70555
rect 253 70543 263 70571
rect 273 70543 293 70577
rect 318 70574 335 70584
rect 303 70558 316 70568
rect 318 70558 324 70574
rect 346 70568 348 70653
rect 400 70645 430 70653
rect 476 70651 480 70719
rect 511 70688 582 70722
rect 544 70681 548 70688
rect 400 70641 436 70645
rect 400 70611 408 70641
rect 420 70611 436 70641
rect 544 70643 548 70651
rect 28 70531 64 70539
rect 127 70538 161 70539
rect 127 70531 182 70538
rect 62 70522 64 70531
rect 282 70485 292 70543
rect 295 70534 324 70558
rect 333 70558 353 70568
rect 428 70564 430 70611
rect 476 70571 480 70639
rect 544 70609 552 70643
rect 578 70609 582 70643
rect 544 70601 548 70609
rect 367 70558 380 70564
rect 333 70534 380 70558
rect 318 70521 324 70534
rect 346 70521 348 70534
rect 367 70530 380 70534
rect 396 70530 408 70564
rect 420 70530 436 70564
rect 544 70561 553 70589
rect 319 70510 346 70521
rect 120 70469 170 70471
rect 76 70463 92 70469
rect 94 70463 110 70469
rect 76 70453 99 70462
rect 60 70443 67 70453
rect 76 70433 77 70453
rect 96 70428 99 70453
rect 109 70433 110 70453
rect 119 70443 126 70453
rect 76 70419 110 70423
rect 170 70419 172 70469
rect 186 70451 190 70485
rect 216 70451 220 70485
rect 182 70413 224 70414
rect 186 70389 220 70406
rect 223 70389 257 70406
rect 182 70372 257 70389
rect 182 70371 224 70372
rect 160 70365 246 70371
rect 288 70365 292 70485
rect 296 70483 368 70491
rect 428 70483 430 70530
rect 476 70493 480 70561
rect 485 70517 495 70551
rect 505 70523 525 70551
rect 505 70517 519 70523
rect 544 70517 555 70561
rect 485 70493 492 70517
rect 579 70502 582 70592
rect 612 70574 624 70575
rect 599 70572 649 70574
rect 612 70571 624 70572
rect 610 70564 632 70571
rect 607 70563 632 70564
rect 586 70556 644 70563
rect 607 70555 644 70556
rect 607 70539 610 70555
rect 616 70539 644 70555
rect 607 70538 644 70539
rect 586 70531 644 70538
rect 607 70530 610 70531
rect 612 70523 632 70531
rect 612 70519 624 70523
rect 649 70522 651 70572
rect 544 70485 548 70493
rect 400 70453 408 70483
rect 420 70453 436 70483
rect 400 70449 436 70453
rect 400 70441 430 70449
rect 428 70425 430 70441
rect 476 70413 480 70481
rect 544 70451 552 70485
rect 578 70451 582 70485
rect 544 70443 548 70451
rect 295 70372 300 70406
rect 324 70372 329 70406
rect 378 70403 450 70411
rect 544 70408 548 70413
rect 544 70404 582 70408
rect 544 70389 552 70404
rect 578 70389 582 70404
rect 544 70371 586 70389
rect 522 70365 608 70371
rect 182 70349 224 70365
rect 544 70349 586 70365
rect 17 70335 67 70337
rect 119 70335 169 70337
rect 186 70335 220 70349
rect 548 70335 582 70349
rect 599 70335 649 70337
rect 42 70293 59 70327
rect 67 70285 69 70335
rect 160 70327 246 70335
rect 522 70327 608 70335
rect 76 70293 110 70327
rect 127 70293 144 70327
rect 152 70293 161 70327
rect 162 70325 195 70327
rect 224 70325 244 70327
rect 162 70293 244 70325
rect 524 70325 548 70327
rect 573 70325 582 70327
rect 586 70325 606 70327
rect 160 70285 246 70293
rect 186 70269 220 70285
rect 182 70255 224 70256
rect 160 70249 182 70255
rect 224 70249 246 70255
rect 186 70214 220 70248
rect 223 70214 257 70248
rect 120 70201 170 70203
rect 76 70197 130 70201
rect 110 70192 130 70197
rect 60 70167 67 70177
rect 76 70167 77 70187
rect 96 70158 99 70192
rect 109 70167 110 70187
rect 119 70167 126 70177
rect 76 70151 92 70157
rect 94 70151 110 70157
rect 170 70151 172 70201
rect 186 70135 190 70169
rect 216 70135 220 70169
rect 288 70135 292 70323
rect 476 70255 480 70323
rect 524 70293 606 70325
rect 607 70293 616 70327
rect 522 70285 608 70293
rect 649 70285 651 70335
rect 548 70269 582 70285
rect 522 70250 548 70255
rect 522 70249 582 70250
rect 586 70249 608 70255
rect 295 70214 300 70248
rect 324 70214 329 70248
rect 544 70246 582 70249
rect 378 70209 450 70217
rect 428 70179 430 70195
rect 400 70171 430 70179
rect 476 70177 480 70245
rect 544 70216 552 70246
rect 578 70216 582 70246
rect 544 70207 548 70216
rect 400 70167 436 70171
rect 400 70137 408 70167
rect 420 70137 436 70167
rect 544 70169 548 70177
rect 12 70098 62 70100
rect 28 70089 59 70097
rect 62 70089 64 70098
rect 28 70081 64 70089
rect 127 70089 158 70097
rect 127 70082 182 70089
rect 215 70087 224 70115
rect 127 70081 161 70082
rect 59 70065 64 70081
rect 158 70065 161 70081
rect 28 70057 64 70065
rect 127 70064 161 70065
rect 127 70057 182 70064
rect 62 70048 64 70057
rect 213 70049 224 70087
rect 282 70077 292 70135
rect 296 70129 368 70137
rect 319 70099 346 70110
rect 318 70086 324 70099
rect 346 70086 348 70099
rect 428 70090 430 70137
rect 443 70127 450 70129
rect 476 70097 480 70165
rect 544 70135 552 70169
rect 578 70135 582 70169
rect 481 70103 517 70131
rect 481 70097 495 70103
rect 367 70086 380 70090
rect 251 70043 263 70077
rect 273 70043 293 70077
rect 295 70062 324 70086
rect 303 70052 316 70062
rect 318 70046 324 70062
rect 333 70062 380 70086
rect 333 70052 353 70062
rect 367 70056 380 70062
rect 396 70056 408 70090
rect 420 70056 436 70090
rect 120 69995 170 69997
rect 76 69989 92 69995
rect 94 69989 110 69995
rect 76 69979 99 69988
rect 60 69969 67 69979
rect 76 69959 77 69979
rect 96 69954 99 69979
rect 109 69959 110 69979
rect 119 69969 126 69979
rect 76 69945 110 69949
rect 170 69945 172 69995
rect 186 69977 190 70011
rect 216 69977 220 70011
rect 186 69900 220 69934
rect 282 69931 292 70043
rect 318 70036 335 70046
rect 318 69967 324 70036
rect 346 69967 348 70052
rect 428 70009 430 70056
rect 476 70019 480 70087
rect 485 70069 495 70097
rect 505 70097 519 70103
rect 544 70097 555 70135
rect 505 70069 525 70097
rect 544 70069 553 70097
rect 544 70049 548 70069
rect 579 70028 582 70118
rect 612 70100 624 70101
rect 599 70098 649 70100
rect 612 70097 624 70098
rect 610 70090 632 70097
rect 607 70089 632 70090
rect 586 70082 644 70089
rect 607 70081 644 70082
rect 607 70065 610 70081
rect 616 70065 644 70081
rect 607 70064 644 70065
rect 586 70057 644 70064
rect 607 70056 610 70057
rect 612 70049 632 70057
rect 612 70045 624 70049
rect 649 70048 651 70098
rect 544 70011 548 70019
rect 400 69979 408 70009
rect 420 69979 436 70009
rect 400 69975 436 69979
rect 400 69967 430 69975
rect 428 69951 430 69967
rect 476 69939 480 70007
rect 544 69977 552 70011
rect 578 69977 582 70011
rect 544 69969 548 69977
rect 544 69939 586 69940
rect 288 69899 292 69931
rect 296 69929 368 69937
rect 378 69929 450 69937
rect 544 69932 548 69939
rect 439 69901 444 69929
rect 120 69885 170 69887
rect 76 69881 130 69885
rect 110 69876 130 69881
rect 60 69851 67 69861
rect 76 69851 77 69871
rect 96 69842 99 69876
rect 109 69851 110 69871
rect 119 69851 126 69861
rect 76 69835 92 69841
rect 94 69835 110 69841
rect 170 69835 172 69885
rect 186 69819 190 69853
rect 216 69819 220 69853
rect 213 69787 224 69819
rect 282 69815 292 69899
rect 296 69893 368 69901
rect 378 69893 450 69901
rect 468 69898 473 69932
rect 428 69863 430 69879
rect 251 69787 292 69815
rect 318 69794 324 69863
rect 12 69782 62 69784
rect 28 69773 59 69781
rect 62 69773 64 69782
rect 251 69781 263 69787
rect 28 69765 64 69773
rect 127 69773 158 69781
rect 127 69766 182 69773
rect 127 69765 161 69766
rect 59 69749 64 69765
rect 158 69749 161 69765
rect 253 69753 263 69781
rect 273 69753 293 69787
rect 318 69784 335 69794
rect 303 69768 316 69778
rect 318 69768 324 69784
rect 346 69778 348 69863
rect 400 69855 430 69863
rect 476 69861 480 69929
rect 511 69898 582 69932
rect 544 69891 548 69898
rect 400 69851 436 69855
rect 400 69821 408 69851
rect 420 69821 436 69851
rect 544 69853 548 69861
rect 28 69741 64 69749
rect 127 69748 161 69749
rect 127 69741 182 69748
rect 62 69732 64 69741
rect 282 69695 292 69753
rect 295 69744 324 69768
rect 333 69768 353 69778
rect 428 69774 430 69821
rect 476 69781 480 69849
rect 544 69819 552 69853
rect 578 69819 582 69853
rect 544 69811 548 69819
rect 367 69768 380 69774
rect 333 69744 380 69768
rect 318 69731 324 69744
rect 346 69731 348 69744
rect 367 69740 380 69744
rect 396 69740 408 69774
rect 420 69740 436 69774
rect 544 69771 553 69799
rect 319 69720 346 69731
rect 120 69679 170 69681
rect 76 69673 92 69679
rect 94 69673 110 69679
rect 76 69663 99 69672
rect 60 69653 67 69663
rect 76 69643 77 69663
rect 96 69638 99 69663
rect 109 69643 110 69663
rect 119 69653 126 69663
rect 76 69629 110 69633
rect 170 69629 172 69679
rect 186 69661 190 69695
rect 216 69661 220 69695
rect 182 69623 224 69624
rect 186 69599 220 69616
rect 223 69599 257 69616
rect 182 69582 257 69599
rect 182 69581 224 69582
rect 160 69575 246 69581
rect 288 69575 292 69695
rect 296 69693 368 69701
rect 428 69693 430 69740
rect 476 69703 480 69771
rect 485 69727 495 69761
rect 505 69733 525 69761
rect 505 69727 519 69733
rect 544 69727 555 69771
rect 485 69703 492 69727
rect 579 69712 582 69802
rect 612 69784 624 69785
rect 599 69782 649 69784
rect 612 69781 624 69782
rect 610 69774 632 69781
rect 607 69773 632 69774
rect 586 69766 644 69773
rect 607 69765 644 69766
rect 607 69749 610 69765
rect 616 69749 644 69765
rect 607 69748 644 69749
rect 586 69741 644 69748
rect 607 69740 610 69741
rect 612 69733 632 69741
rect 612 69729 624 69733
rect 649 69732 651 69782
rect 544 69695 548 69703
rect 400 69663 408 69693
rect 420 69663 436 69693
rect 400 69659 436 69663
rect 400 69651 430 69659
rect 428 69635 430 69651
rect 476 69623 480 69691
rect 544 69661 552 69695
rect 578 69661 582 69695
rect 544 69653 548 69661
rect 295 69582 300 69616
rect 324 69582 329 69616
rect 378 69613 450 69621
rect 544 69618 548 69623
rect 544 69614 582 69618
rect 544 69599 552 69614
rect 578 69599 582 69614
rect 544 69581 586 69599
rect 522 69575 608 69581
rect 182 69559 224 69575
rect 544 69559 586 69575
rect 17 69545 67 69547
rect 119 69545 169 69547
rect 186 69545 220 69559
rect 548 69545 582 69559
rect 599 69545 649 69547
rect 42 69503 59 69537
rect 67 69495 69 69545
rect 160 69537 246 69545
rect 522 69537 608 69545
rect 76 69503 110 69537
rect 127 69503 144 69537
rect 152 69503 161 69537
rect 162 69535 195 69537
rect 224 69535 244 69537
rect 162 69503 244 69535
rect 524 69535 548 69537
rect 573 69535 582 69537
rect 586 69535 606 69537
rect 160 69495 246 69503
rect 186 69479 220 69495
rect 182 69465 224 69466
rect 160 69459 182 69465
rect 224 69459 246 69465
rect 186 69424 220 69458
rect 223 69424 257 69458
rect 120 69411 170 69413
rect 76 69407 130 69411
rect 110 69402 130 69407
rect 60 69377 67 69387
rect 76 69377 77 69397
rect 96 69368 99 69402
rect 109 69377 110 69397
rect 119 69377 126 69387
rect 76 69361 92 69367
rect 94 69361 110 69367
rect 170 69361 172 69411
rect 186 69345 190 69379
rect 216 69345 220 69379
rect 288 69345 292 69533
rect 476 69465 480 69533
rect 524 69503 606 69535
rect 607 69503 616 69537
rect 522 69495 608 69503
rect 649 69495 651 69545
rect 548 69479 582 69495
rect 522 69460 548 69465
rect 522 69459 582 69460
rect 586 69459 608 69465
rect 295 69424 300 69458
rect 324 69424 329 69458
rect 544 69456 582 69459
rect 378 69419 450 69427
rect 428 69389 430 69405
rect 400 69381 430 69389
rect 476 69387 480 69455
rect 544 69426 552 69456
rect 578 69426 582 69456
rect 544 69417 548 69426
rect 400 69377 436 69381
rect 400 69347 408 69377
rect 420 69347 436 69377
rect 544 69379 548 69387
rect 12 69308 62 69310
rect 28 69299 59 69307
rect 62 69299 64 69308
rect 28 69291 64 69299
rect 127 69299 158 69307
rect 127 69292 182 69299
rect 215 69297 224 69325
rect 127 69291 161 69292
rect 59 69275 64 69291
rect 158 69275 161 69291
rect 28 69267 64 69275
rect 127 69274 161 69275
rect 127 69267 182 69274
rect 62 69258 64 69267
rect 213 69259 224 69297
rect 282 69287 292 69345
rect 296 69339 368 69347
rect 319 69309 346 69320
rect 318 69296 324 69309
rect 346 69296 348 69309
rect 428 69300 430 69347
rect 443 69337 450 69339
rect 476 69307 480 69375
rect 544 69345 552 69379
rect 578 69345 582 69379
rect 481 69313 517 69341
rect 481 69307 495 69313
rect 367 69296 380 69300
rect 251 69253 263 69287
rect 273 69253 293 69287
rect 295 69272 324 69296
rect 303 69262 316 69272
rect 318 69256 324 69272
rect 333 69272 380 69296
rect 333 69262 353 69272
rect 367 69266 380 69272
rect 396 69266 408 69300
rect 420 69266 436 69300
rect 120 69205 170 69207
rect 76 69199 92 69205
rect 94 69199 110 69205
rect 76 69189 99 69198
rect 60 69179 67 69189
rect 76 69169 77 69189
rect 96 69164 99 69189
rect 109 69169 110 69189
rect 119 69179 126 69189
rect 76 69155 110 69159
rect 170 69155 172 69205
rect 186 69187 190 69221
rect 216 69187 220 69221
rect 186 69110 220 69144
rect 282 69141 292 69253
rect 318 69246 335 69256
rect 318 69177 324 69246
rect 346 69177 348 69262
rect 428 69219 430 69266
rect 476 69229 480 69297
rect 485 69279 495 69307
rect 505 69307 519 69313
rect 544 69307 555 69345
rect 505 69279 525 69307
rect 544 69279 553 69307
rect 544 69259 548 69279
rect 579 69238 582 69328
rect 612 69310 624 69311
rect 599 69308 649 69310
rect 612 69307 624 69308
rect 610 69300 632 69307
rect 607 69299 632 69300
rect 586 69292 644 69299
rect 607 69291 644 69292
rect 607 69275 610 69291
rect 616 69275 644 69291
rect 607 69274 644 69275
rect 586 69267 644 69274
rect 607 69266 610 69267
rect 612 69259 632 69267
rect 612 69255 624 69259
rect 649 69258 651 69308
rect 544 69221 548 69229
rect 400 69189 408 69219
rect 420 69189 436 69219
rect 400 69185 436 69189
rect 400 69177 430 69185
rect 428 69161 430 69177
rect 476 69149 480 69217
rect 544 69187 552 69221
rect 578 69187 582 69221
rect 544 69179 548 69187
rect 544 69149 586 69150
rect 288 69109 292 69141
rect 296 69139 368 69147
rect 378 69139 450 69147
rect 544 69142 548 69149
rect 439 69111 444 69139
rect 120 69095 170 69097
rect 76 69091 130 69095
rect 110 69086 130 69091
rect 60 69061 67 69071
rect 76 69061 77 69081
rect 96 69052 99 69086
rect 109 69061 110 69081
rect 119 69061 126 69071
rect 76 69045 92 69051
rect 94 69045 110 69051
rect 170 69045 172 69095
rect 186 69029 190 69063
rect 216 69029 220 69063
rect 213 68997 224 69029
rect 282 69025 292 69109
rect 296 69103 368 69111
rect 378 69103 450 69111
rect 468 69108 473 69142
rect 428 69073 430 69089
rect 251 68997 292 69025
rect 318 69004 324 69073
rect 12 68992 62 68994
rect 28 68983 59 68991
rect 62 68983 64 68992
rect 251 68991 263 68997
rect 28 68975 64 68983
rect 127 68983 158 68991
rect 127 68976 182 68983
rect 127 68975 161 68976
rect 59 68959 64 68975
rect 158 68959 161 68975
rect 253 68963 263 68991
rect 273 68963 293 68997
rect 318 68994 335 69004
rect 303 68978 316 68988
rect 318 68978 324 68994
rect 346 68988 348 69073
rect 400 69065 430 69073
rect 476 69071 480 69139
rect 511 69108 582 69142
rect 544 69101 548 69108
rect 400 69061 436 69065
rect 400 69031 408 69061
rect 420 69031 436 69061
rect 544 69063 548 69071
rect 28 68951 64 68959
rect 127 68958 161 68959
rect 127 68951 182 68958
rect 62 68942 64 68951
rect 282 68905 292 68963
rect 295 68954 324 68978
rect 333 68978 353 68988
rect 428 68984 430 69031
rect 476 68991 480 69059
rect 544 69029 552 69063
rect 578 69029 582 69063
rect 544 69021 548 69029
rect 367 68978 380 68984
rect 333 68954 380 68978
rect 318 68941 324 68954
rect 346 68941 348 68954
rect 367 68950 380 68954
rect 396 68950 408 68984
rect 420 68950 436 68984
rect 544 68981 553 69009
rect 319 68930 346 68941
rect 120 68889 170 68891
rect 76 68883 92 68889
rect 94 68883 110 68889
rect 76 68873 99 68882
rect 60 68863 67 68873
rect 76 68853 77 68873
rect 96 68848 99 68873
rect 109 68853 110 68873
rect 119 68863 126 68873
rect 76 68839 110 68843
rect 170 68839 172 68889
rect 186 68871 190 68905
rect 216 68871 220 68905
rect 182 68833 224 68834
rect 186 68809 220 68826
rect 223 68809 257 68826
rect 182 68792 257 68809
rect 182 68791 224 68792
rect 160 68785 246 68791
rect 288 68785 292 68905
rect 296 68903 368 68911
rect 428 68903 430 68950
rect 476 68913 480 68981
rect 485 68937 495 68971
rect 505 68943 525 68971
rect 505 68937 519 68943
rect 544 68937 555 68981
rect 485 68913 492 68937
rect 579 68922 582 69012
rect 612 68994 624 68995
rect 599 68992 649 68994
rect 612 68991 624 68992
rect 610 68984 632 68991
rect 607 68983 632 68984
rect 586 68976 644 68983
rect 607 68975 644 68976
rect 607 68959 610 68975
rect 616 68959 644 68975
rect 607 68958 644 68959
rect 586 68951 644 68958
rect 607 68950 610 68951
rect 612 68943 632 68951
rect 612 68939 624 68943
rect 649 68942 651 68992
rect 544 68905 548 68913
rect 400 68873 408 68903
rect 420 68873 436 68903
rect 400 68869 436 68873
rect 400 68861 430 68869
rect 428 68845 430 68861
rect 476 68833 480 68901
rect 544 68871 552 68905
rect 578 68871 582 68905
rect 544 68863 548 68871
rect 295 68792 300 68826
rect 324 68792 329 68826
rect 378 68823 450 68831
rect 544 68828 548 68833
rect 544 68824 582 68828
rect 544 68809 552 68824
rect 578 68809 582 68824
rect 544 68791 586 68809
rect 522 68785 608 68791
rect 182 68769 224 68785
rect 544 68769 586 68785
rect 17 68755 67 68757
rect 119 68755 169 68757
rect 186 68755 220 68769
rect 548 68755 582 68769
rect 599 68755 649 68757
rect 42 68713 59 68747
rect 67 68705 69 68755
rect 160 68747 246 68755
rect 522 68747 608 68755
rect 76 68713 110 68747
rect 127 68713 144 68747
rect 152 68713 161 68747
rect 162 68745 195 68747
rect 224 68745 244 68747
rect 162 68713 244 68745
rect 524 68745 548 68747
rect 573 68745 582 68747
rect 586 68745 606 68747
rect 160 68705 246 68713
rect 186 68689 220 68705
rect 182 68675 224 68676
rect 160 68669 182 68675
rect 224 68669 246 68675
rect 186 68634 220 68668
rect 223 68634 257 68668
rect 120 68621 170 68623
rect 76 68617 130 68621
rect 110 68612 130 68617
rect 60 68587 67 68597
rect 76 68587 77 68607
rect 96 68578 99 68612
rect 109 68587 110 68607
rect 119 68587 126 68597
rect 76 68571 92 68577
rect 94 68571 110 68577
rect 170 68571 172 68621
rect 186 68555 190 68589
rect 216 68555 220 68589
rect 288 68555 292 68743
rect 476 68675 480 68743
rect 524 68713 606 68745
rect 607 68713 616 68747
rect 522 68705 608 68713
rect 649 68705 651 68755
rect 548 68689 582 68705
rect 522 68670 548 68675
rect 522 68669 582 68670
rect 586 68669 608 68675
rect 295 68634 300 68668
rect 324 68634 329 68668
rect 544 68666 582 68669
rect 378 68629 450 68637
rect 428 68599 430 68615
rect 400 68591 430 68599
rect 476 68597 480 68665
rect 544 68636 552 68666
rect 578 68636 582 68666
rect 544 68627 548 68636
rect 400 68587 436 68591
rect 400 68557 408 68587
rect 420 68557 436 68587
rect 544 68589 548 68597
rect 12 68518 62 68520
rect 28 68509 59 68517
rect 62 68509 64 68518
rect 28 68501 64 68509
rect 127 68509 158 68517
rect 127 68502 182 68509
rect 215 68507 224 68535
rect 127 68501 161 68502
rect 59 68485 64 68501
rect 158 68485 161 68501
rect 28 68477 64 68485
rect 127 68484 161 68485
rect 127 68477 182 68484
rect 62 68468 64 68477
rect 213 68469 224 68507
rect 282 68497 292 68555
rect 296 68549 368 68557
rect 319 68519 346 68530
rect 318 68506 324 68519
rect 346 68506 348 68519
rect 428 68510 430 68557
rect 443 68547 450 68549
rect 476 68517 480 68585
rect 544 68555 552 68589
rect 578 68555 582 68589
rect 481 68523 517 68551
rect 481 68517 495 68523
rect 367 68506 380 68510
rect 251 68463 263 68497
rect 273 68463 293 68497
rect 295 68482 324 68506
rect 303 68472 316 68482
rect 318 68466 324 68482
rect 333 68482 380 68506
rect 333 68472 353 68482
rect 367 68476 380 68482
rect 396 68476 408 68510
rect 420 68476 436 68510
rect 120 68415 170 68417
rect 76 68409 92 68415
rect 94 68409 110 68415
rect 76 68399 99 68408
rect 60 68389 67 68399
rect 76 68379 77 68399
rect 96 68374 99 68399
rect 109 68379 110 68399
rect 119 68389 126 68399
rect 76 68365 110 68369
rect 170 68365 172 68415
rect 186 68397 190 68431
rect 216 68397 220 68431
rect 186 68320 220 68354
rect 282 68351 292 68463
rect 318 68456 335 68466
rect 318 68387 324 68456
rect 346 68387 348 68472
rect 428 68429 430 68476
rect 476 68439 480 68507
rect 485 68489 495 68517
rect 505 68517 519 68523
rect 544 68517 555 68555
rect 505 68489 525 68517
rect 544 68489 553 68517
rect 544 68469 548 68489
rect 579 68448 582 68538
rect 612 68520 624 68521
rect 599 68518 649 68520
rect 612 68517 624 68518
rect 610 68510 632 68517
rect 607 68509 632 68510
rect 586 68502 644 68509
rect 607 68501 644 68502
rect 607 68485 610 68501
rect 616 68485 644 68501
rect 607 68484 644 68485
rect 586 68477 644 68484
rect 607 68476 610 68477
rect 612 68469 632 68477
rect 612 68465 624 68469
rect 649 68468 651 68518
rect 544 68431 548 68439
rect 400 68399 408 68429
rect 420 68399 436 68429
rect 400 68395 436 68399
rect 400 68387 430 68395
rect 428 68371 430 68387
rect 476 68359 480 68427
rect 544 68397 552 68431
rect 578 68397 582 68431
rect 544 68389 548 68397
rect 544 68359 586 68360
rect 288 68319 292 68351
rect 296 68349 368 68357
rect 378 68349 450 68357
rect 544 68352 548 68359
rect 439 68321 444 68349
rect 120 68305 170 68307
rect 76 68301 130 68305
rect 110 68296 130 68301
rect 60 68271 67 68281
rect 76 68271 77 68291
rect 96 68262 99 68296
rect 109 68271 110 68291
rect 119 68271 126 68281
rect 76 68255 92 68261
rect 94 68255 110 68261
rect 170 68255 172 68305
rect 186 68239 190 68273
rect 216 68239 220 68273
rect 213 68207 224 68239
rect 282 68235 292 68319
rect 296 68313 368 68321
rect 378 68313 450 68321
rect 468 68318 473 68352
rect 428 68283 430 68299
rect 251 68207 292 68235
rect 318 68214 324 68283
rect 12 68202 62 68204
rect 28 68193 59 68201
rect 62 68193 64 68202
rect 251 68201 263 68207
rect 28 68185 64 68193
rect 127 68193 158 68201
rect 127 68186 182 68193
rect 127 68185 161 68186
rect 59 68169 64 68185
rect 158 68169 161 68185
rect 253 68173 263 68201
rect 273 68173 293 68207
rect 318 68204 335 68214
rect 303 68188 316 68198
rect 318 68188 324 68204
rect 346 68198 348 68283
rect 400 68275 430 68283
rect 476 68281 480 68349
rect 511 68318 582 68352
rect 544 68311 548 68318
rect 400 68271 436 68275
rect 400 68241 408 68271
rect 420 68241 436 68271
rect 544 68273 548 68281
rect 28 68161 64 68169
rect 127 68168 161 68169
rect 127 68161 182 68168
rect 62 68152 64 68161
rect 282 68115 292 68173
rect 295 68164 324 68188
rect 333 68188 353 68198
rect 428 68194 430 68241
rect 476 68201 480 68269
rect 544 68239 552 68273
rect 578 68239 582 68273
rect 544 68231 548 68239
rect 367 68188 380 68194
rect 333 68164 380 68188
rect 318 68151 324 68164
rect 346 68151 348 68164
rect 367 68160 380 68164
rect 396 68160 408 68194
rect 420 68160 436 68194
rect 544 68191 553 68219
rect 319 68140 346 68151
rect 120 68099 170 68101
rect 76 68093 92 68099
rect 94 68093 110 68099
rect 76 68083 99 68092
rect 60 68073 67 68083
rect 76 68063 77 68083
rect 96 68058 99 68083
rect 109 68063 110 68083
rect 119 68073 126 68083
rect 76 68049 110 68053
rect 170 68049 172 68099
rect 186 68081 190 68115
rect 216 68081 220 68115
rect 182 68043 224 68044
rect 186 68019 220 68036
rect 223 68019 257 68036
rect 182 68002 257 68019
rect 182 68001 224 68002
rect 160 67995 246 68001
rect 288 67995 292 68115
rect 296 68113 368 68121
rect 428 68113 430 68160
rect 476 68123 480 68191
rect 485 68147 495 68181
rect 505 68153 525 68181
rect 505 68147 519 68153
rect 544 68147 555 68191
rect 485 68123 492 68147
rect 579 68132 582 68222
rect 612 68204 624 68205
rect 599 68202 649 68204
rect 612 68201 624 68202
rect 610 68194 632 68201
rect 607 68193 632 68194
rect 586 68186 644 68193
rect 607 68185 644 68186
rect 607 68169 610 68185
rect 616 68169 644 68185
rect 607 68168 644 68169
rect 586 68161 644 68168
rect 607 68160 610 68161
rect 612 68153 632 68161
rect 612 68149 624 68153
rect 649 68152 651 68202
rect 544 68115 548 68123
rect 400 68083 408 68113
rect 420 68083 436 68113
rect 400 68079 436 68083
rect 400 68071 430 68079
rect 428 68055 430 68071
rect 476 68043 480 68111
rect 544 68081 552 68115
rect 578 68081 582 68115
rect 544 68073 548 68081
rect 295 68002 300 68036
rect 324 68002 329 68036
rect 378 68033 450 68041
rect 544 68038 548 68043
rect 544 68034 582 68038
rect 544 68019 552 68034
rect 578 68019 582 68034
rect 544 68001 586 68019
rect 522 67995 608 68001
rect 182 67979 224 67995
rect 544 67979 586 67995
rect 17 67965 67 67967
rect 119 67965 169 67967
rect 186 67965 220 67979
rect 548 67965 582 67979
rect 599 67965 649 67967
rect 42 67923 59 67957
rect 67 67915 69 67965
rect 160 67957 246 67965
rect 522 67957 608 67965
rect 76 67923 110 67957
rect 127 67923 144 67957
rect 152 67923 161 67957
rect 162 67955 195 67957
rect 224 67955 244 67957
rect 162 67923 244 67955
rect 524 67955 548 67957
rect 573 67955 582 67957
rect 586 67955 606 67957
rect 160 67915 246 67923
rect 186 67899 220 67915
rect 182 67885 224 67886
rect 160 67879 182 67885
rect 224 67879 246 67885
rect 186 67844 220 67878
rect 223 67844 257 67878
rect 120 67831 170 67833
rect 76 67827 130 67831
rect 110 67822 130 67827
rect 60 67797 67 67807
rect 76 67797 77 67817
rect 96 67788 99 67822
rect 109 67797 110 67817
rect 119 67797 126 67807
rect 76 67781 92 67787
rect 94 67781 110 67787
rect 170 67781 172 67831
rect 186 67765 190 67799
rect 216 67765 220 67799
rect 288 67765 292 67953
rect 476 67885 480 67953
rect 524 67923 606 67955
rect 607 67923 616 67957
rect 522 67915 608 67923
rect 649 67915 651 67965
rect 548 67899 582 67915
rect 522 67880 548 67885
rect 522 67879 582 67880
rect 586 67879 608 67885
rect 295 67844 300 67878
rect 324 67844 329 67878
rect 544 67876 582 67879
rect 378 67839 450 67847
rect 428 67809 430 67825
rect 400 67801 430 67809
rect 476 67807 480 67875
rect 544 67846 552 67876
rect 578 67846 582 67876
rect 544 67837 548 67846
rect 400 67797 436 67801
rect 400 67767 408 67797
rect 420 67767 436 67797
rect 544 67799 548 67807
rect 12 67728 62 67730
rect 28 67719 59 67727
rect 62 67719 64 67728
rect 28 67711 64 67719
rect 127 67719 158 67727
rect 127 67712 182 67719
rect 215 67717 224 67745
rect 127 67711 161 67712
rect 59 67695 64 67711
rect 158 67695 161 67711
rect 28 67687 64 67695
rect 127 67694 161 67695
rect 127 67687 182 67694
rect 62 67678 64 67687
rect 213 67679 224 67717
rect 282 67707 292 67765
rect 296 67759 368 67767
rect 319 67729 346 67740
rect 318 67716 324 67729
rect 346 67716 348 67729
rect 428 67720 430 67767
rect 443 67757 450 67759
rect 476 67727 480 67795
rect 544 67765 552 67799
rect 578 67765 582 67799
rect 481 67733 517 67761
rect 481 67727 495 67733
rect 367 67716 380 67720
rect 251 67673 263 67707
rect 273 67673 293 67707
rect 295 67692 324 67716
rect 303 67682 316 67692
rect 318 67676 324 67692
rect 333 67692 380 67716
rect 333 67682 353 67692
rect 367 67686 380 67692
rect 396 67686 408 67720
rect 420 67686 436 67720
rect 120 67625 170 67627
rect 76 67619 92 67625
rect 94 67619 110 67625
rect 76 67609 99 67618
rect 60 67599 67 67609
rect 76 67589 77 67609
rect 96 67584 99 67609
rect 109 67589 110 67609
rect 119 67599 126 67609
rect 76 67575 110 67579
rect 170 67575 172 67625
rect 186 67607 190 67641
rect 216 67607 220 67641
rect 186 67530 220 67564
rect 282 67561 292 67673
rect 318 67666 335 67676
rect 318 67597 324 67666
rect 346 67597 348 67682
rect 428 67639 430 67686
rect 476 67649 480 67717
rect 485 67699 495 67727
rect 505 67727 519 67733
rect 544 67727 555 67765
rect 505 67699 525 67727
rect 544 67699 553 67727
rect 544 67679 548 67699
rect 579 67658 582 67748
rect 612 67730 624 67731
rect 599 67728 649 67730
rect 612 67727 624 67728
rect 610 67720 632 67727
rect 607 67719 632 67720
rect 586 67712 644 67719
rect 607 67711 644 67712
rect 607 67695 610 67711
rect 616 67695 644 67711
rect 607 67694 644 67695
rect 586 67687 644 67694
rect 607 67686 610 67687
rect 612 67679 632 67687
rect 612 67675 624 67679
rect 649 67678 651 67728
rect 544 67641 548 67649
rect 400 67609 408 67639
rect 420 67609 436 67639
rect 400 67605 436 67609
rect 400 67597 430 67605
rect 428 67581 430 67597
rect 476 67569 480 67637
rect 544 67607 552 67641
rect 578 67607 582 67641
rect 544 67599 548 67607
rect 544 67569 586 67570
rect 288 67529 292 67561
rect 296 67559 368 67567
rect 378 67559 450 67567
rect 544 67562 548 67569
rect 439 67531 444 67559
rect 120 67515 170 67517
rect 76 67511 130 67515
rect 110 67506 130 67511
rect 60 67481 67 67491
rect 76 67481 77 67501
rect 96 67472 99 67506
rect 109 67481 110 67501
rect 119 67481 126 67491
rect 76 67465 92 67471
rect 94 67465 110 67471
rect 170 67465 172 67515
rect 186 67449 190 67483
rect 216 67449 220 67483
rect 213 67417 224 67449
rect 282 67445 292 67529
rect 296 67523 368 67531
rect 378 67523 450 67531
rect 468 67528 473 67562
rect 428 67493 430 67509
rect 251 67417 292 67445
rect 318 67424 324 67493
rect 12 67412 62 67414
rect 28 67403 59 67411
rect 62 67403 64 67412
rect 251 67411 263 67417
rect 28 67395 64 67403
rect 127 67403 158 67411
rect 127 67396 182 67403
rect 127 67395 161 67396
rect 59 67379 64 67395
rect 158 67379 161 67395
rect 253 67383 263 67411
rect 273 67383 293 67417
rect 318 67414 335 67424
rect 303 67398 316 67408
rect 318 67398 324 67414
rect 346 67408 348 67493
rect 400 67485 430 67493
rect 476 67491 480 67559
rect 511 67528 582 67562
rect 544 67521 548 67528
rect 400 67481 436 67485
rect 400 67451 408 67481
rect 420 67451 436 67481
rect 544 67483 548 67491
rect 28 67371 64 67379
rect 127 67378 161 67379
rect 127 67371 182 67378
rect 62 67362 64 67371
rect 282 67325 292 67383
rect 295 67374 324 67398
rect 333 67398 353 67408
rect 428 67404 430 67451
rect 476 67411 480 67479
rect 544 67449 552 67483
rect 578 67449 582 67483
rect 544 67441 548 67449
rect 367 67398 380 67404
rect 333 67374 380 67398
rect 318 67361 324 67374
rect 346 67361 348 67374
rect 367 67370 380 67374
rect 396 67370 408 67404
rect 420 67370 436 67404
rect 544 67401 553 67429
rect 319 67350 346 67361
rect 120 67309 170 67311
rect 76 67303 92 67309
rect 94 67303 110 67309
rect 76 67293 99 67302
rect 60 67283 67 67293
rect 76 67273 77 67293
rect 96 67268 99 67293
rect 109 67273 110 67293
rect 119 67283 126 67293
rect 76 67259 110 67263
rect 170 67259 172 67309
rect 186 67291 190 67325
rect 216 67291 220 67325
rect 182 67253 224 67254
rect 186 67229 220 67246
rect 223 67229 257 67246
rect 182 67212 257 67229
rect 182 67211 224 67212
rect 160 67205 246 67211
rect 288 67205 292 67325
rect 296 67323 368 67331
rect 428 67323 430 67370
rect 476 67333 480 67401
rect 485 67357 495 67391
rect 505 67363 525 67391
rect 505 67357 519 67363
rect 544 67357 555 67401
rect 485 67333 492 67357
rect 579 67342 582 67432
rect 612 67414 624 67415
rect 599 67412 649 67414
rect 612 67411 624 67412
rect 610 67404 632 67411
rect 607 67403 632 67404
rect 586 67396 644 67403
rect 607 67395 644 67396
rect 607 67379 610 67395
rect 616 67379 644 67395
rect 607 67378 644 67379
rect 586 67371 644 67378
rect 607 67370 610 67371
rect 612 67363 632 67371
rect 612 67359 624 67363
rect 649 67362 651 67412
rect 544 67325 548 67333
rect 400 67293 408 67323
rect 420 67293 436 67323
rect 400 67289 436 67293
rect 400 67281 430 67289
rect 428 67265 430 67281
rect 476 67253 480 67321
rect 544 67291 552 67325
rect 578 67291 582 67325
rect 544 67283 548 67291
rect 295 67212 300 67246
rect 324 67212 329 67246
rect 378 67243 450 67251
rect 544 67248 548 67253
rect 544 67244 582 67248
rect 544 67229 552 67244
rect 578 67229 582 67244
rect 544 67211 586 67229
rect 522 67205 608 67211
rect 182 67189 224 67205
rect 544 67189 586 67205
rect 17 67175 67 67177
rect 119 67175 169 67177
rect 186 67175 220 67189
rect 548 67175 582 67189
rect 599 67175 649 67177
rect 42 67133 59 67167
rect 67 67125 69 67175
rect 160 67167 246 67175
rect 522 67167 608 67175
rect 76 67133 110 67167
rect 127 67133 144 67167
rect 152 67133 161 67167
rect 162 67165 195 67167
rect 224 67165 244 67167
rect 162 67133 244 67165
rect 524 67165 548 67167
rect 573 67165 582 67167
rect 586 67165 606 67167
rect 160 67125 246 67133
rect 186 67109 220 67125
rect 182 67095 224 67096
rect 160 67089 182 67095
rect 224 67089 246 67095
rect 186 67054 220 67088
rect 223 67054 257 67088
rect 120 67041 170 67043
rect 76 67037 130 67041
rect 110 67032 130 67037
rect 60 67007 67 67017
rect 76 67007 77 67027
rect 96 66998 99 67032
rect 109 67007 110 67027
rect 119 67007 126 67017
rect 76 66991 92 66997
rect 94 66991 110 66997
rect 170 66991 172 67041
rect 186 66975 190 67009
rect 216 66975 220 67009
rect 288 66975 292 67163
rect 476 67095 480 67163
rect 524 67133 606 67165
rect 607 67133 616 67167
rect 522 67125 608 67133
rect 649 67125 651 67175
rect 548 67109 582 67125
rect 522 67090 548 67095
rect 522 67089 582 67090
rect 586 67089 608 67095
rect 295 67054 300 67088
rect 324 67054 329 67088
rect 544 67086 582 67089
rect 378 67049 450 67057
rect 428 67019 430 67035
rect 400 67011 430 67019
rect 476 67017 480 67085
rect 544 67056 552 67086
rect 578 67056 582 67086
rect 544 67047 548 67056
rect 400 67007 436 67011
rect 400 66977 408 67007
rect 420 66977 436 67007
rect 544 67009 548 67017
rect 12 66938 62 66940
rect 28 66929 59 66937
rect 62 66929 64 66938
rect 28 66921 64 66929
rect 127 66929 158 66937
rect 127 66922 182 66929
rect 215 66927 224 66955
rect 127 66921 161 66922
rect 59 66905 64 66921
rect 158 66905 161 66921
rect 28 66897 64 66905
rect 127 66904 161 66905
rect 127 66897 182 66904
rect 62 66888 64 66897
rect 213 66889 224 66927
rect 282 66917 292 66975
rect 296 66969 368 66977
rect 319 66939 346 66950
rect 318 66926 324 66939
rect 346 66926 348 66939
rect 428 66930 430 66977
rect 443 66967 450 66969
rect 476 66937 480 67005
rect 544 66975 552 67009
rect 578 66975 582 67009
rect 481 66943 517 66971
rect 481 66937 495 66943
rect 367 66926 380 66930
rect 251 66883 263 66917
rect 273 66883 293 66917
rect 295 66902 324 66926
rect 303 66892 316 66902
rect 318 66886 324 66902
rect 333 66902 380 66926
rect 333 66892 353 66902
rect 367 66896 380 66902
rect 396 66896 408 66930
rect 420 66896 436 66930
rect 120 66835 170 66837
rect 76 66829 92 66835
rect 94 66829 110 66835
rect 76 66819 99 66828
rect 60 66809 67 66819
rect 76 66799 77 66819
rect 96 66794 99 66819
rect 109 66799 110 66819
rect 119 66809 126 66819
rect 76 66785 110 66789
rect 170 66785 172 66835
rect 186 66817 190 66851
rect 216 66817 220 66851
rect 186 66740 220 66774
rect 282 66771 292 66883
rect 318 66876 335 66886
rect 318 66807 324 66876
rect 346 66807 348 66892
rect 428 66849 430 66896
rect 476 66859 480 66927
rect 485 66909 495 66937
rect 505 66937 519 66943
rect 544 66937 555 66975
rect 505 66909 525 66937
rect 544 66909 553 66937
rect 544 66889 548 66909
rect 579 66868 582 66958
rect 612 66940 624 66941
rect 599 66938 649 66940
rect 612 66937 624 66938
rect 610 66930 632 66937
rect 607 66929 632 66930
rect 586 66922 644 66929
rect 607 66921 644 66922
rect 607 66905 610 66921
rect 616 66905 644 66921
rect 607 66904 644 66905
rect 586 66897 644 66904
rect 607 66896 610 66897
rect 612 66889 632 66897
rect 612 66885 624 66889
rect 649 66888 651 66938
rect 544 66851 548 66859
rect 400 66819 408 66849
rect 420 66819 436 66849
rect 400 66815 436 66819
rect 400 66807 430 66815
rect 428 66791 430 66807
rect 476 66779 480 66847
rect 544 66817 552 66851
rect 578 66817 582 66851
rect 544 66809 548 66817
rect 544 66779 586 66780
rect 288 66739 292 66771
rect 296 66769 368 66777
rect 378 66769 450 66777
rect 544 66772 548 66779
rect 439 66741 444 66769
rect 120 66725 170 66727
rect 76 66721 130 66725
rect 110 66716 130 66721
rect 60 66691 67 66701
rect 76 66691 77 66711
rect 96 66682 99 66716
rect 109 66691 110 66711
rect 119 66691 126 66701
rect 76 66675 92 66681
rect 94 66675 110 66681
rect 170 66675 172 66725
rect 186 66659 190 66693
rect 216 66659 220 66693
rect 213 66627 224 66659
rect 282 66655 292 66739
rect 296 66733 368 66741
rect 378 66733 450 66741
rect 468 66738 473 66772
rect 428 66703 430 66719
rect 251 66627 292 66655
rect 318 66634 324 66703
rect 12 66622 62 66624
rect 28 66613 59 66621
rect 62 66613 64 66622
rect 251 66621 263 66627
rect 28 66605 64 66613
rect 127 66613 158 66621
rect 127 66606 182 66613
rect 127 66605 161 66606
rect 59 66589 64 66605
rect 158 66589 161 66605
rect 253 66593 263 66621
rect 273 66593 293 66627
rect 318 66624 335 66634
rect 303 66608 316 66618
rect 318 66608 324 66624
rect 346 66618 348 66703
rect 400 66695 430 66703
rect 476 66701 480 66769
rect 511 66738 582 66772
rect 544 66731 548 66738
rect 400 66691 436 66695
rect 400 66661 408 66691
rect 420 66661 436 66691
rect 544 66693 548 66701
rect 28 66581 64 66589
rect 127 66588 161 66589
rect 127 66581 182 66588
rect 62 66572 64 66581
rect 282 66535 292 66593
rect 295 66584 324 66608
rect 333 66608 353 66618
rect 428 66614 430 66661
rect 476 66621 480 66689
rect 544 66659 552 66693
rect 578 66659 582 66693
rect 544 66651 548 66659
rect 367 66608 380 66614
rect 333 66584 380 66608
rect 318 66571 324 66584
rect 346 66571 348 66584
rect 367 66580 380 66584
rect 396 66580 408 66614
rect 420 66580 436 66614
rect 544 66611 553 66639
rect 319 66560 346 66571
rect 120 66519 170 66521
rect 76 66513 92 66519
rect 94 66513 110 66519
rect 76 66503 99 66512
rect 60 66493 67 66503
rect 76 66483 77 66503
rect 96 66478 99 66503
rect 109 66483 110 66503
rect 119 66493 126 66503
rect 76 66469 110 66473
rect 170 66469 172 66519
rect 186 66501 190 66535
rect 216 66501 220 66535
rect 182 66463 224 66464
rect 186 66439 220 66456
rect 223 66439 257 66456
rect 182 66422 257 66439
rect 182 66421 224 66422
rect 160 66415 246 66421
rect 288 66415 292 66535
rect 296 66533 368 66541
rect 428 66533 430 66580
rect 476 66543 480 66611
rect 485 66567 495 66601
rect 505 66573 525 66601
rect 505 66567 519 66573
rect 544 66567 555 66611
rect 485 66543 492 66567
rect 579 66552 582 66642
rect 612 66624 624 66625
rect 599 66622 649 66624
rect 612 66621 624 66622
rect 610 66614 632 66621
rect 607 66613 632 66614
rect 586 66606 644 66613
rect 607 66605 644 66606
rect 607 66589 610 66605
rect 616 66589 644 66605
rect 607 66588 644 66589
rect 586 66581 644 66588
rect 607 66580 610 66581
rect 612 66573 632 66581
rect 612 66569 624 66573
rect 649 66572 651 66622
rect 544 66535 548 66543
rect 400 66503 408 66533
rect 420 66503 436 66533
rect 400 66499 436 66503
rect 400 66491 430 66499
rect 428 66475 430 66491
rect 476 66463 480 66531
rect 544 66501 552 66535
rect 578 66501 582 66535
rect 544 66493 548 66501
rect 295 66422 300 66456
rect 324 66422 329 66456
rect 378 66453 450 66461
rect 544 66458 548 66463
rect 544 66454 582 66458
rect 544 66439 552 66454
rect 578 66439 582 66454
rect 544 66421 586 66439
rect 522 66415 608 66421
rect 182 66399 224 66415
rect 544 66399 586 66415
rect 17 66385 67 66387
rect 119 66385 169 66387
rect 186 66385 220 66399
rect 548 66385 582 66399
rect 599 66385 649 66387
rect 42 66343 59 66377
rect 67 66335 69 66385
rect 160 66377 246 66385
rect 522 66377 608 66385
rect 76 66343 110 66377
rect 127 66343 144 66377
rect 152 66343 161 66377
rect 162 66375 195 66377
rect 224 66375 244 66377
rect 162 66343 244 66375
rect 524 66375 548 66377
rect 573 66375 582 66377
rect 586 66375 606 66377
rect 160 66335 246 66343
rect 186 66319 220 66335
rect 182 66305 224 66306
rect 160 66299 182 66305
rect 224 66299 246 66305
rect 186 66264 220 66298
rect 223 66264 257 66298
rect 120 66251 170 66253
rect 76 66247 130 66251
rect 110 66242 130 66247
rect 60 66217 67 66227
rect 76 66217 77 66237
rect 96 66208 99 66242
rect 109 66217 110 66237
rect 119 66217 126 66227
rect 76 66201 92 66207
rect 94 66201 110 66207
rect 170 66201 172 66251
rect 186 66185 190 66219
rect 216 66185 220 66219
rect 288 66185 292 66373
rect 476 66305 480 66373
rect 524 66343 606 66375
rect 607 66343 616 66377
rect 522 66335 608 66343
rect 649 66335 651 66385
rect 548 66319 582 66335
rect 522 66300 548 66305
rect 522 66299 582 66300
rect 586 66299 608 66305
rect 295 66264 300 66298
rect 324 66264 329 66298
rect 544 66296 582 66299
rect 378 66259 450 66267
rect 428 66229 430 66245
rect 400 66221 430 66229
rect 476 66227 480 66295
rect 544 66266 552 66296
rect 578 66266 582 66296
rect 544 66257 548 66266
rect 400 66217 436 66221
rect 400 66187 408 66217
rect 420 66187 436 66217
rect 544 66219 548 66227
rect 12 66148 62 66150
rect 28 66139 59 66147
rect 62 66139 64 66148
rect 28 66131 64 66139
rect 127 66139 158 66147
rect 127 66132 182 66139
rect 215 66137 224 66165
rect 127 66131 161 66132
rect 59 66115 64 66131
rect 158 66115 161 66131
rect 28 66107 64 66115
rect 127 66114 161 66115
rect 127 66107 182 66114
rect 62 66098 64 66107
rect 213 66099 224 66137
rect 282 66127 292 66185
rect 296 66179 368 66187
rect 319 66149 346 66160
rect 318 66136 324 66149
rect 346 66136 348 66149
rect 428 66140 430 66187
rect 443 66177 450 66179
rect 476 66147 480 66215
rect 544 66185 552 66219
rect 578 66185 582 66219
rect 481 66153 517 66181
rect 481 66147 495 66153
rect 367 66136 380 66140
rect 251 66093 263 66127
rect 273 66093 293 66127
rect 295 66112 324 66136
rect 303 66102 316 66112
rect 318 66096 324 66112
rect 333 66112 380 66136
rect 333 66102 353 66112
rect 367 66106 380 66112
rect 396 66106 408 66140
rect 420 66106 436 66140
rect 120 66045 170 66047
rect 76 66039 92 66045
rect 94 66039 110 66045
rect 76 66029 99 66038
rect 60 66019 67 66029
rect 76 66009 77 66029
rect 96 66004 99 66029
rect 109 66009 110 66029
rect 119 66019 126 66029
rect 76 65995 110 65999
rect 170 65995 172 66045
rect 186 66027 190 66061
rect 216 66027 220 66061
rect 186 65950 220 65984
rect 282 65981 292 66093
rect 318 66086 335 66096
rect 318 66017 324 66086
rect 346 66017 348 66102
rect 428 66059 430 66106
rect 476 66069 480 66137
rect 485 66119 495 66147
rect 505 66147 519 66153
rect 544 66147 555 66185
rect 505 66119 525 66147
rect 544 66119 553 66147
rect 544 66099 548 66119
rect 579 66078 582 66168
rect 612 66150 624 66151
rect 599 66148 649 66150
rect 612 66147 624 66148
rect 610 66140 632 66147
rect 607 66139 632 66140
rect 586 66132 644 66139
rect 607 66131 644 66132
rect 607 66115 610 66131
rect 616 66115 644 66131
rect 607 66114 644 66115
rect 586 66107 644 66114
rect 607 66106 610 66107
rect 612 66099 632 66107
rect 612 66095 624 66099
rect 649 66098 651 66148
rect 544 66061 548 66069
rect 400 66029 408 66059
rect 420 66029 436 66059
rect 400 66025 436 66029
rect 400 66017 430 66025
rect 428 66001 430 66017
rect 476 65989 480 66057
rect 544 66027 552 66061
rect 578 66027 582 66061
rect 544 66019 548 66027
rect 544 65989 586 65990
rect 288 65949 292 65981
rect 296 65979 368 65987
rect 378 65979 450 65987
rect 544 65982 548 65989
rect 439 65951 444 65979
rect 120 65935 170 65937
rect 76 65931 130 65935
rect 110 65926 130 65931
rect 60 65901 67 65911
rect 76 65901 77 65921
rect 96 65892 99 65926
rect 109 65901 110 65921
rect 119 65901 126 65911
rect 76 65885 92 65891
rect 94 65885 110 65891
rect 170 65885 172 65935
rect 186 65869 190 65903
rect 216 65869 220 65903
rect 213 65837 224 65869
rect 282 65865 292 65949
rect 296 65943 368 65951
rect 378 65943 450 65951
rect 468 65948 473 65982
rect 428 65913 430 65929
rect 251 65837 292 65865
rect 318 65844 324 65913
rect 12 65832 62 65834
rect 28 65823 59 65831
rect 62 65823 64 65832
rect 251 65831 263 65837
rect 28 65815 64 65823
rect 127 65823 158 65831
rect 127 65816 182 65823
rect 127 65815 161 65816
rect 59 65799 64 65815
rect 158 65799 161 65815
rect 253 65803 263 65831
rect 273 65803 293 65837
rect 318 65834 335 65844
rect 303 65818 316 65828
rect 318 65818 324 65834
rect 346 65828 348 65913
rect 400 65905 430 65913
rect 476 65911 480 65979
rect 511 65948 582 65982
rect 544 65941 548 65948
rect 400 65901 436 65905
rect 400 65871 408 65901
rect 420 65871 436 65901
rect 544 65903 548 65911
rect 28 65791 64 65799
rect 127 65798 161 65799
rect 127 65791 182 65798
rect 62 65782 64 65791
rect 282 65745 292 65803
rect 295 65794 324 65818
rect 333 65818 353 65828
rect 428 65824 430 65871
rect 476 65831 480 65899
rect 544 65869 552 65903
rect 578 65869 582 65903
rect 544 65861 548 65869
rect 367 65818 380 65824
rect 333 65794 380 65818
rect 318 65781 324 65794
rect 346 65781 348 65794
rect 367 65790 380 65794
rect 396 65790 408 65824
rect 420 65790 436 65824
rect 544 65821 553 65849
rect 319 65770 346 65781
rect 120 65729 170 65731
rect 76 65723 92 65729
rect 94 65723 110 65729
rect 76 65713 99 65722
rect 60 65703 67 65713
rect 76 65693 77 65713
rect 96 65688 99 65713
rect 109 65693 110 65713
rect 119 65703 126 65713
rect 76 65679 110 65683
rect 170 65679 172 65729
rect 186 65711 190 65745
rect 216 65711 220 65745
rect 182 65673 224 65674
rect 186 65649 220 65666
rect 223 65649 257 65666
rect 182 65632 257 65649
rect 182 65631 224 65632
rect 160 65625 246 65631
rect 288 65625 292 65745
rect 296 65743 368 65751
rect 428 65743 430 65790
rect 476 65753 480 65821
rect 485 65777 495 65811
rect 505 65783 525 65811
rect 505 65777 519 65783
rect 544 65777 555 65821
rect 485 65753 492 65777
rect 579 65762 582 65852
rect 612 65834 624 65835
rect 599 65832 649 65834
rect 612 65831 624 65832
rect 610 65824 632 65831
rect 607 65823 632 65824
rect 586 65816 644 65823
rect 607 65815 644 65816
rect 607 65799 610 65815
rect 616 65799 644 65815
rect 607 65798 644 65799
rect 586 65791 644 65798
rect 607 65790 610 65791
rect 612 65783 632 65791
rect 612 65779 624 65783
rect 649 65782 651 65832
rect 544 65745 548 65753
rect 400 65713 408 65743
rect 420 65713 436 65743
rect 400 65709 436 65713
rect 400 65701 430 65709
rect 428 65685 430 65701
rect 476 65673 480 65741
rect 544 65711 552 65745
rect 578 65711 582 65745
rect 544 65703 548 65711
rect 295 65632 300 65666
rect 324 65632 329 65666
rect 378 65663 450 65671
rect 544 65668 548 65673
rect 544 65664 582 65668
rect 544 65649 552 65664
rect 578 65649 582 65664
rect 544 65631 586 65649
rect 522 65625 608 65631
rect 182 65609 224 65625
rect 544 65609 586 65625
rect 17 65595 67 65597
rect 119 65595 169 65597
rect 186 65595 220 65609
rect 548 65595 582 65609
rect 599 65595 649 65597
rect 42 65553 59 65587
rect 67 65545 69 65595
rect 160 65587 246 65595
rect 522 65587 608 65595
rect 76 65553 110 65587
rect 127 65553 144 65587
rect 152 65553 161 65587
rect 162 65585 195 65587
rect 224 65585 244 65587
rect 162 65553 244 65585
rect 524 65585 548 65587
rect 573 65585 582 65587
rect 586 65585 606 65587
rect 160 65545 246 65553
rect 186 65529 220 65545
rect 182 65515 224 65516
rect 160 65509 182 65515
rect 224 65509 246 65515
rect 186 65474 220 65508
rect 223 65474 257 65508
rect 120 65461 170 65463
rect 76 65457 130 65461
rect 110 65452 130 65457
rect 60 65427 67 65437
rect 76 65427 77 65447
rect 96 65418 99 65452
rect 109 65427 110 65447
rect 119 65427 126 65437
rect 76 65411 92 65417
rect 94 65411 110 65417
rect 170 65411 172 65461
rect 186 65395 190 65429
rect 216 65395 220 65429
rect 288 65395 292 65583
rect 476 65515 480 65583
rect 524 65553 606 65585
rect 607 65553 616 65587
rect 522 65545 608 65553
rect 649 65545 651 65595
rect 548 65529 582 65545
rect 522 65510 548 65515
rect 522 65509 582 65510
rect 586 65509 608 65515
rect 295 65474 300 65508
rect 324 65474 329 65508
rect 544 65506 582 65509
rect 378 65469 450 65477
rect 428 65439 430 65455
rect 400 65431 430 65439
rect 476 65437 480 65505
rect 544 65476 552 65506
rect 578 65476 582 65506
rect 544 65467 548 65476
rect 400 65427 436 65431
rect 400 65397 408 65427
rect 420 65397 436 65427
rect 544 65429 548 65437
rect 12 65358 62 65360
rect 28 65349 59 65357
rect 62 65349 64 65358
rect 28 65341 64 65349
rect 127 65349 158 65357
rect 127 65342 182 65349
rect 215 65347 224 65375
rect 127 65341 161 65342
rect 59 65325 64 65341
rect 158 65325 161 65341
rect 28 65317 64 65325
rect 127 65324 161 65325
rect 127 65317 182 65324
rect 62 65308 64 65317
rect 213 65309 224 65347
rect 282 65337 292 65395
rect 296 65389 368 65397
rect 319 65359 346 65370
rect 318 65346 324 65359
rect 346 65346 348 65359
rect 428 65350 430 65397
rect 443 65387 450 65389
rect 476 65357 480 65425
rect 544 65395 552 65429
rect 578 65395 582 65429
rect 481 65363 517 65391
rect 481 65357 495 65363
rect 367 65346 380 65350
rect 251 65303 263 65337
rect 273 65303 293 65337
rect 295 65322 324 65346
rect 303 65312 316 65322
rect 318 65306 324 65322
rect 333 65322 380 65346
rect 333 65312 353 65322
rect 367 65316 380 65322
rect 396 65316 408 65350
rect 420 65316 436 65350
rect 120 65255 170 65257
rect 76 65249 92 65255
rect 94 65249 110 65255
rect 76 65239 99 65248
rect 60 65229 67 65239
rect 76 65219 77 65239
rect 96 65214 99 65239
rect 109 65219 110 65239
rect 119 65229 126 65239
rect 76 65205 110 65209
rect 170 65205 172 65255
rect 186 65237 190 65271
rect 216 65237 220 65271
rect 186 65160 220 65194
rect 282 65191 292 65303
rect 318 65296 335 65306
rect 318 65227 324 65296
rect 346 65227 348 65312
rect 428 65269 430 65316
rect 476 65279 480 65347
rect 485 65329 495 65357
rect 505 65357 519 65363
rect 544 65357 555 65395
rect 505 65329 525 65357
rect 544 65329 553 65357
rect 544 65309 548 65329
rect 579 65288 582 65378
rect 612 65360 624 65361
rect 599 65358 649 65360
rect 612 65357 624 65358
rect 610 65350 632 65357
rect 607 65349 632 65350
rect 586 65342 644 65349
rect 607 65341 644 65342
rect 607 65325 610 65341
rect 616 65325 644 65341
rect 607 65324 644 65325
rect 586 65317 644 65324
rect 607 65316 610 65317
rect 612 65309 632 65317
rect 612 65305 624 65309
rect 649 65308 651 65358
rect 544 65271 548 65279
rect 400 65239 408 65269
rect 420 65239 436 65269
rect 400 65235 436 65239
rect 400 65227 430 65235
rect 428 65211 430 65227
rect 476 65199 480 65267
rect 544 65237 552 65271
rect 578 65237 582 65271
rect 544 65229 548 65237
rect 544 65199 586 65200
rect 288 65159 292 65191
rect 296 65189 368 65197
rect 378 65189 450 65197
rect 544 65192 548 65199
rect 439 65161 444 65189
rect 120 65145 170 65147
rect 76 65141 130 65145
rect 110 65136 130 65141
rect 60 65111 67 65121
rect 76 65111 77 65131
rect 96 65102 99 65136
rect 109 65111 110 65131
rect 119 65111 126 65121
rect 76 65095 92 65101
rect 94 65095 110 65101
rect 170 65095 172 65145
rect 186 65079 190 65113
rect 216 65079 220 65113
rect 213 65047 224 65079
rect 282 65075 292 65159
rect 296 65153 368 65161
rect 378 65153 450 65161
rect 468 65158 473 65192
rect 428 65123 430 65139
rect 251 65047 292 65075
rect 318 65054 324 65123
rect 12 65042 62 65044
rect 28 65033 59 65041
rect 62 65033 64 65042
rect 251 65041 263 65047
rect 28 65025 64 65033
rect 127 65033 158 65041
rect 127 65026 182 65033
rect 127 65025 161 65026
rect 59 65009 64 65025
rect 158 65009 161 65025
rect 253 65013 263 65041
rect 273 65013 293 65047
rect 318 65044 335 65054
rect 303 65028 316 65038
rect 318 65028 324 65044
rect 346 65038 348 65123
rect 400 65115 430 65123
rect 476 65121 480 65189
rect 511 65158 582 65192
rect 544 65151 548 65158
rect 400 65111 436 65115
rect 400 65081 408 65111
rect 420 65081 436 65111
rect 544 65113 548 65121
rect 28 65001 64 65009
rect 127 65008 161 65009
rect 127 65001 182 65008
rect 62 64992 64 65001
rect 282 64955 292 65013
rect 295 65004 324 65028
rect 333 65028 353 65038
rect 428 65034 430 65081
rect 476 65041 480 65109
rect 544 65079 552 65113
rect 578 65079 582 65113
rect 544 65071 548 65079
rect 367 65028 380 65034
rect 333 65004 380 65028
rect 318 64991 324 65004
rect 346 64991 348 65004
rect 367 65000 380 65004
rect 396 65000 408 65034
rect 420 65000 436 65034
rect 544 65031 553 65059
rect 319 64980 346 64991
rect 120 64939 170 64941
rect 76 64933 92 64939
rect 94 64933 110 64939
rect 76 64923 99 64932
rect 60 64913 67 64923
rect 76 64903 77 64923
rect 96 64898 99 64923
rect 109 64903 110 64923
rect 119 64913 126 64923
rect 76 64889 110 64893
rect 170 64889 172 64939
rect 186 64921 190 64955
rect 216 64921 220 64955
rect 182 64883 224 64884
rect 186 64859 220 64876
rect 223 64859 257 64876
rect 182 64842 257 64859
rect 182 64841 224 64842
rect 160 64835 246 64841
rect 288 64835 292 64955
rect 296 64953 368 64961
rect 428 64953 430 65000
rect 476 64963 480 65031
rect 485 64987 495 65021
rect 505 64993 525 65021
rect 505 64987 519 64993
rect 544 64987 555 65031
rect 485 64963 492 64987
rect 579 64972 582 65062
rect 612 65044 624 65045
rect 599 65042 649 65044
rect 612 65041 624 65042
rect 610 65034 632 65041
rect 607 65033 632 65034
rect 586 65026 644 65033
rect 607 65025 644 65026
rect 607 65009 610 65025
rect 616 65009 644 65025
rect 607 65008 644 65009
rect 586 65001 644 65008
rect 607 65000 610 65001
rect 612 64993 632 65001
rect 612 64989 624 64993
rect 649 64992 651 65042
rect 544 64955 548 64963
rect 400 64923 408 64953
rect 420 64923 436 64953
rect 400 64919 436 64923
rect 400 64911 430 64919
rect 428 64895 430 64911
rect 476 64883 480 64951
rect 544 64921 552 64955
rect 578 64921 582 64955
rect 544 64913 548 64921
rect 295 64842 300 64876
rect 324 64842 329 64876
rect 378 64873 450 64881
rect 544 64878 548 64883
rect 544 64874 582 64878
rect 544 64859 552 64874
rect 578 64859 582 64874
rect 544 64841 586 64859
rect 522 64835 608 64841
rect 182 64819 224 64835
rect 544 64819 586 64835
rect 17 64805 67 64807
rect 119 64805 169 64807
rect 186 64805 220 64819
rect 548 64805 582 64819
rect 599 64805 649 64807
rect 42 64763 59 64797
rect 67 64755 69 64805
rect 160 64797 246 64805
rect 522 64797 608 64805
rect 76 64763 110 64797
rect 127 64763 144 64797
rect 152 64763 161 64797
rect 162 64795 195 64797
rect 224 64795 244 64797
rect 162 64763 244 64795
rect 524 64795 548 64797
rect 573 64795 582 64797
rect 586 64795 606 64797
rect 160 64755 246 64763
rect 186 64739 220 64755
rect 182 64725 224 64726
rect 160 64719 182 64725
rect 224 64719 246 64725
rect 186 64684 220 64718
rect 223 64684 257 64718
rect 120 64671 170 64673
rect 76 64667 130 64671
rect 110 64662 130 64667
rect 60 64637 67 64647
rect 76 64637 77 64657
rect 96 64628 99 64662
rect 109 64637 110 64657
rect 119 64637 126 64647
rect 76 64621 92 64627
rect 94 64621 110 64627
rect 170 64621 172 64671
rect 186 64605 190 64639
rect 216 64605 220 64639
rect 288 64605 292 64793
rect 476 64725 480 64793
rect 524 64763 606 64795
rect 607 64763 616 64797
rect 522 64755 608 64763
rect 649 64755 651 64805
rect 548 64739 582 64755
rect 522 64720 548 64725
rect 522 64719 582 64720
rect 586 64719 608 64725
rect 295 64684 300 64718
rect 324 64684 329 64718
rect 544 64716 582 64719
rect 378 64679 450 64687
rect 428 64649 430 64665
rect 400 64641 430 64649
rect 476 64647 480 64715
rect 544 64686 552 64716
rect 578 64686 582 64716
rect 544 64677 548 64686
rect 400 64637 436 64641
rect 400 64607 408 64637
rect 420 64607 436 64637
rect 544 64639 548 64647
rect 12 64568 62 64570
rect 28 64559 59 64567
rect 62 64559 64 64568
rect 28 64551 64 64559
rect 127 64559 158 64567
rect 127 64552 182 64559
rect 215 64557 224 64585
rect 127 64551 161 64552
rect 59 64535 64 64551
rect 158 64535 161 64551
rect 28 64527 64 64535
rect 127 64534 161 64535
rect 127 64527 182 64534
rect 62 64518 64 64527
rect 213 64519 224 64557
rect 282 64547 292 64605
rect 296 64599 368 64607
rect 319 64569 346 64580
rect 318 64556 324 64569
rect 346 64556 348 64569
rect 428 64560 430 64607
rect 443 64597 450 64599
rect 476 64567 480 64635
rect 544 64605 552 64639
rect 578 64605 582 64639
rect 481 64573 517 64601
rect 481 64567 495 64573
rect 367 64556 380 64560
rect 251 64513 263 64547
rect 273 64513 293 64547
rect 295 64532 324 64556
rect 303 64522 316 64532
rect 318 64516 324 64532
rect 333 64532 380 64556
rect 333 64522 353 64532
rect 367 64526 380 64532
rect 396 64526 408 64560
rect 420 64526 436 64560
rect 120 64465 170 64467
rect 76 64459 92 64465
rect 94 64459 110 64465
rect 76 64449 99 64458
rect 60 64439 67 64449
rect 76 64429 77 64449
rect 96 64424 99 64449
rect 109 64429 110 64449
rect 119 64439 126 64449
rect 76 64415 110 64419
rect 170 64415 172 64465
rect 186 64447 190 64481
rect 216 64447 220 64481
rect 186 64370 220 64404
rect 282 64401 292 64513
rect 318 64506 335 64516
rect 318 64437 324 64506
rect 346 64437 348 64522
rect 428 64479 430 64526
rect 476 64489 480 64557
rect 485 64539 495 64567
rect 505 64567 519 64573
rect 544 64567 555 64605
rect 505 64539 525 64567
rect 544 64539 553 64567
rect 544 64519 548 64539
rect 579 64498 582 64588
rect 612 64570 624 64571
rect 599 64568 649 64570
rect 612 64567 624 64568
rect 610 64560 632 64567
rect 607 64559 632 64560
rect 586 64552 644 64559
rect 607 64551 644 64552
rect 607 64535 610 64551
rect 616 64535 644 64551
rect 607 64534 644 64535
rect 586 64527 644 64534
rect 607 64526 610 64527
rect 612 64519 632 64527
rect 612 64515 624 64519
rect 649 64518 651 64568
rect 544 64481 548 64489
rect 400 64449 408 64479
rect 420 64449 436 64479
rect 400 64445 436 64449
rect 400 64437 430 64445
rect 428 64421 430 64437
rect 476 64409 480 64477
rect 544 64447 552 64481
rect 578 64447 582 64481
rect 544 64439 548 64447
rect 544 64409 586 64410
rect 288 64369 292 64401
rect 296 64399 368 64407
rect 378 64399 450 64407
rect 544 64402 548 64409
rect 439 64371 444 64399
rect 120 64355 170 64357
rect 76 64351 130 64355
rect 110 64346 130 64351
rect 60 64321 67 64331
rect 76 64321 77 64341
rect 96 64312 99 64346
rect 109 64321 110 64341
rect 119 64321 126 64331
rect 76 64305 92 64311
rect 94 64305 110 64311
rect 170 64305 172 64355
rect 186 64289 190 64323
rect 216 64289 220 64323
rect 213 64257 224 64289
rect 282 64285 292 64369
rect 296 64363 368 64371
rect 378 64363 450 64371
rect 468 64368 473 64402
rect 428 64333 430 64349
rect 251 64257 292 64285
rect 318 64264 324 64333
rect 12 64252 62 64254
rect 28 64243 59 64251
rect 62 64243 64 64252
rect 251 64251 263 64257
rect 28 64235 64 64243
rect 127 64243 158 64251
rect 127 64236 182 64243
rect 127 64235 161 64236
rect 59 64219 64 64235
rect 158 64219 161 64235
rect 253 64223 263 64251
rect 273 64223 293 64257
rect 318 64254 335 64264
rect 303 64238 316 64248
rect 318 64238 324 64254
rect 346 64248 348 64333
rect 400 64325 430 64333
rect 476 64331 480 64399
rect 511 64368 582 64402
rect 544 64361 548 64368
rect 400 64321 436 64325
rect 400 64291 408 64321
rect 420 64291 436 64321
rect 544 64323 548 64331
rect 28 64211 64 64219
rect 127 64218 161 64219
rect 127 64211 182 64218
rect 62 64202 64 64211
rect 282 64165 292 64223
rect 295 64214 324 64238
rect 333 64238 353 64248
rect 428 64244 430 64291
rect 476 64251 480 64319
rect 544 64289 552 64323
rect 578 64289 582 64323
rect 544 64281 548 64289
rect 367 64238 380 64244
rect 333 64214 380 64238
rect 318 64201 324 64214
rect 346 64201 348 64214
rect 367 64210 380 64214
rect 396 64210 408 64244
rect 420 64210 436 64244
rect 544 64241 553 64269
rect 319 64190 346 64201
rect 120 64149 170 64151
rect 76 64143 92 64149
rect 94 64143 110 64149
rect 76 64133 99 64142
rect 60 64123 67 64133
rect 76 64113 77 64133
rect 96 64108 99 64133
rect 109 64113 110 64133
rect 119 64123 126 64133
rect 76 64099 110 64103
rect 170 64099 172 64149
rect 186 64131 190 64165
rect 216 64131 220 64165
rect 182 64093 224 64094
rect 186 64069 220 64086
rect 223 64069 257 64086
rect 182 64052 257 64069
rect 182 64051 224 64052
rect 160 64045 246 64051
rect 288 64045 292 64165
rect 296 64163 368 64171
rect 428 64163 430 64210
rect 476 64173 480 64241
rect 485 64197 495 64231
rect 505 64203 525 64231
rect 505 64197 519 64203
rect 544 64197 555 64241
rect 485 64173 492 64197
rect 579 64182 582 64272
rect 612 64254 624 64255
rect 599 64252 649 64254
rect 612 64251 624 64252
rect 610 64244 632 64251
rect 607 64243 632 64244
rect 586 64236 644 64243
rect 607 64235 644 64236
rect 607 64219 610 64235
rect 616 64219 644 64235
rect 607 64218 644 64219
rect 586 64211 644 64218
rect 607 64210 610 64211
rect 612 64203 632 64211
rect 612 64199 624 64203
rect 649 64202 651 64252
rect 544 64165 548 64173
rect 400 64133 408 64163
rect 420 64133 436 64163
rect 400 64129 436 64133
rect 400 64121 430 64129
rect 428 64105 430 64121
rect 476 64093 480 64161
rect 544 64131 552 64165
rect 578 64131 582 64165
rect 544 64123 548 64131
rect 295 64052 300 64086
rect 324 64052 329 64086
rect 378 64083 450 64091
rect 544 64088 548 64093
rect 544 64084 582 64088
rect 544 64069 552 64084
rect 578 64069 582 64084
rect 544 64051 586 64069
rect 522 64045 608 64051
rect 182 64029 224 64045
rect 544 64029 586 64045
rect 17 64015 67 64017
rect 119 64015 169 64017
rect 186 64015 220 64029
rect 548 64015 582 64029
rect 599 64015 649 64017
rect 42 63973 59 64007
rect 67 63965 69 64015
rect 160 64007 246 64015
rect 522 64007 608 64015
rect 76 63973 110 64007
rect 127 63973 144 64007
rect 152 63973 161 64007
rect 162 64005 195 64007
rect 224 64005 244 64007
rect 162 63973 244 64005
rect 524 64005 548 64007
rect 573 64005 582 64007
rect 586 64005 606 64007
rect 160 63965 246 63973
rect 186 63949 220 63965
rect 182 63935 224 63936
rect 160 63929 182 63935
rect 224 63929 246 63935
rect 186 63894 220 63928
rect 223 63894 257 63928
rect 120 63881 170 63883
rect 76 63877 130 63881
rect 110 63872 130 63877
rect 60 63847 67 63857
rect 76 63847 77 63867
rect 96 63838 99 63872
rect 109 63847 110 63867
rect 119 63847 126 63857
rect 76 63831 92 63837
rect 94 63831 110 63837
rect 170 63831 172 63881
rect 186 63815 190 63849
rect 216 63815 220 63849
rect 288 63815 292 64003
rect 476 63935 480 64003
rect 524 63973 606 64005
rect 607 63973 616 64007
rect 522 63965 608 63973
rect 649 63965 651 64015
rect 548 63949 582 63965
rect 522 63930 548 63935
rect 522 63929 582 63930
rect 586 63929 608 63935
rect 295 63894 300 63928
rect 324 63894 329 63928
rect 544 63926 582 63929
rect 378 63889 450 63897
rect 428 63859 430 63875
rect 400 63851 430 63859
rect 476 63857 480 63925
rect 544 63896 552 63926
rect 578 63896 582 63926
rect 544 63887 548 63896
rect 400 63847 436 63851
rect 400 63817 408 63847
rect 420 63817 436 63847
rect 544 63849 548 63857
rect 12 63778 62 63780
rect 28 63769 59 63777
rect 62 63769 64 63778
rect 28 63761 64 63769
rect 127 63769 158 63777
rect 127 63762 182 63769
rect 215 63767 224 63795
rect 127 63761 161 63762
rect 59 63745 64 63761
rect 158 63745 161 63761
rect 28 63737 64 63745
rect 127 63744 161 63745
rect 127 63737 182 63744
rect 62 63728 64 63737
rect 213 63729 224 63767
rect 282 63757 292 63815
rect 296 63809 368 63817
rect 319 63779 346 63790
rect 318 63766 324 63779
rect 346 63766 348 63779
rect 428 63770 430 63817
rect 443 63807 450 63809
rect 476 63777 480 63845
rect 544 63815 552 63849
rect 578 63815 582 63849
rect 481 63783 517 63811
rect 481 63777 495 63783
rect 367 63766 380 63770
rect 251 63723 263 63757
rect 273 63723 293 63757
rect 295 63742 324 63766
rect 303 63732 316 63742
rect 318 63726 324 63742
rect 333 63742 380 63766
rect 333 63732 353 63742
rect 367 63736 380 63742
rect 396 63736 408 63770
rect 420 63736 436 63770
rect 120 63675 170 63677
rect 76 63669 92 63675
rect 94 63669 110 63675
rect 76 63659 99 63668
rect 60 63649 67 63659
rect 76 63639 77 63659
rect 96 63634 99 63659
rect 109 63639 110 63659
rect 119 63649 126 63659
rect 76 63625 110 63629
rect 170 63625 172 63675
rect 186 63657 190 63691
rect 216 63657 220 63691
rect 186 63580 220 63614
rect 282 63611 292 63723
rect 318 63716 335 63726
rect 318 63647 324 63716
rect 346 63647 348 63732
rect 428 63689 430 63736
rect 476 63699 480 63767
rect 485 63749 495 63777
rect 505 63777 519 63783
rect 544 63777 555 63815
rect 505 63749 525 63777
rect 544 63749 553 63777
rect 544 63729 548 63749
rect 579 63708 582 63798
rect 612 63780 624 63781
rect 599 63778 649 63780
rect 612 63777 624 63778
rect 610 63770 632 63777
rect 607 63769 632 63770
rect 586 63762 644 63769
rect 607 63761 644 63762
rect 607 63745 610 63761
rect 616 63745 644 63761
rect 607 63744 644 63745
rect 586 63737 644 63744
rect 607 63736 610 63737
rect 612 63729 632 63737
rect 612 63725 624 63729
rect 649 63728 651 63778
rect 544 63691 548 63699
rect 400 63659 408 63689
rect 420 63659 436 63689
rect 400 63655 436 63659
rect 400 63647 430 63655
rect 428 63631 430 63647
rect 476 63619 480 63687
rect 544 63657 552 63691
rect 578 63657 582 63691
rect 544 63649 548 63657
rect 544 63619 586 63620
rect 288 63579 292 63611
rect 296 63609 368 63617
rect 378 63609 450 63617
rect 544 63612 548 63619
rect 439 63581 444 63609
rect 120 63565 170 63567
rect 76 63561 130 63565
rect 110 63556 130 63561
rect 60 63531 67 63541
rect 76 63531 77 63551
rect 96 63522 99 63556
rect 109 63531 110 63551
rect 119 63531 126 63541
rect 76 63515 92 63521
rect 94 63515 110 63521
rect 170 63515 172 63565
rect 186 63499 190 63533
rect 216 63499 220 63533
rect 213 63467 224 63499
rect 282 63495 292 63579
rect 296 63573 368 63581
rect 378 63573 450 63581
rect 468 63578 473 63612
rect 428 63543 430 63559
rect 251 63467 292 63495
rect 318 63474 324 63543
rect 12 63462 62 63464
rect 28 63453 59 63461
rect 62 63453 64 63462
rect 251 63461 263 63467
rect 28 63445 64 63453
rect 127 63453 158 63461
rect 127 63446 182 63453
rect 127 63445 161 63446
rect 59 63429 64 63445
rect 158 63429 161 63445
rect 253 63433 263 63461
rect 273 63433 293 63467
rect 318 63464 335 63474
rect 303 63448 316 63458
rect 318 63448 324 63464
rect 346 63458 348 63543
rect 400 63535 430 63543
rect 476 63541 480 63609
rect 511 63578 582 63612
rect 544 63571 548 63578
rect 400 63531 436 63535
rect 400 63501 408 63531
rect 420 63501 436 63531
rect 544 63533 548 63541
rect 28 63421 64 63429
rect 127 63428 161 63429
rect 127 63421 182 63428
rect 62 63412 64 63421
rect 282 63375 292 63433
rect 295 63424 324 63448
rect 333 63448 353 63458
rect 428 63454 430 63501
rect 476 63461 480 63529
rect 544 63499 552 63533
rect 578 63499 582 63533
rect 544 63491 548 63499
rect 367 63448 380 63454
rect 333 63424 380 63448
rect 318 63411 324 63424
rect 346 63411 348 63424
rect 367 63420 380 63424
rect 396 63420 408 63454
rect 420 63420 436 63454
rect 544 63451 553 63479
rect 319 63400 346 63411
rect 120 63359 170 63361
rect 76 63353 92 63359
rect 94 63353 110 63359
rect 76 63343 99 63352
rect 60 63333 67 63343
rect 76 63323 77 63343
rect 96 63318 99 63343
rect 109 63323 110 63343
rect 119 63333 126 63343
rect 76 63309 110 63313
rect 170 63309 172 63359
rect 186 63341 190 63375
rect 216 63341 220 63375
rect 182 63303 224 63304
rect 186 63279 220 63296
rect 223 63279 257 63296
rect 182 63262 257 63279
rect 182 63261 224 63262
rect 160 63255 246 63261
rect 288 63255 292 63375
rect 296 63373 368 63381
rect 428 63373 430 63420
rect 476 63383 480 63451
rect 485 63407 495 63441
rect 505 63413 525 63441
rect 505 63407 519 63413
rect 544 63407 555 63451
rect 485 63383 492 63407
rect 579 63392 582 63482
rect 612 63464 624 63465
rect 599 63462 649 63464
rect 612 63461 624 63462
rect 610 63454 632 63461
rect 607 63453 632 63454
rect 586 63446 644 63453
rect 607 63445 644 63446
rect 607 63429 610 63445
rect 616 63429 644 63445
rect 607 63428 644 63429
rect 586 63421 644 63428
rect 607 63420 610 63421
rect 612 63413 632 63421
rect 612 63409 624 63413
rect 649 63412 651 63462
rect 544 63375 548 63383
rect 400 63343 408 63373
rect 420 63343 436 63373
rect 400 63339 436 63343
rect 400 63331 430 63339
rect 428 63315 430 63331
rect 476 63303 480 63371
rect 544 63341 552 63375
rect 578 63341 582 63375
rect 544 63333 548 63341
rect 295 63262 300 63296
rect 324 63262 329 63296
rect 378 63293 450 63301
rect 544 63298 548 63303
rect 544 63294 582 63298
rect 544 63279 552 63294
rect 578 63279 582 63294
rect 544 63261 586 63279
rect 522 63255 608 63261
rect 182 63239 224 63255
rect 544 63239 586 63255
rect 17 63225 67 63227
rect 119 63225 169 63227
rect 186 63225 220 63239
rect 548 63225 582 63239
rect 599 63225 649 63227
rect 42 63183 59 63217
rect 67 63175 69 63225
rect 160 63217 246 63225
rect 522 63217 608 63225
rect 76 63183 110 63217
rect 127 63183 144 63217
rect 152 63183 161 63217
rect 162 63215 195 63217
rect 224 63215 244 63217
rect 162 63183 244 63215
rect 524 63215 548 63217
rect 573 63215 582 63217
rect 586 63215 606 63217
rect 160 63175 246 63183
rect 186 63159 220 63175
rect 182 63145 224 63146
rect 160 63139 182 63145
rect 224 63139 246 63145
rect 186 63104 220 63138
rect 223 63104 257 63138
rect 120 63091 170 63093
rect 76 63087 130 63091
rect 110 63082 130 63087
rect 60 63057 67 63067
rect 76 63057 77 63077
rect 96 63048 99 63082
rect 109 63057 110 63077
rect 119 63057 126 63067
rect 76 63041 92 63047
rect 94 63041 110 63047
rect 170 63041 172 63091
rect 186 63025 190 63059
rect 216 63025 220 63059
rect 288 63025 292 63213
rect 476 63145 480 63213
rect 524 63183 606 63215
rect 607 63183 616 63217
rect 522 63175 608 63183
rect 649 63175 651 63225
rect 548 63159 582 63175
rect 522 63140 548 63145
rect 522 63139 582 63140
rect 586 63139 608 63145
rect 295 63104 300 63138
rect 324 63104 329 63138
rect 544 63136 582 63139
rect 378 63099 450 63107
rect 428 63069 430 63085
rect 400 63061 430 63069
rect 476 63067 480 63135
rect 544 63106 552 63136
rect 578 63106 582 63136
rect 544 63097 548 63106
rect 400 63057 436 63061
rect 400 63027 408 63057
rect 420 63027 436 63057
rect 544 63059 548 63067
rect 12 62988 62 62990
rect 28 62979 59 62987
rect 62 62979 64 62988
rect 28 62971 64 62979
rect 127 62979 158 62987
rect 127 62972 182 62979
rect 215 62977 224 63005
rect 127 62971 161 62972
rect 59 62955 64 62971
rect 158 62955 161 62971
rect 28 62947 64 62955
rect 127 62954 161 62955
rect 127 62947 182 62954
rect 62 62938 64 62947
rect 213 62939 224 62977
rect 282 62967 292 63025
rect 296 63019 368 63027
rect 319 62989 346 63000
rect 318 62976 324 62989
rect 346 62976 348 62989
rect 428 62980 430 63027
rect 443 63017 450 63019
rect 476 62987 480 63055
rect 544 63025 552 63059
rect 578 63025 582 63059
rect 481 62993 517 63021
rect 481 62987 495 62993
rect 367 62976 380 62980
rect 251 62933 263 62967
rect 273 62933 293 62967
rect 295 62952 324 62976
rect 303 62942 316 62952
rect 318 62936 324 62952
rect 333 62952 380 62976
rect 333 62942 353 62952
rect 367 62946 380 62952
rect 396 62946 408 62980
rect 420 62946 436 62980
rect 120 62885 170 62887
rect 76 62879 92 62885
rect 94 62879 110 62885
rect 76 62869 99 62878
rect 60 62859 67 62869
rect 76 62849 77 62869
rect 96 62844 99 62869
rect 109 62849 110 62869
rect 119 62859 126 62869
rect 76 62835 110 62839
rect 170 62835 172 62885
rect 186 62867 190 62901
rect 216 62867 220 62901
rect 186 62790 220 62824
rect 282 62821 292 62933
rect 318 62926 335 62936
rect 318 62857 324 62926
rect 346 62857 348 62942
rect 428 62899 430 62946
rect 476 62909 480 62977
rect 485 62959 495 62987
rect 505 62987 519 62993
rect 544 62987 555 63025
rect 505 62959 525 62987
rect 544 62959 553 62987
rect 544 62939 548 62959
rect 579 62918 582 63008
rect 612 62990 624 62991
rect 599 62988 649 62990
rect 612 62987 624 62988
rect 610 62980 632 62987
rect 607 62979 632 62980
rect 586 62972 644 62979
rect 607 62971 644 62972
rect 607 62955 610 62971
rect 616 62955 644 62971
rect 607 62954 644 62955
rect 586 62947 644 62954
rect 607 62946 610 62947
rect 612 62939 632 62947
rect 612 62935 624 62939
rect 649 62938 651 62988
rect 544 62901 548 62909
rect 400 62869 408 62899
rect 420 62869 436 62899
rect 400 62865 436 62869
rect 400 62857 430 62865
rect 428 62841 430 62857
rect 476 62829 480 62897
rect 544 62867 552 62901
rect 578 62867 582 62901
rect 544 62859 548 62867
rect 544 62829 586 62830
rect 288 62789 292 62821
rect 296 62819 368 62827
rect 378 62819 450 62827
rect 544 62822 548 62829
rect 439 62791 444 62819
rect 120 62775 170 62777
rect 76 62771 130 62775
rect 110 62766 130 62771
rect 60 62741 67 62751
rect 76 62741 77 62761
rect 96 62732 99 62766
rect 109 62741 110 62761
rect 119 62741 126 62751
rect 76 62725 92 62731
rect 94 62725 110 62731
rect 170 62725 172 62775
rect 186 62709 190 62743
rect 216 62709 220 62743
rect 213 62677 224 62709
rect 282 62705 292 62789
rect 296 62783 368 62791
rect 378 62783 450 62791
rect 468 62788 473 62822
rect 428 62753 430 62769
rect 251 62677 292 62705
rect 318 62684 324 62753
rect 12 62672 62 62674
rect 28 62663 59 62671
rect 62 62663 64 62672
rect 251 62671 263 62677
rect 28 62655 64 62663
rect 127 62663 158 62671
rect 127 62656 182 62663
rect 127 62655 161 62656
rect 59 62639 64 62655
rect 158 62639 161 62655
rect 253 62643 263 62671
rect 273 62643 293 62677
rect 318 62674 335 62684
rect 303 62658 316 62668
rect 318 62658 324 62674
rect 346 62668 348 62753
rect 400 62745 430 62753
rect 476 62751 480 62819
rect 511 62788 582 62822
rect 544 62781 548 62788
rect 400 62741 436 62745
rect 400 62711 408 62741
rect 420 62711 436 62741
rect 544 62743 548 62751
rect 28 62631 64 62639
rect 127 62638 161 62639
rect 127 62631 182 62638
rect 62 62622 64 62631
rect 282 62585 292 62643
rect 295 62634 324 62658
rect 333 62658 353 62668
rect 428 62664 430 62711
rect 476 62671 480 62739
rect 544 62709 552 62743
rect 578 62709 582 62743
rect 544 62701 548 62709
rect 367 62658 380 62664
rect 333 62634 380 62658
rect 318 62621 324 62634
rect 346 62621 348 62634
rect 367 62630 380 62634
rect 396 62630 408 62664
rect 420 62630 436 62664
rect 544 62661 553 62689
rect 319 62610 346 62621
rect 120 62569 170 62571
rect 76 62563 92 62569
rect 94 62563 110 62569
rect 76 62553 99 62562
rect 60 62543 67 62553
rect 76 62533 77 62553
rect 96 62528 99 62553
rect 109 62533 110 62553
rect 119 62543 126 62553
rect 76 62519 110 62523
rect 170 62519 172 62569
rect 186 62551 190 62585
rect 216 62551 220 62585
rect 182 62513 224 62514
rect 186 62489 220 62506
rect 223 62489 257 62506
rect 182 62472 257 62489
rect 182 62471 224 62472
rect 160 62465 246 62471
rect 288 62465 292 62585
rect 296 62583 368 62591
rect 428 62583 430 62630
rect 476 62593 480 62661
rect 485 62617 495 62651
rect 505 62623 525 62651
rect 505 62617 519 62623
rect 544 62617 555 62661
rect 485 62593 492 62617
rect 579 62602 582 62692
rect 612 62674 624 62675
rect 599 62672 649 62674
rect 612 62671 624 62672
rect 610 62664 632 62671
rect 607 62663 632 62664
rect 586 62656 644 62663
rect 607 62655 644 62656
rect 607 62639 610 62655
rect 616 62639 644 62655
rect 607 62638 644 62639
rect 586 62631 644 62638
rect 607 62630 610 62631
rect 612 62623 632 62631
rect 612 62619 624 62623
rect 649 62622 651 62672
rect 544 62585 548 62593
rect 400 62553 408 62583
rect 420 62553 436 62583
rect 400 62549 436 62553
rect 400 62541 430 62549
rect 428 62525 430 62541
rect 476 62513 480 62581
rect 544 62551 552 62585
rect 578 62551 582 62585
rect 544 62543 548 62551
rect 295 62472 300 62506
rect 324 62472 329 62506
rect 378 62503 450 62511
rect 544 62508 548 62513
rect 544 62504 582 62508
rect 544 62489 552 62504
rect 578 62489 582 62504
rect 544 62471 586 62489
rect 522 62465 608 62471
rect 182 62449 224 62465
rect 544 62449 586 62465
rect 17 62435 67 62437
rect 119 62435 169 62437
rect 186 62435 220 62449
rect 548 62435 582 62449
rect 599 62435 649 62437
rect 42 62393 59 62427
rect 67 62385 69 62435
rect 160 62427 246 62435
rect 522 62427 608 62435
rect 76 62393 110 62427
rect 127 62393 144 62427
rect 152 62393 161 62427
rect 162 62425 195 62427
rect 224 62425 244 62427
rect 162 62393 244 62425
rect 524 62425 548 62427
rect 573 62425 582 62427
rect 586 62425 606 62427
rect 160 62385 246 62393
rect 186 62369 220 62385
rect 182 62355 224 62356
rect 160 62349 182 62355
rect 224 62349 246 62355
rect 186 62314 220 62348
rect 223 62314 257 62348
rect 120 62301 170 62303
rect 76 62297 130 62301
rect 110 62292 130 62297
rect 60 62267 67 62277
rect 76 62267 77 62287
rect 96 62258 99 62292
rect 109 62267 110 62287
rect 119 62267 126 62277
rect 76 62251 92 62257
rect 94 62251 110 62257
rect 170 62251 172 62301
rect 186 62235 190 62269
rect 216 62235 220 62269
rect 288 62235 292 62423
rect 476 62355 480 62423
rect 524 62393 606 62425
rect 607 62393 616 62427
rect 522 62385 608 62393
rect 649 62385 651 62435
rect 548 62369 582 62385
rect 522 62350 548 62355
rect 522 62349 582 62350
rect 586 62349 608 62355
rect 295 62314 300 62348
rect 324 62314 329 62348
rect 544 62346 582 62349
rect 378 62309 450 62317
rect 428 62279 430 62295
rect 400 62271 430 62279
rect 476 62277 480 62345
rect 544 62316 552 62346
rect 578 62316 582 62346
rect 544 62307 548 62316
rect 400 62267 436 62271
rect 400 62237 408 62267
rect 420 62237 436 62267
rect 544 62269 548 62277
rect 12 62198 62 62200
rect 28 62189 59 62197
rect 62 62189 64 62198
rect 28 62181 64 62189
rect 127 62189 158 62197
rect 127 62182 182 62189
rect 215 62187 224 62215
rect 127 62181 161 62182
rect 59 62165 64 62181
rect 158 62165 161 62181
rect 28 62157 64 62165
rect 127 62164 161 62165
rect 127 62157 182 62164
rect 62 62148 64 62157
rect 213 62149 224 62187
rect 282 62177 292 62235
rect 296 62229 368 62237
rect 319 62199 346 62210
rect 318 62186 324 62199
rect 346 62186 348 62199
rect 428 62190 430 62237
rect 443 62227 450 62229
rect 476 62197 480 62265
rect 544 62235 552 62269
rect 578 62235 582 62269
rect 481 62203 517 62231
rect 481 62197 495 62203
rect 367 62186 380 62190
rect 251 62143 263 62177
rect 273 62143 293 62177
rect 295 62162 324 62186
rect 303 62152 316 62162
rect 318 62146 324 62162
rect 333 62162 380 62186
rect 333 62152 353 62162
rect 367 62156 380 62162
rect 396 62156 408 62190
rect 420 62156 436 62190
rect 120 62095 170 62097
rect 76 62089 92 62095
rect 94 62089 110 62095
rect 76 62079 99 62088
rect 60 62069 67 62079
rect 76 62059 77 62079
rect 96 62054 99 62079
rect 109 62059 110 62079
rect 119 62069 126 62079
rect 76 62045 110 62049
rect 170 62045 172 62095
rect 186 62077 190 62111
rect 216 62077 220 62111
rect 186 62000 220 62034
rect 282 62031 292 62143
rect 318 62136 335 62146
rect 318 62067 324 62136
rect 346 62067 348 62152
rect 428 62109 430 62156
rect 476 62119 480 62187
rect 485 62169 495 62197
rect 505 62197 519 62203
rect 544 62197 555 62235
rect 505 62169 525 62197
rect 544 62169 553 62197
rect 544 62149 548 62169
rect 579 62128 582 62218
rect 612 62200 624 62201
rect 599 62198 649 62200
rect 612 62197 624 62198
rect 610 62190 632 62197
rect 607 62189 632 62190
rect 586 62182 644 62189
rect 607 62181 644 62182
rect 607 62165 610 62181
rect 616 62165 644 62181
rect 607 62164 644 62165
rect 586 62157 644 62164
rect 607 62156 610 62157
rect 612 62149 632 62157
rect 612 62145 624 62149
rect 649 62148 651 62198
rect 544 62111 548 62119
rect 400 62079 408 62109
rect 420 62079 436 62109
rect 400 62075 436 62079
rect 400 62067 430 62075
rect 428 62051 430 62067
rect 476 62039 480 62107
rect 544 62077 552 62111
rect 578 62077 582 62111
rect 544 62069 548 62077
rect 544 62039 586 62040
rect 288 61999 292 62031
rect 296 62029 368 62037
rect 378 62029 450 62037
rect 544 62032 548 62039
rect 439 62001 444 62029
rect 120 61985 170 61987
rect 76 61981 130 61985
rect 110 61976 130 61981
rect 60 61951 67 61961
rect 76 61951 77 61971
rect 96 61942 99 61976
rect 109 61951 110 61971
rect 119 61951 126 61961
rect 76 61935 92 61941
rect 94 61935 110 61941
rect 170 61935 172 61985
rect 186 61919 190 61953
rect 216 61919 220 61953
rect 213 61887 224 61919
rect 282 61915 292 61999
rect 296 61993 368 62001
rect 378 61993 450 62001
rect 468 61998 473 62032
rect 428 61963 430 61979
rect 251 61887 292 61915
rect 318 61894 324 61963
rect 12 61882 62 61884
rect 28 61873 59 61881
rect 62 61873 64 61882
rect 251 61881 263 61887
rect 28 61865 64 61873
rect 127 61873 158 61881
rect 127 61866 182 61873
rect 127 61865 161 61866
rect 59 61849 64 61865
rect 158 61849 161 61865
rect 253 61853 263 61881
rect 273 61853 293 61887
rect 318 61884 335 61894
rect 303 61868 316 61878
rect 318 61868 324 61884
rect 346 61878 348 61963
rect 400 61955 430 61963
rect 476 61961 480 62029
rect 511 61998 582 62032
rect 544 61991 548 61998
rect 400 61951 436 61955
rect 400 61921 408 61951
rect 420 61921 436 61951
rect 544 61953 548 61961
rect 28 61841 64 61849
rect 127 61848 161 61849
rect 127 61841 182 61848
rect 62 61832 64 61841
rect 282 61795 292 61853
rect 295 61844 324 61868
rect 333 61868 353 61878
rect 428 61874 430 61921
rect 476 61881 480 61949
rect 544 61919 552 61953
rect 578 61919 582 61953
rect 544 61911 548 61919
rect 367 61868 380 61874
rect 333 61844 380 61868
rect 318 61831 324 61844
rect 346 61831 348 61844
rect 367 61840 380 61844
rect 396 61840 408 61874
rect 420 61840 436 61874
rect 544 61871 553 61899
rect 319 61820 346 61831
rect 120 61779 170 61781
rect 76 61773 92 61779
rect 94 61773 110 61779
rect 76 61763 99 61772
rect 60 61753 67 61763
rect 76 61743 77 61763
rect 96 61738 99 61763
rect 109 61743 110 61763
rect 119 61753 126 61763
rect 76 61729 110 61733
rect 170 61729 172 61779
rect 186 61761 190 61795
rect 216 61761 220 61795
rect 182 61723 224 61724
rect 186 61699 220 61716
rect 223 61699 257 61716
rect 182 61682 257 61699
rect 182 61681 224 61682
rect 160 61675 246 61681
rect 288 61675 292 61795
rect 296 61793 368 61801
rect 428 61793 430 61840
rect 476 61803 480 61871
rect 485 61827 495 61861
rect 505 61833 525 61861
rect 505 61827 519 61833
rect 544 61827 555 61871
rect 485 61803 492 61827
rect 579 61812 582 61902
rect 612 61884 624 61885
rect 599 61882 649 61884
rect 612 61881 624 61882
rect 610 61874 632 61881
rect 607 61873 632 61874
rect 586 61866 644 61873
rect 607 61865 644 61866
rect 607 61849 610 61865
rect 616 61849 644 61865
rect 607 61848 644 61849
rect 586 61841 644 61848
rect 607 61840 610 61841
rect 612 61833 632 61841
rect 612 61829 624 61833
rect 649 61832 651 61882
rect 544 61795 548 61803
rect 400 61763 408 61793
rect 420 61763 436 61793
rect 400 61759 436 61763
rect 400 61751 430 61759
rect 428 61735 430 61751
rect 476 61723 480 61791
rect 544 61761 552 61795
rect 578 61761 582 61795
rect 544 61753 548 61761
rect 295 61682 300 61716
rect 324 61682 329 61716
rect 378 61713 450 61721
rect 544 61718 548 61723
rect 544 61714 582 61718
rect 544 61699 552 61714
rect 578 61699 582 61714
rect 544 61681 586 61699
rect 522 61675 608 61681
rect 182 61659 224 61675
rect 544 61659 586 61675
rect 17 61645 67 61647
rect 119 61645 169 61647
rect 186 61645 220 61659
rect 548 61645 582 61659
rect 599 61645 649 61647
rect 42 61603 59 61637
rect 67 61595 69 61645
rect 160 61637 246 61645
rect 522 61637 608 61645
rect 76 61603 110 61637
rect 127 61603 144 61637
rect 152 61603 161 61637
rect 162 61635 195 61637
rect 224 61635 244 61637
rect 162 61603 244 61635
rect 524 61635 548 61637
rect 573 61635 582 61637
rect 586 61635 606 61637
rect 160 61595 246 61603
rect 186 61579 220 61595
rect 182 61565 224 61566
rect 160 61559 182 61565
rect 224 61559 246 61565
rect 186 61524 220 61558
rect 223 61524 257 61558
rect 120 61511 170 61513
rect 76 61507 130 61511
rect 110 61502 130 61507
rect 60 61477 67 61487
rect 76 61477 77 61497
rect 96 61468 99 61502
rect 109 61477 110 61497
rect 119 61477 126 61487
rect 76 61461 92 61467
rect 94 61461 110 61467
rect 170 61461 172 61511
rect 186 61445 190 61479
rect 216 61445 220 61479
rect 288 61445 292 61633
rect 476 61565 480 61633
rect 524 61603 606 61635
rect 607 61603 616 61637
rect 522 61595 608 61603
rect 649 61595 651 61645
rect 548 61579 582 61595
rect 522 61560 548 61565
rect 522 61559 582 61560
rect 586 61559 608 61565
rect 295 61524 300 61558
rect 324 61524 329 61558
rect 544 61556 582 61559
rect 378 61519 450 61527
rect 428 61489 430 61505
rect 400 61481 430 61489
rect 476 61487 480 61555
rect 544 61526 552 61556
rect 578 61526 582 61556
rect 544 61517 548 61526
rect 400 61477 436 61481
rect 400 61447 408 61477
rect 420 61447 436 61477
rect 544 61479 548 61487
rect 12 61408 62 61410
rect 28 61399 59 61407
rect 62 61399 64 61408
rect 28 61391 64 61399
rect 127 61399 158 61407
rect 127 61392 182 61399
rect 215 61397 224 61425
rect 127 61391 161 61392
rect 59 61375 64 61391
rect 158 61375 161 61391
rect 28 61367 64 61375
rect 127 61374 161 61375
rect 127 61367 182 61374
rect 62 61358 64 61367
rect 213 61359 224 61397
rect 282 61387 292 61445
rect 296 61439 368 61447
rect 319 61409 346 61420
rect 318 61396 324 61409
rect 346 61396 348 61409
rect 428 61400 430 61447
rect 443 61437 450 61439
rect 476 61407 480 61475
rect 544 61445 552 61479
rect 578 61445 582 61479
rect 481 61413 517 61441
rect 481 61407 495 61413
rect 367 61396 380 61400
rect 251 61353 263 61387
rect 273 61353 293 61387
rect 295 61372 324 61396
rect 303 61362 316 61372
rect 318 61356 324 61372
rect 333 61372 380 61396
rect 333 61362 353 61372
rect 367 61366 380 61372
rect 396 61366 408 61400
rect 420 61366 436 61400
rect 120 61305 170 61307
rect 76 61299 92 61305
rect 94 61299 110 61305
rect 76 61289 99 61298
rect 60 61279 67 61289
rect 76 61269 77 61289
rect 96 61264 99 61289
rect 109 61269 110 61289
rect 119 61279 126 61289
rect 76 61255 110 61259
rect 170 61255 172 61305
rect 186 61287 190 61321
rect 216 61287 220 61321
rect 186 61210 220 61244
rect 282 61241 292 61353
rect 318 61346 335 61356
rect 318 61277 324 61346
rect 346 61277 348 61362
rect 428 61319 430 61366
rect 476 61329 480 61397
rect 485 61379 495 61407
rect 505 61407 519 61413
rect 544 61407 555 61445
rect 505 61379 525 61407
rect 544 61379 553 61407
rect 544 61359 548 61379
rect 579 61338 582 61428
rect 612 61410 624 61411
rect 599 61408 649 61410
rect 612 61407 624 61408
rect 610 61400 632 61407
rect 607 61399 632 61400
rect 586 61392 644 61399
rect 607 61391 644 61392
rect 607 61375 610 61391
rect 616 61375 644 61391
rect 607 61374 644 61375
rect 586 61367 644 61374
rect 607 61366 610 61367
rect 612 61359 632 61367
rect 612 61355 624 61359
rect 649 61358 651 61408
rect 544 61321 548 61329
rect 400 61289 408 61319
rect 420 61289 436 61319
rect 400 61285 436 61289
rect 400 61277 430 61285
rect 428 61261 430 61277
rect 476 61249 480 61317
rect 544 61287 552 61321
rect 578 61287 582 61321
rect 544 61279 548 61287
rect 544 61249 586 61250
rect 288 61209 292 61241
rect 296 61239 368 61247
rect 378 61239 450 61247
rect 544 61242 548 61249
rect 439 61211 444 61239
rect 120 61195 170 61197
rect 76 61191 130 61195
rect 110 61186 130 61191
rect 60 61161 67 61171
rect 76 61161 77 61181
rect 96 61152 99 61186
rect 109 61161 110 61181
rect 119 61161 126 61171
rect 76 61145 92 61151
rect 94 61145 110 61151
rect 170 61145 172 61195
rect 186 61129 190 61163
rect 216 61129 220 61163
rect 213 61097 224 61129
rect 282 61125 292 61209
rect 296 61203 368 61211
rect 378 61203 450 61211
rect 468 61208 473 61242
rect 428 61173 430 61189
rect 251 61097 292 61125
rect 318 61104 324 61173
rect 12 61092 62 61094
rect 28 61083 59 61091
rect 62 61083 64 61092
rect 251 61091 263 61097
rect 28 61075 64 61083
rect 127 61083 158 61091
rect 127 61076 182 61083
rect 127 61075 161 61076
rect 59 61059 64 61075
rect 158 61059 161 61075
rect 253 61063 263 61091
rect 273 61063 293 61097
rect 318 61094 335 61104
rect 303 61078 316 61088
rect 318 61078 324 61094
rect 346 61088 348 61173
rect 400 61165 430 61173
rect 476 61171 480 61239
rect 511 61208 582 61242
rect 544 61201 548 61208
rect 400 61161 436 61165
rect 400 61131 408 61161
rect 420 61131 436 61161
rect 544 61163 548 61171
rect 28 61051 64 61059
rect 127 61058 161 61059
rect 127 61051 182 61058
rect 62 61042 64 61051
rect 282 61005 292 61063
rect 295 61054 324 61078
rect 333 61078 353 61088
rect 428 61084 430 61131
rect 476 61091 480 61159
rect 544 61129 552 61163
rect 578 61129 582 61163
rect 544 61121 548 61129
rect 367 61078 380 61084
rect 333 61054 380 61078
rect 318 61041 324 61054
rect 346 61041 348 61054
rect 367 61050 380 61054
rect 396 61050 408 61084
rect 420 61050 436 61084
rect 544 61081 553 61109
rect 319 61030 346 61041
rect 120 60989 170 60991
rect 76 60983 92 60989
rect 94 60983 110 60989
rect 76 60973 99 60982
rect 60 60963 67 60973
rect 76 60953 77 60973
rect 96 60948 99 60973
rect 109 60953 110 60973
rect 119 60963 126 60973
rect 76 60939 110 60943
rect 170 60939 172 60989
rect 186 60971 190 61005
rect 216 60971 220 61005
rect 182 60933 224 60934
rect 186 60909 220 60926
rect 223 60909 257 60926
rect 182 60892 257 60909
rect 182 60891 224 60892
rect 160 60885 246 60891
rect 288 60885 292 61005
rect 296 61003 368 61011
rect 428 61003 430 61050
rect 476 61013 480 61081
rect 485 61037 495 61071
rect 505 61043 525 61071
rect 505 61037 519 61043
rect 544 61037 555 61081
rect 485 61013 492 61037
rect 579 61022 582 61112
rect 612 61094 624 61095
rect 599 61092 649 61094
rect 612 61091 624 61092
rect 610 61084 632 61091
rect 607 61083 632 61084
rect 586 61076 644 61083
rect 607 61075 644 61076
rect 607 61059 610 61075
rect 616 61059 644 61075
rect 607 61058 644 61059
rect 586 61051 644 61058
rect 607 61050 610 61051
rect 612 61043 632 61051
rect 612 61039 624 61043
rect 649 61042 651 61092
rect 544 61005 548 61013
rect 400 60973 408 61003
rect 420 60973 436 61003
rect 400 60969 436 60973
rect 400 60961 430 60969
rect 428 60945 430 60961
rect 476 60933 480 61001
rect 544 60971 552 61005
rect 578 60971 582 61005
rect 544 60963 548 60971
rect 295 60892 300 60926
rect 324 60892 329 60926
rect 378 60923 450 60931
rect 544 60928 548 60933
rect 544 60924 582 60928
rect 544 60909 552 60924
rect 578 60909 582 60924
rect 544 60891 586 60909
rect 522 60885 608 60891
rect 182 60869 224 60885
rect 544 60869 586 60885
rect 17 60855 67 60857
rect 119 60855 169 60857
rect 186 60855 220 60869
rect 548 60855 582 60869
rect 599 60855 649 60857
rect 42 60813 59 60847
rect 67 60805 69 60855
rect 160 60847 246 60855
rect 522 60847 608 60855
rect 76 60813 110 60847
rect 127 60813 144 60847
rect 152 60813 161 60847
rect 162 60845 195 60847
rect 224 60845 244 60847
rect 162 60813 244 60845
rect 524 60845 548 60847
rect 573 60845 582 60847
rect 586 60845 606 60847
rect 160 60805 246 60813
rect 186 60789 220 60805
rect 182 60775 224 60776
rect 160 60769 182 60775
rect 224 60769 246 60775
rect 186 60734 220 60768
rect 223 60734 257 60768
rect 120 60721 170 60723
rect 76 60717 130 60721
rect 110 60712 130 60717
rect 60 60687 67 60697
rect 76 60687 77 60707
rect 96 60678 99 60712
rect 109 60687 110 60707
rect 119 60687 126 60697
rect 76 60671 92 60677
rect 94 60671 110 60677
rect 170 60671 172 60721
rect 186 60655 190 60689
rect 216 60655 220 60689
rect 288 60655 292 60843
rect 476 60775 480 60843
rect 524 60813 606 60845
rect 607 60813 616 60847
rect 522 60805 608 60813
rect 649 60805 651 60855
rect 548 60789 582 60805
rect 522 60770 548 60775
rect 522 60769 582 60770
rect 586 60769 608 60775
rect 295 60734 300 60768
rect 324 60734 329 60768
rect 544 60766 582 60769
rect 378 60729 450 60737
rect 428 60699 430 60715
rect 400 60691 430 60699
rect 476 60697 480 60765
rect 544 60736 552 60766
rect 578 60736 582 60766
rect 544 60727 548 60736
rect 400 60687 436 60691
rect 400 60657 408 60687
rect 420 60657 436 60687
rect 544 60689 548 60697
rect 12 60618 62 60620
rect 28 60609 59 60617
rect 62 60609 64 60618
rect 28 60601 64 60609
rect 127 60609 158 60617
rect 127 60602 182 60609
rect 215 60607 224 60635
rect 127 60601 161 60602
rect 59 60585 64 60601
rect 158 60585 161 60601
rect 28 60577 64 60585
rect 127 60584 161 60585
rect 127 60577 182 60584
rect 62 60568 64 60577
rect 213 60569 224 60607
rect 282 60597 292 60655
rect 296 60649 368 60657
rect 319 60619 346 60630
rect 318 60606 324 60619
rect 346 60606 348 60619
rect 428 60610 430 60657
rect 443 60647 450 60649
rect 476 60617 480 60685
rect 544 60655 552 60689
rect 578 60655 582 60689
rect 481 60623 517 60651
rect 481 60617 495 60623
rect 367 60606 380 60610
rect 251 60563 263 60597
rect 273 60563 293 60597
rect 295 60582 324 60606
rect 303 60572 316 60582
rect 318 60566 324 60582
rect 333 60582 380 60606
rect 333 60572 353 60582
rect 367 60576 380 60582
rect 396 60576 408 60610
rect 420 60576 436 60610
rect 120 60515 170 60517
rect 76 60509 92 60515
rect 94 60509 110 60515
rect 76 60499 99 60508
rect 60 60489 67 60499
rect 76 60480 77 60499
rect 96 60474 99 60499
rect 109 60480 110 60499
rect 119 60489 126 60499
rect 76 60465 110 60469
rect 170 60465 172 60515
rect 186 60497 190 60531
rect 216 60497 220 60531
rect 186 60420 220 60454
rect 282 60451 292 60563
rect 318 60556 335 60566
rect 318 60487 324 60556
rect 346 60487 348 60572
rect 428 60529 430 60576
rect 476 60539 480 60607
rect 485 60589 495 60617
rect 505 60617 519 60623
rect 544 60617 555 60655
rect 505 60589 525 60617
rect 544 60589 553 60617
rect 544 60569 548 60589
rect 579 60548 582 60638
rect 612 60620 624 60621
rect 599 60618 649 60620
rect 612 60617 624 60618
rect 610 60610 632 60617
rect 607 60609 632 60610
rect 586 60602 644 60609
rect 607 60601 644 60602
rect 607 60585 610 60601
rect 616 60585 644 60601
rect 607 60584 644 60585
rect 586 60577 644 60584
rect 607 60576 610 60577
rect 612 60569 632 60577
rect 612 60565 624 60569
rect 649 60568 651 60618
rect 544 60531 548 60539
rect 400 60499 408 60529
rect 420 60499 436 60529
rect 400 60495 436 60499
rect 400 60487 430 60495
rect 428 60471 430 60487
rect 476 60459 480 60527
rect 544 60497 552 60531
rect 578 60497 582 60531
rect 544 60489 548 60497
rect 544 60459 586 60460
rect 288 60419 292 60451
rect 296 60449 368 60457
rect 378 60449 450 60457
rect 544 60452 548 60459
rect 439 60421 444 60449
rect 120 60405 170 60407
rect 76 60401 130 60405
rect 110 60396 130 60401
rect 60 60371 67 60381
rect 76 60371 77 60391
rect 96 60362 99 60396
rect 109 60371 110 60391
rect 119 60371 126 60381
rect 76 60355 92 60361
rect 94 60355 110 60361
rect 170 60355 172 60405
rect 186 60339 190 60373
rect 216 60339 220 60373
rect 213 60307 224 60339
rect 282 60335 292 60419
rect 296 60413 368 60421
rect 378 60413 450 60421
rect 468 60418 473 60452
rect 428 60383 430 60399
rect 251 60307 292 60335
rect 318 60314 324 60383
rect 12 60302 62 60304
rect 28 60293 59 60301
rect 62 60293 64 60302
rect 251 60301 263 60307
rect 28 60285 64 60293
rect 127 60293 158 60301
rect 127 60286 182 60293
rect 127 60285 161 60286
rect 59 60269 64 60285
rect 158 60269 161 60285
rect 253 60273 263 60301
rect 273 60273 293 60307
rect 318 60304 335 60314
rect 303 60288 316 60298
rect 318 60288 324 60304
rect 346 60298 348 60383
rect 400 60375 430 60383
rect 476 60381 480 60449
rect 511 60418 582 60452
rect 544 60411 548 60418
rect 400 60371 436 60375
rect 400 60341 408 60371
rect 420 60341 436 60371
rect 544 60373 548 60381
rect 28 60261 64 60269
rect 127 60268 161 60269
rect 127 60261 182 60268
rect 62 60252 64 60261
rect 282 60215 292 60273
rect 295 60264 324 60288
rect 333 60288 353 60298
rect 428 60294 430 60341
rect 476 60301 480 60369
rect 544 60339 552 60373
rect 578 60339 582 60373
rect 544 60331 548 60339
rect 367 60288 380 60294
rect 333 60264 380 60288
rect 318 60251 324 60264
rect 346 60251 348 60264
rect 367 60260 380 60264
rect 396 60260 408 60294
rect 420 60260 436 60294
rect 544 60291 553 60319
rect 319 60240 346 60251
rect 120 60199 170 60201
rect 76 60193 92 60199
rect 94 60193 110 60199
rect 76 60183 99 60192
rect 60 60173 67 60183
rect 76 60163 77 60183
rect 96 60158 99 60183
rect 109 60163 110 60183
rect 119 60173 126 60183
rect 76 60149 110 60153
rect 170 60149 172 60199
rect 186 60181 190 60215
rect 216 60181 220 60215
rect 182 60143 224 60144
rect 186 60119 220 60136
rect 223 60119 257 60136
rect 182 60102 257 60119
rect 182 60101 224 60102
rect 160 60095 246 60101
rect 288 60095 292 60215
rect 296 60213 368 60221
rect 428 60213 430 60260
rect 476 60223 480 60291
rect 485 60247 495 60281
rect 505 60253 525 60281
rect 505 60247 519 60253
rect 544 60247 555 60291
rect 485 60223 492 60247
rect 579 60232 582 60322
rect 612 60304 624 60305
rect 599 60302 649 60304
rect 612 60301 624 60302
rect 610 60294 632 60301
rect 607 60293 632 60294
rect 586 60286 644 60293
rect 607 60285 644 60286
rect 607 60269 610 60285
rect 616 60269 644 60285
rect 607 60268 644 60269
rect 586 60261 644 60268
rect 607 60260 610 60261
rect 612 60253 632 60261
rect 612 60249 624 60253
rect 649 60252 651 60302
rect 544 60215 548 60223
rect 400 60183 408 60213
rect 420 60183 436 60213
rect 400 60179 436 60183
rect 400 60171 430 60179
rect 428 60155 430 60171
rect 476 60143 480 60211
rect 544 60181 552 60215
rect 578 60181 582 60215
rect 544 60173 548 60181
rect 295 60102 300 60136
rect 324 60102 329 60136
rect 378 60133 450 60141
rect 544 60138 548 60143
rect 544 60134 582 60138
rect 544 60119 552 60134
rect 578 60119 582 60134
rect 544 60101 586 60119
rect 522 60095 608 60101
rect 182 60079 224 60095
rect 544 60079 586 60095
rect 17 60065 67 60067
rect 119 60065 169 60067
rect 186 60065 220 60079
rect 548 60065 582 60079
rect 599 60065 649 60067
rect 42 60023 59 60057
rect 67 60015 69 60065
rect 160 60057 246 60065
rect 522 60057 608 60065
rect 76 60023 110 60057
rect 127 60023 144 60057
rect 152 60023 161 60057
rect 162 60055 195 60057
rect 224 60055 244 60057
rect 162 60023 244 60055
rect 524 60055 548 60057
rect 573 60055 582 60057
rect 586 60055 606 60057
rect 160 60015 246 60023
rect 186 59999 220 60015
rect 182 59985 224 59986
rect 160 59979 182 59985
rect 224 59979 246 59985
rect 186 59944 220 59978
rect 223 59944 257 59978
rect 120 59931 170 59933
rect 76 59927 130 59931
rect 110 59922 130 59927
rect 60 59897 67 59907
rect 76 59897 77 59917
rect 96 59888 99 59922
rect 109 59897 110 59917
rect 119 59897 126 59907
rect 76 59881 92 59887
rect 94 59881 110 59887
rect 170 59881 172 59931
rect 186 59865 190 59899
rect 216 59865 220 59899
rect 288 59865 292 60053
rect 476 59985 480 60053
rect 524 60023 606 60055
rect 607 60023 616 60057
rect 522 60015 608 60023
rect 649 60015 651 60065
rect 548 59999 582 60015
rect 522 59980 548 59985
rect 522 59979 582 59980
rect 586 59979 608 59985
rect 295 59944 300 59978
rect 324 59944 329 59978
rect 544 59976 582 59979
rect 378 59939 450 59947
rect 428 59909 430 59925
rect 400 59901 430 59909
rect 476 59907 480 59975
rect 544 59946 552 59976
rect 578 59946 582 59976
rect 544 59937 548 59946
rect 400 59897 436 59901
rect 400 59867 408 59897
rect 420 59867 436 59897
rect 544 59899 548 59907
rect 12 59828 62 59830
rect 28 59819 59 59827
rect 62 59819 64 59828
rect 28 59811 64 59819
rect 127 59819 158 59827
rect 127 59812 182 59819
rect 215 59817 224 59845
rect 127 59811 161 59812
rect 59 59795 64 59811
rect 158 59795 161 59811
rect 28 59787 64 59795
rect 127 59794 161 59795
rect 127 59787 182 59794
rect 62 59778 64 59787
rect 213 59779 224 59817
rect 282 59807 292 59865
rect 296 59859 368 59867
rect 319 59829 346 59840
rect 318 59816 324 59829
rect 346 59816 348 59829
rect 428 59820 430 59867
rect 443 59857 450 59859
rect 476 59827 480 59895
rect 544 59865 552 59899
rect 578 59865 582 59899
rect 481 59833 517 59861
rect 481 59827 495 59833
rect 367 59816 380 59820
rect 251 59773 263 59807
rect 273 59773 293 59807
rect 295 59792 324 59816
rect 303 59782 316 59792
rect 318 59776 324 59792
rect 333 59792 380 59816
rect 333 59782 353 59792
rect 367 59786 380 59792
rect 396 59786 408 59820
rect 420 59786 436 59820
rect 120 59725 170 59727
rect 76 59719 92 59725
rect 94 59719 110 59725
rect 76 59709 99 59718
rect 60 59699 67 59709
rect 76 59689 77 59709
rect 96 59684 99 59709
rect 109 59689 110 59709
rect 119 59699 126 59709
rect 76 59675 110 59679
rect 170 59675 172 59725
rect 186 59707 190 59741
rect 216 59707 220 59741
rect 186 59630 220 59664
rect 282 59661 292 59773
rect 318 59766 335 59776
rect 318 59697 324 59766
rect 346 59697 348 59782
rect 428 59739 430 59786
rect 476 59749 480 59817
rect 485 59799 495 59827
rect 505 59827 519 59833
rect 544 59827 555 59865
rect 505 59799 525 59827
rect 544 59799 553 59827
rect 544 59779 548 59799
rect 579 59758 582 59848
rect 612 59830 624 59831
rect 599 59828 649 59830
rect 612 59827 624 59828
rect 610 59820 632 59827
rect 607 59819 632 59820
rect 586 59812 644 59819
rect 607 59811 644 59812
rect 607 59795 610 59811
rect 616 59795 644 59811
rect 607 59794 644 59795
rect 586 59787 644 59794
rect 607 59786 610 59787
rect 612 59779 632 59787
rect 612 59775 624 59779
rect 649 59778 651 59828
rect 544 59741 548 59749
rect 400 59709 408 59739
rect 420 59709 436 59739
rect 400 59705 436 59709
rect 400 59697 430 59705
rect 428 59681 430 59697
rect 476 59669 480 59737
rect 544 59707 552 59741
rect 578 59707 582 59741
rect 544 59699 548 59707
rect 544 59669 586 59670
rect 288 59629 292 59661
rect 296 59659 368 59667
rect 378 59659 450 59667
rect 544 59662 548 59669
rect 439 59631 444 59659
rect 120 59615 170 59617
rect 76 59611 130 59615
rect 110 59606 130 59611
rect 60 59581 67 59591
rect 76 59581 77 59601
rect 96 59572 99 59606
rect 109 59581 110 59601
rect 119 59581 126 59591
rect 76 59565 92 59571
rect 94 59565 110 59571
rect 170 59565 172 59615
rect 186 59549 190 59583
rect 216 59549 220 59583
rect 213 59517 224 59549
rect 282 59545 292 59629
rect 296 59623 368 59631
rect 378 59623 450 59631
rect 468 59628 473 59662
rect 428 59593 430 59609
rect 251 59517 292 59545
rect 318 59524 324 59593
rect 12 59512 62 59514
rect 28 59503 59 59511
rect 62 59503 64 59512
rect 251 59511 263 59517
rect 28 59495 64 59503
rect 127 59503 158 59511
rect 127 59496 182 59503
rect 127 59495 161 59496
rect 59 59479 64 59495
rect 158 59479 161 59495
rect 253 59483 263 59511
rect 273 59483 293 59517
rect 318 59514 335 59524
rect 303 59498 316 59508
rect 318 59498 324 59514
rect 346 59508 348 59593
rect 400 59585 430 59593
rect 476 59591 480 59659
rect 511 59628 582 59662
rect 544 59621 548 59628
rect 400 59581 436 59585
rect 400 59551 408 59581
rect 420 59551 436 59581
rect 544 59583 548 59591
rect 28 59471 64 59479
rect 127 59478 161 59479
rect 127 59471 182 59478
rect 62 59462 64 59471
rect 282 59425 292 59483
rect 295 59474 324 59498
rect 333 59498 353 59508
rect 428 59504 430 59551
rect 476 59511 480 59579
rect 544 59549 552 59583
rect 578 59549 582 59583
rect 544 59541 548 59549
rect 367 59498 380 59504
rect 333 59474 380 59498
rect 318 59461 324 59474
rect 346 59461 348 59474
rect 367 59470 380 59474
rect 396 59470 408 59504
rect 420 59470 436 59504
rect 544 59501 553 59529
rect 319 59450 346 59461
rect 120 59409 170 59411
rect 76 59403 92 59409
rect 94 59403 110 59409
rect 76 59393 99 59402
rect 60 59383 67 59393
rect 76 59373 77 59393
rect 96 59368 99 59393
rect 109 59373 110 59393
rect 119 59383 126 59393
rect 76 59359 110 59363
rect 170 59359 172 59409
rect 186 59391 190 59425
rect 216 59391 220 59425
rect 182 59353 224 59354
rect 186 59329 220 59346
rect 223 59329 257 59346
rect 182 59312 257 59329
rect 182 59311 224 59312
rect 160 59305 246 59311
rect 288 59305 292 59425
rect 296 59423 368 59431
rect 428 59423 430 59470
rect 476 59433 480 59501
rect 485 59457 495 59491
rect 505 59463 525 59491
rect 505 59457 519 59463
rect 544 59457 555 59501
rect 485 59433 492 59457
rect 579 59442 582 59532
rect 612 59514 624 59515
rect 599 59512 649 59514
rect 612 59511 624 59512
rect 610 59504 632 59511
rect 607 59503 632 59504
rect 586 59496 644 59503
rect 607 59495 644 59496
rect 607 59479 610 59495
rect 616 59479 644 59495
rect 607 59478 644 59479
rect 586 59471 644 59478
rect 607 59470 610 59471
rect 612 59463 632 59471
rect 612 59459 624 59463
rect 649 59462 651 59512
rect 544 59425 548 59433
rect 400 59393 408 59423
rect 420 59393 436 59423
rect 400 59389 436 59393
rect 400 59381 430 59389
rect 428 59365 430 59381
rect 476 59353 480 59421
rect 544 59391 552 59425
rect 578 59391 582 59425
rect 544 59383 548 59391
rect 295 59312 300 59346
rect 324 59312 329 59346
rect 378 59343 450 59351
rect 544 59348 548 59353
rect 544 59344 582 59348
rect 544 59329 552 59344
rect 578 59329 582 59344
rect 544 59311 586 59329
rect 522 59305 608 59311
rect 182 59289 224 59305
rect 544 59289 586 59305
rect 17 59275 67 59277
rect 119 59275 169 59277
rect 186 59275 220 59289
rect 548 59275 582 59289
rect 599 59275 649 59277
rect 42 59233 59 59267
rect 67 59225 69 59275
rect 160 59267 246 59275
rect 522 59267 608 59275
rect 76 59233 110 59267
rect 127 59233 144 59267
rect 152 59233 161 59267
rect 162 59265 195 59267
rect 224 59265 244 59267
rect 162 59233 244 59265
rect 524 59265 548 59267
rect 573 59265 582 59267
rect 586 59265 606 59267
rect 160 59225 246 59233
rect 186 59209 220 59225
rect 182 59195 224 59196
rect 160 59189 182 59195
rect 224 59189 246 59195
rect 186 59154 220 59188
rect 223 59154 257 59188
rect 120 59141 170 59143
rect 76 59137 130 59141
rect 110 59132 130 59137
rect 60 59107 67 59117
rect 76 59107 77 59127
rect 96 59098 99 59132
rect 109 59107 110 59127
rect 119 59107 126 59117
rect 76 59091 92 59097
rect 94 59091 110 59097
rect 170 59091 172 59141
rect 186 59075 190 59109
rect 216 59075 220 59109
rect 288 59075 292 59263
rect 476 59195 480 59263
rect 524 59233 606 59265
rect 607 59233 616 59267
rect 522 59225 608 59233
rect 649 59225 651 59275
rect 548 59209 582 59225
rect 522 59190 548 59195
rect 522 59189 582 59190
rect 586 59189 608 59195
rect 295 59154 300 59188
rect 324 59154 329 59188
rect 544 59186 582 59189
rect 378 59149 450 59157
rect 428 59119 430 59135
rect 400 59111 430 59119
rect 476 59117 480 59185
rect 544 59156 552 59186
rect 578 59156 582 59186
rect 544 59147 548 59156
rect 400 59107 436 59111
rect 400 59077 408 59107
rect 420 59077 436 59107
rect 544 59109 548 59117
rect 12 59038 62 59040
rect 28 59029 59 59037
rect 62 59029 64 59038
rect 28 59021 64 59029
rect 127 59029 158 59037
rect 127 59022 182 59029
rect 215 59027 224 59055
rect 127 59021 161 59022
rect 59 59005 64 59021
rect 158 59005 161 59021
rect 28 58997 64 59005
rect 127 59004 161 59005
rect 127 58997 182 59004
rect 62 58988 64 58997
rect 213 58989 224 59027
rect 282 59017 292 59075
rect 296 59069 368 59077
rect 319 59039 346 59050
rect 318 59026 324 59039
rect 346 59026 348 59039
rect 428 59030 430 59077
rect 443 59067 450 59069
rect 476 59037 480 59105
rect 544 59075 552 59109
rect 578 59075 582 59109
rect 481 59043 517 59071
rect 481 59037 495 59043
rect 367 59026 380 59030
rect 251 58983 263 59017
rect 273 58983 293 59017
rect 295 59002 324 59026
rect 303 58992 316 59002
rect 318 58986 324 59002
rect 333 59002 380 59026
rect 333 58992 353 59002
rect 367 58996 380 59002
rect 396 58996 408 59030
rect 420 58996 436 59030
rect 120 58935 170 58937
rect 76 58929 92 58935
rect 94 58929 110 58935
rect 76 58919 99 58928
rect 60 58909 67 58919
rect 76 58899 77 58919
rect 96 58894 99 58919
rect 109 58899 110 58919
rect 119 58909 126 58919
rect 76 58885 110 58889
rect 170 58885 172 58935
rect 186 58917 190 58951
rect 216 58917 220 58951
rect 186 58840 220 58874
rect 282 58871 292 58983
rect 318 58976 335 58986
rect 318 58907 324 58976
rect 346 58907 348 58992
rect 428 58949 430 58996
rect 476 58959 480 59027
rect 485 59009 495 59037
rect 505 59037 519 59043
rect 544 59037 555 59075
rect 505 59009 525 59037
rect 544 59009 553 59037
rect 544 58989 548 59009
rect 579 58968 582 59058
rect 612 59040 624 59041
rect 599 59038 649 59040
rect 612 59037 624 59038
rect 610 59030 632 59037
rect 607 59029 632 59030
rect 586 59022 644 59029
rect 607 59021 644 59022
rect 607 59005 610 59021
rect 616 59005 644 59021
rect 607 59004 644 59005
rect 586 58997 644 59004
rect 607 58996 610 58997
rect 612 58989 632 58997
rect 612 58985 624 58989
rect 649 58988 651 59038
rect 544 58951 548 58959
rect 400 58919 408 58949
rect 420 58919 436 58949
rect 400 58915 436 58919
rect 400 58907 430 58915
rect 428 58891 430 58907
rect 476 58879 480 58947
rect 544 58917 552 58951
rect 578 58917 582 58951
rect 544 58909 548 58917
rect 544 58879 586 58880
rect 288 58839 292 58871
rect 296 58869 368 58877
rect 378 58869 450 58877
rect 544 58872 548 58879
rect 439 58841 444 58869
rect 120 58825 170 58827
rect 76 58821 130 58825
rect 110 58816 130 58821
rect 60 58791 67 58801
rect 76 58791 77 58811
rect 96 58782 99 58816
rect 109 58791 110 58811
rect 119 58791 126 58801
rect 76 58775 92 58781
rect 94 58775 110 58781
rect 170 58775 172 58825
rect 186 58759 190 58793
rect 216 58759 220 58793
rect 213 58727 224 58759
rect 282 58755 292 58839
rect 296 58833 368 58841
rect 378 58833 450 58841
rect 468 58838 473 58872
rect 428 58803 430 58819
rect 251 58727 292 58755
rect 318 58734 324 58803
rect 12 58722 62 58724
rect 28 58713 59 58721
rect 62 58713 64 58722
rect 251 58721 263 58727
rect 28 58705 64 58713
rect 127 58713 158 58721
rect 127 58706 182 58713
rect 127 58705 161 58706
rect 59 58689 64 58705
rect 158 58689 161 58705
rect 253 58693 263 58721
rect 273 58693 293 58727
rect 318 58724 335 58734
rect 303 58708 316 58718
rect 318 58708 324 58724
rect 346 58718 348 58803
rect 400 58795 430 58803
rect 476 58801 480 58869
rect 511 58838 582 58872
rect 544 58831 548 58838
rect 400 58791 436 58795
rect 400 58761 408 58791
rect 420 58761 436 58791
rect 544 58793 548 58801
rect 28 58681 64 58689
rect 127 58688 161 58689
rect 127 58681 182 58688
rect 62 58672 64 58681
rect 282 58635 292 58693
rect 295 58684 324 58708
rect 333 58708 353 58718
rect 428 58714 430 58761
rect 476 58721 480 58789
rect 544 58759 552 58793
rect 578 58759 582 58793
rect 544 58751 548 58759
rect 367 58708 380 58714
rect 333 58684 380 58708
rect 318 58671 324 58684
rect 346 58671 348 58684
rect 367 58680 380 58684
rect 396 58680 408 58714
rect 420 58680 436 58714
rect 544 58711 553 58739
rect 319 58660 346 58671
rect 120 58619 170 58621
rect 76 58613 92 58619
rect 94 58613 110 58619
rect 76 58603 99 58612
rect 60 58593 67 58603
rect 76 58583 77 58603
rect 96 58578 99 58603
rect 109 58583 110 58603
rect 119 58593 126 58603
rect 76 58569 110 58573
rect 170 58569 172 58619
rect 186 58601 190 58635
rect 216 58601 220 58635
rect 182 58563 224 58564
rect 186 58539 220 58556
rect 223 58539 257 58556
rect 182 58522 257 58539
rect 182 58521 224 58522
rect 160 58515 246 58521
rect 288 58515 292 58635
rect 296 58633 368 58641
rect 428 58633 430 58680
rect 476 58643 480 58711
rect 485 58667 495 58701
rect 505 58673 525 58701
rect 505 58667 519 58673
rect 544 58667 555 58711
rect 485 58643 492 58667
rect 579 58652 582 58742
rect 612 58724 624 58725
rect 599 58722 649 58724
rect 612 58721 624 58722
rect 610 58714 632 58721
rect 607 58713 632 58714
rect 586 58706 644 58713
rect 607 58705 644 58706
rect 607 58689 610 58705
rect 616 58689 644 58705
rect 607 58688 644 58689
rect 586 58681 644 58688
rect 607 58680 610 58681
rect 612 58673 632 58681
rect 612 58669 624 58673
rect 649 58672 651 58722
rect 544 58635 548 58643
rect 400 58603 408 58633
rect 420 58603 436 58633
rect 400 58599 436 58603
rect 400 58591 430 58599
rect 428 58575 430 58591
rect 476 58563 480 58631
rect 544 58601 552 58635
rect 578 58601 582 58635
rect 544 58593 548 58601
rect 295 58522 300 58556
rect 324 58522 329 58556
rect 378 58553 450 58561
rect 544 58558 548 58563
rect 544 58554 582 58558
rect 544 58539 552 58554
rect 578 58539 582 58554
rect 544 58521 586 58539
rect 522 58515 608 58521
rect 182 58499 224 58515
rect 544 58499 586 58515
rect 17 58485 67 58487
rect 119 58485 169 58487
rect 186 58485 220 58499
rect 548 58485 582 58499
rect 599 58485 649 58487
rect 42 58443 59 58477
rect 67 58435 69 58485
rect 160 58477 246 58485
rect 522 58477 608 58485
rect 76 58443 110 58477
rect 127 58443 144 58477
rect 152 58443 161 58477
rect 162 58475 195 58477
rect 224 58475 244 58477
rect 162 58443 244 58475
rect 524 58475 548 58477
rect 573 58475 582 58477
rect 586 58475 606 58477
rect 160 58435 246 58443
rect 186 58419 220 58435
rect 182 58405 224 58406
rect 160 58399 182 58405
rect 224 58399 246 58405
rect 186 58364 220 58398
rect 223 58364 257 58398
rect 120 58351 170 58353
rect 76 58347 130 58351
rect 110 58342 130 58347
rect 60 58317 67 58327
rect 76 58317 77 58337
rect 96 58308 99 58342
rect 109 58317 110 58337
rect 119 58317 126 58327
rect 76 58301 92 58307
rect 94 58301 110 58307
rect 170 58301 172 58351
rect 186 58285 190 58319
rect 216 58285 220 58319
rect 288 58285 292 58473
rect 476 58405 480 58473
rect 524 58443 606 58475
rect 607 58443 616 58477
rect 522 58435 608 58443
rect 649 58435 651 58485
rect 548 58419 582 58435
rect 522 58400 548 58405
rect 522 58399 582 58400
rect 586 58399 608 58405
rect 295 58364 300 58398
rect 324 58364 329 58398
rect 544 58396 582 58399
rect 378 58359 450 58367
rect 428 58329 430 58345
rect 400 58321 430 58329
rect 476 58327 480 58395
rect 544 58366 552 58396
rect 578 58366 582 58396
rect 544 58357 548 58366
rect 400 58317 436 58321
rect 400 58287 408 58317
rect 420 58287 436 58317
rect 544 58319 548 58327
rect 12 58248 62 58250
rect 28 58239 59 58247
rect 62 58239 64 58248
rect 28 58231 64 58239
rect 127 58239 158 58247
rect 127 58232 182 58239
rect 215 58237 224 58265
rect 127 58231 161 58232
rect 59 58215 64 58231
rect 158 58215 161 58231
rect 28 58207 64 58215
rect 127 58214 161 58215
rect 127 58207 182 58214
rect 62 58198 64 58207
rect 213 58199 224 58237
rect 282 58227 292 58285
rect 296 58279 368 58287
rect 319 58249 346 58260
rect 318 58236 324 58249
rect 346 58236 348 58249
rect 428 58240 430 58287
rect 443 58277 450 58279
rect 476 58247 480 58315
rect 544 58285 552 58319
rect 578 58285 582 58319
rect 481 58253 517 58281
rect 481 58247 495 58253
rect 367 58236 380 58240
rect 251 58193 263 58227
rect 273 58193 293 58227
rect 295 58212 324 58236
rect 303 58202 316 58212
rect 318 58196 324 58212
rect 333 58212 380 58236
rect 333 58202 353 58212
rect 367 58206 380 58212
rect 396 58206 408 58240
rect 420 58206 436 58240
rect 120 58145 170 58147
rect 76 58139 92 58145
rect 94 58139 110 58145
rect 76 58129 99 58138
rect 60 58119 67 58129
rect 76 58109 77 58129
rect 96 58104 99 58129
rect 109 58109 110 58129
rect 119 58119 126 58129
rect 76 58095 110 58099
rect 170 58095 172 58145
rect 186 58127 190 58161
rect 216 58127 220 58161
rect 186 58050 220 58084
rect 282 58081 292 58193
rect 318 58186 335 58196
rect 318 58117 324 58186
rect 346 58117 348 58202
rect 428 58159 430 58206
rect 476 58169 480 58237
rect 485 58219 495 58247
rect 505 58247 519 58253
rect 544 58247 555 58285
rect 505 58219 525 58247
rect 544 58219 553 58247
rect 544 58199 548 58219
rect 579 58178 582 58268
rect 612 58250 624 58251
rect 599 58248 649 58250
rect 612 58247 624 58248
rect 610 58240 632 58247
rect 607 58239 632 58240
rect 586 58232 644 58239
rect 607 58231 644 58232
rect 607 58215 610 58231
rect 616 58215 644 58231
rect 607 58214 644 58215
rect 586 58207 644 58214
rect 607 58206 610 58207
rect 612 58199 632 58207
rect 612 58195 624 58199
rect 649 58198 651 58248
rect 544 58161 548 58169
rect 400 58129 408 58159
rect 420 58129 436 58159
rect 400 58125 436 58129
rect 400 58117 430 58125
rect 428 58101 430 58117
rect 476 58089 480 58157
rect 544 58127 552 58161
rect 578 58127 582 58161
rect 544 58119 548 58127
rect 544 58089 586 58090
rect 288 58049 292 58081
rect 296 58079 368 58087
rect 378 58079 450 58087
rect 544 58082 548 58089
rect 439 58051 444 58079
rect 120 58035 170 58037
rect 76 58031 130 58035
rect 110 58026 130 58031
rect 60 58001 67 58011
rect 76 58001 77 58021
rect 96 57992 99 58026
rect 109 58001 110 58021
rect 119 58001 126 58011
rect 76 57985 92 57991
rect 94 57985 110 57991
rect 170 57985 172 58035
rect 186 57969 190 58003
rect 216 57969 220 58003
rect 213 57937 224 57969
rect 282 57965 292 58049
rect 296 58043 368 58051
rect 378 58043 450 58051
rect 468 58048 473 58082
rect 428 58013 430 58029
rect 251 57937 292 57965
rect 318 57944 324 58013
rect 12 57932 62 57934
rect 28 57923 59 57931
rect 62 57923 64 57932
rect 251 57931 263 57937
rect 28 57915 64 57923
rect 127 57923 158 57931
rect 127 57916 182 57923
rect 127 57915 161 57916
rect 59 57899 64 57915
rect 158 57899 161 57915
rect 253 57903 263 57931
rect 273 57903 293 57937
rect 318 57934 335 57944
rect 303 57918 316 57928
rect 318 57918 324 57934
rect 346 57928 348 58013
rect 400 58005 430 58013
rect 476 58011 480 58079
rect 511 58048 582 58082
rect 544 58041 548 58048
rect 400 58001 436 58005
rect 400 57971 408 58001
rect 420 57971 436 58001
rect 544 58003 548 58011
rect 28 57891 64 57899
rect 127 57898 161 57899
rect 127 57891 182 57898
rect 62 57882 64 57891
rect 282 57845 292 57903
rect 295 57894 324 57918
rect 333 57918 353 57928
rect 428 57924 430 57971
rect 476 57931 480 57999
rect 544 57969 552 58003
rect 578 57969 582 58003
rect 544 57961 548 57969
rect 367 57918 380 57924
rect 333 57894 380 57918
rect 318 57881 324 57894
rect 346 57881 348 57894
rect 367 57890 380 57894
rect 396 57890 408 57924
rect 420 57890 436 57924
rect 544 57921 553 57949
rect 319 57870 346 57881
rect 120 57829 170 57831
rect 76 57823 92 57829
rect 94 57823 110 57829
rect 76 57813 99 57822
rect 60 57803 67 57813
rect 76 57793 77 57813
rect 96 57788 99 57813
rect 109 57793 110 57813
rect 119 57803 126 57813
rect 76 57779 110 57783
rect 170 57779 172 57829
rect 186 57811 190 57845
rect 216 57811 220 57845
rect 182 57773 224 57774
rect 186 57749 220 57766
rect 223 57749 257 57766
rect 182 57732 257 57749
rect 182 57731 224 57732
rect 160 57725 246 57731
rect 288 57725 292 57845
rect 296 57843 368 57851
rect 428 57843 430 57890
rect 476 57853 480 57921
rect 485 57877 495 57911
rect 505 57883 525 57911
rect 505 57877 519 57883
rect 544 57877 555 57921
rect 485 57853 492 57877
rect 579 57862 582 57952
rect 612 57934 624 57935
rect 599 57932 649 57934
rect 612 57931 624 57932
rect 610 57924 632 57931
rect 607 57923 632 57924
rect 586 57916 644 57923
rect 607 57915 644 57916
rect 607 57899 610 57915
rect 616 57899 644 57915
rect 607 57898 644 57899
rect 586 57891 644 57898
rect 607 57890 610 57891
rect 612 57883 632 57891
rect 612 57879 624 57883
rect 649 57882 651 57932
rect 544 57845 548 57853
rect 400 57813 408 57843
rect 420 57813 436 57843
rect 400 57809 436 57813
rect 400 57801 430 57809
rect 428 57785 430 57801
rect 476 57773 480 57841
rect 544 57811 552 57845
rect 578 57811 582 57845
rect 544 57803 548 57811
rect 295 57732 300 57766
rect 324 57732 329 57766
rect 378 57763 450 57771
rect 544 57768 548 57773
rect 544 57764 582 57768
rect 544 57749 552 57764
rect 578 57749 582 57764
rect 544 57731 586 57749
rect 522 57725 608 57731
rect 182 57709 224 57725
rect 544 57709 586 57725
rect 17 57695 67 57697
rect 119 57695 169 57697
rect 186 57695 220 57709
rect 548 57695 582 57709
rect 599 57695 649 57697
rect 42 57653 59 57687
rect 67 57645 69 57695
rect 160 57687 246 57695
rect 522 57687 608 57695
rect 76 57653 110 57687
rect 127 57653 144 57687
rect 152 57653 161 57687
rect 162 57685 195 57687
rect 224 57685 244 57687
rect 162 57653 244 57685
rect 524 57685 548 57687
rect 573 57685 582 57687
rect 586 57685 606 57687
rect 160 57645 246 57653
rect 186 57629 220 57645
rect 182 57615 224 57616
rect 160 57609 182 57615
rect 224 57609 246 57615
rect 186 57574 220 57608
rect 223 57574 257 57608
rect 120 57561 170 57563
rect 76 57557 130 57561
rect 110 57552 130 57557
rect 60 57527 67 57537
rect 76 57527 77 57547
rect 96 57518 99 57552
rect 109 57527 110 57547
rect 119 57527 126 57537
rect 76 57511 92 57517
rect 94 57511 110 57517
rect 170 57511 172 57561
rect 186 57495 190 57529
rect 216 57495 220 57529
rect 288 57495 292 57683
rect 476 57615 480 57683
rect 524 57653 606 57685
rect 607 57653 616 57687
rect 522 57645 608 57653
rect 649 57645 651 57695
rect 548 57629 582 57645
rect 522 57610 548 57615
rect 522 57609 582 57610
rect 586 57609 608 57615
rect 295 57574 300 57608
rect 324 57574 329 57608
rect 544 57606 582 57609
rect 378 57569 450 57577
rect 428 57539 430 57555
rect 400 57531 430 57539
rect 476 57537 480 57605
rect 544 57576 552 57606
rect 578 57576 582 57606
rect 544 57567 548 57576
rect 400 57527 436 57531
rect 400 57497 408 57527
rect 420 57497 436 57527
rect 544 57529 548 57537
rect 12 57458 62 57460
rect 28 57449 59 57457
rect 62 57449 64 57458
rect 28 57441 64 57449
rect 127 57449 158 57457
rect 127 57442 182 57449
rect 215 57447 224 57475
rect 127 57441 161 57442
rect 59 57425 64 57441
rect 158 57425 161 57441
rect 28 57417 64 57425
rect 127 57424 161 57425
rect 127 57417 182 57424
rect 62 57408 64 57417
rect 213 57409 224 57447
rect 282 57437 292 57495
rect 296 57489 368 57497
rect 319 57459 346 57470
rect 318 57446 324 57459
rect 346 57446 348 57459
rect 428 57450 430 57497
rect 443 57487 450 57489
rect 476 57457 480 57525
rect 544 57495 552 57529
rect 578 57495 582 57529
rect 481 57463 517 57491
rect 481 57457 495 57463
rect 367 57446 380 57450
rect 251 57403 263 57437
rect 273 57403 293 57437
rect 295 57422 324 57446
rect 303 57412 316 57422
rect 318 57406 324 57422
rect 333 57422 380 57446
rect 333 57412 353 57422
rect 367 57416 380 57422
rect 396 57416 408 57450
rect 420 57416 436 57450
rect 120 57355 170 57357
rect 76 57349 92 57355
rect 94 57349 110 57355
rect 76 57339 99 57348
rect 60 57329 67 57339
rect 76 57319 77 57339
rect 96 57314 99 57339
rect 109 57319 110 57339
rect 119 57329 126 57339
rect 76 57305 110 57309
rect 170 57305 172 57355
rect 186 57337 190 57371
rect 216 57337 220 57371
rect 186 57260 220 57294
rect 282 57291 292 57403
rect 318 57396 335 57406
rect 318 57327 324 57396
rect 346 57327 348 57412
rect 428 57369 430 57416
rect 476 57379 480 57447
rect 485 57429 495 57457
rect 505 57457 519 57463
rect 544 57457 555 57495
rect 505 57429 525 57457
rect 544 57429 553 57457
rect 544 57409 548 57429
rect 579 57388 582 57478
rect 612 57460 624 57461
rect 599 57458 649 57460
rect 612 57457 624 57458
rect 610 57450 632 57457
rect 607 57449 632 57450
rect 586 57442 644 57449
rect 607 57441 644 57442
rect 607 57425 610 57441
rect 616 57425 644 57441
rect 607 57424 644 57425
rect 586 57417 644 57424
rect 607 57416 610 57417
rect 612 57409 632 57417
rect 612 57405 624 57409
rect 649 57408 651 57458
rect 544 57371 548 57379
rect 400 57339 408 57369
rect 420 57339 436 57369
rect 400 57335 436 57339
rect 400 57327 430 57335
rect 428 57311 430 57327
rect 476 57299 480 57367
rect 544 57337 552 57371
rect 578 57337 582 57371
rect 544 57329 548 57337
rect 544 57299 586 57300
rect 288 57259 292 57291
rect 296 57289 368 57297
rect 378 57289 450 57297
rect 544 57292 548 57299
rect 439 57261 444 57289
rect 120 57245 170 57247
rect 76 57241 130 57245
rect 110 57236 130 57241
rect 60 57211 67 57221
rect 76 57211 77 57231
rect 96 57202 99 57236
rect 109 57211 110 57231
rect 119 57211 126 57221
rect 76 57195 92 57201
rect 94 57195 110 57201
rect 170 57195 172 57245
rect 186 57179 190 57213
rect 216 57179 220 57213
rect 213 57147 224 57179
rect 282 57175 292 57259
rect 296 57253 368 57261
rect 378 57253 450 57261
rect 468 57258 473 57292
rect 428 57223 430 57239
rect 251 57147 292 57175
rect 318 57154 324 57223
rect 12 57142 62 57144
rect 28 57133 59 57141
rect 62 57133 64 57142
rect 251 57141 263 57147
rect 28 57125 64 57133
rect 127 57133 158 57141
rect 127 57126 182 57133
rect 127 57125 161 57126
rect 59 57109 64 57125
rect 158 57109 161 57125
rect 253 57113 263 57141
rect 273 57113 293 57147
rect 318 57144 335 57154
rect 303 57128 316 57138
rect 318 57128 324 57144
rect 346 57138 348 57223
rect 400 57215 430 57223
rect 476 57221 480 57289
rect 511 57258 582 57292
rect 544 57251 548 57258
rect 400 57211 436 57215
rect 400 57181 408 57211
rect 420 57181 436 57211
rect 544 57213 548 57221
rect 28 57101 64 57109
rect 127 57108 161 57109
rect 127 57101 182 57108
rect 62 57092 64 57101
rect 282 57055 292 57113
rect 295 57104 324 57128
rect 333 57128 353 57138
rect 428 57134 430 57181
rect 476 57141 480 57209
rect 544 57179 552 57213
rect 578 57179 582 57213
rect 544 57171 548 57179
rect 367 57128 380 57134
rect 333 57104 380 57128
rect 318 57091 324 57104
rect 346 57091 348 57104
rect 367 57100 380 57104
rect 396 57100 408 57134
rect 420 57100 436 57134
rect 544 57131 553 57159
rect 319 57080 346 57091
rect 120 57039 170 57041
rect 76 57033 92 57039
rect 94 57033 110 57039
rect 76 57023 99 57032
rect 60 57013 67 57023
rect 76 57003 77 57023
rect 96 56998 99 57023
rect 109 57003 110 57023
rect 119 57013 126 57023
rect 76 56989 110 56993
rect 170 56989 172 57039
rect 186 57021 190 57055
rect 216 57021 220 57055
rect 182 56983 224 56984
rect 186 56959 220 56976
rect 223 56959 257 56976
rect 182 56942 257 56959
rect 182 56941 224 56942
rect 160 56935 246 56941
rect 288 56935 292 57055
rect 296 57053 368 57061
rect 428 57053 430 57100
rect 476 57063 480 57131
rect 485 57087 495 57121
rect 505 57093 525 57121
rect 505 57087 519 57093
rect 544 57087 555 57131
rect 485 57063 492 57087
rect 579 57072 582 57162
rect 612 57144 624 57145
rect 599 57142 649 57144
rect 612 57141 624 57142
rect 610 57134 632 57141
rect 607 57133 632 57134
rect 586 57126 644 57133
rect 607 57125 644 57126
rect 607 57109 610 57125
rect 616 57109 644 57125
rect 607 57108 644 57109
rect 586 57101 644 57108
rect 607 57100 610 57101
rect 612 57093 632 57101
rect 612 57089 624 57093
rect 649 57092 651 57142
rect 544 57055 548 57063
rect 400 57023 408 57053
rect 420 57023 436 57053
rect 400 57019 436 57023
rect 400 57011 430 57019
rect 428 56995 430 57011
rect 476 56983 480 57051
rect 544 57021 552 57055
rect 578 57021 582 57055
rect 544 57013 548 57021
rect 295 56942 300 56976
rect 324 56942 329 56976
rect 378 56973 450 56981
rect 544 56978 548 56983
rect 544 56974 582 56978
rect 544 56959 552 56974
rect 578 56959 582 56974
rect 544 56941 586 56959
rect 522 56935 608 56941
rect 182 56919 224 56935
rect 544 56919 586 56935
rect 17 56905 67 56907
rect 119 56905 169 56907
rect 186 56905 220 56919
rect 548 56905 582 56919
rect 599 56905 649 56907
rect 42 56863 59 56897
rect 67 56855 69 56905
rect 160 56897 246 56905
rect 522 56897 608 56905
rect 76 56863 110 56897
rect 127 56863 144 56897
rect 152 56863 161 56897
rect 162 56895 195 56897
rect 224 56895 244 56897
rect 162 56863 244 56895
rect 524 56895 548 56897
rect 573 56895 582 56897
rect 586 56895 606 56897
rect 160 56855 246 56863
rect 186 56839 220 56855
rect 182 56825 224 56826
rect 160 56819 182 56825
rect 224 56819 246 56825
rect 186 56784 220 56818
rect 223 56784 257 56818
rect 120 56771 170 56773
rect 76 56767 130 56771
rect 110 56762 130 56767
rect 60 56737 67 56747
rect 76 56737 77 56757
rect 96 56728 99 56762
rect 109 56737 110 56757
rect 119 56737 126 56747
rect 76 56721 92 56727
rect 94 56721 110 56727
rect 170 56721 172 56771
rect 186 56705 190 56739
rect 216 56705 220 56739
rect 288 56705 292 56893
rect 476 56825 480 56893
rect 524 56863 606 56895
rect 607 56863 616 56897
rect 522 56855 608 56863
rect 649 56855 651 56905
rect 548 56839 582 56855
rect 522 56820 548 56825
rect 522 56819 582 56820
rect 586 56819 608 56825
rect 295 56784 300 56818
rect 324 56784 329 56818
rect 544 56816 582 56819
rect 378 56779 450 56787
rect 428 56749 430 56765
rect 400 56741 430 56749
rect 476 56747 480 56815
rect 544 56786 552 56816
rect 578 56786 582 56816
rect 544 56777 548 56786
rect 400 56737 436 56741
rect 400 56707 408 56737
rect 420 56707 436 56737
rect 544 56739 548 56747
rect 12 56668 62 56670
rect 28 56659 59 56667
rect 62 56659 64 56668
rect 28 56651 64 56659
rect 127 56659 158 56667
rect 127 56652 182 56659
rect 215 56657 224 56685
rect 127 56651 161 56652
rect 59 56635 64 56651
rect 158 56635 161 56651
rect 28 56627 64 56635
rect 127 56634 161 56635
rect 127 56627 182 56634
rect 62 56618 64 56627
rect 213 56619 224 56657
rect 282 56647 292 56705
rect 296 56699 368 56707
rect 319 56669 346 56680
rect 318 56656 324 56669
rect 346 56656 348 56669
rect 428 56660 430 56707
rect 443 56697 450 56699
rect 476 56667 480 56735
rect 544 56705 552 56739
rect 578 56705 582 56739
rect 481 56673 517 56701
rect 481 56667 495 56673
rect 367 56656 380 56660
rect 251 56613 263 56647
rect 273 56613 293 56647
rect 295 56632 324 56656
rect 303 56622 316 56632
rect 318 56616 324 56632
rect 333 56632 380 56656
rect 333 56622 353 56632
rect 367 56626 380 56632
rect 396 56626 408 56660
rect 420 56626 436 56660
rect 120 56565 170 56567
rect 76 56559 92 56565
rect 94 56559 110 56565
rect 76 56549 99 56558
rect 60 56539 67 56549
rect 76 56529 77 56549
rect 96 56524 99 56549
rect 109 56529 110 56549
rect 119 56539 126 56549
rect 76 56515 110 56519
rect 170 56515 172 56565
rect 186 56547 190 56581
rect 216 56547 220 56581
rect 186 56470 220 56504
rect 282 56501 292 56613
rect 318 56606 335 56616
rect 318 56537 324 56606
rect 346 56537 348 56622
rect 428 56579 430 56626
rect 476 56589 480 56657
rect 485 56639 495 56667
rect 505 56667 519 56673
rect 544 56667 555 56705
rect 505 56639 525 56667
rect 544 56639 553 56667
rect 544 56619 548 56639
rect 579 56598 582 56688
rect 612 56670 624 56671
rect 599 56668 649 56670
rect 612 56667 624 56668
rect 610 56660 632 56667
rect 607 56659 632 56660
rect 586 56652 644 56659
rect 607 56651 644 56652
rect 607 56635 610 56651
rect 616 56635 644 56651
rect 607 56634 644 56635
rect 586 56627 644 56634
rect 607 56626 610 56627
rect 612 56619 632 56627
rect 612 56615 624 56619
rect 649 56618 651 56668
rect 544 56581 548 56589
rect 400 56549 408 56579
rect 420 56549 436 56579
rect 400 56545 436 56549
rect 400 56537 430 56545
rect 428 56521 430 56537
rect 476 56509 480 56577
rect 544 56547 552 56581
rect 578 56547 582 56581
rect 544 56539 548 56547
rect 544 56509 586 56510
rect 288 56469 292 56501
rect 296 56499 368 56507
rect 378 56499 450 56507
rect 544 56502 548 56509
rect 439 56471 444 56499
rect 120 56455 170 56457
rect 76 56451 130 56455
rect 110 56446 130 56451
rect 60 56421 67 56431
rect 76 56421 77 56441
rect 96 56412 99 56446
rect 109 56421 110 56441
rect 119 56421 126 56431
rect 76 56405 92 56411
rect 94 56405 110 56411
rect 170 56405 172 56455
rect 186 56389 190 56423
rect 216 56389 220 56423
rect 213 56357 224 56389
rect 282 56385 292 56469
rect 296 56463 368 56471
rect 378 56463 450 56471
rect 468 56468 473 56502
rect 428 56433 430 56449
rect 251 56357 292 56385
rect 318 56364 324 56433
rect 12 56352 62 56354
rect 28 56343 59 56351
rect 62 56343 64 56352
rect 251 56351 263 56357
rect 28 56335 64 56343
rect 127 56343 158 56351
rect 127 56336 182 56343
rect 127 56335 161 56336
rect 59 56319 64 56335
rect 158 56319 161 56335
rect 253 56323 263 56351
rect 273 56323 293 56357
rect 318 56354 335 56364
rect 303 56338 316 56348
rect 318 56338 324 56354
rect 346 56348 348 56433
rect 400 56425 430 56433
rect 476 56431 480 56499
rect 511 56468 582 56502
rect 544 56461 548 56468
rect 400 56421 436 56425
rect 400 56391 408 56421
rect 420 56391 436 56421
rect 544 56423 548 56431
rect 28 56311 64 56319
rect 127 56318 161 56319
rect 127 56311 182 56318
rect 62 56302 64 56311
rect 282 56265 292 56323
rect 295 56314 324 56338
rect 333 56338 353 56348
rect 428 56344 430 56391
rect 476 56351 480 56419
rect 544 56389 552 56423
rect 578 56389 582 56423
rect 544 56381 548 56389
rect 367 56338 380 56344
rect 333 56314 380 56338
rect 318 56301 324 56314
rect 346 56301 348 56314
rect 367 56310 380 56314
rect 396 56310 408 56344
rect 420 56310 436 56344
rect 544 56341 553 56369
rect 319 56290 346 56301
rect 120 56249 170 56251
rect 76 56243 92 56249
rect 94 56243 110 56249
rect 76 56233 99 56242
rect 60 56223 67 56233
rect 76 56213 77 56233
rect 96 56208 99 56233
rect 109 56213 110 56233
rect 119 56223 126 56233
rect 76 56199 110 56203
rect 170 56199 172 56249
rect 186 56231 190 56265
rect 216 56231 220 56265
rect 182 56193 224 56194
rect 186 56169 220 56186
rect 223 56169 257 56186
rect 182 56152 257 56169
rect 182 56151 224 56152
rect 160 56145 246 56151
rect 288 56145 292 56265
rect 296 56263 368 56271
rect 428 56263 430 56310
rect 476 56273 480 56341
rect 485 56297 495 56331
rect 505 56303 525 56331
rect 505 56297 519 56303
rect 544 56297 555 56341
rect 485 56273 492 56297
rect 579 56282 582 56372
rect 612 56354 624 56355
rect 599 56352 649 56354
rect 612 56351 624 56352
rect 610 56344 632 56351
rect 607 56343 632 56344
rect 586 56336 644 56343
rect 607 56335 644 56336
rect 607 56319 610 56335
rect 616 56319 644 56335
rect 607 56318 644 56319
rect 586 56311 644 56318
rect 607 56310 610 56311
rect 612 56303 632 56311
rect 612 56299 624 56303
rect 649 56302 651 56352
rect 544 56265 548 56273
rect 400 56233 408 56263
rect 420 56233 436 56263
rect 400 56229 436 56233
rect 400 56221 430 56229
rect 428 56205 430 56221
rect 476 56193 480 56261
rect 544 56231 552 56265
rect 578 56231 582 56265
rect 544 56223 548 56231
rect 295 56152 300 56186
rect 324 56152 329 56186
rect 378 56183 450 56191
rect 544 56188 548 56193
rect 544 56184 582 56188
rect 544 56169 552 56184
rect 578 56169 582 56184
rect 544 56151 586 56169
rect 522 56145 608 56151
rect 182 56129 224 56145
rect 544 56129 586 56145
rect 17 56115 67 56117
rect 119 56115 169 56117
rect 186 56115 220 56129
rect 548 56115 582 56129
rect 599 56115 649 56117
rect 42 56073 59 56107
rect 67 56065 69 56115
rect 160 56107 246 56115
rect 522 56107 608 56115
rect 76 56073 110 56107
rect 127 56073 144 56107
rect 152 56073 161 56107
rect 162 56105 195 56107
rect 224 56105 244 56107
rect 162 56073 244 56105
rect 524 56105 548 56107
rect 573 56105 582 56107
rect 586 56105 606 56107
rect 160 56065 246 56073
rect 186 56049 220 56065
rect 182 56035 224 56036
rect 160 56029 182 56035
rect 224 56029 246 56035
rect 186 55994 220 56028
rect 223 55994 257 56028
rect 120 55981 170 55983
rect 76 55977 130 55981
rect 110 55972 130 55977
rect 60 55947 67 55957
rect 76 55947 77 55967
rect 96 55938 99 55972
rect 109 55947 110 55967
rect 119 55947 126 55957
rect 76 55931 92 55937
rect 94 55931 110 55937
rect 170 55931 172 55981
rect 186 55915 190 55949
rect 216 55915 220 55949
rect 288 55915 292 56103
rect 476 56035 480 56103
rect 524 56073 606 56105
rect 607 56073 616 56107
rect 522 56065 608 56073
rect 649 56065 651 56115
rect 548 56049 582 56065
rect 522 56030 548 56035
rect 522 56029 582 56030
rect 586 56029 608 56035
rect 295 55994 300 56028
rect 324 55994 329 56028
rect 544 56026 582 56029
rect 378 55989 450 55997
rect 428 55959 430 55975
rect 400 55951 430 55959
rect 476 55957 480 56025
rect 544 55996 552 56026
rect 578 55996 582 56026
rect 544 55987 548 55996
rect 400 55947 436 55951
rect 400 55917 408 55947
rect 420 55917 436 55947
rect 544 55949 548 55957
rect 12 55878 62 55880
rect 28 55869 59 55877
rect 62 55869 64 55878
rect 28 55861 64 55869
rect 127 55869 158 55877
rect 127 55862 182 55869
rect 215 55867 224 55895
rect 127 55861 161 55862
rect 59 55845 64 55861
rect 158 55845 161 55861
rect 28 55837 64 55845
rect 127 55844 161 55845
rect 127 55837 182 55844
rect 62 55828 64 55837
rect 213 55829 224 55867
rect 282 55857 292 55915
rect 296 55909 368 55917
rect 319 55879 346 55890
rect 318 55866 324 55879
rect 346 55866 348 55879
rect 428 55870 430 55917
rect 443 55907 450 55909
rect 476 55877 480 55945
rect 544 55915 552 55949
rect 578 55915 582 55949
rect 481 55883 517 55911
rect 481 55877 495 55883
rect 367 55866 380 55870
rect 251 55823 263 55857
rect 273 55823 293 55857
rect 295 55842 324 55866
rect 303 55832 316 55842
rect 318 55826 324 55842
rect 333 55842 380 55866
rect 333 55832 353 55842
rect 367 55836 380 55842
rect 396 55836 408 55870
rect 420 55836 436 55870
rect 120 55775 170 55777
rect 76 55769 92 55775
rect 94 55769 110 55775
rect 76 55759 99 55768
rect 60 55749 67 55759
rect 76 55739 77 55759
rect 96 55734 99 55759
rect 109 55739 110 55759
rect 119 55749 126 55759
rect 76 55725 110 55729
rect 170 55725 172 55775
rect 186 55757 190 55791
rect 216 55757 220 55791
rect 186 55680 220 55714
rect 282 55711 292 55823
rect 318 55816 335 55826
rect 318 55747 324 55816
rect 346 55747 348 55832
rect 428 55789 430 55836
rect 476 55799 480 55867
rect 485 55849 495 55877
rect 505 55877 519 55883
rect 544 55877 555 55915
rect 505 55849 525 55877
rect 544 55849 553 55877
rect 544 55829 548 55849
rect 579 55808 582 55898
rect 612 55880 624 55881
rect 599 55878 649 55880
rect 612 55877 624 55878
rect 610 55870 632 55877
rect 607 55869 632 55870
rect 586 55862 644 55869
rect 607 55861 644 55862
rect 607 55845 610 55861
rect 616 55845 644 55861
rect 607 55844 644 55845
rect 586 55837 644 55844
rect 607 55836 610 55837
rect 612 55829 632 55837
rect 612 55825 624 55829
rect 649 55828 651 55878
rect 544 55791 548 55799
rect 400 55759 408 55789
rect 420 55759 436 55789
rect 400 55755 436 55759
rect 400 55747 430 55755
rect 428 55731 430 55747
rect 476 55719 480 55787
rect 544 55757 552 55791
rect 578 55757 582 55791
rect 544 55749 548 55757
rect 544 55719 586 55720
rect 288 55679 292 55711
rect 296 55709 368 55717
rect 378 55709 450 55717
rect 544 55712 548 55719
rect 439 55681 444 55709
rect 120 55665 170 55667
rect 76 55661 130 55665
rect 110 55656 130 55661
rect 60 55631 67 55641
rect 76 55631 77 55651
rect 96 55622 99 55656
rect 109 55631 110 55651
rect 119 55631 126 55641
rect 76 55615 92 55621
rect 94 55615 110 55621
rect 170 55615 172 55665
rect 186 55599 190 55633
rect 216 55599 220 55633
rect 213 55567 224 55599
rect 282 55595 292 55679
rect 296 55673 368 55681
rect 378 55673 450 55681
rect 468 55678 473 55712
rect 428 55643 430 55659
rect 251 55567 292 55595
rect 318 55574 324 55643
rect 12 55562 62 55564
rect 28 55553 59 55561
rect 62 55553 64 55562
rect 251 55561 263 55567
rect 28 55545 64 55553
rect 127 55553 158 55561
rect 127 55546 182 55553
rect 127 55545 161 55546
rect 59 55529 64 55545
rect 158 55529 161 55545
rect 253 55533 263 55561
rect 273 55533 293 55567
rect 318 55564 335 55574
rect 303 55548 316 55558
rect 318 55548 324 55564
rect 346 55558 348 55643
rect 400 55635 430 55643
rect 476 55641 480 55709
rect 511 55678 582 55712
rect 544 55671 548 55678
rect 400 55631 436 55635
rect 400 55601 408 55631
rect 420 55601 436 55631
rect 544 55633 548 55641
rect 28 55521 64 55529
rect 127 55528 161 55529
rect 127 55521 182 55528
rect 62 55512 64 55521
rect 282 55475 292 55533
rect 295 55524 324 55548
rect 333 55548 353 55558
rect 428 55554 430 55601
rect 476 55561 480 55629
rect 544 55599 552 55633
rect 578 55599 582 55633
rect 544 55591 548 55599
rect 367 55548 380 55554
rect 333 55524 380 55548
rect 318 55511 324 55524
rect 346 55511 348 55524
rect 367 55520 380 55524
rect 396 55520 408 55554
rect 420 55520 436 55554
rect 544 55551 553 55579
rect 319 55500 346 55511
rect 120 55459 170 55461
rect 76 55453 92 55459
rect 94 55453 110 55459
rect 76 55443 99 55452
rect 60 55433 67 55443
rect 76 55423 77 55443
rect 96 55418 99 55443
rect 109 55423 110 55443
rect 119 55433 126 55443
rect 76 55409 110 55413
rect 170 55409 172 55459
rect 186 55441 190 55475
rect 216 55441 220 55475
rect 182 55403 224 55404
rect 186 55379 220 55396
rect 223 55379 257 55396
rect 182 55362 257 55379
rect 182 55361 224 55362
rect 160 55355 246 55361
rect 288 55355 292 55475
rect 296 55473 368 55481
rect 428 55473 430 55520
rect 476 55483 480 55551
rect 485 55507 495 55541
rect 505 55513 525 55541
rect 505 55507 519 55513
rect 544 55507 555 55551
rect 485 55483 492 55507
rect 579 55492 582 55582
rect 612 55564 624 55565
rect 599 55562 649 55564
rect 612 55561 624 55562
rect 610 55554 632 55561
rect 607 55553 632 55554
rect 586 55546 644 55553
rect 607 55545 644 55546
rect 607 55529 610 55545
rect 616 55529 644 55545
rect 607 55528 644 55529
rect 586 55521 644 55528
rect 607 55520 610 55521
rect 612 55513 632 55521
rect 612 55509 624 55513
rect 649 55512 651 55562
rect 544 55475 548 55483
rect 400 55443 408 55473
rect 420 55443 436 55473
rect 400 55439 436 55443
rect 400 55431 430 55439
rect 428 55415 430 55431
rect 476 55403 480 55471
rect 544 55441 552 55475
rect 578 55441 582 55475
rect 544 55433 548 55441
rect 295 55362 300 55396
rect 324 55362 329 55396
rect 378 55393 450 55401
rect 544 55398 548 55403
rect 544 55394 582 55398
rect 544 55379 552 55394
rect 578 55379 582 55394
rect 544 55361 586 55379
rect 522 55355 608 55361
rect 182 55339 224 55355
rect 544 55339 586 55355
rect 17 55325 67 55327
rect 119 55325 169 55327
rect 186 55325 220 55339
rect 548 55325 582 55339
rect 599 55325 649 55327
rect 42 55283 59 55317
rect 67 55275 69 55325
rect 160 55317 246 55325
rect 522 55317 608 55325
rect 76 55283 110 55317
rect 127 55283 144 55317
rect 152 55283 161 55317
rect 162 55315 195 55317
rect 224 55315 244 55317
rect 162 55283 244 55315
rect 524 55315 548 55317
rect 573 55315 582 55317
rect 586 55315 606 55317
rect 160 55275 246 55283
rect 186 55259 220 55275
rect 182 55245 224 55246
rect 160 55239 182 55245
rect 224 55239 246 55245
rect 186 55204 220 55238
rect 223 55204 257 55238
rect 120 55191 170 55193
rect 76 55187 130 55191
rect 110 55182 130 55187
rect 60 55157 67 55167
rect 76 55157 77 55177
rect 96 55148 99 55182
rect 109 55157 110 55177
rect 119 55157 126 55167
rect 76 55141 92 55147
rect 94 55141 110 55147
rect 170 55141 172 55191
rect 186 55125 190 55159
rect 216 55125 220 55159
rect 288 55125 292 55313
rect 476 55245 480 55313
rect 524 55283 606 55315
rect 607 55283 616 55317
rect 522 55275 608 55283
rect 649 55275 651 55325
rect 548 55259 582 55275
rect 522 55240 548 55245
rect 522 55239 582 55240
rect 586 55239 608 55245
rect 295 55204 300 55238
rect 324 55204 329 55238
rect 544 55236 582 55239
rect 378 55199 450 55207
rect 428 55169 430 55185
rect 400 55161 430 55169
rect 476 55167 480 55235
rect 544 55206 552 55236
rect 578 55206 582 55236
rect 544 55197 548 55206
rect 400 55157 436 55161
rect 400 55127 408 55157
rect 420 55127 436 55157
rect 544 55159 548 55167
rect 12 55088 62 55090
rect 28 55079 59 55087
rect 62 55079 64 55088
rect 28 55071 64 55079
rect 127 55079 158 55087
rect 127 55072 182 55079
rect 215 55077 224 55105
rect 127 55071 161 55072
rect 59 55055 64 55071
rect 158 55055 161 55071
rect 28 55047 64 55055
rect 127 55054 161 55055
rect 127 55047 182 55054
rect 62 55038 64 55047
rect 213 55039 224 55077
rect 282 55067 292 55125
rect 296 55119 368 55127
rect 319 55089 346 55100
rect 318 55076 324 55089
rect 346 55076 348 55089
rect 428 55080 430 55127
rect 443 55117 450 55119
rect 476 55087 480 55155
rect 544 55125 552 55159
rect 578 55125 582 55159
rect 481 55093 517 55121
rect 481 55087 495 55093
rect 367 55076 380 55080
rect 251 55033 263 55067
rect 273 55033 293 55067
rect 295 55052 324 55076
rect 303 55042 316 55052
rect 318 55036 324 55052
rect 333 55052 380 55076
rect 333 55042 353 55052
rect 367 55046 380 55052
rect 396 55046 408 55080
rect 420 55046 436 55080
rect 120 54985 170 54987
rect 76 54979 92 54985
rect 94 54979 110 54985
rect 76 54969 99 54978
rect 60 54959 67 54969
rect 76 54949 77 54969
rect 96 54944 99 54969
rect 109 54949 110 54969
rect 119 54959 126 54969
rect 76 54935 110 54939
rect 170 54935 172 54985
rect 186 54967 190 55001
rect 216 54967 220 55001
rect 186 54890 220 54924
rect 282 54921 292 55033
rect 318 55026 335 55036
rect 318 54957 324 55026
rect 346 54957 348 55042
rect 428 54999 430 55046
rect 476 55009 480 55077
rect 485 55059 495 55087
rect 505 55087 519 55093
rect 544 55087 555 55125
rect 505 55059 525 55087
rect 544 55059 553 55087
rect 544 55039 548 55059
rect 579 55018 582 55108
rect 612 55090 624 55091
rect 599 55088 649 55090
rect 612 55087 624 55088
rect 610 55080 632 55087
rect 607 55079 632 55080
rect 586 55072 644 55079
rect 607 55071 644 55072
rect 607 55055 610 55071
rect 616 55055 644 55071
rect 607 55054 644 55055
rect 586 55047 644 55054
rect 607 55046 610 55047
rect 612 55039 632 55047
rect 612 55035 624 55039
rect 649 55038 651 55088
rect 544 55001 548 55009
rect 400 54969 408 54999
rect 420 54969 436 54999
rect 400 54965 436 54969
rect 400 54957 430 54965
rect 428 54941 430 54957
rect 476 54929 480 54997
rect 544 54967 552 55001
rect 578 54967 582 55001
rect 544 54959 548 54967
rect 544 54929 586 54930
rect 288 54889 292 54921
rect 296 54919 368 54927
rect 378 54919 450 54927
rect 544 54922 548 54929
rect 439 54891 444 54919
rect 120 54875 170 54877
rect 76 54871 130 54875
rect 110 54866 130 54871
rect 60 54841 67 54851
rect 76 54841 77 54861
rect 96 54832 99 54866
rect 109 54841 110 54861
rect 119 54841 126 54851
rect 76 54825 92 54831
rect 94 54825 110 54831
rect 170 54825 172 54875
rect 186 54809 190 54843
rect 216 54809 220 54843
rect 213 54777 224 54809
rect 282 54805 292 54889
rect 296 54883 368 54891
rect 378 54883 450 54891
rect 468 54888 473 54922
rect 428 54853 430 54869
rect 251 54777 292 54805
rect 318 54784 324 54853
rect 12 54772 62 54774
rect 28 54763 59 54771
rect 62 54763 64 54772
rect 251 54771 263 54777
rect 28 54755 64 54763
rect 127 54763 158 54771
rect 127 54756 182 54763
rect 127 54755 161 54756
rect 59 54739 64 54755
rect 158 54739 161 54755
rect 253 54743 263 54771
rect 273 54743 293 54777
rect 318 54774 335 54784
rect 303 54758 316 54768
rect 318 54758 324 54774
rect 346 54768 348 54853
rect 400 54845 430 54853
rect 476 54851 480 54919
rect 511 54888 582 54922
rect 544 54881 548 54888
rect 400 54841 436 54845
rect 400 54811 408 54841
rect 420 54811 436 54841
rect 544 54843 548 54851
rect 28 54731 64 54739
rect 127 54738 161 54739
rect 127 54731 182 54738
rect 62 54722 64 54731
rect 282 54685 292 54743
rect 295 54734 324 54758
rect 333 54758 353 54768
rect 428 54764 430 54811
rect 476 54771 480 54839
rect 544 54809 552 54843
rect 578 54809 582 54843
rect 544 54801 548 54809
rect 367 54758 380 54764
rect 333 54734 380 54758
rect 318 54721 324 54734
rect 346 54721 348 54734
rect 367 54730 380 54734
rect 396 54730 408 54764
rect 420 54730 436 54764
rect 544 54761 553 54789
rect 319 54710 346 54721
rect 120 54669 170 54671
rect 76 54663 92 54669
rect 94 54663 110 54669
rect 76 54653 99 54662
rect 60 54643 67 54653
rect 76 54633 77 54653
rect 96 54628 99 54653
rect 109 54633 110 54653
rect 119 54643 126 54653
rect 76 54619 110 54623
rect 170 54619 172 54669
rect 186 54651 190 54685
rect 216 54651 220 54685
rect 182 54613 224 54614
rect 186 54589 220 54606
rect 223 54589 257 54606
rect 182 54572 257 54589
rect 182 54571 224 54572
rect 160 54565 246 54571
rect 288 54565 292 54685
rect 296 54683 368 54691
rect 428 54683 430 54730
rect 476 54693 480 54761
rect 485 54717 495 54751
rect 505 54723 525 54751
rect 505 54717 519 54723
rect 544 54717 555 54761
rect 485 54693 492 54717
rect 579 54702 582 54792
rect 612 54774 624 54775
rect 599 54772 649 54774
rect 612 54771 624 54772
rect 610 54764 632 54771
rect 607 54763 632 54764
rect 586 54756 644 54763
rect 607 54755 644 54756
rect 607 54739 610 54755
rect 616 54739 644 54755
rect 607 54738 644 54739
rect 586 54731 644 54738
rect 607 54730 610 54731
rect 612 54723 632 54731
rect 612 54719 624 54723
rect 649 54722 651 54772
rect 544 54685 548 54693
rect 400 54653 408 54683
rect 420 54653 436 54683
rect 400 54649 436 54653
rect 400 54641 430 54649
rect 428 54625 430 54641
rect 476 54613 480 54681
rect 544 54651 552 54685
rect 578 54651 582 54685
rect 544 54643 548 54651
rect 295 54572 300 54606
rect 324 54572 329 54606
rect 378 54603 450 54611
rect 544 54608 548 54613
rect 544 54604 582 54608
rect 544 54589 552 54604
rect 578 54589 582 54604
rect 544 54571 586 54589
rect 522 54565 608 54571
rect 182 54549 224 54565
rect 544 54549 586 54565
rect 17 54535 67 54537
rect 119 54535 169 54537
rect 186 54535 220 54549
rect 548 54535 582 54549
rect 599 54535 649 54537
rect 42 54493 59 54527
rect 67 54485 69 54535
rect 160 54527 246 54535
rect 522 54527 608 54535
rect 76 54493 110 54527
rect 127 54493 144 54527
rect 152 54493 161 54527
rect 162 54525 195 54527
rect 224 54525 244 54527
rect 162 54493 244 54525
rect 524 54525 548 54527
rect 573 54525 582 54527
rect 586 54525 606 54527
rect 160 54485 246 54493
rect 186 54469 220 54485
rect 182 54455 224 54456
rect 160 54449 182 54455
rect 224 54449 246 54455
rect 186 54414 220 54448
rect 223 54414 257 54448
rect 120 54401 170 54403
rect 76 54397 130 54401
rect 110 54392 130 54397
rect 60 54367 67 54377
rect 76 54367 77 54387
rect 96 54358 99 54392
rect 109 54367 110 54387
rect 119 54367 126 54377
rect 76 54351 92 54357
rect 94 54351 110 54357
rect 170 54351 172 54401
rect 186 54335 190 54369
rect 216 54335 220 54369
rect 288 54335 292 54523
rect 476 54455 480 54523
rect 524 54493 606 54525
rect 607 54493 616 54527
rect 522 54485 608 54493
rect 649 54485 651 54535
rect 548 54469 582 54485
rect 522 54450 548 54455
rect 522 54449 582 54450
rect 586 54449 608 54455
rect 295 54414 300 54448
rect 324 54414 329 54448
rect 544 54446 582 54449
rect 378 54409 450 54417
rect 428 54379 430 54395
rect 400 54371 430 54379
rect 476 54377 480 54445
rect 544 54416 552 54446
rect 578 54416 582 54446
rect 544 54407 548 54416
rect 400 54367 436 54371
rect 400 54337 408 54367
rect 420 54337 436 54367
rect 544 54369 548 54377
rect 12 54298 62 54300
rect 28 54289 59 54297
rect 62 54289 64 54298
rect 28 54281 64 54289
rect 127 54289 158 54297
rect 127 54282 182 54289
rect 215 54287 224 54315
rect 127 54281 161 54282
rect 59 54265 64 54281
rect 158 54265 161 54281
rect 28 54257 64 54265
rect 127 54264 161 54265
rect 127 54257 182 54264
rect 62 54248 64 54257
rect 213 54249 224 54287
rect 282 54277 292 54335
rect 296 54329 368 54337
rect 319 54299 346 54310
rect 318 54286 324 54299
rect 346 54286 348 54299
rect 428 54290 430 54337
rect 443 54327 450 54329
rect 476 54297 480 54365
rect 544 54335 552 54369
rect 578 54335 582 54369
rect 481 54303 517 54331
rect 481 54297 495 54303
rect 367 54286 380 54290
rect 251 54243 263 54277
rect 273 54243 293 54277
rect 295 54262 324 54286
rect 303 54252 316 54262
rect 318 54246 324 54262
rect 333 54262 380 54286
rect 333 54252 353 54262
rect 367 54256 380 54262
rect 396 54256 408 54290
rect 420 54256 436 54290
rect 120 54195 170 54197
rect 76 54189 92 54195
rect 94 54189 110 54195
rect 76 54179 99 54188
rect 60 54169 67 54179
rect 76 54159 77 54179
rect 96 54154 99 54179
rect 109 54159 110 54179
rect 119 54169 126 54179
rect 76 54145 110 54149
rect 170 54145 172 54195
rect 186 54177 190 54211
rect 216 54177 220 54211
rect 186 54100 220 54134
rect 282 54131 292 54243
rect 318 54236 335 54246
rect 318 54167 324 54236
rect 346 54167 348 54252
rect 428 54209 430 54256
rect 476 54219 480 54287
rect 485 54269 495 54297
rect 505 54297 519 54303
rect 544 54297 555 54335
rect 505 54269 525 54297
rect 544 54269 553 54297
rect 544 54249 548 54269
rect 579 54228 582 54318
rect 612 54300 624 54301
rect 599 54298 649 54300
rect 612 54297 624 54298
rect 610 54290 632 54297
rect 607 54289 632 54290
rect 586 54282 644 54289
rect 607 54281 644 54282
rect 607 54265 610 54281
rect 616 54265 644 54281
rect 607 54264 644 54265
rect 586 54257 644 54264
rect 607 54256 610 54257
rect 612 54249 632 54257
rect 612 54245 624 54249
rect 649 54248 651 54298
rect 544 54211 548 54219
rect 400 54179 408 54209
rect 420 54179 436 54209
rect 400 54175 436 54179
rect 400 54167 430 54175
rect 428 54151 430 54167
rect 476 54139 480 54207
rect 544 54177 552 54211
rect 578 54177 582 54211
rect 544 54169 548 54177
rect 544 54139 586 54140
rect 288 54099 292 54131
rect 296 54129 368 54137
rect 378 54129 450 54137
rect 544 54132 548 54139
rect 439 54101 444 54129
rect 120 54085 170 54087
rect 76 54081 130 54085
rect 110 54076 130 54081
rect 60 54051 67 54061
rect 76 54051 77 54071
rect 96 54042 99 54076
rect 109 54051 110 54071
rect 119 54051 126 54061
rect 76 54035 92 54041
rect 94 54035 110 54041
rect 170 54035 172 54085
rect 186 54019 190 54053
rect 216 54019 220 54053
rect 213 53987 224 54019
rect 282 54015 292 54099
rect 296 54093 368 54101
rect 378 54093 450 54101
rect 468 54098 473 54132
rect 428 54063 430 54079
rect 251 53987 292 54015
rect 318 53994 324 54063
rect 12 53982 62 53984
rect 28 53973 59 53981
rect 62 53973 64 53982
rect 251 53981 263 53987
rect 28 53965 64 53973
rect 127 53973 158 53981
rect 127 53966 182 53973
rect 127 53965 161 53966
rect 59 53949 64 53965
rect 158 53949 161 53965
rect 253 53953 263 53981
rect 273 53953 293 53987
rect 318 53984 335 53994
rect 303 53968 316 53978
rect 318 53968 324 53984
rect 346 53978 348 54063
rect 400 54055 430 54063
rect 476 54061 480 54129
rect 511 54098 582 54132
rect 544 54091 548 54098
rect 400 54051 436 54055
rect 400 54021 408 54051
rect 420 54021 436 54051
rect 544 54053 548 54061
rect 28 53941 64 53949
rect 127 53948 161 53949
rect 127 53941 182 53948
rect 62 53932 64 53941
rect 282 53895 292 53953
rect 295 53944 324 53968
rect 333 53968 353 53978
rect 428 53974 430 54021
rect 476 53981 480 54049
rect 544 54019 552 54053
rect 578 54019 582 54053
rect 544 54011 548 54019
rect 367 53968 380 53974
rect 333 53944 380 53968
rect 318 53931 324 53944
rect 346 53931 348 53944
rect 367 53940 380 53944
rect 396 53940 408 53974
rect 420 53940 436 53974
rect 544 53971 553 53999
rect 319 53920 346 53931
rect 120 53879 170 53881
rect 76 53873 92 53879
rect 94 53873 110 53879
rect 76 53863 99 53872
rect 60 53853 67 53863
rect 76 53843 77 53863
rect 96 53838 99 53863
rect 109 53843 110 53863
rect 119 53853 126 53863
rect 76 53829 110 53833
rect 170 53829 172 53879
rect 186 53861 190 53895
rect 216 53861 220 53895
rect 182 53823 224 53824
rect 186 53799 220 53816
rect 223 53799 257 53816
rect 182 53782 257 53799
rect 182 53781 224 53782
rect 160 53775 246 53781
rect 288 53775 292 53895
rect 296 53893 368 53901
rect 428 53893 430 53940
rect 476 53903 480 53971
rect 485 53927 495 53961
rect 505 53933 525 53961
rect 505 53927 519 53933
rect 544 53927 555 53971
rect 485 53903 492 53927
rect 579 53912 582 54002
rect 612 53984 624 53985
rect 599 53982 649 53984
rect 612 53981 624 53982
rect 610 53974 632 53981
rect 607 53973 632 53974
rect 586 53966 644 53973
rect 607 53965 644 53966
rect 607 53949 610 53965
rect 616 53949 644 53965
rect 607 53948 644 53949
rect 586 53941 644 53948
rect 607 53940 610 53941
rect 612 53933 632 53941
rect 612 53929 624 53933
rect 649 53932 651 53982
rect 544 53895 548 53903
rect 400 53863 408 53893
rect 420 53863 436 53893
rect 400 53859 436 53863
rect 400 53851 430 53859
rect 428 53835 430 53851
rect 476 53823 480 53891
rect 544 53861 552 53895
rect 578 53861 582 53895
rect 544 53853 548 53861
rect 295 53782 300 53816
rect 324 53782 329 53816
rect 378 53813 450 53821
rect 544 53818 548 53823
rect 544 53814 582 53818
rect 544 53799 552 53814
rect 578 53799 582 53814
rect 544 53781 586 53799
rect 522 53775 608 53781
rect 182 53759 224 53775
rect 544 53759 586 53775
rect 17 53745 67 53747
rect 119 53745 169 53747
rect 186 53745 220 53759
rect 548 53745 582 53759
rect 599 53745 649 53747
rect 42 53703 59 53737
rect 67 53695 69 53745
rect 160 53737 246 53745
rect 522 53737 608 53745
rect 76 53703 110 53737
rect 127 53703 144 53737
rect 152 53703 161 53737
rect 162 53735 195 53737
rect 224 53735 244 53737
rect 162 53703 244 53735
rect 524 53735 548 53737
rect 573 53735 582 53737
rect 586 53735 606 53737
rect 160 53695 246 53703
rect 186 53679 220 53695
rect 182 53665 224 53666
rect 160 53659 182 53665
rect 224 53659 246 53665
rect 186 53624 220 53658
rect 223 53624 257 53658
rect 120 53611 170 53613
rect 76 53607 130 53611
rect 110 53602 130 53607
rect 60 53577 67 53587
rect 76 53577 77 53597
rect 96 53568 99 53602
rect 109 53577 110 53597
rect 119 53577 126 53587
rect 76 53561 92 53567
rect 94 53561 110 53567
rect 170 53561 172 53611
rect 186 53545 190 53579
rect 216 53545 220 53579
rect 288 53545 292 53733
rect 476 53665 480 53733
rect 524 53703 606 53735
rect 607 53703 616 53737
rect 522 53695 608 53703
rect 649 53695 651 53745
rect 548 53679 582 53695
rect 522 53660 548 53665
rect 522 53659 582 53660
rect 586 53659 608 53665
rect 295 53624 300 53658
rect 324 53624 329 53658
rect 544 53656 582 53659
rect 378 53619 450 53627
rect 428 53589 430 53605
rect 400 53581 430 53589
rect 476 53587 480 53655
rect 544 53626 552 53656
rect 578 53626 582 53656
rect 544 53617 548 53626
rect 400 53577 436 53581
rect 400 53547 408 53577
rect 420 53547 436 53577
rect 544 53579 548 53587
rect 12 53508 62 53510
rect 28 53499 59 53507
rect 62 53499 64 53508
rect 28 53491 64 53499
rect 127 53499 158 53507
rect 127 53492 182 53499
rect 215 53497 224 53525
rect 127 53491 161 53492
rect 59 53475 64 53491
rect 158 53475 161 53491
rect 28 53467 64 53475
rect 127 53474 161 53475
rect 127 53467 182 53474
rect 62 53458 64 53467
rect 213 53459 224 53497
rect 282 53487 292 53545
rect 296 53539 368 53547
rect 319 53509 346 53520
rect 318 53496 324 53509
rect 346 53496 348 53509
rect 428 53500 430 53547
rect 443 53537 450 53539
rect 476 53507 480 53575
rect 544 53545 552 53579
rect 578 53545 582 53579
rect 481 53513 517 53541
rect 481 53507 495 53513
rect 367 53496 380 53500
rect 251 53453 263 53487
rect 273 53453 293 53487
rect 295 53472 324 53496
rect 303 53462 316 53472
rect 318 53456 324 53472
rect 333 53472 380 53496
rect 333 53462 353 53472
rect 367 53466 380 53472
rect 396 53466 408 53500
rect 420 53466 436 53500
rect 120 53405 170 53407
rect 76 53399 92 53405
rect 94 53399 110 53405
rect 76 53389 99 53398
rect 60 53379 67 53389
rect 76 53369 77 53389
rect 96 53364 99 53389
rect 109 53369 110 53389
rect 119 53379 126 53389
rect 76 53355 110 53359
rect 170 53355 172 53405
rect 186 53387 190 53421
rect 216 53387 220 53421
rect 186 53310 220 53344
rect 282 53341 292 53453
rect 318 53446 335 53456
rect 318 53377 324 53446
rect 346 53377 348 53462
rect 428 53419 430 53466
rect 476 53429 480 53497
rect 485 53479 495 53507
rect 505 53507 519 53513
rect 544 53507 555 53545
rect 505 53479 525 53507
rect 544 53479 553 53507
rect 544 53459 548 53479
rect 579 53438 582 53528
rect 612 53510 624 53511
rect 599 53508 649 53510
rect 612 53507 624 53508
rect 610 53500 632 53507
rect 607 53499 632 53500
rect 586 53492 644 53499
rect 607 53491 644 53492
rect 607 53475 610 53491
rect 616 53475 644 53491
rect 607 53474 644 53475
rect 586 53467 644 53474
rect 607 53466 610 53467
rect 612 53459 632 53467
rect 612 53455 624 53459
rect 649 53458 651 53508
rect 544 53421 548 53429
rect 400 53389 408 53419
rect 420 53389 436 53419
rect 400 53385 436 53389
rect 400 53377 430 53385
rect 428 53361 430 53377
rect 476 53349 480 53417
rect 544 53387 552 53421
rect 578 53387 582 53421
rect 544 53379 548 53387
rect 544 53349 586 53350
rect 288 53309 292 53341
rect 296 53339 368 53347
rect 378 53339 450 53347
rect 544 53342 548 53349
rect 439 53311 444 53339
rect 120 53295 170 53297
rect 76 53291 130 53295
rect 110 53286 130 53291
rect 60 53261 67 53271
rect 76 53261 77 53281
rect 96 53252 99 53286
rect 109 53261 110 53281
rect 119 53261 126 53271
rect 76 53245 92 53251
rect 94 53245 110 53251
rect 170 53245 172 53295
rect 186 53229 190 53263
rect 216 53229 220 53263
rect 213 53197 224 53229
rect 282 53225 292 53309
rect 296 53303 368 53311
rect 378 53303 450 53311
rect 468 53308 473 53342
rect 428 53273 430 53289
rect 251 53197 292 53225
rect 318 53204 324 53273
rect 12 53192 62 53194
rect 28 53183 59 53191
rect 62 53183 64 53192
rect 251 53191 263 53197
rect 28 53175 64 53183
rect 127 53183 158 53191
rect 127 53176 182 53183
rect 127 53175 161 53176
rect 59 53159 64 53175
rect 158 53159 161 53175
rect 253 53163 263 53191
rect 273 53163 293 53197
rect 318 53194 335 53204
rect 303 53178 316 53188
rect 318 53178 324 53194
rect 346 53188 348 53273
rect 400 53265 430 53273
rect 476 53271 480 53339
rect 511 53308 582 53342
rect 544 53301 548 53308
rect 400 53261 436 53265
rect 400 53231 408 53261
rect 420 53231 436 53261
rect 544 53263 548 53271
rect 28 53151 64 53159
rect 127 53158 161 53159
rect 127 53151 182 53158
rect 62 53142 64 53151
rect 282 53105 292 53163
rect 295 53154 324 53178
rect 333 53178 353 53188
rect 428 53184 430 53231
rect 476 53191 480 53259
rect 544 53229 552 53263
rect 578 53229 582 53263
rect 544 53221 548 53229
rect 367 53178 380 53184
rect 333 53154 380 53178
rect 318 53141 324 53154
rect 346 53141 348 53154
rect 367 53150 380 53154
rect 396 53150 408 53184
rect 420 53150 436 53184
rect 544 53181 553 53209
rect 319 53130 346 53141
rect 120 53089 170 53091
rect 76 53083 92 53089
rect 94 53083 110 53089
rect 76 53073 99 53082
rect 60 53063 67 53073
rect 76 53053 77 53073
rect 96 53048 99 53073
rect 109 53053 110 53073
rect 119 53063 126 53073
rect 76 53039 110 53043
rect 170 53039 172 53089
rect 186 53071 190 53105
rect 216 53071 220 53105
rect 182 53033 224 53034
rect 186 53009 220 53026
rect 223 53009 257 53026
rect 182 52992 257 53009
rect 182 52991 224 52992
rect 160 52985 246 52991
rect 288 52985 292 53105
rect 296 53103 368 53111
rect 428 53103 430 53150
rect 476 53113 480 53181
rect 485 53137 495 53171
rect 505 53143 525 53171
rect 505 53137 519 53143
rect 544 53137 555 53181
rect 485 53113 492 53137
rect 579 53122 582 53212
rect 612 53194 624 53195
rect 599 53192 649 53194
rect 612 53191 624 53192
rect 610 53184 632 53191
rect 607 53183 632 53184
rect 586 53176 644 53183
rect 607 53175 644 53176
rect 607 53159 610 53175
rect 616 53159 644 53175
rect 607 53158 644 53159
rect 586 53151 644 53158
rect 607 53150 610 53151
rect 612 53143 632 53151
rect 612 53139 624 53143
rect 649 53142 651 53192
rect 544 53105 548 53113
rect 400 53073 408 53103
rect 420 53073 436 53103
rect 400 53069 436 53073
rect 400 53061 430 53069
rect 428 53045 430 53061
rect 476 53033 480 53101
rect 544 53071 552 53105
rect 578 53071 582 53105
rect 544 53063 548 53071
rect 295 52992 300 53026
rect 324 52992 329 53026
rect 378 53023 450 53031
rect 544 53028 548 53033
rect 544 53024 582 53028
rect 544 53009 552 53024
rect 578 53009 582 53024
rect 544 52991 586 53009
rect 522 52985 608 52991
rect 182 52969 224 52985
rect 544 52969 586 52985
rect 17 52955 67 52957
rect 119 52955 169 52957
rect 186 52955 220 52969
rect 548 52955 582 52969
rect 599 52955 649 52957
rect 42 52913 59 52947
rect 67 52905 69 52955
rect 160 52947 246 52955
rect 522 52947 608 52955
rect 76 52913 110 52947
rect 127 52913 144 52947
rect 152 52913 161 52947
rect 162 52945 195 52947
rect 224 52945 244 52947
rect 162 52913 244 52945
rect 524 52945 548 52947
rect 573 52945 582 52947
rect 586 52945 606 52947
rect 160 52905 246 52913
rect 186 52889 220 52905
rect 182 52875 224 52876
rect 160 52869 182 52875
rect 224 52869 246 52875
rect 186 52834 220 52868
rect 223 52834 257 52868
rect 120 52821 170 52823
rect 76 52817 130 52821
rect 110 52812 130 52817
rect 60 52787 67 52797
rect 76 52787 77 52807
rect 96 52778 99 52812
rect 109 52787 110 52807
rect 119 52787 126 52797
rect 76 52771 92 52777
rect 94 52771 110 52777
rect 170 52771 172 52821
rect 186 52755 190 52789
rect 216 52755 220 52789
rect 288 52755 292 52943
rect 476 52875 480 52943
rect 524 52913 606 52945
rect 607 52913 616 52947
rect 522 52905 608 52913
rect 649 52905 651 52955
rect 548 52889 582 52905
rect 522 52870 548 52875
rect 522 52869 582 52870
rect 586 52869 608 52875
rect 295 52834 300 52868
rect 324 52834 329 52868
rect 544 52866 582 52869
rect 378 52829 450 52837
rect 428 52799 430 52815
rect 400 52791 430 52799
rect 476 52797 480 52865
rect 544 52836 552 52866
rect 578 52836 582 52866
rect 544 52827 548 52836
rect 400 52787 436 52791
rect 400 52757 408 52787
rect 420 52757 436 52787
rect 544 52789 548 52797
rect 12 52718 62 52720
rect 28 52709 59 52717
rect 62 52709 64 52718
rect 28 52701 64 52709
rect 127 52709 158 52717
rect 127 52702 182 52709
rect 215 52707 224 52735
rect 127 52701 161 52702
rect 59 52685 64 52701
rect 158 52685 161 52701
rect 28 52677 64 52685
rect 127 52684 161 52685
rect 127 52677 182 52684
rect 62 52668 64 52677
rect 213 52669 224 52707
rect 282 52697 292 52755
rect 296 52749 368 52757
rect 319 52719 346 52730
rect 318 52706 324 52719
rect 346 52706 348 52719
rect 428 52710 430 52757
rect 443 52747 450 52749
rect 476 52717 480 52785
rect 544 52755 552 52789
rect 578 52755 582 52789
rect 481 52723 517 52751
rect 481 52717 495 52723
rect 367 52706 380 52710
rect 251 52663 263 52697
rect 273 52663 293 52697
rect 295 52682 324 52706
rect 303 52672 316 52682
rect 318 52666 324 52682
rect 333 52682 380 52706
rect 333 52672 353 52682
rect 367 52676 380 52682
rect 396 52676 408 52710
rect 420 52676 436 52710
rect 120 52615 170 52617
rect 76 52609 92 52615
rect 94 52609 110 52615
rect 76 52599 99 52608
rect 60 52589 67 52599
rect 76 52579 77 52599
rect 96 52574 99 52599
rect 109 52579 110 52599
rect 119 52589 126 52599
rect 76 52565 110 52569
rect 170 52565 172 52615
rect 186 52597 190 52631
rect 216 52597 220 52631
rect 186 52520 220 52554
rect 282 52551 292 52663
rect 318 52656 335 52666
rect 318 52587 324 52656
rect 346 52587 348 52672
rect 428 52629 430 52676
rect 476 52639 480 52707
rect 485 52689 495 52717
rect 505 52717 519 52723
rect 544 52717 555 52755
rect 505 52689 525 52717
rect 544 52689 553 52717
rect 544 52669 548 52689
rect 579 52648 582 52738
rect 612 52720 624 52721
rect 599 52718 649 52720
rect 612 52717 624 52718
rect 610 52710 632 52717
rect 607 52709 632 52710
rect 586 52702 644 52709
rect 607 52701 644 52702
rect 607 52685 610 52701
rect 616 52685 644 52701
rect 607 52684 644 52685
rect 586 52677 644 52684
rect 607 52676 610 52677
rect 612 52669 632 52677
rect 612 52665 624 52669
rect 649 52668 651 52718
rect 544 52631 548 52639
rect 400 52599 408 52629
rect 420 52599 436 52629
rect 400 52595 436 52599
rect 400 52587 430 52595
rect 428 52571 430 52587
rect 476 52559 480 52627
rect 544 52597 552 52631
rect 578 52597 582 52631
rect 544 52589 548 52597
rect 544 52559 586 52560
rect 288 52519 292 52551
rect 296 52549 368 52557
rect 378 52549 450 52557
rect 544 52552 548 52559
rect 439 52521 444 52549
rect 120 52505 170 52507
rect 76 52501 130 52505
rect 110 52496 130 52501
rect 60 52471 67 52481
rect 76 52471 77 52491
rect 96 52462 99 52496
rect 109 52471 110 52491
rect 119 52471 126 52481
rect 76 52455 92 52461
rect 94 52455 110 52461
rect 170 52455 172 52505
rect 186 52439 190 52473
rect 216 52439 220 52473
rect 213 52407 224 52439
rect 282 52435 292 52519
rect 296 52513 368 52521
rect 378 52513 450 52521
rect 468 52518 473 52552
rect 428 52483 430 52499
rect 251 52407 292 52435
rect 318 52414 324 52483
rect 12 52402 62 52404
rect 28 52393 59 52401
rect 62 52393 64 52402
rect 251 52401 263 52407
rect 28 52385 64 52393
rect 127 52393 158 52401
rect 127 52386 182 52393
rect 127 52385 161 52386
rect 59 52369 64 52385
rect 158 52369 161 52385
rect 253 52373 263 52401
rect 273 52373 293 52407
rect 318 52404 335 52414
rect 303 52388 316 52398
rect 318 52388 324 52404
rect 346 52398 348 52483
rect 400 52475 430 52483
rect 476 52481 480 52549
rect 511 52518 582 52552
rect 544 52511 548 52518
rect 400 52471 436 52475
rect 400 52441 408 52471
rect 420 52441 436 52471
rect 544 52473 548 52481
rect 28 52361 64 52369
rect 127 52368 161 52369
rect 127 52361 182 52368
rect 62 52352 64 52361
rect 282 52315 292 52373
rect 295 52364 324 52388
rect 333 52388 353 52398
rect 428 52394 430 52441
rect 476 52401 480 52469
rect 544 52439 552 52473
rect 578 52439 582 52473
rect 544 52431 548 52439
rect 367 52388 380 52394
rect 333 52364 380 52388
rect 318 52351 324 52364
rect 346 52351 348 52364
rect 367 52360 380 52364
rect 396 52360 408 52394
rect 420 52360 436 52394
rect 544 52391 553 52419
rect 319 52340 346 52351
rect 120 52299 170 52301
rect 76 52293 92 52299
rect 94 52293 110 52299
rect 76 52283 99 52292
rect 60 52273 67 52283
rect 76 52263 77 52283
rect 96 52258 99 52283
rect 109 52263 110 52283
rect 119 52273 126 52283
rect 76 52249 110 52253
rect 170 52249 172 52299
rect 186 52281 190 52315
rect 216 52281 220 52315
rect 182 52243 224 52244
rect 186 52219 220 52236
rect 223 52219 257 52236
rect 182 52202 257 52219
rect 182 52201 224 52202
rect 160 52195 246 52201
rect 288 52195 292 52315
rect 296 52313 368 52321
rect 428 52313 430 52360
rect 476 52323 480 52391
rect 485 52347 495 52381
rect 505 52353 525 52381
rect 505 52347 519 52353
rect 544 52347 555 52391
rect 485 52323 492 52347
rect 579 52332 582 52422
rect 612 52404 624 52405
rect 599 52402 649 52404
rect 612 52401 624 52402
rect 610 52394 632 52401
rect 607 52393 632 52394
rect 586 52386 644 52393
rect 607 52385 644 52386
rect 607 52369 610 52385
rect 616 52369 644 52385
rect 607 52368 644 52369
rect 586 52361 644 52368
rect 607 52360 610 52361
rect 612 52353 632 52361
rect 612 52349 624 52353
rect 649 52352 651 52402
rect 544 52315 548 52323
rect 400 52283 408 52313
rect 420 52283 436 52313
rect 400 52279 436 52283
rect 400 52271 430 52279
rect 428 52255 430 52271
rect 476 52243 480 52311
rect 544 52281 552 52315
rect 578 52281 582 52315
rect 544 52273 548 52281
rect 295 52202 300 52236
rect 324 52202 329 52236
rect 378 52233 450 52241
rect 544 52238 548 52243
rect 544 52234 582 52238
rect 544 52219 552 52234
rect 578 52219 582 52234
rect 544 52201 586 52219
rect 522 52195 608 52201
rect 182 52179 224 52195
rect 544 52179 586 52195
rect 17 52165 67 52167
rect 119 52165 169 52167
rect 186 52165 220 52179
rect 548 52165 582 52179
rect 599 52165 649 52167
rect 42 52123 59 52157
rect 67 52115 69 52165
rect 160 52157 246 52165
rect 522 52157 608 52165
rect 76 52123 110 52157
rect 127 52123 144 52157
rect 152 52123 161 52157
rect 162 52155 195 52157
rect 224 52155 244 52157
rect 162 52123 244 52155
rect 524 52155 548 52157
rect 573 52155 582 52157
rect 586 52155 606 52157
rect 160 52115 246 52123
rect 186 52099 220 52115
rect 182 52085 224 52086
rect 160 52079 182 52085
rect 224 52079 246 52085
rect 186 52044 220 52078
rect 223 52044 257 52078
rect 120 52031 170 52033
rect 76 52027 130 52031
rect 110 52022 130 52027
rect 60 51997 67 52007
rect 76 51997 77 52017
rect 96 51988 99 52022
rect 109 51997 110 52017
rect 119 51997 126 52007
rect 76 51981 92 51987
rect 94 51981 110 51987
rect 170 51981 172 52031
rect 186 51965 190 51999
rect 216 51965 220 51999
rect 288 51965 292 52153
rect 476 52085 480 52153
rect 524 52123 606 52155
rect 607 52123 616 52157
rect 522 52115 608 52123
rect 649 52115 651 52165
rect 548 52099 582 52115
rect 522 52080 548 52085
rect 522 52079 582 52080
rect 586 52079 608 52085
rect 295 52044 300 52078
rect 324 52044 329 52078
rect 544 52076 582 52079
rect 378 52039 450 52047
rect 428 52009 430 52025
rect 400 52001 430 52009
rect 476 52007 480 52075
rect 544 52046 552 52076
rect 578 52046 582 52076
rect 544 52037 548 52046
rect 400 51997 436 52001
rect 400 51967 408 51997
rect 420 51967 436 51997
rect 544 51999 548 52007
rect 12 51928 62 51930
rect 28 51919 59 51927
rect 62 51919 64 51928
rect 28 51911 64 51919
rect 127 51919 158 51927
rect 127 51912 182 51919
rect 215 51917 224 51945
rect 127 51911 161 51912
rect 59 51895 64 51911
rect 158 51895 161 51911
rect 28 51887 64 51895
rect 127 51894 161 51895
rect 127 51887 182 51894
rect 62 51878 64 51887
rect 213 51879 224 51917
rect 282 51907 292 51965
rect 296 51959 368 51967
rect 319 51929 346 51940
rect 318 51916 324 51929
rect 346 51916 348 51929
rect 428 51920 430 51967
rect 443 51957 450 51959
rect 476 51927 480 51995
rect 544 51965 552 51999
rect 578 51965 582 51999
rect 481 51933 517 51961
rect 481 51927 495 51933
rect 367 51916 380 51920
rect 251 51873 263 51907
rect 273 51873 293 51907
rect 295 51892 324 51916
rect 303 51882 316 51892
rect 318 51876 324 51892
rect 333 51892 380 51916
rect 333 51882 353 51892
rect 367 51886 380 51892
rect 396 51886 408 51920
rect 420 51886 436 51920
rect 120 51825 170 51827
rect 76 51819 92 51825
rect 94 51819 110 51825
rect 76 51809 99 51818
rect 60 51799 67 51809
rect 76 51789 77 51809
rect 96 51784 99 51809
rect 109 51789 110 51809
rect 119 51799 126 51809
rect 76 51775 110 51779
rect 170 51775 172 51825
rect 186 51807 190 51841
rect 216 51807 220 51841
rect 186 51730 220 51764
rect 282 51761 292 51873
rect 318 51866 335 51876
rect 318 51797 324 51866
rect 346 51797 348 51882
rect 428 51839 430 51886
rect 476 51849 480 51917
rect 485 51899 495 51927
rect 505 51927 519 51933
rect 544 51927 555 51965
rect 505 51899 525 51927
rect 544 51899 553 51927
rect 544 51879 548 51899
rect 579 51858 582 51948
rect 612 51930 624 51931
rect 599 51928 649 51930
rect 612 51927 624 51928
rect 610 51920 632 51927
rect 607 51919 632 51920
rect 586 51912 644 51919
rect 607 51911 644 51912
rect 607 51895 610 51911
rect 616 51895 644 51911
rect 607 51894 644 51895
rect 586 51887 644 51894
rect 607 51886 610 51887
rect 612 51879 632 51887
rect 612 51875 624 51879
rect 649 51878 651 51928
rect 544 51841 548 51849
rect 400 51809 408 51839
rect 420 51809 436 51839
rect 400 51805 436 51809
rect 400 51797 430 51805
rect 428 51781 430 51797
rect 476 51769 480 51837
rect 544 51807 552 51841
rect 578 51807 582 51841
rect 544 51799 548 51807
rect 544 51769 586 51770
rect 288 51729 292 51761
rect 296 51759 368 51767
rect 378 51759 450 51767
rect 544 51762 548 51769
rect 439 51731 444 51759
rect 120 51715 170 51717
rect 76 51711 130 51715
rect 110 51706 130 51711
rect 60 51681 67 51691
rect 76 51681 77 51701
rect 96 51672 99 51706
rect 109 51681 110 51701
rect 119 51681 126 51691
rect 76 51665 92 51671
rect 94 51665 110 51671
rect 170 51665 172 51715
rect 186 51649 190 51683
rect 216 51649 220 51683
rect 213 51617 224 51649
rect 282 51645 292 51729
rect 296 51723 368 51731
rect 378 51723 450 51731
rect 468 51728 473 51762
rect 428 51693 430 51709
rect 251 51617 292 51645
rect 318 51624 324 51693
rect 12 51612 62 51614
rect 28 51603 59 51611
rect 62 51603 64 51612
rect 251 51611 263 51617
rect 28 51595 64 51603
rect 127 51603 158 51611
rect 127 51596 182 51603
rect 127 51595 161 51596
rect 59 51579 64 51595
rect 158 51579 161 51595
rect 253 51583 263 51611
rect 273 51583 293 51617
rect 318 51614 335 51624
rect 303 51598 316 51608
rect 318 51598 324 51614
rect 346 51608 348 51693
rect 400 51685 430 51693
rect 476 51691 480 51759
rect 511 51728 582 51762
rect 544 51721 548 51728
rect 400 51681 436 51685
rect 400 51651 408 51681
rect 420 51651 436 51681
rect 544 51683 548 51691
rect 28 51571 64 51579
rect 127 51578 161 51579
rect 127 51571 182 51578
rect 62 51562 64 51571
rect 282 51525 292 51583
rect 295 51574 324 51598
rect 333 51598 353 51608
rect 428 51604 430 51651
rect 476 51611 480 51679
rect 544 51649 552 51683
rect 578 51649 582 51683
rect 544 51641 548 51649
rect 367 51598 380 51604
rect 333 51574 380 51598
rect 318 51561 324 51574
rect 346 51561 348 51574
rect 367 51570 380 51574
rect 396 51570 408 51604
rect 420 51570 436 51604
rect 544 51601 553 51629
rect 319 51550 346 51561
rect 120 51509 170 51511
rect 76 51503 92 51509
rect 94 51503 110 51509
rect 76 51493 99 51502
rect 60 51483 67 51493
rect 76 51473 77 51493
rect 96 51468 99 51493
rect 109 51473 110 51493
rect 119 51483 126 51493
rect 76 51459 110 51463
rect 170 51459 172 51509
rect 186 51491 190 51525
rect 216 51491 220 51525
rect 182 51453 224 51454
rect 186 51429 220 51446
rect 223 51429 257 51446
rect 182 51412 257 51429
rect 182 51411 224 51412
rect 160 51405 246 51411
rect 288 51405 292 51525
rect 296 51523 368 51531
rect 428 51523 430 51570
rect 476 51533 480 51601
rect 485 51557 495 51591
rect 505 51563 525 51591
rect 505 51557 519 51563
rect 544 51557 555 51601
rect 485 51533 492 51557
rect 579 51542 582 51632
rect 612 51614 624 51615
rect 599 51612 649 51614
rect 612 51611 624 51612
rect 610 51604 632 51611
rect 607 51603 632 51604
rect 586 51596 644 51603
rect 607 51595 644 51596
rect 607 51579 610 51595
rect 616 51579 644 51595
rect 607 51578 644 51579
rect 586 51571 644 51578
rect 607 51570 610 51571
rect 612 51563 632 51571
rect 612 51559 624 51563
rect 649 51562 651 51612
rect 544 51525 548 51533
rect 400 51493 408 51523
rect 420 51493 436 51523
rect 400 51489 436 51493
rect 400 51481 430 51489
rect 428 51465 430 51481
rect 476 51453 480 51521
rect 544 51491 552 51525
rect 578 51491 582 51525
rect 544 51483 548 51491
rect 295 51412 300 51446
rect 324 51412 329 51446
rect 378 51443 450 51451
rect 544 51448 548 51453
rect 544 51444 582 51448
rect 544 51429 552 51444
rect 578 51429 582 51444
rect 544 51411 586 51429
rect 522 51405 608 51411
rect 182 51389 224 51405
rect 544 51389 586 51405
rect 17 51375 67 51377
rect 119 51375 169 51377
rect 186 51375 220 51389
rect 548 51375 582 51389
rect 599 51375 649 51377
rect 42 51333 59 51367
rect 67 51325 69 51375
rect 160 51367 246 51375
rect 522 51367 608 51375
rect 76 51333 110 51367
rect 127 51333 144 51367
rect 152 51333 161 51367
rect 162 51365 195 51367
rect 224 51365 244 51367
rect 162 51333 244 51365
rect 524 51365 548 51367
rect 573 51365 582 51367
rect 586 51365 606 51367
rect 160 51325 246 51333
rect 186 51309 220 51325
rect 182 51295 224 51296
rect 160 51289 182 51295
rect 224 51289 246 51295
rect 186 51254 220 51288
rect 223 51254 257 51288
rect 120 51241 170 51243
rect 76 51237 130 51241
rect 110 51232 130 51237
rect 60 51207 67 51217
rect 76 51207 77 51227
rect 96 51198 99 51232
rect 109 51207 110 51227
rect 119 51207 126 51217
rect 76 51191 92 51197
rect 94 51191 110 51197
rect 170 51191 172 51241
rect 186 51175 190 51209
rect 216 51175 220 51209
rect 288 51175 292 51363
rect 476 51295 480 51363
rect 524 51333 606 51365
rect 607 51333 616 51367
rect 522 51325 608 51333
rect 649 51325 651 51375
rect 548 51309 582 51325
rect 522 51290 548 51295
rect 522 51289 582 51290
rect 586 51289 608 51295
rect 295 51254 300 51288
rect 324 51254 329 51288
rect 544 51286 582 51289
rect 378 51249 450 51257
rect 428 51219 430 51235
rect 400 51211 430 51219
rect 476 51217 480 51285
rect 544 51256 552 51286
rect 578 51256 582 51286
rect 544 51247 548 51256
rect 400 51207 436 51211
rect 400 51177 408 51207
rect 420 51177 436 51207
rect 544 51209 548 51217
rect 12 51138 62 51140
rect 28 51129 59 51137
rect 62 51129 64 51138
rect 28 51121 64 51129
rect 127 51129 158 51137
rect 127 51122 182 51129
rect 215 51127 224 51155
rect 127 51121 161 51122
rect 59 51105 64 51121
rect 158 51105 161 51121
rect 28 51097 64 51105
rect 127 51104 161 51105
rect 127 51097 182 51104
rect 62 51088 64 51097
rect 213 51089 224 51127
rect 282 51117 292 51175
rect 296 51169 368 51177
rect 319 51139 346 51150
rect 318 51126 324 51139
rect 346 51126 348 51139
rect 428 51130 430 51177
rect 443 51167 450 51169
rect 476 51137 480 51205
rect 544 51175 552 51209
rect 578 51175 582 51209
rect 481 51143 517 51171
rect 481 51137 495 51143
rect 367 51126 380 51130
rect 251 51083 263 51117
rect 273 51083 293 51117
rect 295 51102 324 51126
rect 303 51092 316 51102
rect 318 51086 324 51102
rect 333 51102 380 51126
rect 333 51092 353 51102
rect 367 51096 380 51102
rect 396 51096 408 51130
rect 420 51096 436 51130
rect 120 51035 170 51037
rect 76 51029 92 51035
rect 94 51029 110 51035
rect 76 51019 99 51028
rect 60 51009 67 51019
rect 76 50999 77 51019
rect 96 50994 99 51019
rect 109 50999 110 51019
rect 119 51009 126 51019
rect 76 50985 110 50989
rect 170 50985 172 51035
rect 186 51017 190 51051
rect 216 51017 220 51051
rect 186 50940 220 50974
rect 282 50971 292 51083
rect 318 51076 335 51086
rect 318 51007 324 51076
rect 346 51007 348 51092
rect 428 51049 430 51096
rect 476 51059 480 51127
rect 485 51109 495 51137
rect 505 51137 519 51143
rect 544 51137 555 51175
rect 505 51109 525 51137
rect 544 51109 553 51137
rect 544 51089 548 51109
rect 579 51068 582 51158
rect 612 51140 624 51141
rect 599 51138 649 51140
rect 612 51137 624 51138
rect 610 51130 632 51137
rect 607 51129 632 51130
rect 586 51122 644 51129
rect 607 51121 644 51122
rect 607 51105 610 51121
rect 616 51105 644 51121
rect 607 51104 644 51105
rect 586 51097 644 51104
rect 607 51096 610 51097
rect 612 51089 632 51097
rect 612 51085 624 51089
rect 649 51088 651 51138
rect 544 51051 548 51059
rect 400 51019 408 51049
rect 420 51019 436 51049
rect 400 51015 436 51019
rect 400 51007 430 51015
rect 428 50991 430 51007
rect 476 50979 480 51047
rect 544 51017 552 51051
rect 578 51017 582 51051
rect 544 51009 548 51017
rect 544 50979 586 50980
rect 288 50939 292 50971
rect 296 50969 368 50977
rect 378 50969 450 50977
rect 544 50972 548 50979
rect 439 50941 444 50969
rect 120 50925 170 50927
rect 76 50921 130 50925
rect 110 50916 130 50921
rect 60 50891 67 50901
rect 76 50891 77 50911
rect 96 50882 99 50916
rect 109 50891 110 50911
rect 119 50891 126 50901
rect 76 50875 92 50881
rect 94 50875 110 50881
rect 170 50875 172 50925
rect 186 50859 190 50893
rect 216 50859 220 50893
rect 213 50827 224 50859
rect 282 50855 292 50939
rect 296 50933 368 50941
rect 378 50933 450 50941
rect 468 50938 473 50972
rect 428 50903 430 50919
rect 251 50827 292 50855
rect 318 50834 324 50903
rect 12 50822 62 50824
rect 28 50813 59 50821
rect 62 50813 64 50822
rect 251 50821 263 50827
rect 28 50805 64 50813
rect 127 50813 158 50821
rect 127 50806 182 50813
rect 127 50805 161 50806
rect 59 50789 64 50805
rect 158 50789 161 50805
rect 253 50793 263 50821
rect 273 50793 293 50827
rect 318 50824 335 50834
rect 303 50808 316 50818
rect 318 50808 324 50824
rect 346 50818 348 50903
rect 400 50895 430 50903
rect 476 50901 480 50969
rect 511 50938 582 50972
rect 544 50931 548 50938
rect 400 50891 436 50895
rect 400 50861 408 50891
rect 420 50861 436 50891
rect 544 50893 548 50901
rect 28 50781 64 50789
rect 127 50788 161 50789
rect 127 50781 182 50788
rect 62 50772 64 50781
rect 282 50735 292 50793
rect 295 50784 324 50808
rect 333 50808 353 50818
rect 428 50814 430 50861
rect 476 50821 480 50889
rect 544 50859 552 50893
rect 578 50859 582 50893
rect 544 50851 548 50859
rect 367 50808 380 50814
rect 333 50784 380 50808
rect 318 50771 324 50784
rect 346 50771 348 50784
rect 367 50780 380 50784
rect 396 50780 408 50814
rect 420 50780 436 50814
rect 544 50811 553 50839
rect 319 50760 346 50771
rect 120 50719 170 50721
rect 76 50713 92 50719
rect 94 50713 110 50719
rect 76 50703 99 50712
rect 60 50693 67 50703
rect 76 50683 77 50703
rect 96 50678 99 50703
rect 109 50683 110 50703
rect 119 50693 126 50703
rect 76 50669 110 50673
rect 170 50669 172 50719
rect 186 50701 190 50735
rect 216 50701 220 50735
rect 182 50663 224 50664
rect 186 50639 220 50656
rect 223 50639 257 50656
rect 182 50622 257 50639
rect 182 50621 224 50622
rect 160 50615 246 50621
rect 288 50615 292 50735
rect 296 50733 368 50741
rect 428 50733 430 50780
rect 476 50743 480 50811
rect 485 50767 495 50801
rect 505 50773 525 50801
rect 505 50767 519 50773
rect 544 50767 555 50811
rect 485 50743 492 50767
rect 579 50752 582 50842
rect 612 50824 624 50825
rect 599 50822 649 50824
rect 612 50821 624 50822
rect 610 50814 632 50821
rect 607 50813 632 50814
rect 586 50806 644 50813
rect 607 50805 644 50806
rect 607 50789 610 50805
rect 616 50789 644 50805
rect 607 50788 644 50789
rect 586 50781 644 50788
rect 607 50780 610 50781
rect 612 50773 632 50781
rect 612 50769 624 50773
rect 649 50772 651 50822
rect 544 50735 548 50743
rect 400 50703 408 50733
rect 420 50703 436 50733
rect 400 50699 436 50703
rect 400 50691 430 50699
rect 428 50675 430 50691
rect 476 50663 480 50731
rect 544 50701 552 50735
rect 578 50701 582 50735
rect 544 50693 548 50701
rect 295 50622 300 50656
rect 324 50622 329 50656
rect 378 50653 450 50661
rect 544 50658 548 50663
rect 544 50654 582 50658
rect 544 50639 552 50654
rect 578 50639 582 50654
rect 544 50621 586 50639
rect 522 50615 608 50621
rect 182 50599 224 50615
rect 544 50599 586 50615
rect 17 50585 67 50587
rect 119 50585 169 50587
rect 186 50585 220 50599
rect 548 50585 582 50599
rect 599 50585 649 50587
rect 42 50543 59 50577
rect 67 50535 69 50585
rect 160 50577 246 50585
rect 522 50577 608 50585
rect 76 50543 110 50577
rect 127 50543 144 50577
rect 152 50543 161 50577
rect 162 50575 195 50577
rect 224 50575 244 50577
rect 162 50543 244 50575
rect 524 50575 548 50577
rect 573 50575 582 50577
rect 586 50575 606 50577
rect 160 50535 246 50543
rect 186 50519 220 50535
rect 182 50505 224 50506
rect 160 50499 182 50505
rect 224 50499 246 50505
rect 186 50464 220 50498
rect 223 50464 257 50498
rect 120 50451 170 50453
rect 76 50447 130 50451
rect 110 50442 130 50447
rect 60 50417 67 50427
rect 76 50417 77 50437
rect 96 50408 99 50442
rect 109 50417 110 50437
rect 119 50417 126 50427
rect 76 50401 92 50407
rect 94 50401 110 50407
rect 170 50401 172 50451
rect 186 50385 190 50419
rect 216 50385 220 50419
rect 288 50385 292 50573
rect 476 50505 480 50573
rect 524 50543 606 50575
rect 607 50543 616 50577
rect 522 50535 608 50543
rect 649 50535 651 50585
rect 548 50519 582 50535
rect 522 50500 548 50505
rect 522 50499 582 50500
rect 586 50499 608 50505
rect 295 50464 300 50498
rect 324 50464 329 50498
rect 544 50496 582 50499
rect 378 50459 450 50467
rect 428 50429 430 50445
rect 400 50421 430 50429
rect 476 50427 480 50495
rect 544 50466 552 50496
rect 578 50466 582 50496
rect 544 50457 548 50466
rect 400 50417 436 50421
rect 400 50387 408 50417
rect 420 50387 436 50417
rect 544 50419 548 50427
rect 12 50348 62 50350
rect 28 50339 59 50347
rect 62 50339 64 50348
rect 28 50331 64 50339
rect 127 50339 158 50347
rect 127 50332 182 50339
rect 215 50337 224 50365
rect 127 50331 161 50332
rect 59 50315 64 50331
rect 158 50315 161 50331
rect 28 50307 64 50315
rect 127 50314 161 50315
rect 127 50307 182 50314
rect 62 50298 64 50307
rect 213 50299 224 50337
rect 282 50327 292 50385
rect 296 50379 368 50387
rect 319 50349 346 50360
rect 318 50336 324 50349
rect 346 50336 348 50349
rect 428 50340 430 50387
rect 443 50377 450 50379
rect 476 50347 480 50415
rect 544 50385 552 50419
rect 578 50385 582 50419
rect 481 50353 517 50381
rect 481 50347 495 50353
rect 367 50336 380 50340
rect 251 50293 263 50327
rect 273 50293 293 50327
rect 295 50312 324 50336
rect 303 50302 316 50312
rect 318 50296 324 50312
rect 333 50312 380 50336
rect 333 50302 353 50312
rect 367 50306 380 50312
rect 396 50306 408 50340
rect 420 50306 436 50340
rect 120 50245 170 50247
rect 76 50239 92 50245
rect 94 50239 110 50245
rect 76 50229 99 50238
rect 60 50219 67 50229
rect 76 50209 77 50229
rect 96 50204 99 50229
rect 109 50209 110 50229
rect 119 50219 126 50229
rect 76 50195 110 50199
rect 170 50195 172 50245
rect 186 50227 190 50261
rect 216 50227 220 50261
rect 186 50150 220 50184
rect 282 50181 292 50293
rect 318 50286 335 50296
rect 318 50217 324 50286
rect 346 50217 348 50302
rect 428 50259 430 50306
rect 476 50269 480 50337
rect 485 50319 495 50347
rect 505 50347 519 50353
rect 544 50347 555 50385
rect 505 50319 525 50347
rect 544 50319 553 50347
rect 544 50299 548 50319
rect 579 50278 582 50368
rect 612 50350 624 50351
rect 599 50348 649 50350
rect 612 50347 624 50348
rect 610 50340 632 50347
rect 607 50339 632 50340
rect 586 50332 644 50339
rect 607 50331 644 50332
rect 607 50315 610 50331
rect 616 50315 644 50331
rect 607 50314 644 50315
rect 586 50307 644 50314
rect 607 50306 610 50307
rect 612 50299 632 50307
rect 612 50295 624 50299
rect 649 50298 651 50348
rect 544 50261 548 50269
rect 400 50229 408 50259
rect 420 50229 436 50259
rect 400 50225 436 50229
rect 400 50217 430 50225
rect 428 50201 430 50217
rect 476 50189 480 50257
rect 544 50227 552 50261
rect 578 50227 582 50261
rect 544 50219 548 50227
rect 544 50189 586 50190
rect 288 50149 292 50181
rect 296 50179 368 50187
rect 378 50179 450 50187
rect 544 50182 548 50189
rect 439 50151 444 50179
rect 120 50135 170 50137
rect 76 50131 130 50135
rect 110 50126 130 50131
rect 60 50101 67 50111
rect 76 50101 77 50121
rect 96 50092 99 50126
rect 109 50101 110 50121
rect 119 50101 126 50111
rect 76 50085 92 50091
rect 94 50085 110 50091
rect 170 50085 172 50135
rect 186 50069 190 50103
rect 216 50069 220 50103
rect 213 50037 224 50069
rect 282 50065 292 50149
rect 296 50143 368 50151
rect 378 50143 450 50151
rect 468 50148 473 50182
rect 428 50113 430 50129
rect 251 50037 292 50065
rect 318 50044 324 50113
rect 12 50032 62 50034
rect 28 50023 59 50031
rect 62 50023 64 50032
rect 251 50031 263 50037
rect 28 50015 64 50023
rect 127 50023 158 50031
rect 127 50016 182 50023
rect 127 50015 161 50016
rect 59 49999 64 50015
rect 158 49999 161 50015
rect 253 50003 263 50031
rect 273 50003 293 50037
rect 318 50034 335 50044
rect 303 50018 316 50028
rect 318 50018 324 50034
rect 346 50028 348 50113
rect 400 50105 430 50113
rect 476 50111 480 50179
rect 511 50148 582 50182
rect 544 50141 548 50148
rect 400 50101 436 50105
rect 400 50071 408 50101
rect 420 50071 436 50101
rect 544 50103 548 50111
rect 28 49991 64 49999
rect 127 49998 161 49999
rect 127 49991 182 49998
rect 62 49982 64 49991
rect 282 49945 292 50003
rect 295 49994 324 50018
rect 333 50018 353 50028
rect 428 50024 430 50071
rect 476 50031 480 50099
rect 544 50069 552 50103
rect 578 50069 582 50103
rect 544 50061 548 50069
rect 367 50018 380 50024
rect 333 49994 380 50018
rect 318 49981 324 49994
rect 346 49981 348 49994
rect 367 49990 380 49994
rect 396 49990 408 50024
rect 420 49990 436 50024
rect 544 50021 553 50049
rect 319 49970 346 49981
rect 120 49929 170 49931
rect 76 49923 92 49929
rect 94 49923 110 49929
rect 76 49913 99 49922
rect 60 49903 67 49913
rect 76 49893 77 49913
rect 96 49888 99 49913
rect 109 49893 110 49913
rect 119 49903 126 49913
rect 76 49879 110 49883
rect 170 49879 172 49929
rect 186 49911 190 49945
rect 216 49911 220 49945
rect 182 49873 224 49874
rect 186 49849 220 49866
rect 223 49849 257 49866
rect 182 49832 257 49849
rect 182 49831 224 49832
rect 160 49825 246 49831
rect 288 49825 292 49945
rect 296 49943 368 49951
rect 428 49943 430 49990
rect 476 49953 480 50021
rect 485 49977 495 50011
rect 505 49983 525 50011
rect 505 49977 519 49983
rect 544 49977 555 50021
rect 485 49953 492 49977
rect 579 49962 582 50052
rect 612 50034 624 50035
rect 599 50032 649 50034
rect 612 50031 624 50032
rect 610 50024 632 50031
rect 607 50023 632 50024
rect 586 50016 644 50023
rect 607 50015 644 50016
rect 607 49999 610 50015
rect 616 49999 644 50015
rect 607 49998 644 49999
rect 586 49991 644 49998
rect 607 49990 610 49991
rect 612 49983 632 49991
rect 612 49979 624 49983
rect 649 49982 651 50032
rect 544 49945 548 49953
rect 400 49913 408 49943
rect 420 49913 436 49943
rect 400 49909 436 49913
rect 400 49901 430 49909
rect 428 49885 430 49901
rect 476 49873 480 49941
rect 544 49911 552 49945
rect 578 49911 582 49945
rect 544 49903 548 49911
rect 295 49832 300 49866
rect 324 49832 329 49866
rect 378 49863 450 49871
rect 544 49868 548 49873
rect 544 49864 582 49868
rect 544 49849 552 49864
rect 578 49849 582 49864
rect 544 49831 586 49849
rect 522 49825 608 49831
rect 182 49809 224 49825
rect 544 49809 586 49825
rect 17 49795 67 49797
rect 119 49795 169 49797
rect 186 49795 220 49809
rect 548 49795 582 49809
rect 599 49795 649 49797
rect 42 49753 59 49787
rect 67 49745 69 49795
rect 160 49787 246 49795
rect 522 49787 608 49795
rect 76 49753 110 49787
rect 127 49753 144 49787
rect 152 49753 161 49787
rect 162 49785 195 49787
rect 224 49785 244 49787
rect 162 49753 244 49785
rect 524 49785 548 49787
rect 573 49785 582 49787
rect 586 49785 606 49787
rect 160 49745 246 49753
rect 186 49729 220 49745
rect 182 49715 224 49716
rect 160 49709 182 49715
rect 224 49709 246 49715
rect 186 49674 220 49708
rect 223 49674 257 49708
rect 120 49661 170 49663
rect 76 49657 130 49661
rect 110 49652 130 49657
rect 60 49627 67 49637
rect 76 49627 77 49647
rect 96 49618 99 49652
rect 109 49627 110 49647
rect 119 49627 126 49637
rect 76 49611 92 49617
rect 94 49611 110 49617
rect 170 49611 172 49661
rect 186 49595 190 49629
rect 216 49595 220 49629
rect 288 49595 292 49783
rect 476 49715 480 49783
rect 524 49753 606 49785
rect 607 49753 616 49787
rect 522 49745 608 49753
rect 649 49745 651 49795
rect 548 49729 582 49745
rect 522 49710 548 49715
rect 522 49709 582 49710
rect 586 49709 608 49715
rect 295 49674 300 49708
rect 324 49674 329 49708
rect 544 49706 582 49709
rect 378 49669 450 49677
rect 428 49639 430 49655
rect 400 49631 430 49639
rect 476 49637 480 49705
rect 544 49676 552 49706
rect 578 49676 582 49706
rect 544 49667 548 49676
rect 400 49627 436 49631
rect 400 49597 408 49627
rect 420 49597 436 49627
rect 544 49629 548 49637
rect 12 49558 62 49560
rect 28 49549 59 49557
rect 62 49549 64 49558
rect 28 49541 64 49549
rect 127 49549 158 49557
rect 127 49542 182 49549
rect 215 49547 224 49575
rect 127 49541 161 49542
rect 59 49525 64 49541
rect 158 49525 161 49541
rect 28 49517 64 49525
rect 127 49524 161 49525
rect 127 49517 182 49524
rect 62 49508 64 49517
rect 213 49509 224 49547
rect 282 49537 292 49595
rect 296 49589 368 49597
rect 319 49559 346 49570
rect 318 49546 324 49559
rect 346 49546 348 49559
rect 428 49550 430 49597
rect 443 49587 450 49589
rect 476 49557 480 49625
rect 544 49595 552 49629
rect 578 49595 582 49629
rect 481 49563 517 49591
rect 481 49557 495 49563
rect 367 49546 380 49550
rect 251 49503 263 49537
rect 273 49503 293 49537
rect 295 49522 324 49546
rect 303 49512 316 49522
rect 318 49506 324 49522
rect 333 49522 380 49546
rect 333 49512 353 49522
rect 367 49516 380 49522
rect 396 49516 408 49550
rect 420 49516 436 49550
rect 120 49455 170 49457
rect 76 49449 92 49455
rect 94 49449 110 49455
rect 76 49439 99 49448
rect 60 49429 67 49439
rect 76 49419 77 49439
rect 96 49414 99 49439
rect 109 49419 110 49439
rect 119 49429 126 49439
rect 76 49405 110 49409
rect 170 49405 172 49455
rect 186 49437 190 49471
rect 216 49437 220 49471
rect 186 49360 220 49394
rect 282 49391 292 49503
rect 318 49496 335 49506
rect 318 49427 324 49496
rect 346 49427 348 49512
rect 428 49469 430 49516
rect 476 49479 480 49547
rect 485 49529 495 49557
rect 505 49557 519 49563
rect 544 49557 555 49595
rect 505 49529 525 49557
rect 544 49529 553 49557
rect 544 49509 548 49529
rect 579 49488 582 49578
rect 612 49560 624 49561
rect 599 49558 649 49560
rect 612 49557 624 49558
rect 610 49550 632 49557
rect 607 49549 632 49550
rect 586 49542 644 49549
rect 607 49541 644 49542
rect 607 49525 610 49541
rect 616 49525 644 49541
rect 607 49524 644 49525
rect 586 49517 644 49524
rect 607 49516 610 49517
rect 612 49509 632 49517
rect 612 49505 624 49509
rect 649 49508 651 49558
rect 544 49471 548 49479
rect 400 49439 408 49469
rect 420 49439 436 49469
rect 400 49435 436 49439
rect 400 49427 430 49435
rect 428 49411 430 49427
rect 476 49399 480 49467
rect 544 49437 552 49471
rect 578 49437 582 49471
rect 544 49429 548 49437
rect 544 49399 586 49400
rect 288 49359 292 49391
rect 296 49389 368 49397
rect 378 49389 450 49397
rect 544 49392 548 49399
rect 439 49361 444 49389
rect 120 49345 170 49347
rect 76 49341 130 49345
rect 110 49336 130 49341
rect 60 49311 67 49321
rect 76 49311 77 49331
rect 96 49302 99 49336
rect 109 49311 110 49331
rect 119 49311 126 49321
rect 76 49295 92 49301
rect 94 49295 110 49301
rect 170 49295 172 49345
rect 186 49279 190 49313
rect 216 49279 220 49313
rect 213 49247 224 49279
rect 282 49275 292 49359
rect 296 49353 368 49361
rect 378 49353 450 49361
rect 468 49358 473 49392
rect 428 49323 430 49339
rect 251 49247 292 49275
rect 318 49254 324 49323
rect 12 49242 62 49244
rect 28 49233 59 49241
rect 62 49233 64 49242
rect 251 49241 263 49247
rect 28 49225 64 49233
rect 127 49233 158 49241
rect 127 49226 182 49233
rect 127 49225 161 49226
rect 59 49209 64 49225
rect 158 49209 161 49225
rect 253 49213 263 49241
rect 273 49213 293 49247
rect 318 49244 335 49254
rect 303 49228 316 49238
rect 318 49228 324 49244
rect 346 49238 348 49323
rect 400 49315 430 49323
rect 476 49321 480 49389
rect 511 49358 582 49392
rect 544 49351 548 49358
rect 400 49311 436 49315
rect 400 49281 408 49311
rect 420 49281 436 49311
rect 544 49313 548 49321
rect 28 49201 64 49209
rect 127 49208 161 49209
rect 127 49201 182 49208
rect 62 49192 64 49201
rect 282 49155 292 49213
rect 295 49204 324 49228
rect 333 49228 353 49238
rect 428 49234 430 49281
rect 476 49241 480 49309
rect 544 49279 552 49313
rect 578 49279 582 49313
rect 544 49271 548 49279
rect 367 49228 380 49234
rect 333 49204 380 49228
rect 318 49191 324 49204
rect 346 49191 348 49204
rect 367 49200 380 49204
rect 396 49200 408 49234
rect 420 49200 436 49234
rect 544 49231 553 49259
rect 319 49180 346 49191
rect 120 49139 170 49141
rect 76 49133 92 49139
rect 94 49133 110 49139
rect 76 49123 99 49132
rect 60 49113 67 49123
rect 76 49103 77 49123
rect 96 49098 99 49123
rect 109 49103 110 49123
rect 119 49113 126 49123
rect 76 49089 110 49093
rect 170 49089 172 49139
rect 186 49121 190 49155
rect 216 49121 220 49155
rect 182 49083 224 49084
rect 186 49059 220 49076
rect 223 49059 257 49076
rect 182 49042 257 49059
rect 182 49041 224 49042
rect 160 49035 246 49041
rect 288 49035 292 49155
rect 296 49153 368 49161
rect 428 49153 430 49200
rect 476 49163 480 49231
rect 485 49187 495 49221
rect 505 49193 525 49221
rect 505 49187 519 49193
rect 544 49187 555 49231
rect 485 49163 492 49187
rect 579 49172 582 49262
rect 612 49244 624 49245
rect 599 49242 649 49244
rect 612 49241 624 49242
rect 610 49234 632 49241
rect 607 49233 632 49234
rect 586 49226 644 49233
rect 607 49225 644 49226
rect 607 49209 610 49225
rect 616 49209 644 49225
rect 607 49208 644 49209
rect 586 49201 644 49208
rect 607 49200 610 49201
rect 612 49193 632 49201
rect 612 49189 624 49193
rect 649 49192 651 49242
rect 544 49155 548 49163
rect 400 49123 408 49153
rect 420 49123 436 49153
rect 400 49119 436 49123
rect 400 49111 430 49119
rect 428 49095 430 49111
rect 476 49083 480 49151
rect 544 49121 552 49155
rect 578 49121 582 49155
rect 544 49113 548 49121
rect 295 49042 300 49076
rect 324 49042 329 49076
rect 378 49073 450 49081
rect 544 49078 548 49083
rect 544 49074 582 49078
rect 544 49059 552 49074
rect 578 49059 582 49074
rect 544 49041 586 49059
rect 522 49035 608 49041
rect 182 49019 224 49035
rect 544 49019 586 49035
rect 17 49005 67 49007
rect 119 49005 169 49007
rect 186 49005 220 49019
rect 548 49005 582 49019
rect 599 49005 649 49007
rect 42 48963 59 48997
rect 67 48955 69 49005
rect 160 48997 246 49005
rect 522 48997 608 49005
rect 76 48963 110 48997
rect 127 48963 144 48997
rect 152 48963 161 48997
rect 162 48995 195 48997
rect 224 48995 244 48997
rect 162 48963 244 48995
rect 524 48995 548 48997
rect 573 48995 582 48997
rect 586 48995 606 48997
rect 160 48955 246 48963
rect 186 48939 220 48955
rect 182 48925 224 48926
rect 160 48919 182 48925
rect 224 48919 246 48925
rect 186 48884 220 48918
rect 223 48884 257 48918
rect 120 48871 170 48873
rect 76 48867 130 48871
rect 110 48862 130 48867
rect 60 48837 67 48847
rect 76 48837 77 48857
rect 96 48828 99 48862
rect 109 48837 110 48857
rect 119 48837 126 48847
rect 76 48821 92 48827
rect 94 48821 110 48827
rect 170 48821 172 48871
rect 186 48805 190 48839
rect 216 48805 220 48839
rect 288 48805 292 48993
rect 476 48925 480 48993
rect 524 48963 606 48995
rect 607 48963 616 48997
rect 522 48955 608 48963
rect 649 48955 651 49005
rect 548 48939 582 48955
rect 522 48920 548 48925
rect 522 48919 582 48920
rect 586 48919 608 48925
rect 295 48884 300 48918
rect 324 48884 329 48918
rect 544 48916 582 48919
rect 378 48879 450 48887
rect 428 48849 430 48865
rect 400 48841 430 48849
rect 476 48847 480 48915
rect 544 48886 552 48916
rect 578 48886 582 48916
rect 544 48877 548 48886
rect 400 48837 436 48841
rect 400 48807 408 48837
rect 420 48807 436 48837
rect 544 48839 548 48847
rect 12 48768 62 48770
rect 28 48759 59 48767
rect 62 48759 64 48768
rect 28 48751 64 48759
rect 127 48759 158 48767
rect 127 48752 182 48759
rect 215 48757 224 48785
rect 127 48751 161 48752
rect 59 48735 64 48751
rect 158 48735 161 48751
rect 28 48727 64 48735
rect 127 48734 161 48735
rect 127 48727 182 48734
rect 62 48718 64 48727
rect 213 48719 224 48757
rect 282 48747 292 48805
rect 296 48799 368 48807
rect 319 48769 346 48780
rect 318 48756 324 48769
rect 346 48756 348 48769
rect 428 48760 430 48807
rect 443 48797 450 48799
rect 476 48767 480 48835
rect 544 48805 552 48839
rect 578 48805 582 48839
rect 481 48773 517 48801
rect 481 48767 495 48773
rect 367 48756 380 48760
rect 251 48713 263 48747
rect 273 48713 293 48747
rect 295 48732 324 48756
rect 303 48722 316 48732
rect 318 48716 324 48732
rect 333 48732 380 48756
rect 333 48722 353 48732
rect 367 48726 380 48732
rect 396 48726 408 48760
rect 420 48726 436 48760
rect 120 48665 170 48667
rect 76 48659 92 48665
rect 94 48659 110 48665
rect 76 48649 99 48658
rect 60 48639 67 48649
rect 76 48629 77 48649
rect 96 48624 99 48649
rect 109 48629 110 48649
rect 119 48639 126 48649
rect 76 48615 110 48619
rect 170 48615 172 48665
rect 186 48647 190 48681
rect 216 48647 220 48681
rect 186 48570 220 48604
rect 282 48601 292 48713
rect 318 48706 335 48716
rect 318 48637 324 48706
rect 346 48637 348 48722
rect 428 48679 430 48726
rect 476 48689 480 48757
rect 485 48739 495 48767
rect 505 48767 519 48773
rect 544 48767 555 48805
rect 505 48739 525 48767
rect 544 48739 553 48767
rect 544 48719 548 48739
rect 579 48698 582 48788
rect 612 48770 624 48771
rect 599 48768 649 48770
rect 612 48767 624 48768
rect 610 48760 632 48767
rect 607 48759 632 48760
rect 586 48752 644 48759
rect 607 48751 644 48752
rect 607 48735 610 48751
rect 616 48735 644 48751
rect 607 48734 644 48735
rect 586 48727 644 48734
rect 607 48726 610 48727
rect 612 48719 632 48727
rect 612 48715 624 48719
rect 649 48718 651 48768
rect 544 48681 548 48689
rect 400 48649 408 48679
rect 420 48649 436 48679
rect 400 48645 436 48649
rect 400 48637 430 48645
rect 428 48621 430 48637
rect 476 48609 480 48677
rect 544 48647 552 48681
rect 578 48647 582 48681
rect 544 48639 548 48647
rect 544 48609 586 48610
rect 288 48569 292 48601
rect 296 48599 368 48607
rect 378 48599 450 48607
rect 544 48602 548 48609
rect 439 48571 444 48599
rect 120 48555 170 48557
rect 76 48551 130 48555
rect 110 48546 130 48551
rect 60 48521 67 48531
rect 76 48521 77 48541
rect 96 48512 99 48546
rect 109 48521 110 48541
rect 119 48521 126 48531
rect 76 48505 92 48511
rect 94 48505 110 48511
rect 170 48505 172 48555
rect 186 48489 190 48523
rect 216 48489 220 48523
rect 213 48457 224 48489
rect 282 48485 292 48569
rect 296 48563 368 48571
rect 378 48563 450 48571
rect 468 48568 473 48602
rect 428 48533 430 48549
rect 251 48457 292 48485
rect 318 48464 324 48533
rect 12 48452 62 48454
rect 28 48443 59 48451
rect 62 48443 64 48452
rect 251 48451 263 48457
rect 28 48435 64 48443
rect 127 48443 158 48451
rect 127 48436 182 48443
rect 127 48435 161 48436
rect 59 48419 64 48435
rect 158 48419 161 48435
rect 253 48423 263 48451
rect 273 48423 293 48457
rect 318 48454 335 48464
rect 303 48438 316 48448
rect 318 48438 324 48454
rect 346 48448 348 48533
rect 400 48525 430 48533
rect 476 48531 480 48599
rect 511 48568 582 48602
rect 544 48561 548 48568
rect 400 48521 436 48525
rect 400 48491 408 48521
rect 420 48491 436 48521
rect 544 48523 548 48531
rect 28 48411 64 48419
rect 127 48418 161 48419
rect 127 48411 182 48418
rect 62 48402 64 48411
rect 282 48365 292 48423
rect 295 48414 324 48438
rect 333 48438 353 48448
rect 428 48444 430 48491
rect 476 48451 480 48519
rect 544 48489 552 48523
rect 578 48489 582 48523
rect 544 48481 548 48489
rect 367 48438 380 48444
rect 333 48414 380 48438
rect 318 48401 324 48414
rect 346 48401 348 48414
rect 367 48410 380 48414
rect 396 48410 408 48444
rect 420 48410 436 48444
rect 544 48441 553 48469
rect 319 48390 346 48401
rect 120 48349 170 48351
rect 76 48343 92 48349
rect 94 48343 110 48349
rect 76 48333 99 48342
rect 60 48323 67 48333
rect 76 48313 77 48333
rect 96 48308 99 48333
rect 109 48313 110 48333
rect 119 48323 126 48333
rect 76 48299 110 48303
rect 170 48299 172 48349
rect 186 48331 190 48365
rect 216 48331 220 48365
rect 182 48293 224 48294
rect 186 48269 220 48286
rect 223 48269 257 48286
rect 182 48252 257 48269
rect 182 48251 224 48252
rect 160 48245 246 48251
rect 288 48245 292 48365
rect 296 48363 368 48371
rect 428 48363 430 48410
rect 476 48373 480 48441
rect 485 48397 495 48431
rect 505 48403 525 48431
rect 505 48397 519 48403
rect 544 48397 555 48441
rect 485 48373 492 48397
rect 579 48382 582 48472
rect 612 48454 624 48455
rect 599 48452 649 48454
rect 612 48451 624 48452
rect 610 48444 632 48451
rect 607 48443 632 48444
rect 586 48436 644 48443
rect 607 48435 644 48436
rect 607 48419 610 48435
rect 616 48419 644 48435
rect 607 48418 644 48419
rect 586 48411 644 48418
rect 607 48410 610 48411
rect 612 48403 632 48411
rect 612 48399 624 48403
rect 649 48402 651 48452
rect 544 48365 548 48373
rect 400 48333 408 48363
rect 420 48333 436 48363
rect 400 48329 436 48333
rect 400 48321 430 48329
rect 428 48305 430 48321
rect 476 48293 480 48361
rect 544 48331 552 48365
rect 578 48331 582 48365
rect 544 48323 548 48331
rect 295 48252 300 48286
rect 324 48252 329 48286
rect 378 48283 450 48291
rect 544 48288 548 48293
rect 544 48284 582 48288
rect 544 48269 552 48284
rect 578 48269 582 48284
rect 544 48251 586 48269
rect 522 48245 608 48251
rect 182 48229 224 48245
rect 544 48229 586 48245
rect 17 48215 67 48217
rect 119 48215 169 48217
rect 186 48215 220 48229
rect 548 48215 582 48229
rect 599 48215 649 48217
rect 42 48173 59 48207
rect 67 48165 69 48215
rect 160 48207 246 48215
rect 522 48207 608 48215
rect 76 48173 110 48207
rect 127 48173 144 48207
rect 152 48173 161 48207
rect 162 48205 195 48207
rect 224 48205 244 48207
rect 162 48173 244 48205
rect 524 48205 548 48207
rect 573 48205 582 48207
rect 586 48205 606 48207
rect 160 48165 246 48173
rect 186 48149 220 48165
rect 182 48135 224 48136
rect 160 48129 182 48135
rect 224 48129 246 48135
rect 186 48094 220 48128
rect 223 48094 257 48128
rect 120 48081 170 48083
rect 76 48077 130 48081
rect 110 48072 130 48077
rect 60 48047 67 48057
rect 76 48047 77 48067
rect 96 48038 99 48072
rect 109 48047 110 48067
rect 119 48047 126 48057
rect 76 48031 92 48037
rect 94 48031 110 48037
rect 170 48031 172 48081
rect 186 48015 190 48049
rect 216 48015 220 48049
rect 288 48015 292 48203
rect 476 48135 480 48203
rect 524 48173 606 48205
rect 607 48173 616 48207
rect 522 48165 608 48173
rect 649 48165 651 48215
rect 548 48149 582 48165
rect 522 48130 548 48135
rect 522 48129 582 48130
rect 586 48129 608 48135
rect 295 48094 300 48128
rect 324 48094 329 48128
rect 544 48126 582 48129
rect 378 48089 450 48097
rect 428 48059 430 48075
rect 400 48051 430 48059
rect 476 48057 480 48125
rect 544 48096 552 48126
rect 578 48096 582 48126
rect 544 48087 548 48096
rect 400 48047 436 48051
rect 400 48017 408 48047
rect 420 48017 436 48047
rect 544 48049 548 48057
rect 12 47978 62 47980
rect 28 47969 59 47977
rect 62 47969 64 47978
rect 28 47961 64 47969
rect 127 47969 158 47977
rect 127 47962 182 47969
rect 215 47967 224 47995
rect 127 47961 161 47962
rect 59 47945 64 47961
rect 158 47945 161 47961
rect 28 47937 64 47945
rect 127 47944 161 47945
rect 127 47937 182 47944
rect 62 47928 64 47937
rect 213 47929 224 47967
rect 282 47957 292 48015
rect 296 48009 368 48017
rect 319 47979 346 47990
rect 318 47966 324 47979
rect 346 47966 348 47979
rect 428 47970 430 48017
rect 443 48007 450 48009
rect 476 47977 480 48045
rect 544 48015 552 48049
rect 578 48015 582 48049
rect 481 47983 517 48011
rect 481 47977 495 47983
rect 367 47966 380 47970
rect 251 47923 263 47957
rect 273 47923 293 47957
rect 295 47942 324 47966
rect 303 47932 316 47942
rect 318 47926 324 47942
rect 333 47942 380 47966
rect 333 47932 353 47942
rect 367 47936 380 47942
rect 396 47936 408 47970
rect 420 47936 436 47970
rect 120 47875 170 47877
rect 76 47869 92 47875
rect 94 47869 110 47875
rect 76 47859 99 47868
rect 60 47849 67 47859
rect 76 47839 77 47859
rect 96 47834 99 47859
rect 109 47839 110 47859
rect 119 47849 126 47859
rect 76 47825 110 47829
rect 170 47825 172 47875
rect 186 47857 190 47891
rect 216 47857 220 47891
rect 186 47780 220 47814
rect 282 47811 292 47923
rect 318 47916 335 47926
rect 318 47847 324 47916
rect 346 47847 348 47932
rect 428 47889 430 47936
rect 476 47899 480 47967
rect 485 47949 495 47977
rect 505 47977 519 47983
rect 544 47977 555 48015
rect 505 47949 525 47977
rect 544 47949 553 47977
rect 544 47929 548 47949
rect 579 47908 582 47998
rect 612 47980 624 47981
rect 599 47978 649 47980
rect 612 47977 624 47978
rect 610 47970 632 47977
rect 607 47969 632 47970
rect 586 47962 644 47969
rect 607 47961 644 47962
rect 607 47945 610 47961
rect 616 47945 644 47961
rect 607 47944 644 47945
rect 586 47937 644 47944
rect 607 47936 610 47937
rect 612 47929 632 47937
rect 612 47925 624 47929
rect 649 47928 651 47978
rect 544 47891 548 47899
rect 400 47859 408 47889
rect 420 47859 436 47889
rect 400 47855 436 47859
rect 400 47847 430 47855
rect 428 47831 430 47847
rect 476 47819 480 47887
rect 544 47857 552 47891
rect 578 47857 582 47891
rect 544 47849 548 47857
rect 544 47819 586 47820
rect 288 47779 292 47811
rect 296 47809 368 47817
rect 378 47809 450 47817
rect 544 47812 548 47819
rect 439 47781 444 47809
rect 120 47765 170 47767
rect 76 47761 130 47765
rect 110 47756 130 47761
rect 60 47731 67 47741
rect 76 47731 77 47751
rect 96 47722 99 47756
rect 109 47731 110 47751
rect 119 47731 126 47741
rect 76 47715 92 47721
rect 94 47715 110 47721
rect 170 47715 172 47765
rect 186 47699 190 47733
rect 216 47699 220 47733
rect 213 47667 224 47699
rect 282 47695 292 47779
rect 296 47773 368 47781
rect 378 47773 450 47781
rect 468 47778 473 47812
rect 428 47743 430 47759
rect 251 47667 292 47695
rect 318 47674 324 47743
rect 12 47662 62 47664
rect 28 47653 59 47661
rect 62 47653 64 47662
rect 251 47661 263 47667
rect 28 47645 64 47653
rect 127 47653 158 47661
rect 127 47646 182 47653
rect 127 47645 161 47646
rect 59 47629 64 47645
rect 158 47629 161 47645
rect 253 47633 263 47661
rect 273 47633 293 47667
rect 318 47664 335 47674
rect 303 47648 316 47658
rect 318 47648 324 47664
rect 346 47658 348 47743
rect 400 47735 430 47743
rect 476 47741 480 47809
rect 511 47778 582 47812
rect 544 47771 548 47778
rect 400 47731 436 47735
rect 400 47701 408 47731
rect 420 47701 436 47731
rect 544 47733 548 47741
rect 28 47621 64 47629
rect 127 47628 161 47629
rect 127 47621 182 47628
rect 62 47612 64 47621
rect 282 47575 292 47633
rect 295 47624 324 47648
rect 333 47648 353 47658
rect 428 47654 430 47701
rect 476 47661 480 47729
rect 544 47699 552 47733
rect 578 47699 582 47733
rect 544 47691 548 47699
rect 367 47648 380 47654
rect 333 47624 380 47648
rect 318 47611 324 47624
rect 346 47611 348 47624
rect 367 47620 380 47624
rect 396 47620 408 47654
rect 420 47620 436 47654
rect 544 47651 553 47679
rect 319 47600 346 47611
rect 120 47559 170 47561
rect 76 47553 92 47559
rect 94 47553 110 47559
rect 76 47543 99 47552
rect 60 47533 67 47543
rect 76 47523 77 47543
rect 96 47518 99 47543
rect 109 47523 110 47543
rect 119 47533 126 47543
rect 76 47509 110 47513
rect 170 47509 172 47559
rect 186 47541 190 47575
rect 216 47541 220 47575
rect 182 47503 224 47504
rect 186 47479 220 47496
rect 223 47479 257 47496
rect 182 47462 257 47479
rect 182 47461 224 47462
rect 160 47455 246 47461
rect 288 47455 292 47575
rect 296 47573 368 47581
rect 428 47573 430 47620
rect 476 47583 480 47651
rect 485 47607 495 47641
rect 505 47613 525 47641
rect 505 47607 519 47613
rect 544 47607 555 47651
rect 485 47583 492 47607
rect 579 47592 582 47682
rect 612 47664 624 47665
rect 599 47662 649 47664
rect 612 47661 624 47662
rect 610 47654 632 47661
rect 607 47653 632 47654
rect 586 47646 644 47653
rect 607 47645 644 47646
rect 607 47629 610 47645
rect 616 47629 644 47645
rect 607 47628 644 47629
rect 586 47621 644 47628
rect 607 47620 610 47621
rect 612 47613 632 47621
rect 612 47609 624 47613
rect 649 47612 651 47662
rect 544 47575 548 47583
rect 400 47543 408 47573
rect 420 47543 436 47573
rect 400 47539 436 47543
rect 400 47531 430 47539
rect 428 47515 430 47531
rect 476 47503 480 47571
rect 544 47541 552 47575
rect 578 47541 582 47575
rect 544 47533 548 47541
rect 295 47462 300 47496
rect 324 47462 329 47496
rect 378 47493 450 47501
rect 544 47498 548 47503
rect 544 47494 582 47498
rect 544 47479 552 47494
rect 578 47479 582 47494
rect 544 47461 586 47479
rect 522 47455 608 47461
rect 182 47439 224 47455
rect 544 47439 586 47455
rect 17 47425 67 47427
rect 119 47425 169 47427
rect 186 47425 220 47439
rect 548 47425 582 47439
rect 599 47425 649 47427
rect 42 47383 59 47417
rect 67 47375 69 47425
rect 160 47417 246 47425
rect 522 47417 608 47425
rect 76 47383 110 47417
rect 127 47383 144 47417
rect 152 47383 161 47417
rect 162 47415 195 47417
rect 224 47415 244 47417
rect 162 47383 244 47415
rect 524 47415 548 47417
rect 573 47415 582 47417
rect 586 47415 606 47417
rect 160 47375 246 47383
rect 186 47359 220 47375
rect 182 47345 224 47346
rect 160 47339 182 47345
rect 224 47339 246 47345
rect 186 47304 220 47338
rect 223 47304 257 47338
rect 120 47291 170 47293
rect 76 47287 130 47291
rect 110 47282 130 47287
rect 60 47257 67 47267
rect 76 47257 77 47277
rect 96 47248 99 47282
rect 109 47257 110 47277
rect 119 47257 126 47267
rect 76 47241 92 47247
rect 94 47241 110 47247
rect 170 47241 172 47291
rect 186 47225 190 47259
rect 216 47225 220 47259
rect 288 47225 292 47413
rect 476 47345 480 47413
rect 524 47383 606 47415
rect 607 47383 616 47417
rect 522 47375 608 47383
rect 649 47375 651 47425
rect 548 47359 582 47375
rect 522 47340 548 47345
rect 522 47339 582 47340
rect 586 47339 608 47345
rect 295 47304 300 47338
rect 324 47304 329 47338
rect 544 47336 582 47339
rect 378 47299 450 47307
rect 428 47269 430 47285
rect 400 47261 430 47269
rect 476 47267 480 47335
rect 544 47306 552 47336
rect 578 47306 582 47336
rect 544 47297 548 47306
rect 400 47257 436 47261
rect 400 47227 408 47257
rect 420 47227 436 47257
rect 544 47259 548 47267
rect 12 47188 62 47190
rect 28 47179 59 47187
rect 62 47179 64 47188
rect 28 47171 64 47179
rect 127 47179 158 47187
rect 127 47172 182 47179
rect 215 47177 224 47205
rect 127 47171 161 47172
rect 59 47155 64 47171
rect 158 47155 161 47171
rect 28 47147 64 47155
rect 127 47154 161 47155
rect 127 47147 182 47154
rect 62 47138 64 47147
rect 213 47139 224 47177
rect 282 47167 292 47225
rect 296 47219 368 47227
rect 319 47189 346 47200
rect 318 47176 324 47189
rect 346 47176 348 47189
rect 428 47180 430 47227
rect 443 47217 450 47219
rect 476 47187 480 47255
rect 544 47225 552 47259
rect 578 47225 582 47259
rect 481 47193 517 47221
rect 481 47187 495 47193
rect 367 47176 380 47180
rect 251 47133 263 47167
rect 273 47133 293 47167
rect 295 47152 324 47176
rect 303 47142 316 47152
rect 318 47136 324 47152
rect 333 47152 380 47176
rect 333 47142 353 47152
rect 367 47146 380 47152
rect 396 47146 408 47180
rect 420 47146 436 47180
rect 120 47085 170 47087
rect 76 47079 92 47085
rect 94 47079 110 47085
rect 76 47069 99 47078
rect 60 47059 67 47069
rect 76 47049 77 47069
rect 96 47044 99 47069
rect 109 47049 110 47069
rect 119 47059 126 47069
rect 76 47035 110 47039
rect 170 47035 172 47085
rect 186 47067 190 47101
rect 216 47067 220 47101
rect 186 46990 220 47024
rect 282 47021 292 47133
rect 318 47126 335 47136
rect 318 47057 324 47126
rect 346 47057 348 47142
rect 428 47099 430 47146
rect 476 47109 480 47177
rect 485 47159 495 47187
rect 505 47187 519 47193
rect 544 47187 555 47225
rect 505 47159 525 47187
rect 544 47159 553 47187
rect 544 47139 548 47159
rect 579 47118 582 47208
rect 612 47190 624 47191
rect 599 47188 649 47190
rect 612 47187 624 47188
rect 610 47180 632 47187
rect 607 47179 632 47180
rect 586 47172 644 47179
rect 607 47171 644 47172
rect 607 47155 610 47171
rect 616 47155 644 47171
rect 607 47154 644 47155
rect 586 47147 644 47154
rect 607 47146 610 47147
rect 612 47139 632 47147
rect 612 47135 624 47139
rect 649 47138 651 47188
rect 544 47101 548 47109
rect 400 47069 408 47099
rect 420 47069 436 47099
rect 400 47065 436 47069
rect 400 47057 430 47065
rect 428 47041 430 47057
rect 476 47029 480 47097
rect 544 47067 552 47101
rect 578 47067 582 47101
rect 544 47059 548 47067
rect 544 47029 586 47030
rect 288 46989 292 47021
rect 296 47019 368 47027
rect 378 47019 450 47027
rect 544 47022 548 47029
rect 439 46991 444 47019
rect 120 46975 170 46977
rect 76 46971 130 46975
rect 110 46966 130 46971
rect 60 46941 67 46951
rect 76 46941 77 46961
rect 96 46932 99 46966
rect 109 46941 110 46961
rect 119 46941 126 46951
rect 76 46925 92 46931
rect 94 46925 110 46931
rect 170 46925 172 46975
rect 186 46909 190 46943
rect 216 46909 220 46943
rect 213 46877 224 46909
rect 282 46905 292 46989
rect 296 46983 368 46991
rect 378 46983 450 46991
rect 468 46988 473 47022
rect 428 46953 430 46969
rect 251 46877 292 46905
rect 318 46884 324 46953
rect 12 46872 62 46874
rect 28 46863 59 46871
rect 62 46863 64 46872
rect 251 46871 263 46877
rect 28 46855 64 46863
rect 127 46863 158 46871
rect 127 46856 182 46863
rect 127 46855 161 46856
rect 59 46839 64 46855
rect 158 46839 161 46855
rect 253 46843 263 46871
rect 273 46843 293 46877
rect 318 46874 335 46884
rect 303 46858 316 46868
rect 318 46858 324 46874
rect 346 46868 348 46953
rect 400 46945 430 46953
rect 476 46951 480 47019
rect 511 46988 582 47022
rect 544 46981 548 46988
rect 400 46941 436 46945
rect 400 46911 408 46941
rect 420 46911 436 46941
rect 544 46943 548 46951
rect 28 46831 64 46839
rect 127 46838 161 46839
rect 127 46831 182 46838
rect 62 46822 64 46831
rect 282 46785 292 46843
rect 295 46834 324 46858
rect 333 46858 353 46868
rect 428 46864 430 46911
rect 476 46871 480 46939
rect 544 46909 552 46943
rect 578 46909 582 46943
rect 544 46901 548 46909
rect 367 46858 380 46864
rect 333 46834 380 46858
rect 318 46821 324 46834
rect 346 46821 348 46834
rect 367 46830 380 46834
rect 396 46830 408 46864
rect 420 46830 436 46864
rect 544 46861 553 46889
rect 319 46810 346 46821
rect 120 46769 170 46771
rect 76 46763 92 46769
rect 94 46763 110 46769
rect 76 46753 99 46762
rect 60 46743 67 46753
rect 76 46733 77 46753
rect 96 46728 99 46753
rect 109 46733 110 46753
rect 119 46743 126 46753
rect 76 46719 110 46723
rect 170 46719 172 46769
rect 186 46751 190 46785
rect 216 46751 220 46785
rect 182 46713 224 46714
rect 186 46689 220 46706
rect 223 46689 257 46706
rect 182 46672 257 46689
rect 182 46671 224 46672
rect 160 46665 246 46671
rect 288 46665 292 46785
rect 296 46783 368 46791
rect 428 46783 430 46830
rect 476 46793 480 46861
rect 485 46817 495 46851
rect 505 46823 525 46851
rect 505 46817 519 46823
rect 544 46817 555 46861
rect 485 46793 492 46817
rect 579 46802 582 46892
rect 612 46874 624 46875
rect 599 46872 649 46874
rect 612 46871 624 46872
rect 610 46864 632 46871
rect 607 46863 632 46864
rect 586 46856 644 46863
rect 607 46855 644 46856
rect 607 46839 610 46855
rect 616 46839 644 46855
rect 607 46838 644 46839
rect 586 46831 644 46838
rect 607 46830 610 46831
rect 612 46823 632 46831
rect 612 46819 624 46823
rect 649 46822 651 46872
rect 544 46785 548 46793
rect 400 46753 408 46783
rect 420 46753 436 46783
rect 400 46749 436 46753
rect 400 46741 430 46749
rect 428 46725 430 46741
rect 476 46713 480 46781
rect 544 46751 552 46785
rect 578 46751 582 46785
rect 544 46743 548 46751
rect 295 46672 300 46706
rect 324 46672 329 46706
rect 378 46703 450 46711
rect 544 46708 548 46713
rect 544 46704 582 46708
rect 544 46689 552 46704
rect 578 46689 582 46704
rect 544 46671 586 46689
rect 522 46665 608 46671
rect 182 46649 224 46665
rect 544 46649 586 46665
rect 17 46635 67 46637
rect 119 46635 169 46637
rect 186 46635 220 46649
rect 548 46635 582 46649
rect 599 46635 649 46637
rect 42 46593 59 46627
rect 67 46585 69 46635
rect 160 46627 246 46635
rect 522 46627 608 46635
rect 76 46593 110 46627
rect 127 46593 144 46627
rect 152 46593 161 46627
rect 162 46625 195 46627
rect 224 46625 244 46627
rect 162 46593 244 46625
rect 524 46625 548 46627
rect 573 46625 582 46627
rect 586 46625 606 46627
rect 160 46585 246 46593
rect 186 46569 220 46585
rect 182 46555 224 46556
rect 160 46549 182 46555
rect 224 46549 246 46555
rect 186 46514 220 46548
rect 223 46514 257 46548
rect 120 46501 170 46503
rect 76 46497 130 46501
rect 110 46492 130 46497
rect 60 46467 67 46477
rect 76 46467 77 46487
rect 96 46458 99 46492
rect 109 46467 110 46487
rect 119 46467 126 46477
rect 76 46451 92 46457
rect 94 46451 110 46457
rect 170 46451 172 46501
rect 186 46435 190 46469
rect 216 46435 220 46469
rect 288 46435 292 46623
rect 476 46555 480 46623
rect 524 46593 606 46625
rect 607 46593 616 46627
rect 522 46585 608 46593
rect 649 46585 651 46635
rect 548 46569 582 46585
rect 522 46550 548 46555
rect 522 46549 582 46550
rect 586 46549 608 46555
rect 295 46514 300 46548
rect 324 46514 329 46548
rect 544 46546 582 46549
rect 378 46509 450 46517
rect 428 46479 430 46495
rect 400 46471 430 46479
rect 476 46477 480 46545
rect 544 46516 552 46546
rect 578 46516 582 46546
rect 544 46507 548 46516
rect 400 46467 436 46471
rect 400 46437 408 46467
rect 420 46437 436 46467
rect 544 46469 548 46477
rect 12 46398 62 46400
rect 28 46389 59 46397
rect 62 46389 64 46398
rect 28 46381 64 46389
rect 127 46389 158 46397
rect 127 46382 182 46389
rect 215 46387 224 46415
rect 127 46381 161 46382
rect 59 46365 64 46381
rect 158 46365 161 46381
rect 28 46357 64 46365
rect 127 46364 161 46365
rect 127 46357 182 46364
rect 62 46348 64 46357
rect 213 46349 224 46387
rect 282 46377 292 46435
rect 296 46429 368 46437
rect 319 46399 346 46410
rect 318 46386 324 46399
rect 346 46386 348 46399
rect 428 46390 430 46437
rect 443 46427 450 46429
rect 476 46397 480 46465
rect 544 46435 552 46469
rect 578 46435 582 46469
rect 481 46403 517 46431
rect 481 46397 495 46403
rect 367 46386 380 46390
rect 251 46343 263 46377
rect 273 46343 293 46377
rect 295 46362 324 46386
rect 303 46352 316 46362
rect 318 46346 324 46362
rect 333 46362 380 46386
rect 333 46352 353 46362
rect 367 46356 380 46362
rect 396 46356 408 46390
rect 420 46356 436 46390
rect 120 46295 170 46297
rect 76 46289 92 46295
rect 94 46289 110 46295
rect 76 46279 99 46288
rect 60 46269 67 46279
rect 76 46259 77 46279
rect 96 46254 99 46279
rect 109 46259 110 46279
rect 119 46269 126 46279
rect 76 46245 110 46249
rect 170 46245 172 46295
rect 186 46277 190 46311
rect 216 46277 220 46311
rect 186 46200 220 46234
rect 282 46231 292 46343
rect 318 46336 335 46346
rect 318 46267 324 46336
rect 346 46267 348 46352
rect 428 46309 430 46356
rect 476 46319 480 46387
rect 485 46369 495 46397
rect 505 46397 519 46403
rect 544 46397 555 46435
rect 505 46369 525 46397
rect 544 46369 553 46397
rect 544 46349 548 46369
rect 579 46328 582 46418
rect 612 46400 624 46401
rect 599 46398 649 46400
rect 612 46397 624 46398
rect 610 46390 632 46397
rect 607 46389 632 46390
rect 586 46382 644 46389
rect 607 46381 644 46382
rect 607 46365 610 46381
rect 616 46365 644 46381
rect 607 46364 644 46365
rect 586 46357 644 46364
rect 607 46356 610 46357
rect 612 46349 632 46357
rect 612 46345 624 46349
rect 649 46348 651 46398
rect 544 46311 548 46319
rect 400 46279 408 46309
rect 420 46279 436 46309
rect 400 46275 436 46279
rect 400 46267 430 46275
rect 428 46251 430 46267
rect 476 46239 480 46307
rect 544 46277 552 46311
rect 578 46277 582 46311
rect 544 46269 548 46277
rect 544 46239 586 46240
rect 288 46199 292 46231
rect 296 46229 368 46237
rect 378 46229 450 46237
rect 544 46232 548 46239
rect 439 46201 444 46229
rect 120 46185 170 46187
rect 76 46181 130 46185
rect 110 46176 130 46181
rect 60 46151 67 46161
rect 76 46151 77 46171
rect 96 46142 99 46176
rect 109 46151 110 46171
rect 119 46151 126 46161
rect 76 46135 92 46141
rect 94 46135 110 46141
rect 170 46135 172 46185
rect 186 46119 190 46153
rect 216 46119 220 46153
rect 213 46087 224 46119
rect 282 46115 292 46199
rect 296 46193 368 46201
rect 378 46193 450 46201
rect 468 46198 473 46232
rect 428 46163 430 46179
rect 251 46087 292 46115
rect 318 46094 324 46163
rect 12 46082 62 46084
rect 28 46073 59 46081
rect 62 46073 64 46082
rect 251 46081 263 46087
rect 28 46065 64 46073
rect 127 46073 158 46081
rect 127 46066 182 46073
rect 127 46065 161 46066
rect 59 46049 64 46065
rect 158 46049 161 46065
rect 253 46053 263 46081
rect 273 46053 293 46087
rect 318 46084 335 46094
rect 303 46068 316 46078
rect 318 46068 324 46084
rect 346 46078 348 46163
rect 400 46155 430 46163
rect 476 46161 480 46229
rect 511 46198 582 46232
rect 544 46191 548 46198
rect 400 46151 436 46155
rect 400 46121 408 46151
rect 420 46121 436 46151
rect 544 46153 548 46161
rect 28 46041 64 46049
rect 127 46048 161 46049
rect 127 46041 182 46048
rect 62 46032 64 46041
rect 282 45995 292 46053
rect 295 46044 324 46068
rect 333 46068 353 46078
rect 428 46074 430 46121
rect 476 46081 480 46149
rect 544 46119 552 46153
rect 578 46119 582 46153
rect 544 46111 548 46119
rect 367 46068 380 46074
rect 333 46044 380 46068
rect 318 46031 324 46044
rect 346 46031 348 46044
rect 367 46040 380 46044
rect 396 46040 408 46074
rect 420 46040 436 46074
rect 544 46071 553 46099
rect 319 46020 346 46031
rect 120 45979 170 45981
rect 76 45973 92 45979
rect 94 45973 110 45979
rect 76 45963 99 45972
rect 60 45953 67 45963
rect 76 45943 77 45963
rect 96 45938 99 45963
rect 109 45943 110 45963
rect 119 45953 126 45963
rect 76 45929 110 45933
rect 170 45929 172 45979
rect 186 45961 190 45995
rect 216 45961 220 45995
rect 182 45923 224 45924
rect 186 45899 220 45916
rect 223 45899 257 45916
rect 182 45882 257 45899
rect 182 45881 224 45882
rect 160 45875 246 45881
rect 288 45875 292 45995
rect 296 45993 368 46001
rect 428 45993 430 46040
rect 476 46003 480 46071
rect 485 46027 495 46061
rect 505 46033 525 46061
rect 505 46027 519 46033
rect 544 46027 555 46071
rect 485 46003 492 46027
rect 579 46012 582 46102
rect 612 46084 624 46085
rect 599 46082 649 46084
rect 612 46081 624 46082
rect 610 46074 632 46081
rect 607 46073 632 46074
rect 586 46066 644 46073
rect 607 46065 644 46066
rect 607 46049 610 46065
rect 616 46049 644 46065
rect 607 46048 644 46049
rect 586 46041 644 46048
rect 607 46040 610 46041
rect 612 46033 632 46041
rect 612 46029 624 46033
rect 649 46032 651 46082
rect 544 45995 548 46003
rect 400 45963 408 45993
rect 420 45963 436 45993
rect 400 45959 436 45963
rect 400 45951 430 45959
rect 428 45935 430 45951
rect 476 45923 480 45991
rect 544 45961 552 45995
rect 578 45961 582 45995
rect 544 45953 548 45961
rect 295 45882 300 45916
rect 324 45882 329 45916
rect 378 45913 450 45921
rect 544 45918 548 45923
rect 544 45914 582 45918
rect 544 45899 552 45914
rect 578 45899 582 45914
rect 544 45881 586 45899
rect 522 45875 608 45881
rect 182 45859 224 45875
rect 544 45859 586 45875
rect 17 45845 67 45847
rect 119 45845 169 45847
rect 186 45845 220 45859
rect 548 45845 582 45859
rect 599 45845 649 45847
rect 42 45803 59 45837
rect 67 45795 69 45845
rect 160 45837 246 45845
rect 522 45837 608 45845
rect 76 45803 110 45837
rect 127 45803 144 45837
rect 152 45803 161 45837
rect 162 45835 195 45837
rect 224 45835 244 45837
rect 162 45803 244 45835
rect 524 45835 548 45837
rect 573 45835 582 45837
rect 586 45835 606 45837
rect 160 45795 246 45803
rect 186 45779 220 45795
rect 182 45765 224 45766
rect 160 45759 182 45765
rect 224 45759 246 45765
rect 186 45724 220 45758
rect 223 45724 257 45758
rect 120 45711 170 45713
rect 76 45707 130 45711
rect 110 45702 130 45707
rect 60 45677 67 45687
rect 76 45677 77 45697
rect 96 45668 99 45702
rect 109 45677 110 45697
rect 119 45677 126 45687
rect 76 45661 92 45667
rect 94 45661 110 45667
rect 170 45661 172 45711
rect 186 45645 190 45679
rect 216 45645 220 45679
rect 288 45645 292 45833
rect 476 45765 480 45833
rect 524 45803 606 45835
rect 607 45803 616 45837
rect 522 45795 608 45803
rect 649 45795 651 45845
rect 548 45779 582 45795
rect 522 45760 548 45765
rect 522 45759 582 45760
rect 586 45759 608 45765
rect 295 45724 300 45758
rect 324 45724 329 45758
rect 544 45756 582 45759
rect 378 45719 450 45727
rect 428 45689 430 45705
rect 400 45681 430 45689
rect 476 45687 480 45755
rect 544 45726 552 45756
rect 578 45726 582 45756
rect 544 45717 548 45726
rect 400 45677 436 45681
rect 400 45647 408 45677
rect 420 45647 436 45677
rect 544 45679 548 45687
rect 12 45608 62 45610
rect 28 45599 59 45607
rect 62 45599 64 45608
rect 28 45591 64 45599
rect 127 45599 158 45607
rect 127 45592 182 45599
rect 215 45597 224 45625
rect 127 45591 161 45592
rect 59 45575 64 45591
rect 158 45575 161 45591
rect 28 45567 64 45575
rect 127 45574 161 45575
rect 127 45567 182 45574
rect 62 45558 64 45567
rect 213 45559 224 45597
rect 282 45587 292 45645
rect 296 45639 368 45647
rect 319 45609 346 45620
rect 318 45596 324 45609
rect 346 45596 348 45609
rect 428 45600 430 45647
rect 443 45637 450 45639
rect 476 45607 480 45675
rect 544 45645 552 45679
rect 578 45645 582 45679
rect 481 45613 517 45641
rect 481 45607 495 45613
rect 367 45596 380 45600
rect 251 45553 263 45587
rect 273 45553 293 45587
rect 295 45572 324 45596
rect 303 45562 316 45572
rect 318 45556 324 45572
rect 333 45572 380 45596
rect 333 45562 353 45572
rect 367 45566 380 45572
rect 396 45566 408 45600
rect 420 45566 436 45600
rect 120 45505 170 45507
rect 76 45499 92 45505
rect 94 45499 110 45505
rect 76 45489 99 45498
rect 60 45479 67 45489
rect 76 45469 77 45489
rect 96 45464 99 45489
rect 109 45469 110 45489
rect 119 45479 126 45489
rect 76 45455 110 45459
rect 170 45455 172 45505
rect 186 45487 190 45521
rect 216 45487 220 45521
rect 186 45410 220 45444
rect 282 45441 292 45553
rect 318 45546 335 45556
rect 318 45477 324 45546
rect 346 45477 348 45562
rect 428 45519 430 45566
rect 476 45529 480 45597
rect 485 45579 495 45607
rect 505 45607 519 45613
rect 544 45607 555 45645
rect 505 45579 525 45607
rect 544 45579 553 45607
rect 544 45559 548 45579
rect 579 45538 582 45628
rect 612 45610 624 45611
rect 599 45608 649 45610
rect 612 45607 624 45608
rect 610 45600 632 45607
rect 607 45599 632 45600
rect 586 45592 644 45599
rect 607 45591 644 45592
rect 607 45575 610 45591
rect 616 45575 644 45591
rect 607 45574 644 45575
rect 586 45567 644 45574
rect 607 45566 610 45567
rect 612 45559 632 45567
rect 612 45555 624 45559
rect 649 45558 651 45608
rect 544 45521 548 45529
rect 400 45489 408 45519
rect 420 45489 436 45519
rect 400 45485 436 45489
rect 400 45477 430 45485
rect 428 45461 430 45477
rect 476 45449 480 45517
rect 544 45487 552 45521
rect 578 45487 582 45521
rect 544 45479 548 45487
rect 544 45449 586 45450
rect 288 45409 292 45441
rect 296 45439 368 45447
rect 378 45439 450 45447
rect 544 45442 548 45449
rect 439 45411 444 45439
rect 120 45395 170 45397
rect 76 45391 130 45395
rect 110 45386 130 45391
rect 60 45361 67 45371
rect 76 45361 77 45381
rect 96 45352 99 45386
rect 109 45361 110 45381
rect 119 45361 126 45371
rect 76 45345 92 45351
rect 94 45345 110 45351
rect 170 45345 172 45395
rect 186 45329 190 45363
rect 216 45329 220 45363
rect 213 45297 224 45329
rect 282 45325 292 45409
rect 296 45403 368 45411
rect 378 45403 450 45411
rect 468 45408 473 45442
rect 428 45373 430 45389
rect 251 45297 292 45325
rect 318 45304 324 45373
rect 12 45292 62 45294
rect 28 45283 59 45291
rect 62 45283 64 45292
rect 251 45291 263 45297
rect 28 45275 64 45283
rect 127 45283 158 45291
rect 127 45276 182 45283
rect 127 45275 161 45276
rect 59 45259 64 45275
rect 158 45259 161 45275
rect 253 45263 263 45291
rect 273 45263 293 45297
rect 318 45294 335 45304
rect 303 45278 316 45288
rect 318 45278 324 45294
rect 346 45288 348 45373
rect 400 45365 430 45373
rect 476 45371 480 45439
rect 511 45408 582 45442
rect 544 45401 548 45408
rect 400 45361 436 45365
rect 400 45331 408 45361
rect 420 45331 436 45361
rect 544 45363 548 45371
rect 28 45251 64 45259
rect 127 45258 161 45259
rect 127 45251 182 45258
rect 62 45242 64 45251
rect 282 45205 292 45263
rect 295 45254 324 45278
rect 333 45278 353 45288
rect 428 45284 430 45331
rect 476 45291 480 45359
rect 544 45329 552 45363
rect 578 45329 582 45363
rect 544 45321 548 45329
rect 367 45278 380 45284
rect 333 45254 380 45278
rect 318 45241 324 45254
rect 346 45241 348 45254
rect 367 45250 380 45254
rect 396 45250 408 45284
rect 420 45250 436 45284
rect 544 45281 553 45309
rect 319 45230 346 45241
rect 120 45189 170 45191
rect 76 45183 92 45189
rect 94 45183 110 45189
rect 76 45173 99 45182
rect 60 45163 67 45173
rect 76 45153 77 45173
rect 96 45148 99 45173
rect 109 45153 110 45173
rect 119 45163 126 45173
rect 76 45139 110 45143
rect 170 45139 172 45189
rect 186 45171 190 45205
rect 216 45171 220 45205
rect 182 45133 224 45134
rect 186 45109 220 45126
rect 223 45109 257 45126
rect 182 45092 257 45109
rect 182 45091 224 45092
rect 160 45085 246 45091
rect 288 45085 292 45205
rect 296 45203 368 45211
rect 428 45203 430 45250
rect 476 45213 480 45281
rect 485 45237 495 45271
rect 505 45243 525 45271
rect 505 45237 519 45243
rect 544 45237 555 45281
rect 485 45213 492 45237
rect 579 45222 582 45312
rect 612 45294 624 45295
rect 599 45292 649 45294
rect 612 45291 624 45292
rect 610 45284 632 45291
rect 607 45283 632 45284
rect 586 45276 644 45283
rect 607 45275 644 45276
rect 607 45259 610 45275
rect 616 45259 644 45275
rect 607 45258 644 45259
rect 586 45251 644 45258
rect 607 45250 610 45251
rect 612 45243 632 45251
rect 612 45239 624 45243
rect 649 45242 651 45292
rect 544 45205 548 45213
rect 400 45173 408 45203
rect 420 45173 436 45203
rect 400 45169 436 45173
rect 400 45161 430 45169
rect 428 45145 430 45161
rect 476 45133 480 45201
rect 544 45171 552 45205
rect 578 45171 582 45205
rect 544 45163 548 45171
rect 295 45092 300 45126
rect 324 45092 329 45126
rect 378 45123 450 45131
rect 544 45128 548 45133
rect 544 45124 582 45128
rect 544 45109 552 45124
rect 578 45109 582 45124
rect 544 45091 586 45109
rect 522 45085 608 45091
rect 182 45069 224 45085
rect 544 45069 586 45085
rect 17 45055 67 45057
rect 119 45055 169 45057
rect 186 45055 220 45069
rect 548 45055 582 45069
rect 599 45055 649 45057
rect 42 45013 59 45047
rect 67 45005 69 45055
rect 160 45047 246 45055
rect 522 45047 608 45055
rect 76 45013 110 45047
rect 127 45013 144 45047
rect 152 45013 161 45047
rect 162 45045 195 45047
rect 224 45045 244 45047
rect 162 45013 244 45045
rect 524 45045 548 45047
rect 573 45045 582 45047
rect 586 45045 606 45047
rect 160 45005 246 45013
rect 186 44989 220 45005
rect 182 44975 224 44976
rect 160 44969 182 44975
rect 224 44969 246 44975
rect 186 44934 220 44968
rect 223 44934 257 44968
rect 120 44921 170 44923
rect 76 44917 130 44921
rect 110 44912 130 44917
rect 60 44887 67 44897
rect 76 44887 77 44907
rect 96 44878 99 44912
rect 109 44887 110 44907
rect 119 44887 126 44897
rect 76 44871 92 44877
rect 94 44871 110 44877
rect 170 44871 172 44921
rect 186 44855 190 44889
rect 216 44855 220 44889
rect 288 44855 292 45043
rect 476 44975 480 45043
rect 524 45013 606 45045
rect 607 45013 616 45047
rect 522 45005 608 45013
rect 649 45005 651 45055
rect 548 44989 582 45005
rect 522 44970 548 44975
rect 522 44969 582 44970
rect 586 44969 608 44975
rect 295 44934 300 44968
rect 324 44934 329 44968
rect 544 44966 582 44969
rect 378 44929 450 44937
rect 428 44899 430 44915
rect 400 44891 430 44899
rect 476 44897 480 44965
rect 544 44936 552 44966
rect 578 44936 582 44966
rect 544 44927 548 44936
rect 400 44887 436 44891
rect 400 44857 408 44887
rect 420 44857 436 44887
rect 544 44889 548 44897
rect 12 44818 62 44820
rect 28 44809 59 44817
rect 62 44809 64 44818
rect 28 44801 64 44809
rect 127 44809 158 44817
rect 127 44802 182 44809
rect 215 44807 224 44835
rect 127 44801 161 44802
rect 59 44785 64 44801
rect 158 44785 161 44801
rect 28 44777 64 44785
rect 127 44784 161 44785
rect 127 44777 182 44784
rect 62 44768 64 44777
rect 213 44769 224 44807
rect 282 44797 292 44855
rect 296 44849 368 44857
rect 319 44819 346 44830
rect 318 44806 324 44819
rect 346 44806 348 44819
rect 428 44810 430 44857
rect 443 44847 450 44849
rect 476 44817 480 44885
rect 544 44855 552 44889
rect 578 44855 582 44889
rect 481 44823 517 44851
rect 481 44817 495 44823
rect 367 44806 380 44810
rect 251 44763 263 44797
rect 273 44763 293 44797
rect 295 44782 324 44806
rect 303 44772 316 44782
rect 318 44766 324 44782
rect 333 44782 380 44806
rect 333 44772 353 44782
rect 367 44776 380 44782
rect 396 44776 408 44810
rect 420 44776 436 44810
rect 120 44715 170 44717
rect 76 44709 92 44715
rect 94 44709 110 44715
rect 76 44699 99 44708
rect 60 44689 67 44699
rect 76 44679 77 44699
rect 96 44674 99 44699
rect 109 44679 110 44699
rect 119 44689 126 44699
rect 76 44665 110 44669
rect 170 44665 172 44715
rect 186 44697 190 44731
rect 216 44697 220 44731
rect 186 44620 220 44654
rect 282 44651 292 44763
rect 318 44756 335 44766
rect 318 44687 324 44756
rect 346 44687 348 44772
rect 428 44729 430 44776
rect 476 44739 480 44807
rect 485 44789 495 44817
rect 505 44817 519 44823
rect 544 44817 555 44855
rect 505 44789 525 44817
rect 544 44789 553 44817
rect 544 44769 548 44789
rect 579 44748 582 44838
rect 612 44820 624 44821
rect 599 44818 649 44820
rect 612 44817 624 44818
rect 610 44810 632 44817
rect 607 44809 632 44810
rect 586 44802 644 44809
rect 607 44801 644 44802
rect 607 44785 610 44801
rect 616 44785 644 44801
rect 607 44784 644 44785
rect 586 44777 644 44784
rect 607 44776 610 44777
rect 612 44769 632 44777
rect 612 44765 624 44769
rect 649 44768 651 44818
rect 544 44731 548 44739
rect 400 44699 408 44729
rect 420 44699 436 44729
rect 400 44695 436 44699
rect 400 44687 430 44695
rect 428 44671 430 44687
rect 476 44659 480 44727
rect 544 44697 552 44731
rect 578 44697 582 44731
rect 544 44689 548 44697
rect 544 44659 586 44660
rect 288 44619 292 44651
rect 296 44649 368 44657
rect 378 44649 450 44657
rect 544 44652 548 44659
rect 439 44621 444 44649
rect 120 44605 170 44607
rect 76 44601 130 44605
rect 110 44596 130 44601
rect 60 44571 67 44581
rect 76 44571 77 44591
rect 96 44562 99 44596
rect 109 44571 110 44591
rect 119 44571 126 44581
rect 76 44555 92 44561
rect 94 44555 110 44561
rect 170 44555 172 44605
rect 186 44539 190 44573
rect 216 44539 220 44573
rect 213 44507 224 44539
rect 282 44535 292 44619
rect 296 44613 368 44621
rect 378 44613 450 44621
rect 468 44618 473 44652
rect 428 44583 430 44599
rect 251 44507 292 44535
rect 318 44514 324 44583
rect 12 44502 62 44504
rect 28 44493 59 44501
rect 62 44493 64 44502
rect 251 44501 263 44507
rect 28 44485 64 44493
rect 127 44493 158 44501
rect 127 44486 182 44493
rect 127 44485 161 44486
rect 59 44469 64 44485
rect 158 44469 161 44485
rect 253 44473 263 44501
rect 273 44473 293 44507
rect 318 44504 335 44514
rect 303 44488 316 44498
rect 318 44488 324 44504
rect 346 44498 348 44583
rect 400 44575 430 44583
rect 476 44581 480 44649
rect 511 44618 582 44652
rect 544 44611 548 44618
rect 400 44571 436 44575
rect 400 44541 408 44571
rect 420 44541 436 44571
rect 544 44573 548 44581
rect 28 44461 64 44469
rect 127 44468 161 44469
rect 127 44461 182 44468
rect 62 44452 64 44461
rect 282 44415 292 44473
rect 295 44464 324 44488
rect 333 44488 353 44498
rect 428 44494 430 44541
rect 476 44501 480 44569
rect 544 44539 552 44573
rect 578 44539 582 44573
rect 544 44531 548 44539
rect 367 44488 380 44494
rect 333 44464 380 44488
rect 318 44451 324 44464
rect 346 44451 348 44464
rect 367 44460 380 44464
rect 396 44460 408 44494
rect 420 44460 436 44494
rect 544 44491 553 44519
rect 319 44440 346 44451
rect 120 44399 170 44401
rect 76 44393 92 44399
rect 94 44393 110 44399
rect 76 44383 99 44392
rect 60 44373 67 44383
rect 76 44363 77 44383
rect 96 44358 99 44383
rect 109 44363 110 44383
rect 119 44373 126 44383
rect 76 44349 110 44353
rect 170 44349 172 44399
rect 186 44381 190 44415
rect 216 44381 220 44415
rect 182 44343 224 44344
rect 186 44319 220 44336
rect 223 44319 257 44336
rect 182 44302 257 44319
rect 182 44301 224 44302
rect 160 44295 246 44301
rect 288 44295 292 44415
rect 296 44413 368 44421
rect 428 44413 430 44460
rect 476 44423 480 44491
rect 485 44447 495 44481
rect 505 44453 525 44481
rect 505 44447 519 44453
rect 544 44447 555 44491
rect 485 44423 492 44447
rect 579 44432 582 44522
rect 612 44504 624 44505
rect 599 44502 649 44504
rect 612 44501 624 44502
rect 610 44494 632 44501
rect 607 44493 632 44494
rect 586 44486 644 44493
rect 607 44485 644 44486
rect 607 44469 610 44485
rect 616 44469 644 44485
rect 607 44468 644 44469
rect 586 44461 644 44468
rect 607 44460 610 44461
rect 612 44453 632 44461
rect 612 44449 624 44453
rect 649 44452 651 44502
rect 544 44415 548 44423
rect 400 44383 408 44413
rect 420 44383 436 44413
rect 400 44379 436 44383
rect 400 44371 430 44379
rect 428 44355 430 44371
rect 476 44343 480 44411
rect 544 44381 552 44415
rect 578 44381 582 44415
rect 544 44373 548 44381
rect 295 44302 300 44336
rect 324 44302 329 44336
rect 378 44333 450 44341
rect 544 44338 548 44343
rect 544 44334 582 44338
rect 544 44319 552 44334
rect 578 44319 582 44334
rect 544 44301 586 44319
rect 522 44295 608 44301
rect 182 44279 224 44295
rect 544 44279 586 44295
rect 17 44265 67 44267
rect 119 44265 169 44267
rect 186 44265 220 44279
rect 548 44265 582 44279
rect 599 44265 649 44267
rect 42 44223 59 44257
rect 67 44215 69 44265
rect 160 44257 246 44265
rect 522 44257 608 44265
rect 76 44223 110 44257
rect 127 44223 144 44257
rect 152 44223 161 44257
rect 162 44255 195 44257
rect 224 44255 244 44257
rect 162 44223 244 44255
rect 524 44255 548 44257
rect 573 44255 582 44257
rect 586 44255 606 44257
rect 160 44215 246 44223
rect 186 44199 220 44215
rect 182 44185 224 44186
rect 160 44179 182 44185
rect 224 44179 246 44185
rect 186 44144 220 44178
rect 223 44144 257 44178
rect 120 44131 170 44133
rect 76 44127 130 44131
rect 110 44122 130 44127
rect 60 44097 67 44107
rect 76 44097 77 44117
rect 96 44088 99 44122
rect 109 44097 110 44117
rect 119 44097 126 44107
rect 76 44081 92 44087
rect 94 44081 110 44087
rect 170 44081 172 44131
rect 186 44065 190 44099
rect 216 44065 220 44099
rect 288 44065 292 44253
rect 476 44185 480 44253
rect 524 44223 606 44255
rect 607 44223 616 44257
rect 522 44215 608 44223
rect 649 44215 651 44265
rect 548 44199 582 44215
rect 522 44180 548 44185
rect 522 44179 582 44180
rect 586 44179 608 44185
rect 295 44144 300 44178
rect 324 44144 329 44178
rect 544 44176 582 44179
rect 378 44139 450 44147
rect 428 44109 430 44125
rect 400 44101 430 44109
rect 476 44107 480 44175
rect 544 44146 552 44176
rect 578 44146 582 44176
rect 544 44137 548 44146
rect 400 44097 436 44101
rect 400 44067 408 44097
rect 420 44067 436 44097
rect 544 44099 548 44107
rect 12 44028 62 44030
rect 28 44019 59 44027
rect 62 44019 64 44028
rect 28 44011 64 44019
rect 127 44019 158 44027
rect 127 44012 182 44019
rect 215 44017 224 44045
rect 127 44011 161 44012
rect 59 43995 64 44011
rect 158 43995 161 44011
rect 28 43987 64 43995
rect 127 43994 161 43995
rect 127 43987 182 43994
rect 62 43978 64 43987
rect 213 43979 224 44017
rect 282 44007 292 44065
rect 296 44059 368 44067
rect 319 44029 346 44040
rect 318 44016 324 44029
rect 346 44016 348 44029
rect 428 44020 430 44067
rect 443 44057 450 44059
rect 476 44027 480 44095
rect 544 44065 552 44099
rect 578 44065 582 44099
rect 481 44033 517 44061
rect 481 44027 495 44033
rect 367 44016 380 44020
rect 251 43973 263 44007
rect 273 43973 293 44007
rect 295 43992 324 44016
rect 303 43982 316 43992
rect 318 43976 324 43992
rect 333 43992 380 44016
rect 333 43982 353 43992
rect 367 43986 380 43992
rect 396 43986 408 44020
rect 420 43986 436 44020
rect 120 43925 170 43927
rect 76 43919 92 43925
rect 94 43919 110 43925
rect 76 43909 99 43918
rect 60 43899 67 43909
rect 76 43889 77 43909
rect 96 43884 99 43909
rect 109 43889 110 43909
rect 119 43899 126 43909
rect 76 43875 110 43879
rect 170 43875 172 43925
rect 186 43907 190 43941
rect 216 43907 220 43941
rect 186 43830 220 43864
rect 282 43861 292 43973
rect 318 43966 335 43976
rect 318 43897 324 43966
rect 346 43897 348 43982
rect 428 43939 430 43986
rect 476 43949 480 44017
rect 485 43999 495 44027
rect 505 44027 519 44033
rect 544 44027 555 44065
rect 505 43999 525 44027
rect 544 43999 553 44027
rect 544 43979 548 43999
rect 579 43958 582 44048
rect 612 44030 624 44031
rect 599 44028 649 44030
rect 612 44027 624 44028
rect 610 44020 632 44027
rect 607 44019 632 44020
rect 586 44012 644 44019
rect 607 44011 644 44012
rect 607 43995 610 44011
rect 616 43995 644 44011
rect 607 43994 644 43995
rect 586 43987 644 43994
rect 607 43986 610 43987
rect 612 43979 632 43987
rect 612 43975 624 43979
rect 649 43978 651 44028
rect 544 43941 548 43949
rect 400 43909 408 43939
rect 420 43909 436 43939
rect 400 43905 436 43909
rect 400 43897 430 43905
rect 428 43881 430 43897
rect 476 43869 480 43937
rect 544 43907 552 43941
rect 578 43907 582 43941
rect 544 43899 548 43907
rect 544 43869 586 43870
rect 288 43829 292 43861
rect 296 43859 368 43867
rect 378 43859 450 43867
rect 544 43862 548 43869
rect 439 43831 444 43859
rect 120 43815 170 43817
rect 76 43811 130 43815
rect 110 43806 130 43811
rect 60 43781 67 43791
rect 76 43781 77 43801
rect 96 43772 99 43806
rect 109 43781 110 43801
rect 119 43781 126 43791
rect 76 43765 92 43771
rect 94 43765 110 43771
rect 170 43765 172 43815
rect 186 43749 190 43783
rect 216 43749 220 43783
rect 213 43717 224 43749
rect 282 43745 292 43829
rect 296 43823 368 43831
rect 378 43823 450 43831
rect 468 43828 473 43862
rect 428 43793 430 43809
rect 251 43717 292 43745
rect 318 43724 324 43793
rect 12 43712 62 43714
rect 28 43703 59 43711
rect 62 43703 64 43712
rect 251 43711 263 43717
rect 28 43695 64 43703
rect 127 43703 158 43711
rect 127 43696 182 43703
rect 127 43695 161 43696
rect 59 43679 64 43695
rect 158 43679 161 43695
rect 253 43683 263 43711
rect 273 43683 293 43717
rect 318 43714 335 43724
rect 303 43698 316 43708
rect 318 43698 324 43714
rect 346 43708 348 43793
rect 400 43785 430 43793
rect 476 43791 480 43859
rect 511 43828 582 43862
rect 544 43821 548 43828
rect 400 43781 436 43785
rect 400 43751 408 43781
rect 420 43751 436 43781
rect 544 43783 548 43791
rect 28 43671 64 43679
rect 127 43678 161 43679
rect 127 43671 182 43678
rect 62 43662 64 43671
rect 282 43625 292 43683
rect 295 43674 324 43698
rect 333 43698 353 43708
rect 428 43704 430 43751
rect 476 43711 480 43779
rect 544 43749 552 43783
rect 578 43749 582 43783
rect 544 43741 548 43749
rect 367 43698 380 43704
rect 333 43674 380 43698
rect 318 43661 324 43674
rect 346 43661 348 43674
rect 367 43670 380 43674
rect 396 43670 408 43704
rect 420 43670 436 43704
rect 544 43701 553 43729
rect 319 43650 346 43661
rect 120 43609 170 43611
rect 76 43603 92 43609
rect 94 43603 110 43609
rect 76 43593 99 43602
rect 60 43583 67 43593
rect 76 43573 77 43593
rect 96 43568 99 43593
rect 109 43573 110 43593
rect 119 43583 126 43593
rect 76 43559 110 43563
rect 170 43559 172 43609
rect 186 43591 190 43625
rect 216 43591 220 43625
rect 182 43553 224 43554
rect 186 43529 220 43546
rect 223 43529 257 43546
rect 182 43512 257 43529
rect 182 43511 224 43512
rect 160 43505 246 43511
rect 288 43505 292 43625
rect 296 43623 368 43631
rect 428 43623 430 43670
rect 476 43633 480 43701
rect 485 43657 495 43691
rect 505 43663 525 43691
rect 505 43657 519 43663
rect 544 43657 555 43701
rect 485 43633 492 43657
rect 579 43642 582 43732
rect 612 43714 624 43715
rect 599 43712 649 43714
rect 612 43711 624 43712
rect 610 43704 632 43711
rect 607 43703 632 43704
rect 586 43696 644 43703
rect 607 43695 644 43696
rect 607 43679 610 43695
rect 616 43679 644 43695
rect 607 43678 644 43679
rect 586 43671 644 43678
rect 607 43670 610 43671
rect 612 43663 632 43671
rect 612 43659 624 43663
rect 649 43662 651 43712
rect 544 43625 548 43633
rect 400 43593 408 43623
rect 420 43593 436 43623
rect 400 43589 436 43593
rect 400 43581 430 43589
rect 428 43565 430 43581
rect 476 43553 480 43621
rect 544 43591 552 43625
rect 578 43591 582 43625
rect 544 43583 548 43591
rect 295 43512 300 43546
rect 324 43512 329 43546
rect 378 43543 450 43551
rect 544 43548 548 43553
rect 544 43544 582 43548
rect 544 43529 552 43544
rect 578 43529 582 43544
rect 544 43511 586 43529
rect 522 43505 608 43511
rect 182 43489 224 43505
rect 544 43489 586 43505
rect 17 43475 67 43477
rect 119 43475 169 43477
rect 186 43475 220 43489
rect 548 43475 582 43489
rect 599 43475 649 43477
rect 42 43433 59 43467
rect 67 43425 69 43475
rect 160 43467 246 43475
rect 522 43467 608 43475
rect 76 43433 110 43467
rect 127 43433 144 43467
rect 152 43433 161 43467
rect 162 43465 195 43467
rect 224 43465 244 43467
rect 162 43433 244 43465
rect 524 43465 548 43467
rect 573 43465 582 43467
rect 586 43465 606 43467
rect 160 43425 246 43433
rect 186 43409 220 43425
rect 182 43395 224 43396
rect 160 43389 182 43395
rect 224 43389 246 43395
rect 186 43354 220 43388
rect 223 43354 257 43388
rect 120 43341 170 43343
rect 76 43337 130 43341
rect 110 43332 130 43337
rect 60 43307 67 43317
rect 76 43307 77 43327
rect 96 43298 99 43332
rect 109 43307 110 43327
rect 119 43307 126 43317
rect 76 43291 92 43297
rect 94 43291 110 43297
rect 170 43291 172 43341
rect 186 43275 190 43309
rect 216 43275 220 43309
rect 288 43275 292 43463
rect 476 43395 480 43463
rect 524 43433 606 43465
rect 607 43433 616 43467
rect 522 43425 608 43433
rect 649 43425 651 43475
rect 548 43409 582 43425
rect 522 43390 548 43395
rect 522 43389 582 43390
rect 586 43389 608 43395
rect 295 43354 300 43388
rect 324 43354 329 43388
rect 544 43386 582 43389
rect 378 43349 450 43357
rect 428 43319 430 43335
rect 400 43311 430 43319
rect 476 43317 480 43385
rect 544 43356 552 43386
rect 578 43356 582 43386
rect 544 43347 548 43356
rect 400 43307 436 43311
rect 400 43277 408 43307
rect 420 43277 436 43307
rect 544 43309 548 43317
rect 12 43238 62 43240
rect 28 43229 59 43237
rect 62 43229 64 43238
rect 28 43221 64 43229
rect 127 43229 158 43237
rect 127 43222 182 43229
rect 215 43227 224 43255
rect 127 43221 161 43222
rect 59 43205 64 43221
rect 158 43205 161 43221
rect 28 43197 64 43205
rect 127 43204 161 43205
rect 127 43197 182 43204
rect 62 43188 64 43197
rect 213 43189 224 43227
rect 282 43217 292 43275
rect 296 43269 368 43277
rect 319 43239 346 43250
rect 318 43226 324 43239
rect 346 43226 348 43239
rect 428 43230 430 43277
rect 443 43267 450 43269
rect 476 43237 480 43305
rect 544 43275 552 43309
rect 578 43275 582 43309
rect 481 43243 517 43271
rect 481 43237 495 43243
rect 367 43226 380 43230
rect 251 43183 263 43217
rect 273 43183 293 43217
rect 295 43202 324 43226
rect 303 43192 316 43202
rect 318 43186 324 43202
rect 333 43202 380 43226
rect 333 43192 353 43202
rect 367 43196 380 43202
rect 396 43196 408 43230
rect 420 43196 436 43230
rect 120 43135 170 43137
rect 76 43129 92 43135
rect 94 43129 110 43135
rect 76 43119 99 43128
rect 60 43109 67 43119
rect 76 43099 77 43119
rect 96 43094 99 43119
rect 109 43099 110 43119
rect 119 43109 126 43119
rect 76 43085 110 43089
rect 170 43085 172 43135
rect 186 43117 190 43151
rect 216 43117 220 43151
rect 186 43040 220 43074
rect 282 43071 292 43183
rect 318 43176 335 43186
rect 318 43107 324 43176
rect 346 43107 348 43192
rect 428 43149 430 43196
rect 476 43159 480 43227
rect 485 43209 495 43237
rect 505 43237 519 43243
rect 544 43237 555 43275
rect 505 43209 525 43237
rect 544 43209 553 43237
rect 544 43189 548 43209
rect 579 43168 582 43258
rect 612 43240 624 43241
rect 599 43238 649 43240
rect 612 43237 624 43238
rect 610 43230 632 43237
rect 607 43229 632 43230
rect 586 43222 644 43229
rect 607 43221 644 43222
rect 607 43205 610 43221
rect 616 43205 644 43221
rect 607 43204 644 43205
rect 586 43197 644 43204
rect 607 43196 610 43197
rect 612 43189 632 43197
rect 612 43185 624 43189
rect 649 43188 651 43238
rect 544 43151 548 43159
rect 400 43119 408 43149
rect 420 43119 436 43149
rect 400 43115 436 43119
rect 400 43107 430 43115
rect 428 43091 430 43107
rect 476 43079 480 43147
rect 544 43117 552 43151
rect 578 43117 582 43151
rect 544 43109 548 43117
rect 544 43079 586 43080
rect 288 43039 292 43071
rect 296 43069 368 43077
rect 378 43069 450 43077
rect 544 43072 548 43079
rect 439 43041 444 43069
rect 120 43025 170 43027
rect 76 43021 130 43025
rect 110 43016 130 43021
rect 60 42991 67 43001
rect 76 42991 77 43011
rect 96 42982 99 43016
rect 109 42991 110 43011
rect 119 42991 126 43001
rect 76 42975 92 42981
rect 94 42975 110 42981
rect 170 42975 172 43025
rect 186 42959 190 42993
rect 216 42959 220 42993
rect 213 42927 224 42959
rect 282 42955 292 43039
rect 296 43033 368 43041
rect 378 43033 450 43041
rect 468 43038 473 43072
rect 428 43003 430 43019
rect 251 42927 292 42955
rect 318 42934 324 43003
rect 12 42922 62 42924
rect 28 42913 59 42921
rect 62 42913 64 42922
rect 251 42921 263 42927
rect 28 42905 64 42913
rect 127 42913 158 42921
rect 127 42906 182 42913
rect 127 42905 161 42906
rect 59 42889 64 42905
rect 158 42889 161 42905
rect 253 42893 263 42921
rect 273 42893 293 42927
rect 318 42924 335 42934
rect 303 42908 316 42918
rect 318 42908 324 42924
rect 346 42918 348 43003
rect 400 42995 430 43003
rect 476 43001 480 43069
rect 511 43038 582 43072
rect 544 43031 548 43038
rect 400 42991 436 42995
rect 400 42961 408 42991
rect 420 42961 436 42991
rect 544 42993 548 43001
rect 28 42881 64 42889
rect 127 42888 161 42889
rect 127 42881 182 42888
rect 62 42872 64 42881
rect 282 42835 292 42893
rect 295 42884 324 42908
rect 333 42908 353 42918
rect 428 42914 430 42961
rect 476 42921 480 42989
rect 544 42959 552 42993
rect 578 42959 582 42993
rect 544 42951 548 42959
rect 367 42908 380 42914
rect 333 42884 380 42908
rect 318 42871 324 42884
rect 346 42871 348 42884
rect 367 42880 380 42884
rect 396 42880 408 42914
rect 420 42880 436 42914
rect 544 42911 553 42939
rect 319 42860 346 42871
rect 120 42819 170 42821
rect 76 42813 92 42819
rect 94 42813 110 42819
rect 76 42803 99 42812
rect 60 42793 67 42803
rect 76 42783 77 42803
rect 96 42778 99 42803
rect 109 42783 110 42803
rect 119 42793 126 42803
rect 76 42769 110 42773
rect 170 42769 172 42819
rect 186 42801 190 42835
rect 216 42801 220 42835
rect 182 42763 224 42764
rect 186 42739 220 42756
rect 223 42739 257 42756
rect 182 42722 257 42739
rect 182 42721 224 42722
rect 160 42715 246 42721
rect 288 42715 292 42835
rect 296 42833 368 42841
rect 428 42833 430 42880
rect 476 42843 480 42911
rect 485 42867 495 42901
rect 505 42873 525 42901
rect 505 42867 519 42873
rect 544 42867 555 42911
rect 485 42843 492 42867
rect 579 42852 582 42942
rect 612 42924 624 42925
rect 599 42922 649 42924
rect 612 42921 624 42922
rect 610 42914 632 42921
rect 607 42913 632 42914
rect 586 42906 644 42913
rect 607 42905 644 42906
rect 607 42889 610 42905
rect 616 42889 644 42905
rect 607 42888 644 42889
rect 586 42881 644 42888
rect 607 42880 610 42881
rect 612 42873 632 42881
rect 612 42869 624 42873
rect 649 42872 651 42922
rect 544 42835 548 42843
rect 400 42803 408 42833
rect 420 42803 436 42833
rect 400 42799 436 42803
rect 400 42791 430 42799
rect 428 42775 430 42791
rect 476 42763 480 42831
rect 544 42801 552 42835
rect 578 42801 582 42835
rect 544 42793 548 42801
rect 295 42722 300 42756
rect 324 42722 329 42756
rect 378 42753 450 42761
rect 544 42758 548 42763
rect 544 42754 582 42758
rect 544 42739 552 42754
rect 578 42739 582 42754
rect 544 42721 586 42739
rect 522 42715 608 42721
rect 182 42699 224 42715
rect 544 42699 586 42715
rect 17 42685 67 42687
rect 119 42685 169 42687
rect 186 42685 220 42699
rect 548 42685 582 42699
rect 599 42685 649 42687
rect 42 42643 59 42677
rect 67 42635 69 42685
rect 160 42677 246 42685
rect 522 42677 608 42685
rect 76 42643 110 42677
rect 127 42643 144 42677
rect 152 42643 161 42677
rect 162 42675 195 42677
rect 224 42675 244 42677
rect 162 42643 244 42675
rect 524 42675 548 42677
rect 573 42675 582 42677
rect 586 42675 606 42677
rect 160 42635 246 42643
rect 186 42619 220 42635
rect 182 42605 224 42606
rect 160 42599 182 42605
rect 224 42599 246 42605
rect 186 42564 220 42598
rect 223 42564 257 42598
rect 120 42551 170 42553
rect 76 42547 130 42551
rect 110 42542 130 42547
rect 60 42517 67 42527
rect 76 42517 77 42537
rect 96 42508 99 42542
rect 109 42517 110 42537
rect 119 42517 126 42527
rect 76 42501 92 42507
rect 94 42501 110 42507
rect 170 42501 172 42551
rect 186 42485 190 42519
rect 216 42485 220 42519
rect 288 42485 292 42673
rect 476 42605 480 42673
rect 524 42643 606 42675
rect 607 42643 616 42677
rect 522 42635 608 42643
rect 649 42635 651 42685
rect 548 42619 582 42635
rect 522 42600 548 42605
rect 522 42599 582 42600
rect 586 42599 608 42605
rect 295 42564 300 42598
rect 324 42564 329 42598
rect 544 42596 582 42599
rect 378 42559 450 42567
rect 428 42529 430 42545
rect 400 42521 430 42529
rect 476 42527 480 42595
rect 544 42566 552 42596
rect 578 42566 582 42596
rect 544 42557 548 42566
rect 400 42517 436 42521
rect 400 42487 408 42517
rect 420 42487 436 42517
rect 544 42519 548 42527
rect 12 42448 62 42450
rect 28 42439 59 42447
rect 62 42439 64 42448
rect 28 42431 64 42439
rect 127 42439 158 42447
rect 127 42432 182 42439
rect 215 42437 224 42465
rect 127 42431 161 42432
rect 59 42415 64 42431
rect 158 42415 161 42431
rect 28 42407 64 42415
rect 127 42414 161 42415
rect 127 42407 182 42414
rect 62 42398 64 42407
rect 213 42399 224 42437
rect 282 42427 292 42485
rect 296 42479 368 42487
rect 319 42449 346 42460
rect 318 42436 324 42449
rect 346 42436 348 42449
rect 428 42440 430 42487
rect 443 42477 450 42479
rect 476 42447 480 42515
rect 544 42485 552 42519
rect 578 42485 582 42519
rect 481 42453 517 42481
rect 481 42447 495 42453
rect 367 42436 380 42440
rect 251 42393 263 42427
rect 273 42393 293 42427
rect 295 42412 324 42436
rect 303 42402 316 42412
rect 318 42396 324 42412
rect 333 42412 380 42436
rect 333 42402 353 42412
rect 367 42406 380 42412
rect 396 42406 408 42440
rect 420 42406 436 42440
rect 120 42345 170 42347
rect 76 42339 92 42345
rect 94 42339 110 42345
rect 76 42329 99 42338
rect 60 42319 67 42329
rect 76 42309 77 42329
rect 96 42304 99 42329
rect 109 42309 110 42329
rect 119 42319 126 42329
rect 76 42295 110 42299
rect 170 42295 172 42345
rect 186 42327 190 42361
rect 216 42327 220 42361
rect 186 42250 220 42284
rect 282 42281 292 42393
rect 318 42386 335 42396
rect 318 42317 324 42386
rect 346 42317 348 42402
rect 428 42359 430 42406
rect 476 42369 480 42437
rect 485 42419 495 42447
rect 505 42447 519 42453
rect 544 42447 555 42485
rect 505 42419 525 42447
rect 544 42419 553 42447
rect 544 42399 548 42419
rect 579 42378 582 42468
rect 612 42450 624 42451
rect 599 42448 649 42450
rect 612 42447 624 42448
rect 610 42440 632 42447
rect 607 42439 632 42440
rect 586 42432 644 42439
rect 607 42431 644 42432
rect 607 42415 610 42431
rect 616 42415 644 42431
rect 607 42414 644 42415
rect 586 42407 644 42414
rect 607 42406 610 42407
rect 612 42399 632 42407
rect 612 42395 624 42399
rect 649 42398 651 42448
rect 544 42361 548 42369
rect 400 42329 408 42359
rect 420 42329 436 42359
rect 400 42325 436 42329
rect 400 42317 430 42325
rect 428 42301 430 42317
rect 476 42289 480 42357
rect 544 42327 552 42361
rect 578 42327 582 42361
rect 544 42319 548 42327
rect 544 42289 586 42290
rect 288 42249 292 42281
rect 296 42279 368 42287
rect 378 42279 450 42287
rect 544 42282 548 42289
rect 439 42251 444 42279
rect 120 42235 170 42237
rect 76 42231 130 42235
rect 110 42226 130 42231
rect 60 42201 67 42211
rect 76 42201 77 42221
rect 96 42192 99 42226
rect 109 42201 110 42221
rect 119 42201 126 42211
rect 76 42185 92 42191
rect 94 42185 110 42191
rect 170 42185 172 42235
rect 186 42169 190 42203
rect 216 42169 220 42203
rect 213 42137 224 42169
rect 282 42165 292 42249
rect 296 42243 368 42251
rect 378 42243 450 42251
rect 468 42248 473 42282
rect 428 42213 430 42229
rect 251 42137 292 42165
rect 318 42144 324 42213
rect 12 42132 62 42134
rect 28 42123 59 42131
rect 62 42123 64 42132
rect 251 42131 263 42137
rect 28 42115 64 42123
rect 127 42123 158 42131
rect 127 42116 182 42123
rect 127 42115 161 42116
rect 59 42099 64 42115
rect 158 42099 161 42115
rect 253 42103 263 42131
rect 273 42103 293 42137
rect 318 42134 335 42144
rect 303 42118 316 42128
rect 318 42118 324 42134
rect 346 42128 348 42213
rect 400 42205 430 42213
rect 476 42211 480 42279
rect 511 42248 582 42282
rect 544 42241 548 42248
rect 400 42201 436 42205
rect 400 42171 408 42201
rect 420 42171 436 42201
rect 544 42203 548 42211
rect 28 42091 64 42099
rect 127 42098 161 42099
rect 127 42091 182 42098
rect 62 42082 64 42091
rect 282 42045 292 42103
rect 295 42094 324 42118
rect 333 42118 353 42128
rect 428 42124 430 42171
rect 476 42131 480 42199
rect 544 42169 552 42203
rect 578 42169 582 42203
rect 544 42161 548 42169
rect 367 42118 380 42124
rect 333 42094 380 42118
rect 318 42081 324 42094
rect 346 42081 348 42094
rect 367 42090 380 42094
rect 396 42090 408 42124
rect 420 42090 436 42124
rect 544 42121 553 42149
rect 319 42070 346 42081
rect 120 42029 170 42031
rect 76 42023 92 42029
rect 94 42023 110 42029
rect 76 42013 99 42022
rect 60 42003 67 42013
rect 76 41993 77 42013
rect 96 41988 99 42013
rect 109 41993 110 42013
rect 119 42003 126 42013
rect 76 41979 110 41983
rect 170 41979 172 42029
rect 186 42011 190 42045
rect 216 42011 220 42045
rect 182 41973 224 41974
rect 186 41949 220 41966
rect 223 41949 257 41966
rect 182 41932 257 41949
rect 182 41931 224 41932
rect 160 41925 246 41931
rect 288 41925 292 42045
rect 296 42043 368 42051
rect 428 42043 430 42090
rect 476 42053 480 42121
rect 485 42077 495 42111
rect 505 42083 525 42111
rect 505 42077 519 42083
rect 544 42077 555 42121
rect 485 42053 492 42077
rect 579 42062 582 42152
rect 612 42134 624 42135
rect 599 42132 649 42134
rect 612 42131 624 42132
rect 610 42124 632 42131
rect 607 42123 632 42124
rect 586 42116 644 42123
rect 607 42115 644 42116
rect 607 42099 610 42115
rect 616 42099 644 42115
rect 607 42098 644 42099
rect 586 42091 644 42098
rect 607 42090 610 42091
rect 612 42083 632 42091
rect 612 42079 624 42083
rect 649 42082 651 42132
rect 544 42045 548 42053
rect 400 42013 408 42043
rect 420 42013 436 42043
rect 400 42009 436 42013
rect 400 42001 430 42009
rect 428 41985 430 42001
rect 476 41973 480 42041
rect 544 42011 552 42045
rect 578 42011 582 42045
rect 544 42003 548 42011
rect 295 41932 300 41966
rect 324 41932 329 41966
rect 378 41963 450 41971
rect 544 41968 548 41973
rect 544 41964 582 41968
rect 544 41949 552 41964
rect 578 41949 582 41964
rect 544 41931 586 41949
rect 522 41925 608 41931
rect 182 41909 224 41925
rect 544 41909 586 41925
rect 17 41895 67 41897
rect 119 41895 169 41897
rect 186 41895 220 41909
rect 548 41895 582 41909
rect 599 41895 649 41897
rect 42 41853 59 41887
rect 67 41845 69 41895
rect 160 41887 246 41895
rect 522 41887 608 41895
rect 76 41853 110 41887
rect 127 41853 144 41887
rect 152 41853 161 41887
rect 162 41885 195 41887
rect 224 41885 244 41887
rect 162 41853 244 41885
rect 524 41885 548 41887
rect 573 41885 582 41887
rect 586 41885 606 41887
rect 160 41845 246 41853
rect 186 41829 220 41845
rect 182 41815 224 41816
rect 160 41809 182 41815
rect 224 41809 246 41815
rect 186 41774 220 41808
rect 223 41774 257 41808
rect 120 41761 170 41763
rect 76 41757 130 41761
rect 110 41752 130 41757
rect 60 41727 67 41737
rect 76 41727 77 41747
rect 96 41718 99 41752
rect 109 41727 110 41747
rect 119 41727 126 41737
rect 76 41711 92 41717
rect 94 41711 110 41717
rect 170 41711 172 41761
rect 186 41695 190 41729
rect 216 41695 220 41729
rect 288 41695 292 41883
rect 476 41815 480 41883
rect 524 41853 606 41885
rect 607 41853 616 41887
rect 522 41845 608 41853
rect 649 41845 651 41895
rect 548 41829 582 41845
rect 522 41810 548 41815
rect 522 41809 582 41810
rect 586 41809 608 41815
rect 295 41774 300 41808
rect 324 41774 329 41808
rect 544 41806 582 41809
rect 378 41769 450 41777
rect 428 41739 430 41755
rect 400 41731 430 41739
rect 476 41737 480 41805
rect 544 41776 552 41806
rect 578 41776 582 41806
rect 544 41767 548 41776
rect 400 41727 436 41731
rect 400 41697 408 41727
rect 420 41697 436 41727
rect 544 41729 548 41737
rect 12 41658 62 41660
rect 28 41649 59 41657
rect 62 41649 64 41658
rect 28 41641 64 41649
rect 127 41649 158 41657
rect 127 41642 182 41649
rect 215 41647 224 41675
rect 127 41641 161 41642
rect 59 41625 64 41641
rect 158 41625 161 41641
rect 28 41617 64 41625
rect 127 41624 161 41625
rect 127 41617 182 41624
rect 62 41608 64 41617
rect 213 41609 224 41647
rect 282 41637 292 41695
rect 296 41689 368 41697
rect 319 41659 346 41670
rect 318 41646 324 41659
rect 346 41646 348 41659
rect 428 41650 430 41697
rect 443 41687 450 41689
rect 476 41657 480 41725
rect 544 41695 552 41729
rect 578 41695 582 41729
rect 481 41663 517 41691
rect 481 41657 495 41663
rect 367 41646 380 41650
rect 251 41603 263 41637
rect 273 41603 293 41637
rect 295 41622 324 41646
rect 303 41612 316 41622
rect 318 41606 324 41622
rect 333 41622 380 41646
rect 333 41612 353 41622
rect 367 41616 380 41622
rect 396 41616 408 41650
rect 420 41616 436 41650
rect 120 41555 170 41557
rect 76 41549 92 41555
rect 94 41549 110 41555
rect 76 41539 99 41548
rect 60 41529 67 41539
rect 76 41519 77 41539
rect 96 41514 99 41539
rect 109 41519 110 41539
rect 119 41529 126 41539
rect 76 41505 110 41509
rect 170 41505 172 41555
rect 186 41537 190 41571
rect 216 41537 220 41571
rect 186 41460 220 41494
rect 282 41491 292 41603
rect 318 41596 335 41606
rect 318 41527 324 41596
rect 346 41527 348 41612
rect 428 41569 430 41616
rect 476 41579 480 41647
rect 485 41629 495 41657
rect 505 41657 519 41663
rect 544 41657 555 41695
rect 505 41629 525 41657
rect 544 41629 553 41657
rect 544 41609 548 41629
rect 579 41588 582 41678
rect 612 41660 624 41661
rect 599 41658 649 41660
rect 612 41657 624 41658
rect 610 41650 632 41657
rect 607 41649 632 41650
rect 586 41642 644 41649
rect 607 41641 644 41642
rect 607 41625 610 41641
rect 616 41625 644 41641
rect 607 41624 644 41625
rect 586 41617 644 41624
rect 607 41616 610 41617
rect 612 41609 632 41617
rect 612 41605 624 41609
rect 649 41608 651 41658
rect 544 41571 548 41579
rect 400 41539 408 41569
rect 420 41539 436 41569
rect 400 41535 436 41539
rect 400 41527 430 41535
rect 428 41511 430 41527
rect 476 41499 480 41567
rect 544 41537 552 41571
rect 578 41537 582 41571
rect 544 41529 548 41537
rect 544 41499 586 41500
rect 288 41459 292 41491
rect 296 41489 368 41497
rect 378 41489 450 41497
rect 544 41492 548 41499
rect 439 41461 444 41489
rect 120 41445 170 41447
rect 76 41441 130 41445
rect 110 41436 130 41441
rect 60 41411 67 41421
rect 76 41411 77 41431
rect 96 41402 99 41436
rect 109 41411 110 41431
rect 119 41411 126 41421
rect 76 41395 92 41401
rect 94 41395 110 41401
rect 170 41395 172 41445
rect 186 41379 190 41413
rect 216 41379 220 41413
rect 213 41347 224 41379
rect 282 41375 292 41459
rect 296 41453 368 41461
rect 378 41453 450 41461
rect 468 41458 473 41492
rect 428 41423 430 41439
rect 251 41347 292 41375
rect 318 41354 324 41423
rect 12 41342 62 41344
rect 28 41333 59 41341
rect 62 41333 64 41342
rect 251 41341 263 41347
rect 28 41325 64 41333
rect 127 41333 158 41341
rect 127 41326 182 41333
rect 127 41325 161 41326
rect 59 41309 64 41325
rect 158 41309 161 41325
rect 253 41313 263 41341
rect 273 41313 293 41347
rect 318 41344 335 41354
rect 303 41328 316 41338
rect 318 41328 324 41344
rect 346 41338 348 41423
rect 400 41415 430 41423
rect 476 41421 480 41489
rect 511 41458 582 41492
rect 544 41451 548 41458
rect 400 41411 436 41415
rect 400 41381 408 41411
rect 420 41381 436 41411
rect 544 41413 548 41421
rect 28 41301 64 41309
rect 127 41308 161 41309
rect 127 41301 182 41308
rect 62 41292 64 41301
rect 282 41255 292 41313
rect 295 41304 324 41328
rect 333 41328 353 41338
rect 428 41334 430 41381
rect 476 41341 480 41409
rect 544 41379 552 41413
rect 578 41379 582 41413
rect 544 41371 548 41379
rect 367 41328 380 41334
rect 333 41304 380 41328
rect 318 41291 324 41304
rect 346 41291 348 41304
rect 367 41300 380 41304
rect 396 41300 408 41334
rect 420 41300 436 41334
rect 544 41331 553 41359
rect 319 41280 346 41291
rect 120 41239 170 41241
rect 76 41233 92 41239
rect 94 41233 110 41239
rect 76 41223 99 41232
rect 60 41213 67 41223
rect 76 41203 77 41223
rect 96 41198 99 41223
rect 109 41203 110 41223
rect 119 41213 126 41223
rect 76 41189 110 41193
rect 170 41189 172 41239
rect 186 41221 190 41255
rect 216 41221 220 41255
rect 182 41183 224 41184
rect 186 41159 220 41176
rect 223 41159 257 41176
rect 182 41142 257 41159
rect 182 41141 224 41142
rect 160 41135 246 41141
rect 288 41135 292 41255
rect 296 41253 368 41261
rect 428 41253 430 41300
rect 476 41263 480 41331
rect 485 41287 495 41321
rect 505 41293 525 41321
rect 505 41287 519 41293
rect 544 41287 555 41331
rect 485 41263 492 41287
rect 579 41272 582 41362
rect 612 41344 624 41345
rect 599 41342 649 41344
rect 612 41341 624 41342
rect 610 41334 632 41341
rect 607 41333 632 41334
rect 586 41326 644 41333
rect 607 41325 644 41326
rect 607 41309 610 41325
rect 616 41309 644 41325
rect 607 41308 644 41309
rect 586 41301 644 41308
rect 607 41300 610 41301
rect 612 41293 632 41301
rect 612 41289 624 41293
rect 649 41292 651 41342
rect 544 41255 548 41263
rect 400 41223 408 41253
rect 420 41223 436 41253
rect 400 41219 436 41223
rect 400 41211 430 41219
rect 428 41195 430 41211
rect 476 41183 480 41251
rect 544 41221 552 41255
rect 578 41221 582 41255
rect 544 41213 548 41221
rect 295 41142 300 41176
rect 324 41142 329 41176
rect 378 41173 450 41181
rect 544 41178 548 41183
rect 544 41174 582 41178
rect 544 41159 552 41174
rect 578 41159 582 41174
rect 544 41141 586 41159
rect 522 41135 608 41141
rect 182 41119 224 41135
rect 544 41119 586 41135
rect 17 41105 67 41107
rect 119 41105 169 41107
rect 186 41105 220 41119
rect 548 41105 582 41119
rect 599 41105 649 41107
rect 42 41063 59 41097
rect 67 41055 69 41105
rect 160 41097 246 41105
rect 522 41097 608 41105
rect 76 41063 110 41097
rect 127 41063 144 41097
rect 152 41063 161 41097
rect 162 41095 195 41097
rect 224 41095 244 41097
rect 162 41063 244 41095
rect 524 41095 548 41097
rect 573 41095 582 41097
rect 586 41095 606 41097
rect 160 41055 246 41063
rect 186 41039 220 41055
rect 182 41025 224 41026
rect 160 41019 182 41025
rect 224 41019 246 41025
rect 186 40984 220 41018
rect 223 40984 257 41018
rect 120 40971 170 40973
rect 76 40967 130 40971
rect 110 40962 130 40967
rect 60 40937 67 40947
rect 76 40937 77 40957
rect 96 40928 99 40962
rect 109 40937 110 40957
rect 119 40937 126 40947
rect 76 40921 92 40927
rect 94 40921 110 40927
rect 170 40921 172 40971
rect 186 40905 190 40939
rect 216 40905 220 40939
rect 288 40905 292 41093
rect 476 41025 480 41093
rect 524 41063 606 41095
rect 607 41063 616 41097
rect 522 41055 608 41063
rect 649 41055 651 41105
rect 548 41039 582 41055
rect 522 41020 548 41025
rect 522 41019 582 41020
rect 586 41019 608 41025
rect 295 40984 300 41018
rect 324 40984 329 41018
rect 544 41016 582 41019
rect 378 40979 450 40987
rect 428 40949 430 40965
rect 400 40941 430 40949
rect 476 40947 480 41015
rect 544 40986 552 41016
rect 578 40986 582 41016
rect 544 40977 548 40986
rect 400 40937 436 40941
rect 400 40907 408 40937
rect 420 40907 436 40937
rect 544 40939 548 40947
rect 12 40868 62 40870
rect 28 40859 59 40867
rect 62 40859 64 40868
rect 28 40851 64 40859
rect 127 40859 158 40867
rect 127 40852 182 40859
rect 215 40857 224 40885
rect 127 40851 161 40852
rect 59 40835 64 40851
rect 158 40835 161 40851
rect 28 40827 64 40835
rect 127 40834 161 40835
rect 127 40827 182 40834
rect 62 40818 64 40827
rect 213 40819 224 40857
rect 282 40847 292 40905
rect 296 40899 368 40907
rect 319 40869 346 40880
rect 318 40856 324 40869
rect 346 40856 348 40869
rect 428 40860 430 40907
rect 443 40897 450 40899
rect 476 40867 480 40935
rect 544 40905 552 40939
rect 578 40905 582 40939
rect 481 40873 517 40901
rect 481 40867 495 40873
rect 367 40856 380 40860
rect 251 40813 263 40847
rect 273 40813 293 40847
rect 295 40832 324 40856
rect 303 40822 316 40832
rect 318 40816 324 40832
rect 333 40832 380 40856
rect 333 40822 353 40832
rect 367 40826 380 40832
rect 396 40826 408 40860
rect 420 40826 436 40860
rect 120 40765 170 40767
rect 76 40759 92 40765
rect 94 40759 110 40765
rect 76 40749 99 40758
rect 60 40739 67 40749
rect 76 40729 77 40749
rect 96 40724 99 40749
rect 109 40729 110 40749
rect 119 40739 126 40749
rect 76 40715 110 40719
rect 170 40715 172 40765
rect 186 40747 190 40781
rect 216 40747 220 40781
rect 186 40670 220 40704
rect 282 40701 292 40813
rect 318 40806 335 40816
rect 318 40737 324 40806
rect 346 40737 348 40822
rect 428 40779 430 40826
rect 476 40789 480 40857
rect 485 40839 495 40867
rect 505 40867 519 40873
rect 544 40867 555 40905
rect 505 40839 525 40867
rect 544 40839 553 40867
rect 544 40819 548 40839
rect 579 40798 582 40888
rect 612 40870 624 40871
rect 599 40868 649 40870
rect 612 40867 624 40868
rect 610 40860 632 40867
rect 607 40859 632 40860
rect 586 40852 644 40859
rect 607 40851 644 40852
rect 607 40835 610 40851
rect 616 40835 644 40851
rect 607 40834 644 40835
rect 586 40827 644 40834
rect 607 40826 610 40827
rect 612 40819 632 40827
rect 612 40815 624 40819
rect 649 40818 651 40868
rect 544 40781 548 40789
rect 400 40749 408 40779
rect 420 40749 436 40779
rect 400 40745 436 40749
rect 400 40737 430 40745
rect 428 40721 430 40737
rect 476 40709 480 40777
rect 544 40747 552 40781
rect 578 40747 582 40781
rect 544 40739 548 40747
rect 544 40709 586 40710
rect 288 40669 292 40701
rect 296 40699 368 40707
rect 378 40699 450 40707
rect 544 40702 548 40709
rect 439 40671 444 40699
rect 120 40655 170 40657
rect 76 40651 130 40655
rect 110 40646 130 40651
rect 60 40621 67 40631
rect 76 40621 77 40641
rect 96 40612 99 40646
rect 109 40621 110 40641
rect 119 40621 126 40631
rect 76 40605 92 40611
rect 94 40605 110 40611
rect 170 40605 172 40655
rect 186 40589 190 40623
rect 216 40589 220 40623
rect 213 40557 224 40589
rect 282 40585 292 40669
rect 296 40663 368 40671
rect 378 40663 450 40671
rect 468 40668 473 40702
rect 428 40633 430 40649
rect 251 40557 292 40585
rect 318 40564 324 40633
rect 12 40552 62 40554
rect 28 40543 59 40551
rect 62 40543 64 40552
rect 251 40551 263 40557
rect 28 40535 64 40543
rect 127 40543 158 40551
rect 127 40536 182 40543
rect 127 40535 161 40536
rect 59 40519 64 40535
rect 158 40519 161 40535
rect 253 40523 263 40551
rect 273 40523 293 40557
rect 318 40554 335 40564
rect 303 40538 316 40548
rect 318 40538 324 40554
rect 346 40548 348 40633
rect 400 40625 430 40633
rect 476 40631 480 40699
rect 511 40668 582 40702
rect 544 40661 548 40668
rect 400 40621 436 40625
rect 400 40591 408 40621
rect 420 40591 436 40621
rect 544 40623 548 40631
rect 28 40511 64 40519
rect 127 40518 161 40519
rect 127 40511 182 40518
rect 62 40502 64 40511
rect 282 40465 292 40523
rect 295 40514 324 40538
rect 333 40538 353 40548
rect 428 40544 430 40591
rect 476 40551 480 40619
rect 544 40589 552 40623
rect 578 40589 582 40623
rect 544 40581 548 40589
rect 367 40538 380 40544
rect 333 40514 380 40538
rect 318 40501 324 40514
rect 346 40501 348 40514
rect 367 40510 380 40514
rect 396 40510 408 40544
rect 420 40510 436 40544
rect 544 40541 553 40569
rect 319 40490 346 40501
rect 120 40449 170 40451
rect 76 40443 92 40449
rect 94 40443 110 40449
rect 76 40433 99 40442
rect 60 40423 67 40433
rect 76 40413 77 40433
rect 96 40408 99 40433
rect 109 40413 110 40433
rect 119 40423 126 40433
rect 76 40399 110 40403
rect 170 40399 172 40449
rect 186 40431 190 40465
rect 216 40431 220 40465
rect 182 40393 224 40394
rect 186 40369 220 40386
rect 223 40369 257 40386
rect 182 40352 257 40369
rect 182 40351 224 40352
rect 160 40345 246 40351
rect 288 40345 292 40465
rect 296 40463 368 40471
rect 428 40463 430 40510
rect 476 40473 480 40541
rect 485 40497 495 40531
rect 505 40503 525 40531
rect 505 40497 519 40503
rect 544 40497 555 40541
rect 485 40473 492 40497
rect 579 40482 582 40572
rect 612 40554 624 40555
rect 599 40552 649 40554
rect 612 40551 624 40552
rect 610 40544 632 40551
rect 607 40543 632 40544
rect 586 40536 644 40543
rect 607 40535 644 40536
rect 607 40519 610 40535
rect 616 40519 644 40535
rect 607 40518 644 40519
rect 586 40511 644 40518
rect 607 40510 610 40511
rect 612 40503 632 40511
rect 612 40499 624 40503
rect 649 40502 651 40552
rect 544 40465 548 40473
rect 400 40433 408 40463
rect 420 40433 436 40463
rect 400 40429 436 40433
rect 400 40421 430 40429
rect 428 40405 430 40421
rect 476 40393 480 40461
rect 544 40431 552 40465
rect 578 40431 582 40465
rect 544 40423 548 40431
rect 295 40352 300 40386
rect 324 40352 329 40386
rect 378 40383 450 40391
rect 544 40388 548 40393
rect 544 40384 582 40388
rect 544 40369 552 40384
rect 578 40369 582 40384
rect 544 40351 586 40369
rect 522 40345 608 40351
rect 182 40329 224 40345
rect 544 40329 586 40345
rect 17 40315 67 40317
rect 119 40315 169 40317
rect 186 40315 220 40329
rect 548 40315 582 40329
rect 599 40315 649 40317
rect 42 40273 59 40307
rect 67 40265 69 40315
rect 160 40307 246 40315
rect 522 40307 608 40315
rect 76 40273 110 40307
rect 127 40273 144 40307
rect 152 40273 161 40307
rect 162 40305 195 40307
rect 224 40305 244 40307
rect 162 40273 244 40305
rect 524 40305 548 40307
rect 573 40305 582 40307
rect 586 40305 606 40307
rect 160 40265 246 40273
rect 186 40249 220 40265
rect 182 40235 224 40236
rect 160 40229 182 40235
rect 224 40229 246 40235
rect 186 40194 220 40228
rect 223 40194 257 40228
rect 120 40181 170 40183
rect 76 40177 130 40181
rect 110 40172 130 40177
rect 60 40147 67 40157
rect 76 40147 77 40167
rect 96 40138 99 40172
rect 109 40147 110 40167
rect 119 40147 126 40157
rect 76 40131 92 40137
rect 94 40131 110 40137
rect 170 40131 172 40181
rect 186 40115 190 40149
rect 216 40115 220 40149
rect 288 40115 292 40303
rect 476 40235 480 40303
rect 524 40273 606 40305
rect 607 40273 616 40307
rect 522 40265 608 40273
rect 649 40265 651 40315
rect 548 40249 582 40265
rect 522 40230 548 40235
rect 522 40229 582 40230
rect 586 40229 608 40235
rect 295 40194 300 40228
rect 324 40194 329 40228
rect 544 40226 582 40229
rect 378 40189 450 40197
rect 428 40159 430 40175
rect 400 40151 430 40159
rect 476 40157 480 40225
rect 544 40196 552 40226
rect 578 40196 582 40226
rect 544 40187 548 40196
rect 400 40147 436 40151
rect 400 40117 408 40147
rect 420 40117 436 40147
rect 544 40149 548 40157
rect 12 40078 62 40080
rect 28 40069 59 40077
rect 62 40069 64 40078
rect 28 40061 64 40069
rect 127 40069 158 40077
rect 127 40062 182 40069
rect 215 40067 224 40095
rect 127 40061 161 40062
rect 59 40045 64 40061
rect 158 40045 161 40061
rect 28 40037 64 40045
rect 127 40044 161 40045
rect 127 40037 182 40044
rect 62 40028 64 40037
rect 213 40029 224 40067
rect 282 40057 292 40115
rect 296 40109 368 40117
rect 319 40079 346 40090
rect 318 40066 324 40079
rect 346 40066 348 40079
rect 428 40070 430 40117
rect 443 40107 450 40109
rect 476 40077 480 40145
rect 544 40115 552 40149
rect 578 40115 582 40149
rect 481 40083 517 40111
rect 481 40077 495 40083
rect 367 40066 380 40070
rect 251 40023 263 40057
rect 273 40023 293 40057
rect 295 40042 324 40066
rect 303 40032 316 40042
rect 318 40026 324 40042
rect 333 40042 380 40066
rect 333 40032 353 40042
rect 367 40036 380 40042
rect 396 40036 408 40070
rect 420 40036 436 40070
rect 120 39975 170 39977
rect 76 39969 92 39975
rect 94 39969 110 39975
rect 76 39959 99 39968
rect 60 39949 67 39959
rect 76 39939 77 39959
rect 96 39934 99 39959
rect 109 39939 110 39959
rect 119 39949 126 39959
rect 76 39925 110 39929
rect 170 39925 172 39975
rect 186 39957 190 39991
rect 216 39957 220 39991
rect 186 39880 220 39914
rect 282 39911 292 40023
rect 318 40016 335 40026
rect 318 39947 324 40016
rect 346 39947 348 40032
rect 428 39989 430 40036
rect 476 39999 480 40067
rect 485 40049 495 40077
rect 505 40077 519 40083
rect 544 40077 555 40115
rect 505 40049 525 40077
rect 544 40049 553 40077
rect 544 40029 548 40049
rect 579 40008 582 40098
rect 612 40080 624 40081
rect 599 40078 649 40080
rect 612 40077 624 40078
rect 610 40070 632 40077
rect 607 40069 632 40070
rect 586 40062 644 40069
rect 607 40061 644 40062
rect 607 40045 610 40061
rect 616 40045 644 40061
rect 607 40044 644 40045
rect 586 40037 644 40044
rect 607 40036 610 40037
rect 612 40029 632 40037
rect 612 40025 624 40029
rect 649 40028 651 40078
rect 544 39991 548 39999
rect 400 39959 408 39989
rect 420 39959 436 39989
rect 400 39955 436 39959
rect 400 39947 430 39955
rect 428 39931 430 39947
rect 476 39919 480 39987
rect 544 39957 552 39991
rect 578 39957 582 39991
rect 544 39949 548 39957
rect 544 39919 586 39920
rect 288 39879 292 39911
rect 296 39909 368 39917
rect 378 39909 450 39917
rect 544 39912 548 39919
rect 439 39881 444 39909
rect 120 39865 170 39867
rect 76 39861 130 39865
rect 110 39856 130 39861
rect 60 39831 67 39841
rect 76 39831 77 39851
rect 96 39822 99 39856
rect 109 39831 110 39851
rect 119 39831 126 39841
rect 76 39815 92 39821
rect 94 39815 110 39821
rect 170 39815 172 39865
rect 186 39799 190 39833
rect 216 39799 220 39833
rect 213 39767 224 39799
rect 282 39795 292 39879
rect 296 39873 368 39881
rect 378 39873 450 39881
rect 468 39878 473 39912
rect 428 39843 430 39859
rect 251 39767 292 39795
rect 318 39774 324 39843
rect 12 39762 62 39764
rect 28 39753 59 39761
rect 62 39753 64 39762
rect 251 39761 263 39767
rect 28 39745 64 39753
rect 127 39753 158 39761
rect 127 39746 182 39753
rect 127 39745 161 39746
rect 59 39729 64 39745
rect 158 39729 161 39745
rect 253 39733 263 39761
rect 273 39733 293 39767
rect 318 39764 335 39774
rect 303 39748 316 39758
rect 318 39748 324 39764
rect 346 39758 348 39843
rect 400 39835 430 39843
rect 476 39841 480 39909
rect 511 39878 582 39912
rect 544 39871 548 39878
rect 400 39831 436 39835
rect 400 39801 408 39831
rect 420 39801 436 39831
rect 544 39833 548 39841
rect 28 39721 64 39729
rect 127 39728 161 39729
rect 127 39721 182 39728
rect 62 39712 64 39721
rect 282 39675 292 39733
rect 295 39724 324 39748
rect 333 39748 353 39758
rect 428 39754 430 39801
rect 476 39761 480 39829
rect 544 39799 552 39833
rect 578 39799 582 39833
rect 544 39791 548 39799
rect 367 39748 380 39754
rect 333 39724 380 39748
rect 318 39711 324 39724
rect 346 39711 348 39724
rect 367 39720 380 39724
rect 396 39720 408 39754
rect 420 39720 436 39754
rect 544 39751 553 39779
rect 319 39700 346 39711
rect 120 39659 170 39661
rect 76 39653 92 39659
rect 94 39653 110 39659
rect 76 39643 99 39652
rect 60 39633 67 39643
rect 76 39623 77 39643
rect 96 39618 99 39643
rect 109 39623 110 39643
rect 119 39633 126 39643
rect 76 39609 110 39613
rect 170 39609 172 39659
rect 186 39641 190 39675
rect 216 39641 220 39675
rect 182 39603 224 39604
rect 186 39579 220 39596
rect 223 39579 257 39596
rect 182 39562 257 39579
rect 182 39561 224 39562
rect 160 39555 246 39561
rect 288 39555 292 39675
rect 296 39673 368 39681
rect 428 39673 430 39720
rect 476 39683 480 39751
rect 485 39707 495 39741
rect 505 39713 525 39741
rect 505 39707 519 39713
rect 544 39707 555 39751
rect 485 39683 492 39707
rect 579 39692 582 39782
rect 612 39764 624 39765
rect 599 39762 649 39764
rect 612 39761 624 39762
rect 610 39754 632 39761
rect 607 39753 632 39754
rect 586 39746 644 39753
rect 607 39745 644 39746
rect 607 39729 610 39745
rect 616 39729 644 39745
rect 607 39728 644 39729
rect 586 39721 644 39728
rect 607 39720 610 39721
rect 612 39713 632 39721
rect 612 39709 624 39713
rect 649 39712 651 39762
rect 544 39675 548 39683
rect 400 39643 408 39673
rect 420 39643 436 39673
rect 400 39639 436 39643
rect 400 39631 430 39639
rect 428 39615 430 39631
rect 476 39603 480 39671
rect 544 39641 552 39675
rect 578 39641 582 39675
rect 544 39633 548 39641
rect 295 39562 300 39596
rect 324 39562 329 39596
rect 378 39593 450 39601
rect 544 39598 548 39603
rect 544 39594 582 39598
rect 544 39579 552 39594
rect 578 39579 582 39594
rect 544 39561 586 39579
rect 522 39555 608 39561
rect 182 39539 224 39555
rect 544 39539 586 39555
rect 17 39525 67 39527
rect 119 39525 169 39527
rect 186 39525 220 39539
rect 548 39525 582 39539
rect 599 39525 649 39527
rect 42 39483 59 39517
rect 67 39475 69 39525
rect 160 39517 246 39525
rect 522 39517 608 39525
rect 76 39483 110 39517
rect 127 39483 144 39517
rect 152 39483 161 39517
rect 162 39515 195 39517
rect 224 39515 244 39517
rect 162 39483 244 39515
rect 524 39515 548 39517
rect 573 39515 582 39517
rect 586 39515 606 39517
rect 160 39475 246 39483
rect 186 39459 220 39475
rect 182 39445 224 39446
rect 160 39439 182 39445
rect 224 39439 246 39445
rect 186 39404 220 39438
rect 223 39404 257 39438
rect 120 39391 170 39393
rect 76 39387 130 39391
rect 110 39382 130 39387
rect 60 39357 67 39367
rect 76 39357 77 39377
rect 96 39348 99 39382
rect 109 39357 110 39377
rect 119 39357 126 39367
rect 76 39341 92 39347
rect 94 39341 110 39347
rect 170 39341 172 39391
rect 186 39325 190 39359
rect 216 39325 220 39359
rect 288 39325 292 39513
rect 476 39445 480 39513
rect 524 39483 606 39515
rect 607 39483 616 39517
rect 522 39475 608 39483
rect 649 39475 651 39525
rect 548 39459 582 39475
rect 522 39440 548 39445
rect 522 39439 582 39440
rect 586 39439 608 39445
rect 295 39404 300 39438
rect 324 39404 329 39438
rect 544 39436 582 39439
rect 378 39399 450 39407
rect 428 39369 430 39385
rect 400 39361 430 39369
rect 476 39367 480 39435
rect 544 39406 552 39436
rect 578 39406 582 39436
rect 544 39397 548 39406
rect 400 39357 436 39361
rect 400 39327 408 39357
rect 420 39327 436 39357
rect 544 39359 548 39367
rect 12 39288 62 39290
rect 28 39279 59 39287
rect 62 39279 64 39288
rect 28 39271 64 39279
rect 127 39279 158 39287
rect 127 39272 182 39279
rect 215 39277 224 39305
rect 127 39271 161 39272
rect 59 39255 64 39271
rect 158 39255 161 39271
rect 28 39247 64 39255
rect 127 39254 161 39255
rect 127 39247 182 39254
rect 62 39238 64 39247
rect 213 39239 224 39277
rect 282 39267 292 39325
rect 296 39319 368 39327
rect 319 39289 346 39300
rect 318 39276 324 39289
rect 346 39276 348 39289
rect 428 39280 430 39327
rect 443 39317 450 39319
rect 476 39287 480 39355
rect 544 39325 552 39359
rect 578 39325 582 39359
rect 481 39293 517 39321
rect 481 39287 495 39293
rect 367 39276 380 39280
rect 251 39233 263 39267
rect 273 39233 293 39267
rect 295 39252 324 39276
rect 303 39242 316 39252
rect 318 39236 324 39252
rect 333 39252 380 39276
rect 333 39242 353 39252
rect 367 39246 380 39252
rect 396 39246 408 39280
rect 420 39246 436 39280
rect 120 39185 170 39187
rect 76 39179 92 39185
rect 94 39179 110 39185
rect 76 39169 99 39178
rect 60 39159 67 39169
rect 76 39149 77 39169
rect 96 39144 99 39169
rect 109 39149 110 39169
rect 119 39159 126 39169
rect 76 39135 110 39139
rect 170 39135 172 39185
rect 186 39167 190 39201
rect 216 39167 220 39201
rect 186 39090 220 39124
rect 282 39121 292 39233
rect 318 39226 335 39236
rect 318 39157 324 39226
rect 346 39157 348 39242
rect 428 39199 430 39246
rect 476 39209 480 39277
rect 485 39259 495 39287
rect 505 39287 519 39293
rect 544 39287 555 39325
rect 505 39259 525 39287
rect 544 39259 553 39287
rect 544 39239 548 39259
rect 579 39218 582 39308
rect 612 39290 624 39291
rect 599 39288 649 39290
rect 612 39287 624 39288
rect 610 39280 632 39287
rect 607 39279 632 39280
rect 586 39272 644 39279
rect 607 39271 644 39272
rect 607 39255 610 39271
rect 616 39255 644 39271
rect 607 39254 644 39255
rect 586 39247 644 39254
rect 607 39246 610 39247
rect 612 39239 632 39247
rect 612 39235 624 39239
rect 649 39238 651 39288
rect 544 39201 548 39209
rect 400 39169 408 39199
rect 420 39169 436 39199
rect 400 39165 436 39169
rect 400 39157 430 39165
rect 428 39141 430 39157
rect 476 39129 480 39197
rect 544 39167 552 39201
rect 578 39167 582 39201
rect 544 39159 548 39167
rect 544 39129 586 39130
rect 288 39089 292 39121
rect 296 39119 368 39127
rect 378 39119 450 39127
rect 544 39122 548 39129
rect 439 39091 444 39119
rect 120 39075 170 39077
rect 76 39071 130 39075
rect 110 39066 130 39071
rect 60 39041 67 39051
rect 76 39041 77 39061
rect 96 39032 99 39066
rect 109 39041 110 39061
rect 119 39041 126 39051
rect 76 39025 92 39031
rect 94 39025 110 39031
rect 170 39025 172 39075
rect 186 39009 190 39043
rect 216 39009 220 39043
rect 213 38977 224 39009
rect 282 39005 292 39089
rect 296 39083 368 39091
rect 378 39083 450 39091
rect 468 39088 473 39122
rect 428 39053 430 39069
rect 251 38977 292 39005
rect 318 38984 324 39053
rect 12 38972 62 38974
rect 28 38963 59 38971
rect 62 38963 64 38972
rect 251 38971 263 38977
rect 28 38955 64 38963
rect 127 38963 158 38971
rect 127 38956 182 38963
rect 127 38955 161 38956
rect 59 38939 64 38955
rect 158 38939 161 38955
rect 253 38943 263 38971
rect 273 38943 293 38977
rect 318 38974 335 38984
rect 303 38958 316 38968
rect 318 38958 324 38974
rect 346 38968 348 39053
rect 400 39045 430 39053
rect 476 39051 480 39119
rect 511 39088 582 39122
rect 544 39081 548 39088
rect 400 39041 436 39045
rect 400 39011 408 39041
rect 420 39011 436 39041
rect 544 39043 548 39051
rect 28 38931 64 38939
rect 127 38938 161 38939
rect 127 38931 182 38938
rect 62 38922 64 38931
rect 282 38885 292 38943
rect 295 38934 324 38958
rect 333 38958 353 38968
rect 428 38964 430 39011
rect 476 38971 480 39039
rect 544 39009 552 39043
rect 578 39009 582 39043
rect 544 39001 548 39009
rect 367 38958 380 38964
rect 333 38934 380 38958
rect 318 38921 324 38934
rect 346 38921 348 38934
rect 367 38930 380 38934
rect 396 38930 408 38964
rect 420 38930 436 38964
rect 544 38961 553 38989
rect 319 38910 346 38921
rect 120 38869 170 38871
rect 76 38863 92 38869
rect 94 38863 110 38869
rect 76 38853 99 38862
rect 60 38843 67 38853
rect 76 38833 77 38853
rect 96 38828 99 38853
rect 109 38833 110 38853
rect 119 38843 126 38853
rect 76 38819 110 38823
rect 170 38819 172 38869
rect 186 38851 190 38885
rect 216 38851 220 38885
rect 182 38813 224 38814
rect 186 38789 220 38806
rect 223 38789 257 38806
rect 182 38772 257 38789
rect 182 38771 224 38772
rect 160 38765 246 38771
rect 288 38765 292 38885
rect 296 38883 368 38891
rect 428 38883 430 38930
rect 476 38893 480 38961
rect 485 38917 495 38951
rect 505 38923 525 38951
rect 505 38917 519 38923
rect 544 38917 555 38961
rect 485 38893 492 38917
rect 579 38902 582 38992
rect 612 38974 624 38975
rect 599 38972 649 38974
rect 612 38971 624 38972
rect 610 38964 632 38971
rect 607 38963 632 38964
rect 586 38956 644 38963
rect 607 38955 644 38956
rect 607 38939 610 38955
rect 616 38939 644 38955
rect 607 38938 644 38939
rect 586 38931 644 38938
rect 607 38930 610 38931
rect 612 38923 632 38931
rect 612 38919 624 38923
rect 649 38922 651 38972
rect 544 38885 548 38893
rect 400 38853 408 38883
rect 420 38853 436 38883
rect 400 38849 436 38853
rect 400 38841 430 38849
rect 428 38825 430 38841
rect 476 38813 480 38881
rect 544 38851 552 38885
rect 578 38851 582 38885
rect 544 38843 548 38851
rect 295 38772 300 38806
rect 324 38772 329 38806
rect 378 38803 450 38811
rect 544 38808 548 38813
rect 544 38804 582 38808
rect 544 38789 552 38804
rect 578 38789 582 38804
rect 544 38771 586 38789
rect 522 38765 608 38771
rect 182 38749 224 38765
rect 544 38749 586 38765
rect 17 38735 67 38737
rect 119 38735 169 38737
rect 186 38735 220 38749
rect 548 38735 582 38749
rect 599 38735 649 38737
rect 42 38693 59 38727
rect 67 38685 69 38735
rect 160 38727 246 38735
rect 522 38727 608 38735
rect 76 38693 110 38727
rect 127 38693 144 38727
rect 152 38693 161 38727
rect 162 38725 195 38727
rect 224 38725 244 38727
rect 162 38693 244 38725
rect 524 38725 548 38727
rect 573 38725 582 38727
rect 586 38725 606 38727
rect 160 38685 246 38693
rect 186 38669 220 38685
rect 182 38655 224 38656
rect 160 38649 182 38655
rect 224 38649 246 38655
rect 186 38614 220 38648
rect 223 38614 257 38648
rect 120 38601 170 38603
rect 76 38597 130 38601
rect 110 38592 130 38597
rect 60 38567 67 38577
rect 76 38567 77 38587
rect 96 38558 99 38592
rect 109 38567 110 38587
rect 119 38567 126 38577
rect 76 38551 92 38557
rect 94 38551 110 38557
rect 170 38551 172 38601
rect 186 38535 190 38569
rect 216 38535 220 38569
rect 288 38535 292 38723
rect 476 38655 480 38723
rect 524 38693 606 38725
rect 607 38693 616 38727
rect 522 38685 608 38693
rect 649 38685 651 38735
rect 548 38669 582 38685
rect 522 38650 548 38655
rect 522 38649 582 38650
rect 586 38649 608 38655
rect 295 38614 300 38648
rect 324 38614 329 38648
rect 544 38646 582 38649
rect 378 38609 450 38617
rect 428 38579 430 38595
rect 400 38571 430 38579
rect 476 38577 480 38645
rect 544 38616 552 38646
rect 578 38616 582 38646
rect 544 38607 548 38616
rect 400 38567 436 38571
rect 400 38537 408 38567
rect 420 38537 436 38567
rect 544 38569 548 38577
rect 12 38498 62 38500
rect 28 38489 59 38497
rect 62 38489 64 38498
rect 28 38481 64 38489
rect 127 38489 158 38497
rect 127 38482 182 38489
rect 215 38487 224 38515
rect 127 38481 161 38482
rect 59 38465 64 38481
rect 158 38465 161 38481
rect 28 38457 64 38465
rect 127 38464 161 38465
rect 127 38457 182 38464
rect 62 38448 64 38457
rect 213 38449 224 38487
rect 282 38477 292 38535
rect 296 38529 368 38537
rect 319 38499 346 38510
rect 318 38486 324 38499
rect 346 38486 348 38499
rect 428 38490 430 38537
rect 443 38527 450 38529
rect 476 38497 480 38565
rect 544 38535 552 38569
rect 578 38535 582 38569
rect 481 38503 517 38531
rect 481 38497 495 38503
rect 367 38486 380 38490
rect 251 38443 263 38477
rect 273 38443 293 38477
rect 295 38462 324 38486
rect 303 38452 316 38462
rect 318 38446 324 38462
rect 333 38462 380 38486
rect 333 38452 353 38462
rect 367 38456 380 38462
rect 396 38456 408 38490
rect 420 38456 436 38490
rect 120 38395 170 38397
rect 76 38389 92 38395
rect 94 38389 110 38395
rect 76 38379 99 38388
rect 60 38369 67 38379
rect 76 38359 77 38379
rect 96 38354 99 38379
rect 109 38359 110 38379
rect 119 38369 126 38379
rect 76 38345 110 38349
rect 170 38345 172 38395
rect 186 38377 190 38411
rect 216 38377 220 38411
rect 186 38300 220 38334
rect 282 38331 292 38443
rect 318 38436 335 38446
rect 318 38367 324 38436
rect 346 38367 348 38452
rect 428 38409 430 38456
rect 476 38419 480 38487
rect 485 38469 495 38497
rect 505 38497 519 38503
rect 544 38497 555 38535
rect 505 38469 525 38497
rect 544 38469 553 38497
rect 544 38449 548 38469
rect 579 38428 582 38518
rect 612 38500 624 38501
rect 599 38498 649 38500
rect 612 38497 624 38498
rect 610 38490 632 38497
rect 607 38489 632 38490
rect 586 38482 644 38489
rect 607 38481 644 38482
rect 607 38465 610 38481
rect 616 38465 644 38481
rect 607 38464 644 38465
rect 586 38457 644 38464
rect 607 38456 610 38457
rect 612 38449 632 38457
rect 612 38445 624 38449
rect 649 38448 651 38498
rect 544 38411 548 38419
rect 400 38379 408 38409
rect 420 38379 436 38409
rect 400 38375 436 38379
rect 400 38367 430 38375
rect 428 38351 430 38367
rect 476 38339 480 38407
rect 544 38377 552 38411
rect 578 38377 582 38411
rect 544 38369 548 38377
rect 544 38339 586 38340
rect 288 38299 292 38331
rect 296 38329 368 38337
rect 378 38329 450 38337
rect 544 38332 548 38339
rect 439 38301 444 38329
rect 120 38285 170 38287
rect 76 38281 130 38285
rect 110 38276 130 38281
rect 60 38251 67 38261
rect 76 38251 77 38271
rect 96 38242 99 38276
rect 109 38251 110 38271
rect 119 38251 126 38261
rect 76 38235 92 38241
rect 94 38235 110 38241
rect 170 38235 172 38285
rect 186 38219 190 38253
rect 216 38219 220 38253
rect 213 38187 224 38219
rect 282 38215 292 38299
rect 296 38293 368 38301
rect 378 38293 450 38301
rect 468 38298 473 38332
rect 428 38263 430 38279
rect 251 38187 292 38215
rect 318 38194 324 38263
rect 12 38182 62 38184
rect 28 38173 59 38181
rect 62 38173 64 38182
rect 251 38181 263 38187
rect 28 38165 64 38173
rect 127 38173 158 38181
rect 127 38166 182 38173
rect 127 38165 161 38166
rect 59 38149 64 38165
rect 158 38149 161 38165
rect 253 38153 263 38181
rect 273 38153 293 38187
rect 318 38184 335 38194
rect 303 38168 316 38178
rect 318 38168 324 38184
rect 346 38178 348 38263
rect 400 38255 430 38263
rect 476 38261 480 38329
rect 511 38298 582 38332
rect 544 38291 548 38298
rect 400 38251 436 38255
rect 400 38221 408 38251
rect 420 38221 436 38251
rect 544 38253 548 38261
rect 28 38141 64 38149
rect 127 38148 161 38149
rect 127 38141 182 38148
rect 62 38132 64 38141
rect 282 38095 292 38153
rect 295 38144 324 38168
rect 333 38168 353 38178
rect 428 38174 430 38221
rect 476 38181 480 38249
rect 544 38219 552 38253
rect 578 38219 582 38253
rect 544 38211 548 38219
rect 367 38168 380 38174
rect 333 38144 380 38168
rect 318 38131 324 38144
rect 346 38131 348 38144
rect 367 38140 380 38144
rect 396 38140 408 38174
rect 420 38140 436 38174
rect 544 38171 553 38199
rect 319 38120 346 38131
rect 120 38079 170 38081
rect 76 38073 92 38079
rect 94 38073 110 38079
rect 76 38063 99 38072
rect 60 38053 67 38063
rect 76 38043 77 38063
rect 96 38038 99 38063
rect 109 38043 110 38063
rect 119 38053 126 38063
rect 76 38029 110 38033
rect 170 38029 172 38079
rect 186 38061 190 38095
rect 216 38061 220 38095
rect 182 38023 224 38024
rect 186 37999 220 38016
rect 223 37999 257 38016
rect 182 37982 257 37999
rect 182 37981 224 37982
rect 160 37975 246 37981
rect 288 37975 292 38095
rect 296 38093 368 38101
rect 428 38093 430 38140
rect 476 38103 480 38171
rect 485 38127 495 38161
rect 505 38133 525 38161
rect 505 38127 519 38133
rect 544 38127 555 38171
rect 485 38103 492 38127
rect 579 38112 582 38202
rect 612 38184 624 38185
rect 599 38182 649 38184
rect 612 38181 624 38182
rect 610 38174 632 38181
rect 607 38173 632 38174
rect 586 38166 644 38173
rect 607 38165 644 38166
rect 607 38149 610 38165
rect 616 38149 644 38165
rect 607 38148 644 38149
rect 586 38141 644 38148
rect 607 38140 610 38141
rect 612 38133 632 38141
rect 612 38129 624 38133
rect 649 38132 651 38182
rect 544 38095 548 38103
rect 400 38063 408 38093
rect 420 38063 436 38093
rect 400 38059 436 38063
rect 400 38051 430 38059
rect 428 38035 430 38051
rect 476 38023 480 38091
rect 544 38061 552 38095
rect 578 38061 582 38095
rect 544 38053 548 38061
rect 295 37982 300 38016
rect 324 37982 329 38016
rect 378 38013 450 38021
rect 544 38018 548 38023
rect 544 38014 582 38018
rect 544 37999 552 38014
rect 578 37999 582 38014
rect 544 37981 586 37999
rect 522 37975 608 37981
rect 182 37959 224 37975
rect 544 37959 586 37975
rect 17 37945 67 37947
rect 119 37945 169 37947
rect 186 37945 220 37959
rect 548 37945 582 37959
rect 599 37945 649 37947
rect 42 37903 59 37937
rect 67 37895 69 37945
rect 160 37937 246 37945
rect 522 37937 608 37945
rect 76 37903 110 37937
rect 127 37903 144 37937
rect 152 37903 161 37937
rect 162 37935 195 37937
rect 224 37935 244 37937
rect 162 37903 244 37935
rect 524 37935 548 37937
rect 573 37935 582 37937
rect 586 37935 606 37937
rect 160 37895 246 37903
rect 186 37879 220 37895
rect 182 37865 224 37866
rect 160 37859 182 37865
rect 224 37859 246 37865
rect 186 37824 220 37858
rect 223 37824 257 37858
rect 120 37811 170 37813
rect 76 37807 130 37811
rect 110 37802 130 37807
rect 60 37777 67 37787
rect 76 37777 77 37797
rect 96 37768 99 37802
rect 109 37777 110 37797
rect 119 37777 126 37787
rect 76 37761 92 37767
rect 94 37761 110 37767
rect 170 37761 172 37811
rect 186 37745 190 37779
rect 216 37745 220 37779
rect 288 37745 292 37933
rect 476 37865 480 37933
rect 524 37903 606 37935
rect 607 37903 616 37937
rect 522 37895 608 37903
rect 649 37895 651 37945
rect 548 37879 582 37895
rect 522 37860 548 37865
rect 522 37859 582 37860
rect 586 37859 608 37865
rect 295 37824 300 37858
rect 324 37824 329 37858
rect 544 37856 582 37859
rect 378 37819 450 37827
rect 428 37789 430 37805
rect 400 37781 430 37789
rect 476 37787 480 37855
rect 544 37826 552 37856
rect 578 37826 582 37856
rect 544 37817 548 37826
rect 400 37777 436 37781
rect 400 37747 408 37777
rect 420 37747 436 37777
rect 544 37779 548 37787
rect 12 37708 62 37710
rect 28 37699 59 37707
rect 62 37699 64 37708
rect 28 37691 64 37699
rect 127 37699 158 37707
rect 127 37692 182 37699
rect 215 37697 224 37725
rect 127 37691 161 37692
rect 59 37675 64 37691
rect 158 37675 161 37691
rect 28 37667 64 37675
rect 127 37674 161 37675
rect 127 37667 182 37674
rect 62 37658 64 37667
rect 213 37659 224 37697
rect 282 37687 292 37745
rect 296 37739 368 37747
rect 319 37709 346 37720
rect 318 37696 324 37709
rect 346 37696 348 37709
rect 428 37700 430 37747
rect 443 37737 450 37739
rect 476 37707 480 37775
rect 544 37745 552 37779
rect 578 37745 582 37779
rect 481 37713 517 37741
rect 481 37707 495 37713
rect 367 37696 380 37700
rect 251 37653 263 37687
rect 273 37653 293 37687
rect 295 37672 324 37696
rect 303 37662 316 37672
rect 318 37656 324 37672
rect 333 37672 380 37696
rect 333 37662 353 37672
rect 367 37666 380 37672
rect 396 37666 408 37700
rect 420 37666 436 37700
rect 120 37605 170 37607
rect 76 37599 92 37605
rect 94 37599 110 37605
rect 76 37589 99 37598
rect 60 37579 67 37589
rect 76 37569 77 37589
rect 96 37564 99 37589
rect 109 37569 110 37589
rect 119 37579 126 37589
rect 76 37555 110 37559
rect 170 37555 172 37605
rect 186 37587 190 37621
rect 216 37587 220 37621
rect 186 37510 220 37544
rect 282 37541 292 37653
rect 318 37646 335 37656
rect 318 37577 324 37646
rect 346 37577 348 37662
rect 428 37619 430 37666
rect 476 37629 480 37697
rect 485 37679 495 37707
rect 505 37707 519 37713
rect 544 37707 555 37745
rect 505 37679 525 37707
rect 544 37679 553 37707
rect 544 37659 548 37679
rect 579 37638 582 37728
rect 612 37710 624 37711
rect 599 37708 649 37710
rect 612 37707 624 37708
rect 610 37700 632 37707
rect 607 37699 632 37700
rect 586 37692 644 37699
rect 607 37691 644 37692
rect 607 37675 610 37691
rect 616 37675 644 37691
rect 607 37674 644 37675
rect 586 37667 644 37674
rect 607 37666 610 37667
rect 612 37659 632 37667
rect 612 37655 624 37659
rect 649 37658 651 37708
rect 544 37621 548 37629
rect 400 37589 408 37619
rect 420 37589 436 37619
rect 400 37585 436 37589
rect 400 37577 430 37585
rect 428 37561 430 37577
rect 476 37549 480 37617
rect 544 37587 552 37621
rect 578 37587 582 37621
rect 544 37579 548 37587
rect 544 37549 586 37550
rect 288 37509 292 37541
rect 296 37539 368 37547
rect 378 37539 450 37547
rect 544 37542 548 37549
rect 439 37511 444 37539
rect 120 37495 170 37497
rect 76 37491 130 37495
rect 110 37486 130 37491
rect 60 37461 67 37471
rect 76 37461 77 37481
rect 96 37452 99 37486
rect 109 37461 110 37481
rect 119 37461 126 37471
rect 76 37445 92 37451
rect 94 37445 110 37451
rect 170 37445 172 37495
rect 186 37429 190 37463
rect 216 37429 220 37463
rect 213 37397 224 37429
rect 282 37425 292 37509
rect 296 37503 368 37511
rect 378 37503 450 37511
rect 468 37508 473 37542
rect 428 37473 430 37489
rect 251 37397 292 37425
rect 318 37404 324 37473
rect 12 37392 62 37394
rect 28 37383 59 37391
rect 62 37383 64 37392
rect 251 37391 263 37397
rect 28 37375 64 37383
rect 127 37383 158 37391
rect 127 37376 182 37383
rect 127 37375 161 37376
rect 59 37359 64 37375
rect 158 37359 161 37375
rect 253 37363 263 37391
rect 273 37363 293 37397
rect 318 37394 335 37404
rect 303 37378 316 37388
rect 318 37378 324 37394
rect 346 37388 348 37473
rect 400 37465 430 37473
rect 476 37471 480 37539
rect 511 37508 582 37542
rect 544 37501 548 37508
rect 400 37461 436 37465
rect 400 37431 408 37461
rect 420 37431 436 37461
rect 544 37463 548 37471
rect 28 37351 64 37359
rect 127 37358 161 37359
rect 127 37351 182 37358
rect 62 37342 64 37351
rect 282 37305 292 37363
rect 295 37354 324 37378
rect 333 37378 353 37388
rect 428 37384 430 37431
rect 476 37391 480 37459
rect 544 37429 552 37463
rect 578 37429 582 37463
rect 544 37421 548 37429
rect 367 37378 380 37384
rect 333 37354 380 37378
rect 318 37341 324 37354
rect 346 37341 348 37354
rect 367 37350 380 37354
rect 396 37350 408 37384
rect 420 37350 436 37384
rect 544 37381 553 37409
rect 319 37330 346 37341
rect 120 37289 170 37291
rect 76 37283 92 37289
rect 94 37283 110 37289
rect 76 37273 99 37282
rect 60 37263 67 37273
rect 76 37253 77 37273
rect 96 37248 99 37273
rect 109 37253 110 37273
rect 119 37263 126 37273
rect 76 37239 110 37243
rect 170 37239 172 37289
rect 186 37271 190 37305
rect 216 37271 220 37305
rect 182 37233 224 37234
rect 186 37209 220 37226
rect 223 37209 257 37226
rect 182 37192 257 37209
rect 182 37191 224 37192
rect 160 37185 246 37191
rect 288 37185 292 37305
rect 296 37303 368 37311
rect 428 37303 430 37350
rect 476 37313 480 37381
rect 485 37337 495 37371
rect 505 37343 525 37371
rect 505 37337 519 37343
rect 544 37337 555 37381
rect 485 37313 492 37337
rect 579 37322 582 37412
rect 612 37394 624 37395
rect 599 37392 649 37394
rect 612 37391 624 37392
rect 610 37384 632 37391
rect 607 37383 632 37384
rect 586 37376 644 37383
rect 607 37375 644 37376
rect 607 37359 610 37375
rect 616 37359 644 37375
rect 607 37358 644 37359
rect 586 37351 644 37358
rect 607 37350 610 37351
rect 612 37343 632 37351
rect 612 37339 624 37343
rect 649 37342 651 37392
rect 544 37305 548 37313
rect 400 37273 408 37303
rect 420 37273 436 37303
rect 400 37269 436 37273
rect 400 37261 430 37269
rect 428 37245 430 37261
rect 476 37233 480 37301
rect 544 37271 552 37305
rect 578 37271 582 37305
rect 544 37263 548 37271
rect 295 37192 300 37226
rect 324 37192 329 37226
rect 378 37223 450 37231
rect 544 37228 548 37233
rect 544 37224 582 37228
rect 544 37209 552 37224
rect 578 37209 582 37224
rect 544 37191 586 37209
rect 522 37185 608 37191
rect 182 37169 224 37185
rect 544 37169 586 37185
rect 17 37155 67 37157
rect 119 37155 169 37157
rect 186 37155 220 37169
rect 548 37155 582 37169
rect 599 37155 649 37157
rect 42 37113 59 37147
rect 67 37105 69 37155
rect 160 37147 246 37155
rect 522 37147 608 37155
rect 76 37113 110 37147
rect 127 37113 144 37147
rect 152 37113 161 37147
rect 162 37145 195 37147
rect 224 37145 244 37147
rect 162 37113 244 37145
rect 524 37145 548 37147
rect 573 37145 582 37147
rect 586 37145 606 37147
rect 160 37105 246 37113
rect 186 37089 220 37105
rect 182 37075 224 37076
rect 160 37069 182 37075
rect 224 37069 246 37075
rect 186 37034 220 37068
rect 223 37034 257 37068
rect 120 37021 170 37023
rect 76 37017 130 37021
rect 110 37012 130 37017
rect 60 36987 67 36997
rect 76 36987 77 37007
rect 96 36978 99 37012
rect 109 36987 110 37007
rect 119 36987 126 36997
rect 76 36971 92 36977
rect 94 36971 110 36977
rect 170 36971 172 37021
rect 186 36955 190 36989
rect 216 36955 220 36989
rect 288 36955 292 37143
rect 476 37075 480 37143
rect 524 37113 606 37145
rect 607 37113 616 37147
rect 522 37105 608 37113
rect 649 37105 651 37155
rect 548 37089 582 37105
rect 522 37070 548 37075
rect 522 37069 582 37070
rect 586 37069 608 37075
rect 295 37034 300 37068
rect 324 37034 329 37068
rect 544 37066 582 37069
rect 378 37029 450 37037
rect 428 36999 430 37015
rect 400 36991 430 36999
rect 476 36997 480 37065
rect 544 37036 552 37066
rect 578 37036 582 37066
rect 544 37027 548 37036
rect 400 36987 436 36991
rect 400 36957 408 36987
rect 420 36957 436 36987
rect 544 36989 548 36997
rect 12 36918 62 36920
rect 28 36909 59 36917
rect 62 36909 64 36918
rect 28 36901 64 36909
rect 127 36909 158 36917
rect 127 36902 182 36909
rect 215 36907 224 36935
rect 127 36901 161 36902
rect 59 36885 64 36901
rect 158 36885 161 36901
rect 28 36877 64 36885
rect 127 36884 161 36885
rect 127 36877 182 36884
rect 62 36868 64 36877
rect 213 36869 224 36907
rect 282 36897 292 36955
rect 296 36949 368 36957
rect 319 36919 346 36930
rect 318 36906 324 36919
rect 346 36906 348 36919
rect 428 36910 430 36957
rect 443 36947 450 36949
rect 476 36917 480 36985
rect 544 36955 552 36989
rect 578 36955 582 36989
rect 481 36923 517 36951
rect 481 36917 495 36923
rect 367 36906 380 36910
rect 251 36863 263 36897
rect 273 36863 293 36897
rect 295 36882 324 36906
rect 303 36872 316 36882
rect 318 36866 324 36882
rect 333 36882 380 36906
rect 333 36872 353 36882
rect 367 36876 380 36882
rect 396 36876 408 36910
rect 420 36876 436 36910
rect 120 36815 170 36817
rect 76 36809 92 36815
rect 94 36809 110 36815
rect 76 36799 99 36808
rect 60 36789 67 36799
rect 76 36779 77 36799
rect 96 36774 99 36799
rect 109 36779 110 36799
rect 119 36789 126 36799
rect 76 36765 110 36769
rect 170 36765 172 36815
rect 186 36797 190 36831
rect 216 36797 220 36831
rect 186 36720 220 36754
rect 282 36751 292 36863
rect 318 36856 335 36866
rect 318 36787 324 36856
rect 346 36787 348 36872
rect 428 36829 430 36876
rect 476 36839 480 36907
rect 485 36889 495 36917
rect 505 36917 519 36923
rect 544 36917 555 36955
rect 505 36889 525 36917
rect 544 36889 553 36917
rect 544 36869 548 36889
rect 579 36848 582 36938
rect 612 36920 624 36921
rect 599 36918 649 36920
rect 612 36917 624 36918
rect 610 36910 632 36917
rect 607 36909 632 36910
rect 586 36902 644 36909
rect 607 36901 644 36902
rect 607 36885 610 36901
rect 616 36885 644 36901
rect 607 36884 644 36885
rect 586 36877 644 36884
rect 607 36876 610 36877
rect 612 36869 632 36877
rect 612 36865 624 36869
rect 649 36868 651 36918
rect 544 36831 548 36839
rect 400 36799 408 36829
rect 420 36799 436 36829
rect 400 36795 436 36799
rect 400 36787 430 36795
rect 428 36771 430 36787
rect 476 36759 480 36827
rect 544 36797 552 36831
rect 578 36797 582 36831
rect 544 36789 548 36797
rect 544 36759 586 36760
rect 288 36719 292 36751
rect 296 36749 368 36757
rect 378 36749 450 36757
rect 544 36752 548 36759
rect 439 36721 444 36749
rect 120 36705 170 36707
rect 76 36701 130 36705
rect 110 36696 130 36701
rect 60 36671 67 36681
rect 76 36671 77 36691
rect 96 36662 99 36696
rect 109 36671 110 36691
rect 119 36671 126 36681
rect 76 36655 92 36661
rect 94 36655 110 36661
rect 170 36655 172 36705
rect 186 36639 190 36673
rect 216 36639 220 36673
rect 213 36607 224 36639
rect 282 36635 292 36719
rect 296 36713 368 36721
rect 378 36713 450 36721
rect 468 36718 473 36752
rect 428 36683 430 36699
rect 251 36607 292 36635
rect 318 36614 324 36683
rect 12 36602 62 36604
rect 28 36593 59 36601
rect 62 36593 64 36602
rect 251 36601 263 36607
rect 28 36585 64 36593
rect 127 36593 158 36601
rect 127 36586 182 36593
rect 127 36585 161 36586
rect 59 36569 64 36585
rect 158 36569 161 36585
rect 253 36573 263 36601
rect 273 36573 293 36607
rect 318 36604 335 36614
rect 303 36588 316 36598
rect 318 36588 324 36604
rect 346 36598 348 36683
rect 400 36675 430 36683
rect 476 36681 480 36749
rect 511 36718 582 36752
rect 544 36711 548 36718
rect 400 36671 436 36675
rect 400 36641 408 36671
rect 420 36641 436 36671
rect 544 36673 548 36681
rect 28 36561 64 36569
rect 127 36568 161 36569
rect 127 36561 182 36568
rect 62 36552 64 36561
rect 282 36515 292 36573
rect 295 36564 324 36588
rect 333 36588 353 36598
rect 428 36594 430 36641
rect 476 36601 480 36669
rect 544 36639 552 36673
rect 578 36639 582 36673
rect 544 36631 548 36639
rect 367 36588 380 36594
rect 333 36564 380 36588
rect 318 36551 324 36564
rect 346 36551 348 36564
rect 367 36560 380 36564
rect 396 36560 408 36594
rect 420 36560 436 36594
rect 544 36591 553 36619
rect 319 36540 346 36551
rect 120 36499 170 36501
rect 76 36493 92 36499
rect 94 36493 110 36499
rect 76 36483 99 36492
rect 60 36473 67 36483
rect 76 36463 77 36483
rect 96 36458 99 36483
rect 109 36463 110 36483
rect 119 36473 126 36483
rect 76 36449 110 36453
rect 170 36449 172 36499
rect 186 36481 190 36515
rect 216 36481 220 36515
rect 182 36443 224 36444
rect 186 36419 220 36436
rect 223 36419 257 36436
rect 182 36402 257 36419
rect 182 36401 224 36402
rect 160 36395 246 36401
rect 288 36395 292 36515
rect 296 36513 368 36521
rect 428 36513 430 36560
rect 476 36523 480 36591
rect 485 36547 495 36581
rect 505 36553 525 36581
rect 505 36547 519 36553
rect 544 36547 555 36591
rect 485 36523 492 36547
rect 579 36532 582 36622
rect 612 36604 624 36605
rect 599 36602 649 36604
rect 612 36601 624 36602
rect 610 36594 632 36601
rect 607 36593 632 36594
rect 586 36586 644 36593
rect 607 36585 644 36586
rect 607 36569 610 36585
rect 616 36569 644 36585
rect 607 36568 644 36569
rect 586 36561 644 36568
rect 607 36560 610 36561
rect 612 36553 632 36561
rect 612 36549 624 36553
rect 649 36552 651 36602
rect 544 36515 548 36523
rect 400 36483 408 36513
rect 420 36483 436 36513
rect 400 36479 436 36483
rect 400 36471 430 36479
rect 428 36455 430 36471
rect 476 36443 480 36511
rect 544 36481 552 36515
rect 578 36481 582 36515
rect 544 36473 548 36481
rect 295 36402 300 36436
rect 324 36402 329 36436
rect 378 36433 450 36441
rect 544 36438 548 36443
rect 544 36434 582 36438
rect 544 36419 552 36434
rect 578 36419 582 36434
rect 544 36401 586 36419
rect 522 36395 608 36401
rect 182 36379 224 36395
rect 544 36379 586 36395
rect 17 36365 67 36367
rect 119 36365 169 36367
rect 186 36365 220 36379
rect 548 36365 582 36379
rect 599 36365 649 36367
rect 42 36323 59 36357
rect 67 36315 69 36365
rect 160 36357 246 36365
rect 522 36357 608 36365
rect 76 36323 110 36357
rect 127 36323 144 36357
rect 152 36323 161 36357
rect 162 36355 195 36357
rect 224 36355 244 36357
rect 162 36323 244 36355
rect 524 36355 548 36357
rect 573 36355 582 36357
rect 586 36355 606 36357
rect 160 36315 246 36323
rect 186 36299 220 36315
rect 182 36285 224 36286
rect 160 36279 182 36285
rect 224 36279 246 36285
rect 186 36244 220 36278
rect 223 36244 257 36278
rect 120 36231 170 36233
rect 76 36227 130 36231
rect 110 36222 130 36227
rect 60 36197 67 36207
rect 76 36197 77 36217
rect 96 36188 99 36222
rect 109 36197 110 36217
rect 119 36197 126 36207
rect 76 36181 92 36187
rect 94 36181 110 36187
rect 170 36181 172 36231
rect 186 36165 190 36199
rect 216 36165 220 36199
rect 288 36165 292 36353
rect 476 36285 480 36353
rect 524 36323 606 36355
rect 607 36323 616 36357
rect 522 36315 608 36323
rect 649 36315 651 36365
rect 548 36299 582 36315
rect 522 36280 548 36285
rect 522 36279 582 36280
rect 586 36279 608 36285
rect 295 36244 300 36278
rect 324 36244 329 36278
rect 544 36276 582 36279
rect 378 36239 450 36247
rect 428 36209 430 36225
rect 400 36201 430 36209
rect 476 36207 480 36275
rect 544 36246 552 36276
rect 578 36246 582 36276
rect 544 36237 548 36246
rect 400 36197 436 36201
rect 400 36167 408 36197
rect 420 36167 436 36197
rect 544 36199 548 36207
rect 12 36128 62 36130
rect 28 36119 59 36127
rect 62 36119 64 36128
rect 28 36111 64 36119
rect 127 36119 158 36127
rect 127 36112 182 36119
rect 215 36117 224 36145
rect 127 36111 161 36112
rect 59 36095 64 36111
rect 158 36095 161 36111
rect 28 36087 64 36095
rect 127 36094 161 36095
rect 127 36087 182 36094
rect 62 36078 64 36087
rect 213 36079 224 36117
rect 282 36107 292 36165
rect 296 36159 368 36167
rect 319 36129 346 36140
rect 318 36116 324 36129
rect 346 36116 348 36129
rect 428 36120 430 36167
rect 443 36157 450 36159
rect 476 36127 480 36195
rect 544 36165 552 36199
rect 578 36165 582 36199
rect 481 36133 517 36161
rect 481 36127 495 36133
rect 367 36116 380 36120
rect 251 36073 263 36107
rect 273 36073 293 36107
rect 295 36092 324 36116
rect 303 36082 316 36092
rect 318 36076 324 36092
rect 333 36092 380 36116
rect 333 36082 353 36092
rect 367 36086 380 36092
rect 396 36086 408 36120
rect 420 36086 436 36120
rect 120 36025 170 36027
rect 76 36019 92 36025
rect 94 36019 110 36025
rect 76 36009 99 36018
rect 60 35999 67 36009
rect 76 35989 77 36009
rect 96 35984 99 36009
rect 109 35989 110 36009
rect 119 35999 126 36009
rect 76 35975 110 35979
rect 170 35975 172 36025
rect 186 36007 190 36041
rect 216 36007 220 36041
rect 186 35930 220 35964
rect 282 35961 292 36073
rect 318 36066 335 36076
rect 318 35997 324 36066
rect 346 35997 348 36082
rect 428 36039 430 36086
rect 476 36049 480 36117
rect 485 36099 495 36127
rect 505 36127 519 36133
rect 544 36127 555 36165
rect 505 36099 525 36127
rect 544 36099 553 36127
rect 544 36079 548 36099
rect 579 36058 582 36148
rect 612 36130 624 36131
rect 599 36128 649 36130
rect 612 36127 624 36128
rect 610 36120 632 36127
rect 607 36119 632 36120
rect 586 36112 644 36119
rect 607 36111 644 36112
rect 607 36095 610 36111
rect 616 36095 644 36111
rect 607 36094 644 36095
rect 586 36087 644 36094
rect 607 36086 610 36087
rect 612 36079 632 36087
rect 612 36075 624 36079
rect 649 36078 651 36128
rect 544 36041 548 36049
rect 400 36009 408 36039
rect 420 36009 436 36039
rect 400 36005 436 36009
rect 400 35997 430 36005
rect 428 35981 430 35997
rect 476 35969 480 36037
rect 544 36007 552 36041
rect 578 36007 582 36041
rect 544 35999 548 36007
rect 544 35969 586 35970
rect 288 35929 292 35961
rect 296 35959 368 35967
rect 378 35959 450 35967
rect 544 35962 548 35969
rect 439 35931 444 35959
rect 120 35915 170 35917
rect 76 35911 130 35915
rect 110 35906 130 35911
rect 60 35881 67 35891
rect 76 35881 77 35901
rect 96 35872 99 35906
rect 109 35881 110 35901
rect 119 35881 126 35891
rect 76 35865 92 35871
rect 94 35865 110 35871
rect 170 35865 172 35915
rect 186 35849 190 35883
rect 216 35849 220 35883
rect 213 35817 224 35849
rect 282 35845 292 35929
rect 296 35923 368 35931
rect 378 35923 450 35931
rect 468 35928 473 35962
rect 428 35893 430 35909
rect 251 35817 292 35845
rect 318 35824 324 35893
rect 12 35812 62 35814
rect 28 35803 59 35811
rect 62 35803 64 35812
rect 251 35811 263 35817
rect 28 35795 64 35803
rect 127 35803 158 35811
rect 127 35796 182 35803
rect 127 35795 161 35796
rect 59 35779 64 35795
rect 158 35779 161 35795
rect 253 35783 263 35811
rect 273 35783 293 35817
rect 318 35814 335 35824
rect 303 35798 316 35808
rect 318 35798 324 35814
rect 346 35808 348 35893
rect 400 35885 430 35893
rect 476 35891 480 35959
rect 511 35928 582 35962
rect 544 35921 548 35928
rect 400 35881 436 35885
rect 400 35851 408 35881
rect 420 35851 436 35881
rect 544 35883 548 35891
rect 28 35771 64 35779
rect 127 35778 161 35779
rect 127 35771 182 35778
rect 62 35762 64 35771
rect 282 35725 292 35783
rect 295 35774 324 35798
rect 333 35798 353 35808
rect 428 35804 430 35851
rect 476 35811 480 35879
rect 544 35849 552 35883
rect 578 35849 582 35883
rect 544 35841 548 35849
rect 367 35798 380 35804
rect 333 35774 380 35798
rect 318 35761 324 35774
rect 346 35761 348 35774
rect 367 35770 380 35774
rect 396 35770 408 35804
rect 420 35770 436 35804
rect 544 35801 553 35829
rect 319 35750 346 35761
rect 120 35709 170 35711
rect 76 35703 92 35709
rect 94 35703 110 35709
rect 76 35693 99 35702
rect 60 35683 67 35693
rect 76 35673 77 35693
rect 96 35668 99 35693
rect 109 35673 110 35693
rect 119 35683 126 35693
rect 76 35659 110 35663
rect 170 35659 172 35709
rect 186 35691 190 35725
rect 216 35691 220 35725
rect 182 35653 224 35654
rect 186 35629 220 35646
rect 223 35629 257 35646
rect 182 35612 257 35629
rect 182 35611 224 35612
rect 160 35605 246 35611
rect 288 35605 292 35725
rect 296 35723 368 35731
rect 428 35723 430 35770
rect 476 35733 480 35801
rect 485 35757 495 35791
rect 505 35763 525 35791
rect 505 35757 519 35763
rect 544 35757 555 35801
rect 485 35733 492 35757
rect 579 35742 582 35832
rect 612 35814 624 35815
rect 599 35812 649 35814
rect 612 35811 624 35812
rect 610 35804 632 35811
rect 607 35803 632 35804
rect 586 35796 644 35803
rect 607 35795 644 35796
rect 607 35779 610 35795
rect 616 35779 644 35795
rect 607 35778 644 35779
rect 586 35771 644 35778
rect 607 35770 610 35771
rect 612 35763 632 35771
rect 612 35759 624 35763
rect 649 35762 651 35812
rect 544 35725 548 35733
rect 400 35693 408 35723
rect 420 35693 436 35723
rect 400 35689 436 35693
rect 400 35681 430 35689
rect 428 35665 430 35681
rect 476 35653 480 35721
rect 544 35691 552 35725
rect 578 35691 582 35725
rect 544 35683 548 35691
rect 295 35612 300 35646
rect 324 35612 329 35646
rect 378 35643 450 35651
rect 544 35648 548 35653
rect 544 35644 582 35648
rect 544 35629 552 35644
rect 578 35629 582 35644
rect 544 35611 586 35629
rect 522 35605 608 35611
rect 182 35589 224 35605
rect 544 35589 586 35605
rect 17 35575 67 35577
rect 119 35575 169 35577
rect 186 35575 220 35589
rect 548 35575 582 35589
rect 599 35575 649 35577
rect 42 35533 59 35567
rect 67 35525 69 35575
rect 160 35567 246 35575
rect 522 35567 608 35575
rect 76 35533 110 35567
rect 127 35533 144 35567
rect 152 35533 161 35567
rect 162 35565 195 35567
rect 224 35565 244 35567
rect 162 35533 244 35565
rect 524 35565 548 35567
rect 573 35565 582 35567
rect 586 35565 606 35567
rect 160 35525 246 35533
rect 186 35509 220 35525
rect 182 35495 224 35496
rect 160 35489 182 35495
rect 224 35489 246 35495
rect 186 35454 220 35488
rect 223 35454 257 35488
rect 120 35441 170 35443
rect 76 35437 130 35441
rect 110 35432 130 35437
rect 60 35407 67 35417
rect 76 35407 77 35427
rect 96 35398 99 35432
rect 109 35407 110 35427
rect 119 35407 126 35417
rect 76 35391 92 35397
rect 94 35391 110 35397
rect 170 35391 172 35441
rect 186 35375 190 35409
rect 216 35375 220 35409
rect 288 35375 292 35563
rect 476 35495 480 35563
rect 524 35533 606 35565
rect 607 35533 616 35567
rect 522 35525 608 35533
rect 649 35525 651 35575
rect 548 35509 582 35525
rect 522 35490 548 35495
rect 522 35489 582 35490
rect 586 35489 608 35495
rect 295 35454 300 35488
rect 324 35454 329 35488
rect 544 35486 582 35489
rect 378 35449 450 35457
rect 428 35419 430 35435
rect 400 35411 430 35419
rect 476 35417 480 35485
rect 544 35456 552 35486
rect 578 35456 582 35486
rect 544 35447 548 35456
rect 400 35407 436 35411
rect 400 35377 408 35407
rect 420 35377 436 35407
rect 544 35409 548 35417
rect 12 35338 62 35340
rect 28 35329 59 35337
rect 62 35329 64 35338
rect 28 35321 64 35329
rect 127 35329 158 35337
rect 127 35322 182 35329
rect 215 35327 224 35355
rect 127 35321 161 35322
rect 59 35305 64 35321
rect 158 35305 161 35321
rect 28 35297 64 35305
rect 127 35304 161 35305
rect 127 35297 182 35304
rect 62 35288 64 35297
rect 213 35289 224 35327
rect 282 35317 292 35375
rect 296 35369 368 35377
rect 319 35339 346 35350
rect 318 35326 324 35339
rect 346 35326 348 35339
rect 428 35330 430 35377
rect 443 35367 450 35369
rect 476 35337 480 35405
rect 544 35375 552 35409
rect 578 35375 582 35409
rect 481 35343 517 35371
rect 481 35337 495 35343
rect 367 35326 380 35330
rect 251 35283 263 35317
rect 273 35283 293 35317
rect 295 35302 324 35326
rect 303 35292 316 35302
rect 318 35286 324 35302
rect 333 35302 380 35326
rect 333 35292 353 35302
rect 367 35296 380 35302
rect 396 35296 408 35330
rect 420 35296 436 35330
rect 120 35235 170 35237
rect 76 35229 92 35235
rect 94 35229 110 35235
rect 76 35219 99 35228
rect 60 35209 67 35219
rect 76 35199 77 35219
rect 96 35194 99 35219
rect 109 35199 110 35219
rect 119 35209 126 35219
rect 76 35185 110 35189
rect 170 35185 172 35235
rect 186 35217 190 35251
rect 216 35217 220 35251
rect 186 35140 220 35174
rect 282 35171 292 35283
rect 318 35276 335 35286
rect 318 35207 324 35276
rect 346 35207 348 35292
rect 428 35249 430 35296
rect 476 35259 480 35327
rect 485 35309 495 35337
rect 505 35337 519 35343
rect 544 35337 555 35375
rect 505 35309 525 35337
rect 544 35309 553 35337
rect 544 35289 548 35309
rect 579 35268 582 35358
rect 612 35340 624 35341
rect 599 35338 649 35340
rect 612 35337 624 35338
rect 610 35330 632 35337
rect 607 35329 632 35330
rect 586 35322 644 35329
rect 607 35321 644 35322
rect 607 35305 610 35321
rect 616 35305 644 35321
rect 607 35304 644 35305
rect 586 35297 644 35304
rect 607 35296 610 35297
rect 612 35289 632 35297
rect 612 35285 624 35289
rect 649 35288 651 35338
rect 544 35251 548 35259
rect 400 35219 408 35249
rect 420 35219 436 35249
rect 400 35215 436 35219
rect 400 35207 430 35215
rect 428 35191 430 35207
rect 476 35179 480 35247
rect 544 35217 552 35251
rect 578 35217 582 35251
rect 544 35209 548 35217
rect 544 35179 586 35180
rect 288 35139 292 35171
rect 296 35169 368 35177
rect 378 35169 450 35177
rect 544 35172 548 35179
rect 439 35141 444 35169
rect 120 35125 170 35127
rect 76 35121 130 35125
rect 110 35116 130 35121
rect 60 35091 67 35101
rect 76 35091 77 35111
rect 96 35082 99 35116
rect 109 35091 110 35111
rect 119 35091 126 35101
rect 76 35075 92 35081
rect 94 35075 110 35081
rect 170 35075 172 35125
rect 186 35059 190 35093
rect 216 35059 220 35093
rect 213 35027 224 35059
rect 282 35055 292 35139
rect 296 35133 368 35141
rect 378 35133 450 35141
rect 468 35138 473 35172
rect 428 35103 430 35119
rect 251 35027 292 35055
rect 318 35034 324 35103
rect 12 35022 62 35024
rect 28 35013 59 35021
rect 62 35013 64 35022
rect 251 35021 263 35027
rect 28 35005 64 35013
rect 127 35013 158 35021
rect 127 35006 182 35013
rect 127 35005 161 35006
rect 59 34989 64 35005
rect 158 34989 161 35005
rect 253 34993 263 35021
rect 273 34993 293 35027
rect 318 35024 335 35034
rect 303 35008 316 35018
rect 318 35008 324 35024
rect 346 35018 348 35103
rect 400 35095 430 35103
rect 476 35101 480 35169
rect 511 35138 582 35172
rect 544 35131 548 35138
rect 400 35091 436 35095
rect 400 35061 408 35091
rect 420 35061 436 35091
rect 544 35093 548 35101
rect 28 34981 64 34989
rect 127 34988 161 34989
rect 127 34981 182 34988
rect 62 34972 64 34981
rect 282 34935 292 34993
rect 295 34984 324 35008
rect 333 35008 353 35018
rect 428 35014 430 35061
rect 476 35021 480 35089
rect 544 35059 552 35093
rect 578 35059 582 35093
rect 544 35051 548 35059
rect 367 35008 380 35014
rect 333 34984 380 35008
rect 318 34971 324 34984
rect 346 34971 348 34984
rect 367 34980 380 34984
rect 396 34980 408 35014
rect 420 34980 436 35014
rect 544 35011 553 35039
rect 319 34960 346 34971
rect 120 34919 170 34921
rect 76 34913 92 34919
rect 94 34913 110 34919
rect 76 34903 99 34912
rect 60 34893 67 34903
rect 76 34883 77 34903
rect 96 34878 99 34903
rect 109 34883 110 34903
rect 119 34893 126 34903
rect 76 34869 110 34873
rect 170 34869 172 34919
rect 186 34901 190 34935
rect 216 34901 220 34935
rect 182 34863 224 34864
rect 186 34839 220 34856
rect 223 34839 257 34856
rect 182 34822 257 34839
rect 182 34821 224 34822
rect 160 34815 246 34821
rect 288 34815 292 34935
rect 296 34933 368 34941
rect 428 34933 430 34980
rect 476 34943 480 35011
rect 485 34967 495 35001
rect 505 34973 525 35001
rect 505 34967 519 34973
rect 544 34967 555 35011
rect 485 34943 492 34967
rect 579 34952 582 35042
rect 612 35024 624 35025
rect 599 35022 649 35024
rect 612 35021 624 35022
rect 610 35014 632 35021
rect 607 35013 632 35014
rect 586 35006 644 35013
rect 607 35005 644 35006
rect 607 34989 610 35005
rect 616 34989 644 35005
rect 607 34988 644 34989
rect 586 34981 644 34988
rect 607 34980 610 34981
rect 612 34973 632 34981
rect 612 34969 624 34973
rect 649 34972 651 35022
rect 544 34935 548 34943
rect 400 34903 408 34933
rect 420 34903 436 34933
rect 400 34899 436 34903
rect 400 34891 430 34899
rect 428 34875 430 34891
rect 476 34863 480 34931
rect 544 34901 552 34935
rect 578 34901 582 34935
rect 544 34893 548 34901
rect 295 34822 300 34856
rect 324 34822 329 34856
rect 378 34853 450 34861
rect 544 34858 548 34863
rect 544 34854 582 34858
rect 544 34839 552 34854
rect 578 34839 582 34854
rect 544 34821 586 34839
rect 522 34815 608 34821
rect 182 34799 224 34815
rect 544 34799 586 34815
rect 17 34785 67 34787
rect 119 34785 169 34787
rect 186 34785 220 34799
rect 548 34785 582 34799
rect 599 34785 649 34787
rect 42 34743 59 34777
rect 67 34735 69 34785
rect 160 34777 246 34785
rect 522 34777 608 34785
rect 76 34743 110 34777
rect 127 34743 144 34777
rect 152 34743 161 34777
rect 162 34775 195 34777
rect 224 34775 244 34777
rect 162 34743 244 34775
rect 524 34775 548 34777
rect 573 34775 582 34777
rect 586 34775 606 34777
rect 160 34735 246 34743
rect 186 34719 220 34735
rect 182 34705 224 34706
rect 160 34699 182 34705
rect 224 34699 246 34705
rect 186 34664 220 34698
rect 223 34664 257 34698
rect 120 34651 170 34653
rect 76 34647 130 34651
rect 110 34642 130 34647
rect 60 34617 67 34627
rect 76 34617 77 34637
rect 96 34608 99 34642
rect 109 34617 110 34637
rect 119 34617 126 34627
rect 76 34601 92 34607
rect 94 34601 110 34607
rect 170 34601 172 34651
rect 186 34585 190 34619
rect 216 34585 220 34619
rect 288 34585 292 34773
rect 476 34705 480 34773
rect 524 34743 606 34775
rect 607 34743 616 34777
rect 522 34735 608 34743
rect 649 34735 651 34785
rect 548 34719 582 34735
rect 522 34700 548 34705
rect 522 34699 582 34700
rect 586 34699 608 34705
rect 295 34664 300 34698
rect 324 34664 329 34698
rect 544 34696 582 34699
rect 378 34659 450 34667
rect 428 34629 430 34645
rect 400 34621 430 34629
rect 476 34627 480 34695
rect 544 34666 552 34696
rect 578 34666 582 34696
rect 544 34657 548 34666
rect 400 34617 436 34621
rect 400 34587 408 34617
rect 420 34587 436 34617
rect 544 34619 548 34627
rect 12 34548 62 34550
rect 28 34539 59 34547
rect 62 34539 64 34548
rect 28 34531 64 34539
rect 127 34539 158 34547
rect 127 34532 182 34539
rect 215 34537 224 34565
rect 127 34531 161 34532
rect 59 34515 64 34531
rect 158 34515 161 34531
rect 28 34507 64 34515
rect 127 34514 161 34515
rect 127 34507 182 34514
rect 62 34498 64 34507
rect 213 34499 224 34537
rect 282 34527 292 34585
rect 296 34579 368 34587
rect 319 34549 346 34560
rect 318 34536 324 34549
rect 346 34536 348 34549
rect 428 34540 430 34587
rect 443 34577 450 34579
rect 476 34547 480 34615
rect 544 34585 552 34619
rect 578 34585 582 34619
rect 481 34553 517 34581
rect 481 34547 495 34553
rect 367 34536 380 34540
rect 251 34493 263 34527
rect 273 34493 293 34527
rect 295 34512 324 34536
rect 303 34502 316 34512
rect 318 34496 324 34512
rect 333 34512 380 34536
rect 333 34502 353 34512
rect 367 34506 380 34512
rect 396 34506 408 34540
rect 420 34506 436 34540
rect 120 34445 170 34447
rect 76 34439 92 34445
rect 94 34439 110 34445
rect 76 34429 99 34438
rect 60 34419 67 34429
rect 76 34409 77 34429
rect 96 34404 99 34429
rect 109 34409 110 34429
rect 119 34419 126 34429
rect 76 34395 110 34399
rect 170 34395 172 34445
rect 186 34427 190 34461
rect 216 34427 220 34461
rect 186 34350 220 34384
rect 282 34381 292 34493
rect 318 34486 335 34496
rect 318 34417 324 34486
rect 346 34417 348 34502
rect 428 34459 430 34506
rect 476 34469 480 34537
rect 485 34519 495 34547
rect 505 34547 519 34553
rect 544 34547 555 34585
rect 505 34519 525 34547
rect 544 34519 553 34547
rect 544 34499 548 34519
rect 579 34478 582 34568
rect 612 34550 624 34551
rect 599 34548 649 34550
rect 612 34547 624 34548
rect 610 34540 632 34547
rect 607 34539 632 34540
rect 586 34532 644 34539
rect 607 34531 644 34532
rect 607 34515 610 34531
rect 616 34515 644 34531
rect 607 34514 644 34515
rect 586 34507 644 34514
rect 607 34506 610 34507
rect 612 34499 632 34507
rect 612 34495 624 34499
rect 649 34498 651 34548
rect 544 34461 548 34469
rect 400 34429 408 34459
rect 420 34429 436 34459
rect 400 34425 436 34429
rect 400 34417 430 34425
rect 428 34401 430 34417
rect 476 34389 480 34457
rect 544 34427 552 34461
rect 578 34427 582 34461
rect 544 34419 548 34427
rect 544 34389 586 34390
rect 288 34349 292 34381
rect 296 34379 368 34387
rect 378 34379 450 34387
rect 544 34382 548 34389
rect 439 34351 444 34379
rect 120 34335 170 34337
rect 76 34331 130 34335
rect 110 34326 130 34331
rect 60 34301 67 34311
rect 76 34301 77 34321
rect 96 34292 99 34326
rect 109 34301 110 34321
rect 119 34301 126 34311
rect 76 34285 92 34291
rect 94 34285 110 34291
rect 170 34285 172 34335
rect 186 34269 190 34303
rect 216 34269 220 34303
rect 213 34237 224 34269
rect 282 34265 292 34349
rect 296 34343 368 34351
rect 378 34343 450 34351
rect 468 34348 473 34382
rect 428 34313 430 34329
rect 251 34237 292 34265
rect 318 34244 324 34313
rect 12 34232 62 34234
rect 28 34223 59 34231
rect 62 34223 64 34232
rect 251 34231 263 34237
rect 28 34215 64 34223
rect 127 34223 158 34231
rect 127 34216 182 34223
rect 127 34215 161 34216
rect 59 34199 64 34215
rect 158 34199 161 34215
rect 253 34203 263 34231
rect 273 34203 293 34237
rect 318 34234 335 34244
rect 303 34218 316 34228
rect 318 34218 324 34234
rect 346 34228 348 34313
rect 400 34305 430 34313
rect 476 34311 480 34379
rect 511 34348 582 34382
rect 544 34341 548 34348
rect 400 34301 436 34305
rect 400 34271 408 34301
rect 420 34271 436 34301
rect 544 34303 548 34311
rect 28 34191 64 34199
rect 127 34198 161 34199
rect 127 34191 182 34198
rect 62 34182 64 34191
rect 282 34145 292 34203
rect 295 34194 324 34218
rect 333 34218 353 34228
rect 428 34224 430 34271
rect 476 34231 480 34299
rect 544 34269 552 34303
rect 578 34269 582 34303
rect 544 34261 548 34269
rect 367 34218 380 34224
rect 333 34194 380 34218
rect 318 34181 324 34194
rect 346 34181 348 34194
rect 367 34190 380 34194
rect 396 34190 408 34224
rect 420 34190 436 34224
rect 544 34221 553 34249
rect 319 34170 346 34181
rect 120 34129 170 34131
rect 76 34123 92 34129
rect 94 34123 110 34129
rect 76 34113 99 34122
rect 60 34103 67 34113
rect 76 34093 77 34113
rect 96 34088 99 34113
rect 109 34093 110 34113
rect 119 34103 126 34113
rect 76 34079 110 34083
rect 170 34079 172 34129
rect 186 34111 190 34145
rect 216 34111 220 34145
rect 182 34073 224 34074
rect 186 34049 220 34066
rect 223 34049 257 34066
rect 182 34032 257 34049
rect 182 34031 224 34032
rect 160 34025 246 34031
rect 288 34025 292 34145
rect 296 34143 368 34151
rect 428 34143 430 34190
rect 476 34153 480 34221
rect 485 34177 495 34211
rect 505 34183 525 34211
rect 505 34177 519 34183
rect 544 34177 555 34221
rect 485 34153 492 34177
rect 579 34162 582 34252
rect 612 34234 624 34235
rect 599 34232 649 34234
rect 612 34231 624 34232
rect 610 34224 632 34231
rect 607 34223 632 34224
rect 586 34216 644 34223
rect 607 34215 644 34216
rect 607 34199 610 34215
rect 616 34199 644 34215
rect 607 34198 644 34199
rect 586 34191 644 34198
rect 607 34190 610 34191
rect 612 34183 632 34191
rect 612 34179 624 34183
rect 649 34182 651 34232
rect 544 34145 548 34153
rect 400 34113 408 34143
rect 420 34113 436 34143
rect 400 34109 436 34113
rect 400 34101 430 34109
rect 428 34085 430 34101
rect 476 34073 480 34141
rect 544 34111 552 34145
rect 578 34111 582 34145
rect 544 34103 548 34111
rect 295 34032 300 34066
rect 324 34032 329 34066
rect 378 34063 450 34071
rect 544 34068 548 34073
rect 544 34064 582 34068
rect 544 34049 552 34064
rect 578 34049 582 34064
rect 544 34031 586 34049
rect 522 34025 608 34031
rect 182 34009 224 34025
rect 544 34009 586 34025
rect 17 33995 67 33997
rect 119 33995 169 33997
rect 186 33995 220 34009
rect 548 33995 582 34009
rect 599 33995 649 33997
rect 42 33953 59 33987
rect 67 33945 69 33995
rect 160 33987 246 33995
rect 522 33987 608 33995
rect 76 33953 110 33987
rect 127 33953 144 33987
rect 152 33953 161 33987
rect 162 33985 195 33987
rect 224 33985 244 33987
rect 162 33953 244 33985
rect 524 33985 548 33987
rect 573 33985 582 33987
rect 586 33985 606 33987
rect 160 33945 246 33953
rect 186 33929 220 33945
rect 182 33915 224 33916
rect 160 33909 182 33915
rect 224 33909 246 33915
rect 186 33874 220 33908
rect 223 33874 257 33908
rect 120 33861 170 33863
rect 76 33857 130 33861
rect 110 33852 130 33857
rect 60 33827 67 33837
rect 76 33827 77 33847
rect 96 33818 99 33852
rect 109 33827 110 33847
rect 119 33827 126 33837
rect 76 33811 92 33817
rect 94 33811 110 33817
rect 170 33811 172 33861
rect 186 33795 190 33829
rect 216 33795 220 33829
rect 288 33795 292 33983
rect 476 33915 480 33983
rect 524 33953 606 33985
rect 607 33953 616 33987
rect 522 33945 608 33953
rect 649 33945 651 33995
rect 548 33929 582 33945
rect 522 33910 548 33915
rect 522 33909 582 33910
rect 586 33909 608 33915
rect 295 33874 300 33908
rect 324 33874 329 33908
rect 544 33906 582 33909
rect 378 33869 450 33877
rect 428 33839 430 33855
rect 400 33831 430 33839
rect 476 33837 480 33905
rect 544 33876 552 33906
rect 578 33876 582 33906
rect 544 33867 548 33876
rect 400 33827 436 33831
rect 400 33797 408 33827
rect 420 33797 436 33827
rect 544 33829 548 33837
rect 12 33758 62 33760
rect 28 33749 59 33757
rect 62 33749 64 33758
rect 28 33741 64 33749
rect 127 33749 158 33757
rect 127 33742 182 33749
rect 215 33747 224 33775
rect 127 33741 161 33742
rect 59 33725 64 33741
rect 158 33725 161 33741
rect 28 33717 64 33725
rect 127 33724 161 33725
rect 127 33717 182 33724
rect 62 33708 64 33717
rect 213 33709 224 33747
rect 282 33737 292 33795
rect 296 33789 368 33797
rect 319 33759 346 33770
rect 318 33746 324 33759
rect 346 33746 348 33759
rect 428 33750 430 33797
rect 443 33787 450 33789
rect 476 33757 480 33825
rect 544 33795 552 33829
rect 578 33795 582 33829
rect 481 33763 517 33791
rect 481 33757 495 33763
rect 367 33746 380 33750
rect 251 33703 263 33737
rect 273 33703 293 33737
rect 295 33722 324 33746
rect 303 33712 316 33722
rect 318 33706 324 33722
rect 333 33722 380 33746
rect 333 33712 353 33722
rect 367 33716 380 33722
rect 396 33716 408 33750
rect 420 33716 436 33750
rect 120 33655 170 33657
rect 76 33649 92 33655
rect 94 33649 110 33655
rect 76 33639 99 33648
rect 60 33629 67 33639
rect 76 33619 77 33639
rect 96 33614 99 33639
rect 109 33619 110 33639
rect 119 33629 126 33639
rect 76 33605 110 33609
rect 170 33605 172 33655
rect 186 33637 190 33671
rect 216 33637 220 33671
rect 186 33560 220 33594
rect 282 33591 292 33703
rect 318 33696 335 33706
rect 318 33627 324 33696
rect 346 33627 348 33712
rect 428 33669 430 33716
rect 476 33679 480 33747
rect 485 33729 495 33757
rect 505 33757 519 33763
rect 544 33757 555 33795
rect 505 33729 525 33757
rect 544 33729 553 33757
rect 544 33709 548 33729
rect 579 33688 582 33778
rect 612 33760 624 33761
rect 599 33758 649 33760
rect 612 33757 624 33758
rect 610 33750 632 33757
rect 607 33749 632 33750
rect 586 33742 644 33749
rect 607 33741 644 33742
rect 607 33725 610 33741
rect 616 33725 644 33741
rect 607 33724 644 33725
rect 586 33717 644 33724
rect 607 33716 610 33717
rect 612 33709 632 33717
rect 612 33705 624 33709
rect 649 33708 651 33758
rect 544 33671 548 33679
rect 400 33639 408 33669
rect 420 33639 436 33669
rect 400 33635 436 33639
rect 400 33627 430 33635
rect 428 33611 430 33627
rect 476 33599 480 33667
rect 544 33637 552 33671
rect 578 33637 582 33671
rect 544 33629 548 33637
rect 544 33599 586 33600
rect 288 33559 292 33591
rect 296 33589 368 33597
rect 378 33589 450 33597
rect 544 33592 548 33599
rect 439 33561 444 33589
rect 120 33545 170 33547
rect 76 33541 130 33545
rect 110 33536 130 33541
rect 60 33511 67 33521
rect 76 33511 77 33531
rect 96 33502 99 33536
rect 109 33511 110 33531
rect 119 33511 126 33521
rect 76 33495 92 33501
rect 94 33495 110 33501
rect 170 33495 172 33545
rect 186 33479 190 33513
rect 216 33479 220 33513
rect 213 33447 224 33479
rect 282 33475 292 33559
rect 296 33553 368 33561
rect 378 33553 450 33561
rect 468 33558 473 33592
rect 428 33523 430 33539
rect 251 33447 292 33475
rect 318 33454 324 33523
rect 12 33442 62 33444
rect 28 33433 59 33441
rect 62 33433 64 33442
rect 251 33441 263 33447
rect 28 33425 64 33433
rect 127 33433 158 33441
rect 127 33426 182 33433
rect 127 33425 161 33426
rect 59 33409 64 33425
rect 158 33409 161 33425
rect 253 33413 263 33441
rect 273 33413 293 33447
rect 318 33444 335 33454
rect 303 33428 316 33438
rect 318 33428 324 33444
rect 346 33438 348 33523
rect 400 33515 430 33523
rect 476 33521 480 33589
rect 511 33558 582 33592
rect 544 33551 548 33558
rect 400 33511 436 33515
rect 400 33481 408 33511
rect 420 33481 436 33511
rect 544 33513 548 33521
rect 28 33401 64 33409
rect 127 33408 161 33409
rect 127 33401 182 33408
rect 62 33392 64 33401
rect 282 33355 292 33413
rect 295 33404 324 33428
rect 333 33428 353 33438
rect 428 33434 430 33481
rect 476 33441 480 33509
rect 544 33479 552 33513
rect 578 33479 582 33513
rect 544 33471 548 33479
rect 367 33428 380 33434
rect 333 33404 380 33428
rect 318 33391 324 33404
rect 346 33391 348 33404
rect 367 33400 380 33404
rect 396 33400 408 33434
rect 420 33400 436 33434
rect 544 33431 553 33459
rect 319 33380 346 33391
rect 120 33339 170 33341
rect 76 33333 92 33339
rect 94 33333 110 33339
rect 76 33323 99 33332
rect 60 33313 67 33323
rect 76 33303 77 33323
rect 96 33298 99 33323
rect 109 33303 110 33323
rect 119 33313 126 33323
rect 76 33289 110 33293
rect 170 33289 172 33339
rect 186 33321 190 33355
rect 216 33321 220 33355
rect 182 33283 224 33284
rect 186 33259 220 33276
rect 223 33259 257 33276
rect 182 33242 257 33259
rect 182 33241 224 33242
rect 160 33235 246 33241
rect 288 33235 292 33355
rect 296 33353 368 33361
rect 428 33353 430 33400
rect 476 33363 480 33431
rect 485 33387 495 33421
rect 505 33393 525 33421
rect 505 33387 519 33393
rect 544 33387 555 33431
rect 485 33363 492 33387
rect 579 33372 582 33462
rect 612 33444 624 33445
rect 599 33442 649 33444
rect 612 33441 624 33442
rect 610 33434 632 33441
rect 607 33433 632 33434
rect 586 33426 644 33433
rect 607 33425 644 33426
rect 607 33409 610 33425
rect 616 33409 644 33425
rect 607 33408 644 33409
rect 586 33401 644 33408
rect 607 33400 610 33401
rect 612 33393 632 33401
rect 612 33389 624 33393
rect 649 33392 651 33442
rect 544 33355 548 33363
rect 400 33323 408 33353
rect 420 33323 436 33353
rect 400 33319 436 33323
rect 400 33311 430 33319
rect 428 33295 430 33311
rect 476 33283 480 33351
rect 544 33321 552 33355
rect 578 33321 582 33355
rect 544 33313 548 33321
rect 295 33242 300 33276
rect 324 33242 329 33276
rect 378 33273 450 33281
rect 544 33278 548 33283
rect 544 33274 582 33278
rect 544 33259 552 33274
rect 578 33259 582 33274
rect 544 33241 586 33259
rect 522 33235 608 33241
rect 182 33219 224 33235
rect 544 33219 586 33235
rect 17 33205 67 33207
rect 119 33205 169 33207
rect 186 33205 220 33219
rect 548 33205 582 33219
rect 599 33205 649 33207
rect 42 33163 59 33197
rect 67 33155 69 33205
rect 160 33197 246 33205
rect 522 33197 608 33205
rect 76 33163 110 33197
rect 127 33163 144 33197
rect 152 33163 161 33197
rect 162 33195 195 33197
rect 224 33195 244 33197
rect 162 33163 244 33195
rect 524 33195 548 33197
rect 573 33195 582 33197
rect 586 33195 606 33197
rect 160 33155 246 33163
rect 186 33139 220 33155
rect 182 33125 224 33126
rect 160 33119 182 33125
rect 224 33119 246 33125
rect 186 33084 220 33118
rect 223 33084 257 33118
rect 120 33071 170 33073
rect 76 33067 130 33071
rect 110 33062 130 33067
rect 60 33037 67 33047
rect 76 33037 77 33057
rect 96 33028 99 33062
rect 109 33037 110 33057
rect 119 33037 126 33047
rect 76 33021 92 33027
rect 94 33021 110 33027
rect 170 33021 172 33071
rect 186 33005 190 33039
rect 216 33005 220 33039
rect 288 33005 292 33193
rect 476 33125 480 33193
rect 524 33163 606 33195
rect 607 33163 616 33197
rect 522 33155 608 33163
rect 649 33155 651 33205
rect 548 33139 582 33155
rect 522 33120 548 33125
rect 522 33119 582 33120
rect 586 33119 608 33125
rect 295 33084 300 33118
rect 324 33084 329 33118
rect 544 33116 582 33119
rect 378 33079 450 33087
rect 428 33049 430 33065
rect 400 33041 430 33049
rect 476 33047 480 33115
rect 544 33086 552 33116
rect 578 33086 582 33116
rect 544 33077 548 33086
rect 400 33037 436 33041
rect 400 33007 408 33037
rect 420 33007 436 33037
rect 544 33039 548 33047
rect 12 32968 62 32970
rect 28 32959 59 32967
rect 62 32959 64 32968
rect 28 32951 64 32959
rect 127 32959 158 32967
rect 127 32952 182 32959
rect 215 32957 224 32985
rect 127 32951 161 32952
rect 59 32935 64 32951
rect 158 32935 161 32951
rect 28 32927 64 32935
rect 127 32934 161 32935
rect 127 32927 182 32934
rect 62 32918 64 32927
rect 213 32919 224 32957
rect 282 32947 292 33005
rect 296 32999 368 33007
rect 319 32969 346 32980
rect 318 32956 324 32969
rect 346 32956 348 32969
rect 428 32960 430 33007
rect 443 32997 450 32999
rect 476 32967 480 33035
rect 544 33005 552 33039
rect 578 33005 582 33039
rect 481 32973 517 33001
rect 481 32967 495 32973
rect 367 32956 380 32960
rect 251 32913 263 32947
rect 273 32913 293 32947
rect 295 32932 324 32956
rect 303 32922 316 32932
rect 318 32916 324 32932
rect 333 32932 380 32956
rect 333 32922 353 32932
rect 367 32926 380 32932
rect 396 32926 408 32960
rect 420 32926 436 32960
rect 120 32865 170 32867
rect 76 32859 92 32865
rect 94 32859 110 32865
rect 76 32849 99 32858
rect 60 32839 67 32849
rect 76 32829 77 32849
rect 96 32824 99 32849
rect 109 32829 110 32849
rect 119 32839 126 32849
rect 76 32815 110 32819
rect 170 32815 172 32865
rect 186 32847 190 32881
rect 216 32847 220 32881
rect 186 32770 220 32804
rect 282 32801 292 32913
rect 318 32906 335 32916
rect 318 32837 324 32906
rect 346 32837 348 32922
rect 428 32879 430 32926
rect 476 32889 480 32957
rect 485 32939 495 32967
rect 505 32967 519 32973
rect 544 32967 555 33005
rect 505 32939 525 32967
rect 544 32939 553 32967
rect 544 32919 548 32939
rect 579 32898 582 32988
rect 612 32970 624 32971
rect 599 32968 649 32970
rect 612 32967 624 32968
rect 610 32960 632 32967
rect 607 32959 632 32960
rect 586 32952 644 32959
rect 607 32951 644 32952
rect 607 32935 610 32951
rect 616 32935 644 32951
rect 607 32934 644 32935
rect 586 32927 644 32934
rect 607 32926 610 32927
rect 612 32919 632 32927
rect 612 32915 624 32919
rect 649 32918 651 32968
rect 544 32881 548 32889
rect 400 32849 408 32879
rect 420 32849 436 32879
rect 400 32845 436 32849
rect 400 32837 430 32845
rect 428 32821 430 32837
rect 476 32809 480 32877
rect 544 32847 552 32881
rect 578 32847 582 32881
rect 544 32839 548 32847
rect 544 32809 586 32810
rect 288 32769 292 32801
rect 296 32799 368 32807
rect 378 32799 450 32807
rect 544 32802 548 32809
rect 439 32771 444 32799
rect 120 32755 170 32757
rect 76 32751 130 32755
rect 110 32746 130 32751
rect 60 32721 67 32731
rect 76 32721 77 32741
rect 96 32712 99 32746
rect 109 32721 110 32741
rect 119 32721 126 32731
rect 76 32705 92 32711
rect 94 32705 110 32711
rect 170 32705 172 32755
rect 186 32689 190 32723
rect 216 32689 220 32723
rect 213 32657 224 32689
rect 282 32685 292 32769
rect 296 32763 368 32771
rect 378 32763 450 32771
rect 468 32768 473 32802
rect 428 32733 430 32749
rect 251 32657 292 32685
rect 318 32664 324 32733
rect 12 32652 62 32654
rect 28 32643 59 32651
rect 62 32643 64 32652
rect 251 32651 263 32657
rect 28 32635 64 32643
rect 127 32643 158 32651
rect 127 32636 182 32643
rect 127 32635 161 32636
rect 59 32619 64 32635
rect 158 32619 161 32635
rect 253 32623 263 32651
rect 273 32623 293 32657
rect 318 32654 335 32664
rect 303 32638 316 32648
rect 318 32638 324 32654
rect 346 32648 348 32733
rect 400 32725 430 32733
rect 476 32731 480 32799
rect 511 32768 582 32802
rect 544 32761 548 32768
rect 400 32721 436 32725
rect 400 32691 408 32721
rect 420 32691 436 32721
rect 544 32723 548 32731
rect 28 32611 64 32619
rect 127 32618 161 32619
rect 127 32611 182 32618
rect 62 32602 64 32611
rect 282 32565 292 32623
rect 295 32614 324 32638
rect 333 32638 353 32648
rect 428 32644 430 32691
rect 476 32651 480 32719
rect 544 32689 552 32723
rect 578 32689 582 32723
rect 544 32681 548 32689
rect 367 32638 380 32644
rect 333 32614 380 32638
rect 318 32601 324 32614
rect 346 32601 348 32614
rect 367 32610 380 32614
rect 396 32610 408 32644
rect 420 32610 436 32644
rect 544 32641 553 32669
rect 319 32590 346 32601
rect 120 32549 170 32551
rect 76 32543 92 32549
rect 94 32543 110 32549
rect 76 32533 99 32542
rect 60 32523 67 32533
rect 76 32513 77 32533
rect 96 32508 99 32533
rect 109 32513 110 32533
rect 119 32523 126 32533
rect 76 32499 110 32503
rect 170 32499 172 32549
rect 186 32531 190 32565
rect 216 32531 220 32565
rect 182 32493 224 32494
rect 186 32469 220 32486
rect 223 32469 257 32486
rect 182 32452 257 32469
rect 182 32451 224 32452
rect 160 32445 246 32451
rect 288 32445 292 32565
rect 296 32563 368 32571
rect 428 32563 430 32610
rect 476 32573 480 32641
rect 485 32597 495 32631
rect 505 32603 525 32631
rect 505 32597 519 32603
rect 544 32597 555 32641
rect 485 32573 492 32597
rect 579 32582 582 32672
rect 612 32654 624 32655
rect 599 32652 649 32654
rect 612 32651 624 32652
rect 610 32644 632 32651
rect 607 32643 632 32644
rect 586 32636 644 32643
rect 607 32635 644 32636
rect 607 32619 610 32635
rect 616 32619 644 32635
rect 607 32618 644 32619
rect 586 32611 644 32618
rect 607 32610 610 32611
rect 612 32603 632 32611
rect 612 32599 624 32603
rect 649 32602 651 32652
rect 544 32565 548 32573
rect 400 32533 408 32563
rect 420 32533 436 32563
rect 400 32529 436 32533
rect 400 32521 430 32529
rect 428 32505 430 32521
rect 476 32493 480 32561
rect 544 32531 552 32565
rect 578 32531 582 32565
rect 544 32523 548 32531
rect 295 32452 300 32486
rect 324 32452 329 32486
rect 378 32483 450 32491
rect 544 32488 548 32493
rect 544 32484 582 32488
rect 544 32469 552 32484
rect 578 32469 582 32484
rect 544 32451 586 32469
rect 522 32445 608 32451
rect 182 32429 224 32445
rect 544 32429 586 32445
rect 17 32415 67 32417
rect 119 32415 169 32417
rect 186 32415 220 32429
rect 548 32415 582 32429
rect 599 32415 649 32417
rect 42 32373 59 32407
rect 67 32365 69 32415
rect 160 32407 246 32415
rect 522 32407 608 32415
rect 76 32373 110 32407
rect 127 32373 144 32407
rect 152 32373 161 32407
rect 162 32405 195 32407
rect 224 32405 244 32407
rect 162 32373 244 32405
rect 524 32405 548 32407
rect 573 32405 582 32407
rect 586 32405 606 32407
rect 160 32365 246 32373
rect 186 32349 220 32365
rect 182 32335 224 32336
rect 160 32329 182 32335
rect 224 32329 246 32335
rect 186 32294 220 32328
rect 223 32294 257 32328
rect 120 32281 170 32283
rect 76 32277 130 32281
rect 110 32272 130 32277
rect 60 32247 67 32257
rect 76 32247 77 32267
rect 96 32238 99 32272
rect 109 32247 110 32267
rect 119 32247 126 32257
rect 76 32231 92 32237
rect 94 32231 110 32237
rect 170 32231 172 32281
rect 186 32215 190 32249
rect 216 32215 220 32249
rect 288 32215 292 32403
rect 476 32335 480 32403
rect 524 32373 606 32405
rect 607 32373 616 32407
rect 522 32365 608 32373
rect 649 32365 651 32415
rect 548 32349 582 32365
rect 522 32330 548 32335
rect 522 32329 582 32330
rect 586 32329 608 32335
rect 295 32294 300 32328
rect 324 32294 329 32328
rect 544 32326 582 32329
rect 378 32289 450 32297
rect 428 32259 430 32275
rect 400 32251 430 32259
rect 476 32257 480 32325
rect 544 32296 552 32326
rect 578 32296 582 32326
rect 544 32287 548 32296
rect 400 32247 436 32251
rect 400 32217 408 32247
rect 420 32217 436 32247
rect 544 32249 548 32257
rect 12 32178 62 32180
rect 28 32169 59 32177
rect 62 32169 64 32178
rect 28 32161 64 32169
rect 127 32169 158 32177
rect 127 32162 182 32169
rect 215 32167 224 32195
rect 127 32161 161 32162
rect 59 32145 64 32161
rect 158 32145 161 32161
rect 28 32137 64 32145
rect 127 32144 161 32145
rect 127 32137 182 32144
rect 62 32128 64 32137
rect 213 32129 224 32167
rect 282 32157 292 32215
rect 296 32209 368 32217
rect 319 32179 346 32190
rect 318 32166 324 32179
rect 346 32166 348 32179
rect 428 32170 430 32217
rect 443 32207 450 32209
rect 476 32177 480 32245
rect 544 32215 552 32249
rect 578 32215 582 32249
rect 481 32183 517 32211
rect 481 32177 495 32183
rect 367 32166 380 32170
rect 251 32123 263 32157
rect 273 32123 293 32157
rect 295 32142 324 32166
rect 303 32132 316 32142
rect 318 32126 324 32142
rect 333 32142 380 32166
rect 333 32132 353 32142
rect 367 32136 380 32142
rect 396 32136 408 32170
rect 420 32136 436 32170
rect 120 32075 170 32077
rect 76 32069 92 32075
rect 94 32069 110 32075
rect 76 32059 99 32068
rect 60 32049 67 32059
rect 76 32039 77 32059
rect 96 32034 99 32059
rect 109 32039 110 32059
rect 119 32049 126 32059
rect 76 32025 110 32029
rect 170 32025 172 32075
rect 186 32057 190 32091
rect 216 32057 220 32091
rect 186 31980 220 32014
rect 282 32011 292 32123
rect 318 32116 335 32126
rect 318 32047 324 32116
rect 346 32047 348 32132
rect 428 32089 430 32136
rect 476 32099 480 32167
rect 485 32149 495 32177
rect 505 32177 519 32183
rect 544 32177 555 32215
rect 505 32149 525 32177
rect 544 32149 553 32177
rect 544 32129 548 32149
rect 579 32108 582 32198
rect 612 32180 624 32181
rect 599 32178 649 32180
rect 612 32177 624 32178
rect 610 32170 632 32177
rect 607 32169 632 32170
rect 586 32162 644 32169
rect 607 32161 644 32162
rect 607 32145 610 32161
rect 616 32145 644 32161
rect 607 32144 644 32145
rect 586 32137 644 32144
rect 607 32136 610 32137
rect 612 32129 632 32137
rect 612 32125 624 32129
rect 649 32128 651 32178
rect 544 32091 548 32099
rect 400 32059 408 32089
rect 420 32059 436 32089
rect 400 32055 436 32059
rect 400 32047 430 32055
rect 428 32031 430 32047
rect 476 32019 480 32087
rect 544 32057 552 32091
rect 578 32057 582 32091
rect 544 32049 548 32057
rect 544 32019 586 32020
rect 288 31979 292 32011
rect 296 32009 368 32017
rect 378 32009 450 32017
rect 544 32012 548 32019
rect 439 31981 444 32009
rect 120 31965 170 31967
rect 76 31961 130 31965
rect 110 31956 130 31961
rect 60 31931 67 31941
rect 76 31931 77 31951
rect 96 31922 99 31956
rect 109 31931 110 31951
rect 119 31931 126 31941
rect 76 31915 92 31921
rect 94 31915 110 31921
rect 170 31915 172 31965
rect 186 31899 190 31933
rect 216 31899 220 31933
rect 213 31867 224 31899
rect 282 31895 292 31979
rect 296 31973 368 31981
rect 378 31973 450 31981
rect 468 31978 473 32012
rect 428 31943 430 31959
rect 251 31867 292 31895
rect 318 31874 324 31943
rect 12 31862 62 31864
rect 28 31853 59 31861
rect 62 31853 64 31862
rect 251 31861 263 31867
rect 28 31845 64 31853
rect 127 31853 158 31861
rect 127 31846 182 31853
rect 127 31845 161 31846
rect 59 31829 64 31845
rect 158 31829 161 31845
rect 253 31833 263 31861
rect 273 31833 293 31867
rect 318 31864 335 31874
rect 303 31848 316 31858
rect 318 31848 324 31864
rect 346 31858 348 31943
rect 400 31935 430 31943
rect 476 31941 480 32009
rect 511 31978 582 32012
rect 544 31971 548 31978
rect 400 31931 436 31935
rect 400 31901 408 31931
rect 420 31901 436 31931
rect 544 31933 548 31941
rect 28 31821 64 31829
rect 127 31828 161 31829
rect 127 31821 182 31828
rect 62 31812 64 31821
rect 282 31775 292 31833
rect 295 31824 324 31848
rect 333 31848 353 31858
rect 428 31854 430 31901
rect 476 31861 480 31929
rect 544 31899 552 31933
rect 578 31899 582 31933
rect 544 31891 548 31899
rect 367 31848 380 31854
rect 333 31824 380 31848
rect 318 31811 324 31824
rect 346 31811 348 31824
rect 367 31820 380 31824
rect 396 31820 408 31854
rect 420 31820 436 31854
rect 544 31851 553 31879
rect 319 31800 346 31811
rect 120 31759 170 31761
rect 76 31753 92 31759
rect 94 31753 110 31759
rect 76 31743 99 31752
rect 60 31733 67 31743
rect 76 31723 77 31743
rect 96 31718 99 31743
rect 109 31723 110 31743
rect 119 31733 126 31743
rect 76 31709 110 31713
rect 170 31709 172 31759
rect 186 31741 190 31775
rect 216 31741 220 31775
rect 182 31703 224 31704
rect 186 31679 220 31696
rect 223 31679 257 31696
rect 182 31662 257 31679
rect 182 31661 224 31662
rect 160 31655 246 31661
rect 288 31655 292 31775
rect 296 31773 368 31781
rect 428 31773 430 31820
rect 476 31783 480 31851
rect 485 31807 495 31841
rect 505 31813 525 31841
rect 505 31807 519 31813
rect 544 31807 555 31851
rect 485 31783 492 31807
rect 579 31792 582 31882
rect 612 31864 624 31865
rect 599 31862 649 31864
rect 612 31861 624 31862
rect 610 31854 632 31861
rect 607 31853 632 31854
rect 586 31846 644 31853
rect 607 31845 644 31846
rect 607 31829 610 31845
rect 616 31829 644 31845
rect 607 31828 644 31829
rect 586 31821 644 31828
rect 607 31820 610 31821
rect 612 31813 632 31821
rect 612 31809 624 31813
rect 649 31812 651 31862
rect 544 31775 548 31783
rect 400 31743 408 31773
rect 420 31743 436 31773
rect 400 31739 436 31743
rect 400 31731 430 31739
rect 428 31715 430 31731
rect 476 31703 480 31771
rect 544 31741 552 31775
rect 578 31741 582 31775
rect 544 31733 548 31741
rect 295 31662 300 31696
rect 324 31662 329 31696
rect 378 31693 450 31701
rect 544 31698 548 31703
rect 544 31694 582 31698
rect 544 31679 552 31694
rect 578 31679 582 31694
rect 544 31661 586 31679
rect 522 31655 608 31661
rect 182 31639 224 31655
rect 544 31639 586 31655
rect 17 31625 67 31627
rect 119 31625 169 31627
rect 186 31625 220 31639
rect 548 31625 582 31639
rect 599 31625 649 31627
rect 42 31583 59 31617
rect 67 31575 69 31625
rect 160 31617 246 31625
rect 522 31617 608 31625
rect 76 31583 110 31617
rect 127 31583 144 31617
rect 152 31583 161 31617
rect 162 31615 195 31617
rect 224 31615 244 31617
rect 162 31583 244 31615
rect 524 31615 548 31617
rect 573 31615 582 31617
rect 586 31615 606 31617
rect 160 31575 246 31583
rect 186 31559 220 31575
rect 182 31545 224 31546
rect 160 31539 182 31545
rect 224 31539 246 31545
rect 186 31504 220 31538
rect 223 31504 257 31538
rect 120 31491 170 31493
rect 76 31487 130 31491
rect 110 31482 130 31487
rect 60 31457 67 31467
rect 76 31457 77 31477
rect 96 31448 99 31482
rect 109 31457 110 31477
rect 119 31457 126 31467
rect 76 31441 92 31447
rect 94 31441 110 31447
rect 170 31441 172 31491
rect 186 31425 190 31459
rect 216 31425 220 31459
rect 288 31425 292 31613
rect 476 31545 480 31613
rect 524 31583 606 31615
rect 607 31583 616 31617
rect 522 31575 608 31583
rect 649 31575 651 31625
rect 548 31559 582 31575
rect 522 31540 548 31545
rect 522 31539 582 31540
rect 586 31539 608 31545
rect 295 31504 300 31538
rect 324 31504 329 31538
rect 544 31536 582 31539
rect 378 31499 450 31507
rect 428 31469 430 31485
rect 400 31461 430 31469
rect 476 31467 480 31535
rect 544 31506 552 31536
rect 578 31506 582 31536
rect 544 31497 548 31506
rect 400 31457 436 31461
rect 400 31427 408 31457
rect 420 31427 436 31457
rect 544 31459 548 31467
rect 12 31388 62 31390
rect 28 31379 59 31387
rect 62 31379 64 31388
rect 28 31371 64 31379
rect 127 31379 158 31387
rect 127 31372 182 31379
rect 215 31377 224 31405
rect 127 31371 161 31372
rect 59 31355 64 31371
rect 158 31355 161 31371
rect 28 31347 64 31355
rect 127 31354 161 31355
rect 127 31347 182 31354
rect 62 31338 64 31347
rect 213 31339 224 31377
rect 282 31367 292 31425
rect 296 31419 368 31427
rect 319 31389 346 31400
rect 318 31376 324 31389
rect 346 31376 348 31389
rect 428 31380 430 31427
rect 443 31417 450 31419
rect 476 31387 480 31455
rect 544 31425 552 31459
rect 578 31425 582 31459
rect 481 31393 517 31421
rect 481 31387 495 31393
rect 367 31376 380 31380
rect 251 31333 263 31367
rect 273 31333 293 31367
rect 295 31352 324 31376
rect 303 31342 316 31352
rect 318 31336 324 31352
rect 333 31352 380 31376
rect 333 31342 353 31352
rect 367 31346 380 31352
rect 396 31346 408 31380
rect 420 31346 436 31380
rect 120 31285 170 31287
rect 76 31279 92 31285
rect 94 31279 110 31285
rect 76 31269 99 31278
rect 60 31259 67 31269
rect 76 31249 77 31269
rect 96 31244 99 31269
rect 109 31249 110 31269
rect 119 31259 126 31269
rect 76 31235 110 31239
rect 170 31235 172 31285
rect 186 31267 190 31301
rect 216 31267 220 31301
rect 186 31190 220 31224
rect 282 31221 292 31333
rect 318 31326 335 31336
rect 318 31257 324 31326
rect 346 31257 348 31342
rect 428 31299 430 31346
rect 476 31309 480 31377
rect 485 31359 495 31387
rect 505 31387 519 31393
rect 544 31387 555 31425
rect 505 31359 525 31387
rect 544 31359 553 31387
rect 544 31339 548 31359
rect 579 31318 582 31408
rect 612 31390 624 31391
rect 599 31388 649 31390
rect 612 31387 624 31388
rect 610 31380 632 31387
rect 607 31379 632 31380
rect 586 31372 644 31379
rect 607 31371 644 31372
rect 607 31355 610 31371
rect 616 31355 644 31371
rect 607 31354 644 31355
rect 586 31347 644 31354
rect 607 31346 610 31347
rect 612 31339 632 31347
rect 612 31335 624 31339
rect 649 31338 651 31388
rect 544 31301 548 31309
rect 400 31269 408 31299
rect 420 31269 436 31299
rect 400 31265 436 31269
rect 400 31257 430 31265
rect 428 31241 430 31257
rect 476 31229 480 31297
rect 544 31267 552 31301
rect 578 31267 582 31301
rect 544 31259 548 31267
rect 544 31229 586 31230
rect 288 31189 292 31221
rect 296 31219 368 31227
rect 378 31219 450 31227
rect 544 31222 548 31229
rect 439 31191 444 31219
rect 120 31175 170 31177
rect 76 31171 130 31175
rect 110 31166 130 31171
rect 60 31141 67 31151
rect 76 31141 77 31161
rect 96 31132 99 31166
rect 109 31141 110 31161
rect 119 31141 126 31151
rect 76 31125 92 31131
rect 94 31125 110 31131
rect 170 31125 172 31175
rect 186 31109 190 31143
rect 216 31109 220 31143
rect 213 31077 224 31109
rect 282 31105 292 31189
rect 296 31183 368 31191
rect 378 31183 450 31191
rect 468 31188 473 31222
rect 428 31153 430 31169
rect 251 31077 292 31105
rect 318 31084 324 31153
rect 12 31072 62 31074
rect 28 31063 59 31071
rect 62 31063 64 31072
rect 251 31071 263 31077
rect 28 31055 64 31063
rect 127 31063 158 31071
rect 127 31056 182 31063
rect 127 31055 161 31056
rect 59 31039 64 31055
rect 158 31039 161 31055
rect 253 31043 263 31071
rect 273 31043 293 31077
rect 318 31074 335 31084
rect 303 31058 316 31068
rect 318 31058 324 31074
rect 346 31068 348 31153
rect 400 31145 430 31153
rect 476 31151 480 31219
rect 511 31188 582 31222
rect 544 31181 548 31188
rect 400 31141 436 31145
rect 400 31111 408 31141
rect 420 31111 436 31141
rect 544 31143 548 31151
rect 28 31031 64 31039
rect 127 31038 161 31039
rect 127 31031 182 31038
rect 62 31022 64 31031
rect 282 30985 292 31043
rect 295 31034 324 31058
rect 333 31058 353 31068
rect 428 31064 430 31111
rect 476 31071 480 31139
rect 544 31109 552 31143
rect 578 31109 582 31143
rect 544 31101 548 31109
rect 367 31058 380 31064
rect 333 31034 380 31058
rect 318 31021 324 31034
rect 346 31021 348 31034
rect 367 31030 380 31034
rect 396 31030 408 31064
rect 420 31030 436 31064
rect 544 31061 553 31089
rect 319 31010 346 31021
rect 120 30969 170 30971
rect 76 30963 92 30969
rect 94 30963 110 30969
rect 76 30953 99 30962
rect 60 30943 67 30953
rect 76 30933 77 30953
rect 96 30928 99 30953
rect 109 30933 110 30953
rect 119 30943 126 30953
rect 76 30919 110 30923
rect 170 30919 172 30969
rect 186 30951 190 30985
rect 216 30951 220 30985
rect 182 30913 224 30914
rect 186 30889 220 30906
rect 223 30889 257 30906
rect 182 30872 257 30889
rect 182 30871 224 30872
rect 160 30865 246 30871
rect 288 30865 292 30985
rect 296 30983 368 30991
rect 428 30983 430 31030
rect 476 30993 480 31061
rect 485 31017 495 31051
rect 505 31023 525 31051
rect 505 31017 519 31023
rect 544 31017 555 31061
rect 485 30993 492 31017
rect 579 31002 582 31092
rect 612 31074 624 31075
rect 599 31072 649 31074
rect 612 31071 624 31072
rect 610 31064 632 31071
rect 607 31063 632 31064
rect 586 31056 644 31063
rect 607 31055 644 31056
rect 607 31039 610 31055
rect 616 31039 644 31055
rect 607 31038 644 31039
rect 586 31031 644 31038
rect 607 31030 610 31031
rect 612 31023 632 31031
rect 612 31019 624 31023
rect 649 31022 651 31072
rect 544 30985 548 30993
rect 400 30953 408 30983
rect 420 30953 436 30983
rect 400 30949 436 30953
rect 400 30941 430 30949
rect 428 30925 430 30941
rect 476 30913 480 30981
rect 544 30951 552 30985
rect 578 30951 582 30985
rect 544 30943 548 30951
rect 295 30872 300 30906
rect 324 30872 329 30906
rect 378 30903 450 30911
rect 544 30908 548 30913
rect 544 30904 582 30908
rect 544 30889 552 30904
rect 578 30889 582 30904
rect 544 30871 586 30889
rect 522 30865 608 30871
rect 182 30849 224 30865
rect 544 30849 586 30865
rect 17 30835 67 30837
rect 119 30835 169 30837
rect 186 30835 220 30849
rect 548 30835 582 30849
rect 599 30835 649 30837
rect 42 30793 59 30827
rect 67 30785 69 30835
rect 160 30827 246 30835
rect 522 30827 608 30835
rect 76 30793 110 30827
rect 127 30793 144 30827
rect 152 30793 161 30827
rect 162 30825 195 30827
rect 224 30825 244 30827
rect 162 30793 244 30825
rect 524 30825 548 30827
rect 573 30825 582 30827
rect 586 30825 606 30827
rect 160 30785 246 30793
rect 186 30769 220 30785
rect 182 30755 224 30756
rect 160 30749 182 30755
rect 224 30749 246 30755
rect 186 30714 220 30748
rect 223 30714 257 30748
rect 120 30701 170 30703
rect 76 30697 130 30701
rect 110 30692 130 30697
rect 60 30667 67 30677
rect 76 30667 77 30687
rect 96 30658 99 30692
rect 109 30667 110 30687
rect 119 30667 126 30677
rect 76 30651 92 30657
rect 94 30651 110 30657
rect 170 30651 172 30701
rect 186 30635 190 30669
rect 216 30635 220 30669
rect 288 30635 292 30823
rect 476 30755 480 30823
rect 524 30793 606 30825
rect 607 30793 616 30827
rect 522 30785 608 30793
rect 649 30785 651 30835
rect 548 30769 582 30785
rect 522 30750 548 30755
rect 522 30749 582 30750
rect 586 30749 608 30755
rect 295 30714 300 30748
rect 324 30714 329 30748
rect 544 30746 582 30749
rect 378 30709 450 30717
rect 428 30679 430 30695
rect 400 30671 430 30679
rect 476 30677 480 30745
rect 544 30716 552 30746
rect 578 30716 582 30746
rect 544 30707 548 30716
rect 400 30667 436 30671
rect 400 30637 408 30667
rect 420 30637 436 30667
rect 544 30669 548 30677
rect 12 30598 62 30600
rect 28 30589 59 30597
rect 62 30589 64 30598
rect 28 30581 64 30589
rect 127 30589 158 30597
rect 127 30582 182 30589
rect 215 30587 224 30615
rect 127 30581 161 30582
rect 59 30565 64 30581
rect 158 30565 161 30581
rect 28 30557 64 30565
rect 127 30564 161 30565
rect 127 30557 182 30564
rect 62 30548 64 30557
rect 213 30549 224 30587
rect 282 30577 292 30635
rect 296 30629 368 30637
rect 319 30599 346 30610
rect 318 30586 324 30599
rect 346 30586 348 30599
rect 428 30590 430 30637
rect 443 30627 450 30629
rect 476 30597 480 30665
rect 544 30635 552 30669
rect 578 30635 582 30669
rect 481 30603 517 30631
rect 481 30597 495 30603
rect 367 30586 380 30590
rect 251 30543 263 30577
rect 273 30543 293 30577
rect 295 30562 324 30586
rect 303 30552 316 30562
rect 318 30546 324 30562
rect 333 30562 380 30586
rect 333 30552 353 30562
rect 367 30556 380 30562
rect 396 30556 408 30590
rect 420 30556 436 30590
rect 120 30495 170 30497
rect 76 30489 92 30495
rect 94 30489 110 30495
rect 76 30479 99 30488
rect 60 30469 67 30479
rect 76 30459 77 30479
rect 96 30454 99 30479
rect 109 30459 110 30479
rect 119 30469 126 30479
rect 76 30445 110 30449
rect 170 30445 172 30495
rect 186 30477 190 30511
rect 216 30477 220 30511
rect 186 30400 220 30434
rect 282 30431 292 30543
rect 318 30536 335 30546
rect 318 30467 324 30536
rect 346 30467 348 30552
rect 428 30509 430 30556
rect 476 30519 480 30587
rect 485 30569 495 30597
rect 505 30597 519 30603
rect 544 30597 555 30635
rect 505 30569 525 30597
rect 544 30569 553 30597
rect 544 30549 548 30569
rect 579 30528 582 30618
rect 612 30600 624 30601
rect 599 30598 649 30600
rect 612 30597 624 30598
rect 610 30590 632 30597
rect 607 30589 632 30590
rect 586 30582 644 30589
rect 607 30581 644 30582
rect 607 30565 610 30581
rect 616 30565 644 30581
rect 607 30564 644 30565
rect 586 30557 644 30564
rect 607 30556 610 30557
rect 612 30549 632 30557
rect 612 30545 624 30549
rect 649 30548 651 30598
rect 544 30511 548 30519
rect 400 30479 408 30509
rect 420 30479 436 30509
rect 400 30475 436 30479
rect 400 30467 430 30475
rect 428 30451 430 30467
rect 476 30439 480 30507
rect 544 30477 552 30511
rect 578 30477 582 30511
rect 544 30469 548 30477
rect 544 30439 586 30440
rect 288 30399 292 30431
rect 296 30429 368 30437
rect 378 30429 450 30437
rect 544 30432 548 30439
rect 439 30401 444 30429
rect 120 30385 170 30387
rect 76 30381 130 30385
rect 110 30376 130 30381
rect 60 30351 67 30361
rect 76 30351 77 30371
rect 96 30342 99 30376
rect 109 30351 110 30371
rect 119 30351 126 30361
rect 76 30335 92 30341
rect 94 30335 110 30341
rect 170 30335 172 30385
rect 186 30319 190 30353
rect 216 30319 220 30353
rect 213 30287 224 30319
rect 282 30315 292 30399
rect 296 30393 368 30401
rect 378 30393 450 30401
rect 468 30398 473 30432
rect 428 30363 430 30379
rect 251 30287 292 30315
rect 318 30294 324 30363
rect 12 30282 62 30284
rect 28 30273 59 30281
rect 62 30273 64 30282
rect 251 30281 263 30287
rect 28 30265 64 30273
rect 127 30273 158 30281
rect 127 30266 182 30273
rect 127 30265 161 30266
rect 59 30249 64 30265
rect 158 30249 161 30265
rect 253 30253 263 30281
rect 273 30253 293 30287
rect 318 30284 335 30294
rect 303 30268 316 30278
rect 318 30268 324 30284
rect 346 30278 348 30363
rect 400 30355 430 30363
rect 476 30361 480 30429
rect 511 30398 582 30432
rect 544 30391 548 30398
rect 400 30351 436 30355
rect 400 30321 408 30351
rect 420 30321 436 30351
rect 544 30353 548 30361
rect 28 30241 64 30249
rect 127 30248 161 30249
rect 127 30241 182 30248
rect 62 30232 64 30241
rect 282 30195 292 30253
rect 295 30244 324 30268
rect 333 30268 353 30278
rect 428 30274 430 30321
rect 476 30281 480 30349
rect 544 30319 552 30353
rect 578 30319 582 30353
rect 544 30311 548 30319
rect 367 30268 380 30274
rect 333 30244 380 30268
rect 318 30231 324 30244
rect 346 30231 348 30244
rect 367 30240 380 30244
rect 396 30240 408 30274
rect 420 30240 436 30274
rect 544 30271 553 30299
rect 319 30220 346 30231
rect 120 30179 170 30181
rect 76 30173 92 30179
rect 94 30173 110 30179
rect 76 30163 99 30172
rect 60 30153 67 30163
rect 76 30143 77 30163
rect 96 30138 99 30163
rect 109 30143 110 30163
rect 119 30153 126 30163
rect 76 30129 110 30133
rect 170 30129 172 30179
rect 186 30161 190 30195
rect 216 30161 220 30195
rect 182 30123 224 30124
rect 186 30099 220 30116
rect 223 30099 257 30116
rect 182 30082 257 30099
rect 182 30081 224 30082
rect 160 30075 246 30081
rect 288 30075 292 30195
rect 296 30193 368 30201
rect 428 30193 430 30240
rect 476 30203 480 30271
rect 485 30227 495 30261
rect 505 30233 525 30261
rect 505 30227 519 30233
rect 544 30227 555 30271
rect 485 30203 492 30227
rect 579 30212 582 30302
rect 612 30284 624 30285
rect 599 30282 649 30284
rect 612 30281 624 30282
rect 610 30274 632 30281
rect 607 30273 632 30274
rect 586 30266 644 30273
rect 607 30265 644 30266
rect 607 30249 610 30265
rect 616 30249 644 30265
rect 607 30248 644 30249
rect 586 30241 644 30248
rect 607 30240 610 30241
rect 612 30233 632 30241
rect 612 30229 624 30233
rect 649 30232 651 30282
rect 544 30195 548 30203
rect 400 30163 408 30193
rect 420 30163 436 30193
rect 400 30159 436 30163
rect 400 30151 430 30159
rect 428 30135 430 30151
rect 476 30123 480 30191
rect 544 30161 552 30195
rect 578 30161 582 30195
rect 544 30153 548 30161
rect 295 30082 300 30116
rect 324 30082 329 30116
rect 378 30113 450 30121
rect 544 30118 548 30123
rect 544 30114 582 30118
rect 544 30099 552 30114
rect 578 30099 582 30114
rect 544 30081 586 30099
rect 522 30075 608 30081
rect 182 30059 224 30075
rect 544 30059 586 30075
rect 17 30045 67 30047
rect 119 30045 169 30047
rect 186 30045 220 30059
rect 548 30045 582 30059
rect 599 30045 649 30047
rect 42 30003 59 30037
rect 67 29995 69 30045
rect 160 30037 246 30045
rect 522 30037 608 30045
rect 76 30003 110 30037
rect 127 30003 144 30037
rect 152 30003 161 30037
rect 162 30035 195 30037
rect 224 30035 244 30037
rect 162 30003 244 30035
rect 524 30035 548 30037
rect 573 30035 582 30037
rect 586 30035 606 30037
rect 160 29995 246 30003
rect 186 29979 220 29995
rect 182 29965 224 29966
rect 160 29959 182 29965
rect 224 29959 246 29965
rect 186 29924 220 29958
rect 223 29924 257 29958
rect 120 29911 170 29913
rect 76 29907 130 29911
rect 110 29902 130 29907
rect 60 29877 67 29887
rect 76 29877 77 29897
rect 96 29868 99 29902
rect 109 29877 110 29897
rect 119 29877 126 29887
rect 76 29861 92 29867
rect 94 29861 110 29867
rect 170 29861 172 29911
rect 186 29845 190 29879
rect 216 29845 220 29879
rect 288 29845 292 30033
rect 476 29965 480 30033
rect 524 30003 606 30035
rect 607 30003 616 30037
rect 522 29995 608 30003
rect 649 29995 651 30045
rect 548 29979 582 29995
rect 522 29960 548 29965
rect 522 29959 582 29960
rect 586 29959 608 29965
rect 295 29924 300 29958
rect 324 29924 329 29958
rect 544 29956 582 29959
rect 378 29919 450 29927
rect 428 29889 430 29905
rect 400 29881 430 29889
rect 476 29887 480 29955
rect 544 29926 552 29956
rect 578 29926 582 29956
rect 544 29917 548 29926
rect 400 29877 436 29881
rect 400 29847 408 29877
rect 420 29847 436 29877
rect 544 29879 548 29887
rect 12 29808 62 29810
rect 28 29799 59 29807
rect 62 29799 64 29808
rect 28 29791 64 29799
rect 127 29799 158 29807
rect 127 29792 182 29799
rect 215 29797 224 29825
rect 127 29791 161 29792
rect 59 29775 64 29791
rect 158 29775 161 29791
rect 28 29767 64 29775
rect 127 29774 161 29775
rect 127 29767 182 29774
rect 62 29758 64 29767
rect 213 29759 224 29797
rect 282 29787 292 29845
rect 296 29839 368 29847
rect 319 29809 346 29820
rect 318 29796 324 29809
rect 346 29796 348 29809
rect 428 29800 430 29847
rect 443 29837 450 29839
rect 476 29807 480 29875
rect 544 29845 552 29879
rect 578 29845 582 29879
rect 481 29813 517 29841
rect 481 29807 495 29813
rect 367 29796 380 29800
rect 251 29753 263 29787
rect 273 29753 293 29787
rect 295 29772 324 29796
rect 303 29762 316 29772
rect 318 29756 324 29772
rect 333 29772 380 29796
rect 333 29762 353 29772
rect 367 29766 380 29772
rect 396 29766 408 29800
rect 420 29766 436 29800
rect 120 29705 170 29707
rect 76 29699 92 29705
rect 94 29699 110 29705
rect 76 29689 99 29698
rect 60 29679 67 29689
rect 76 29669 77 29689
rect 96 29664 99 29689
rect 109 29669 110 29689
rect 119 29679 126 29689
rect 76 29655 110 29659
rect 170 29655 172 29705
rect 186 29687 190 29721
rect 216 29687 220 29721
rect 186 29610 220 29644
rect 282 29641 292 29753
rect 318 29746 335 29756
rect 318 29677 324 29746
rect 346 29677 348 29762
rect 428 29719 430 29766
rect 476 29729 480 29797
rect 485 29779 495 29807
rect 505 29807 519 29813
rect 544 29807 555 29845
rect 505 29779 525 29807
rect 544 29779 553 29807
rect 544 29759 548 29779
rect 579 29738 582 29828
rect 612 29810 624 29811
rect 599 29808 649 29810
rect 612 29807 624 29808
rect 610 29800 632 29807
rect 607 29799 632 29800
rect 586 29792 644 29799
rect 607 29791 644 29792
rect 607 29775 610 29791
rect 616 29775 644 29791
rect 607 29774 644 29775
rect 586 29767 644 29774
rect 607 29766 610 29767
rect 612 29759 632 29767
rect 612 29755 624 29759
rect 649 29758 651 29808
rect 544 29721 548 29729
rect 400 29689 408 29719
rect 420 29689 436 29719
rect 400 29685 436 29689
rect 400 29677 430 29685
rect 428 29661 430 29677
rect 476 29649 480 29717
rect 544 29687 552 29721
rect 578 29687 582 29721
rect 544 29679 548 29687
rect 544 29649 586 29650
rect 288 29609 292 29641
rect 296 29639 368 29647
rect 378 29639 450 29647
rect 544 29642 548 29649
rect 439 29611 444 29639
rect 120 29595 170 29597
rect 76 29591 130 29595
rect 110 29586 130 29591
rect 60 29561 67 29571
rect 76 29561 77 29581
rect 96 29552 99 29586
rect 109 29561 110 29581
rect 119 29561 126 29571
rect 76 29545 92 29551
rect 94 29545 110 29551
rect 170 29545 172 29595
rect 186 29529 190 29563
rect 216 29529 220 29563
rect 213 29497 224 29529
rect 282 29525 292 29609
rect 296 29603 368 29611
rect 378 29603 450 29611
rect 468 29608 473 29642
rect 428 29573 430 29589
rect 251 29497 292 29525
rect 318 29504 324 29573
rect 12 29492 62 29494
rect 28 29483 59 29491
rect 62 29483 64 29492
rect 251 29491 263 29497
rect 28 29475 64 29483
rect 127 29483 158 29491
rect 127 29476 182 29483
rect 127 29475 161 29476
rect 59 29459 64 29475
rect 158 29459 161 29475
rect 253 29463 263 29491
rect 273 29463 293 29497
rect 318 29494 335 29504
rect 303 29478 316 29488
rect 318 29478 324 29494
rect 346 29488 348 29573
rect 400 29565 430 29573
rect 476 29571 480 29639
rect 511 29608 582 29642
rect 544 29601 548 29608
rect 400 29561 436 29565
rect 400 29531 408 29561
rect 420 29531 436 29561
rect 544 29563 548 29571
rect 28 29451 64 29459
rect 127 29458 161 29459
rect 127 29451 182 29458
rect 62 29442 64 29451
rect 282 29405 292 29463
rect 295 29454 324 29478
rect 333 29478 353 29488
rect 428 29484 430 29531
rect 476 29491 480 29559
rect 544 29529 552 29563
rect 578 29529 582 29563
rect 544 29521 548 29529
rect 367 29478 380 29484
rect 333 29454 380 29478
rect 318 29441 324 29454
rect 346 29441 348 29454
rect 367 29450 380 29454
rect 396 29450 408 29484
rect 420 29450 436 29484
rect 544 29481 553 29509
rect 319 29430 346 29441
rect 120 29389 170 29391
rect 76 29383 92 29389
rect 94 29383 110 29389
rect 76 29373 99 29382
rect 60 29363 67 29373
rect 76 29353 77 29373
rect 96 29348 99 29373
rect 109 29353 110 29373
rect 119 29363 126 29373
rect 76 29339 110 29343
rect 170 29339 172 29389
rect 186 29371 190 29405
rect 216 29371 220 29405
rect 182 29333 224 29334
rect 186 29309 220 29326
rect 223 29309 257 29326
rect 182 29292 257 29309
rect 182 29291 224 29292
rect 160 29285 246 29291
rect 288 29285 292 29405
rect 296 29403 368 29411
rect 428 29403 430 29450
rect 476 29413 480 29481
rect 485 29437 495 29471
rect 505 29443 525 29471
rect 505 29437 519 29443
rect 544 29437 555 29481
rect 485 29413 492 29437
rect 579 29422 582 29512
rect 612 29494 624 29495
rect 599 29492 649 29494
rect 612 29491 624 29492
rect 610 29484 632 29491
rect 607 29483 632 29484
rect 586 29476 644 29483
rect 607 29475 644 29476
rect 607 29459 610 29475
rect 616 29459 644 29475
rect 607 29458 644 29459
rect 586 29451 644 29458
rect 607 29450 610 29451
rect 612 29443 632 29451
rect 612 29439 624 29443
rect 649 29442 651 29492
rect 544 29405 548 29413
rect 400 29373 408 29403
rect 420 29373 436 29403
rect 400 29369 436 29373
rect 400 29361 430 29369
rect 428 29345 430 29361
rect 476 29333 480 29401
rect 544 29371 552 29405
rect 578 29371 582 29405
rect 544 29363 548 29371
rect 295 29292 300 29326
rect 324 29292 329 29326
rect 378 29323 450 29331
rect 544 29328 548 29333
rect 544 29324 582 29328
rect 544 29309 552 29324
rect 578 29309 582 29324
rect 544 29291 586 29309
rect 522 29285 608 29291
rect 182 29269 224 29285
rect 544 29269 586 29285
rect 17 29255 67 29257
rect 119 29255 169 29257
rect 186 29255 220 29269
rect 548 29255 582 29269
rect 599 29255 649 29257
rect 42 29213 59 29247
rect 67 29205 69 29255
rect 160 29247 246 29255
rect 522 29247 608 29255
rect 76 29213 110 29247
rect 127 29213 144 29247
rect 152 29213 161 29247
rect 162 29245 195 29247
rect 224 29245 244 29247
rect 162 29213 244 29245
rect 524 29245 548 29247
rect 573 29245 582 29247
rect 586 29245 606 29247
rect 160 29205 246 29213
rect 186 29189 220 29205
rect 182 29175 224 29176
rect 160 29169 182 29175
rect 224 29169 246 29175
rect 186 29134 220 29168
rect 223 29134 257 29168
rect 120 29121 170 29123
rect 76 29117 130 29121
rect 110 29112 130 29117
rect 60 29087 67 29097
rect 76 29087 77 29107
rect 96 29078 99 29112
rect 109 29087 110 29107
rect 119 29087 126 29097
rect 76 29071 92 29077
rect 94 29071 110 29077
rect 170 29071 172 29121
rect 186 29055 190 29089
rect 216 29055 220 29089
rect 288 29055 292 29243
rect 476 29175 480 29243
rect 524 29213 606 29245
rect 607 29213 616 29247
rect 522 29205 608 29213
rect 649 29205 651 29255
rect 548 29189 582 29205
rect 522 29170 548 29175
rect 522 29169 582 29170
rect 586 29169 608 29175
rect 295 29134 300 29168
rect 324 29134 329 29168
rect 544 29166 582 29169
rect 378 29129 450 29137
rect 428 29099 430 29115
rect 400 29091 430 29099
rect 476 29097 480 29165
rect 544 29136 552 29166
rect 578 29136 582 29166
rect 544 29127 548 29136
rect 400 29087 436 29091
rect 400 29057 408 29087
rect 420 29057 436 29087
rect 544 29089 548 29097
rect 12 29018 62 29020
rect 28 29009 59 29017
rect 62 29009 64 29018
rect 28 29001 64 29009
rect 127 29009 158 29017
rect 127 29002 182 29009
rect 215 29007 224 29035
rect 127 29001 161 29002
rect 59 28985 64 29001
rect 158 28985 161 29001
rect 28 28977 64 28985
rect 127 28984 161 28985
rect 127 28977 182 28984
rect 62 28968 64 28977
rect 213 28969 224 29007
rect 282 28997 292 29055
rect 296 29049 368 29057
rect 319 29019 346 29030
rect 318 29006 324 29019
rect 346 29006 348 29019
rect 428 29010 430 29057
rect 443 29047 450 29049
rect 476 29017 480 29085
rect 544 29055 552 29089
rect 578 29055 582 29089
rect 481 29023 517 29051
rect 481 29017 495 29023
rect 367 29006 380 29010
rect 251 28963 263 28997
rect 273 28963 293 28997
rect 295 28982 324 29006
rect 303 28972 316 28982
rect 318 28966 324 28982
rect 333 28982 380 29006
rect 333 28972 353 28982
rect 367 28976 380 28982
rect 396 28976 408 29010
rect 420 28976 436 29010
rect 120 28915 170 28917
rect 76 28909 92 28915
rect 94 28909 110 28915
rect 76 28899 99 28908
rect 60 28889 67 28899
rect 76 28879 77 28899
rect 96 28874 99 28899
rect 109 28879 110 28899
rect 119 28889 126 28899
rect 76 28865 110 28869
rect 170 28865 172 28915
rect 186 28897 190 28931
rect 216 28897 220 28931
rect 186 28820 220 28854
rect 282 28851 292 28963
rect 318 28956 335 28966
rect 318 28887 324 28956
rect 346 28887 348 28972
rect 428 28929 430 28976
rect 476 28939 480 29007
rect 485 28989 495 29017
rect 505 29017 519 29023
rect 544 29017 555 29055
rect 505 28989 525 29017
rect 544 28989 553 29017
rect 544 28969 548 28989
rect 579 28948 582 29038
rect 612 29020 624 29021
rect 599 29018 649 29020
rect 612 29017 624 29018
rect 610 29010 632 29017
rect 607 29009 632 29010
rect 586 29002 644 29009
rect 607 29001 644 29002
rect 607 28985 610 29001
rect 616 28985 644 29001
rect 607 28984 644 28985
rect 586 28977 644 28984
rect 607 28976 610 28977
rect 612 28969 632 28977
rect 612 28965 624 28969
rect 649 28968 651 29018
rect 544 28931 548 28939
rect 400 28899 408 28929
rect 420 28899 436 28929
rect 400 28895 436 28899
rect 400 28887 430 28895
rect 428 28871 430 28887
rect 476 28859 480 28927
rect 544 28897 552 28931
rect 578 28897 582 28931
rect 544 28889 548 28897
rect 544 28859 586 28860
rect 288 28819 292 28851
rect 296 28849 368 28857
rect 378 28849 450 28857
rect 544 28852 548 28859
rect 439 28821 444 28849
rect 120 28805 170 28807
rect 76 28801 130 28805
rect 110 28796 130 28801
rect 60 28771 67 28781
rect 76 28771 77 28791
rect 96 28762 99 28796
rect 109 28771 110 28791
rect 119 28771 126 28781
rect 76 28755 92 28761
rect 94 28755 110 28761
rect 170 28755 172 28805
rect 186 28739 190 28773
rect 216 28739 220 28773
rect 213 28707 224 28739
rect 282 28735 292 28819
rect 296 28813 368 28821
rect 378 28813 450 28821
rect 468 28818 473 28852
rect 428 28783 430 28799
rect 251 28707 292 28735
rect 318 28714 324 28783
rect 12 28702 62 28704
rect 28 28693 59 28701
rect 62 28693 64 28702
rect 251 28701 263 28707
rect 28 28685 64 28693
rect 127 28693 158 28701
rect 127 28686 182 28693
rect 127 28685 161 28686
rect 59 28669 64 28685
rect 158 28669 161 28685
rect 253 28673 263 28701
rect 273 28673 293 28707
rect 318 28704 335 28714
rect 303 28688 316 28698
rect 318 28688 324 28704
rect 346 28698 348 28783
rect 400 28775 430 28783
rect 476 28781 480 28849
rect 511 28818 582 28852
rect 544 28811 548 28818
rect 400 28771 436 28775
rect 400 28741 408 28771
rect 420 28741 436 28771
rect 544 28773 548 28781
rect 28 28661 64 28669
rect 127 28668 161 28669
rect 127 28661 182 28668
rect 62 28652 64 28661
rect 282 28615 292 28673
rect 295 28664 324 28688
rect 333 28688 353 28698
rect 428 28694 430 28741
rect 476 28701 480 28769
rect 544 28739 552 28773
rect 578 28739 582 28773
rect 544 28731 548 28739
rect 367 28688 380 28694
rect 333 28664 380 28688
rect 318 28651 324 28664
rect 346 28651 348 28664
rect 367 28660 380 28664
rect 396 28660 408 28694
rect 420 28660 436 28694
rect 544 28691 553 28719
rect 319 28640 346 28651
rect 120 28599 170 28601
rect 76 28593 92 28599
rect 94 28593 110 28599
rect 76 28583 99 28592
rect 60 28573 67 28583
rect 76 28563 77 28583
rect 96 28558 99 28583
rect 109 28563 110 28583
rect 119 28573 126 28583
rect 76 28549 110 28553
rect 170 28549 172 28599
rect 186 28581 190 28615
rect 216 28581 220 28615
rect 182 28543 224 28544
rect 186 28519 220 28536
rect 223 28519 257 28536
rect 182 28502 257 28519
rect 182 28501 224 28502
rect 160 28495 246 28501
rect 288 28495 292 28615
rect 296 28613 368 28621
rect 428 28613 430 28660
rect 476 28623 480 28691
rect 485 28647 495 28681
rect 505 28653 525 28681
rect 505 28647 519 28653
rect 544 28647 555 28691
rect 485 28623 492 28647
rect 579 28632 582 28722
rect 612 28704 624 28705
rect 599 28702 649 28704
rect 612 28701 624 28702
rect 610 28694 632 28701
rect 607 28693 632 28694
rect 586 28686 644 28693
rect 607 28685 644 28686
rect 607 28669 610 28685
rect 616 28669 644 28685
rect 607 28668 644 28669
rect 586 28661 644 28668
rect 607 28660 610 28661
rect 612 28653 632 28661
rect 612 28649 624 28653
rect 649 28652 651 28702
rect 544 28615 548 28623
rect 400 28583 408 28613
rect 420 28583 436 28613
rect 400 28579 436 28583
rect 400 28571 430 28579
rect 428 28555 430 28571
rect 476 28543 480 28611
rect 544 28581 552 28615
rect 578 28581 582 28615
rect 544 28573 548 28581
rect 295 28502 300 28536
rect 324 28502 329 28536
rect 378 28533 450 28541
rect 544 28538 548 28543
rect 544 28534 582 28538
rect 544 28519 552 28534
rect 578 28519 582 28534
rect 544 28501 586 28519
rect 522 28495 608 28501
rect 182 28479 224 28495
rect 544 28479 586 28495
rect 17 28465 67 28467
rect 119 28465 169 28467
rect 186 28465 220 28479
rect 548 28465 582 28479
rect 599 28465 649 28467
rect 42 28423 59 28457
rect 67 28415 69 28465
rect 160 28457 246 28465
rect 522 28457 608 28465
rect 76 28423 110 28457
rect 127 28423 144 28457
rect 152 28423 161 28457
rect 162 28455 195 28457
rect 224 28455 244 28457
rect 162 28423 244 28455
rect 524 28455 548 28457
rect 573 28455 582 28457
rect 586 28455 606 28457
rect 160 28415 246 28423
rect 186 28399 220 28415
rect 182 28385 224 28386
rect 160 28379 182 28385
rect 224 28379 246 28385
rect 186 28344 220 28378
rect 223 28344 257 28378
rect 120 28331 170 28333
rect 76 28327 130 28331
rect 110 28322 130 28327
rect 60 28297 67 28307
rect 76 28297 77 28317
rect 96 28288 99 28322
rect 109 28297 110 28317
rect 119 28297 126 28307
rect 76 28281 92 28287
rect 94 28281 110 28287
rect 170 28281 172 28331
rect 186 28265 190 28299
rect 216 28265 220 28299
rect 288 28265 292 28453
rect 476 28385 480 28453
rect 524 28423 606 28455
rect 607 28423 616 28457
rect 522 28415 608 28423
rect 649 28415 651 28465
rect 548 28399 582 28415
rect 522 28380 548 28385
rect 522 28379 582 28380
rect 586 28379 608 28385
rect 295 28344 300 28378
rect 324 28344 329 28378
rect 544 28376 582 28379
rect 378 28339 450 28347
rect 428 28309 430 28325
rect 400 28301 430 28309
rect 476 28307 480 28375
rect 544 28346 552 28376
rect 578 28346 582 28376
rect 544 28337 548 28346
rect 400 28297 436 28301
rect 400 28267 408 28297
rect 420 28267 436 28297
rect 544 28299 548 28307
rect 12 28228 62 28230
rect 28 28219 59 28227
rect 62 28219 64 28228
rect 28 28211 64 28219
rect 127 28219 158 28227
rect 127 28212 182 28219
rect 215 28217 224 28245
rect 127 28211 161 28212
rect 59 28195 64 28211
rect 158 28195 161 28211
rect 28 28187 64 28195
rect 127 28194 161 28195
rect 127 28187 182 28194
rect 62 28178 64 28187
rect 213 28179 224 28217
rect 282 28207 292 28265
rect 296 28259 368 28267
rect 319 28229 346 28240
rect 318 28216 324 28229
rect 346 28216 348 28229
rect 428 28220 430 28267
rect 443 28257 450 28259
rect 476 28227 480 28295
rect 544 28265 552 28299
rect 578 28265 582 28299
rect 481 28233 517 28261
rect 481 28227 495 28233
rect 367 28216 380 28220
rect 251 28173 263 28207
rect 273 28173 293 28207
rect 295 28192 324 28216
rect 303 28182 316 28192
rect 318 28176 324 28192
rect 333 28192 380 28216
rect 333 28182 353 28192
rect 367 28186 380 28192
rect 396 28186 408 28220
rect 420 28186 436 28220
rect 120 28125 170 28127
rect 76 28119 92 28125
rect 94 28119 110 28125
rect 76 28109 99 28118
rect 60 28099 67 28109
rect 76 28089 77 28109
rect 96 28084 99 28109
rect 109 28089 110 28109
rect 119 28099 126 28109
rect 76 28075 110 28079
rect 170 28075 172 28125
rect 186 28107 190 28141
rect 216 28107 220 28141
rect 186 28030 220 28064
rect 282 28061 292 28173
rect 318 28166 335 28176
rect 318 28097 324 28166
rect 346 28097 348 28182
rect 428 28139 430 28186
rect 476 28149 480 28217
rect 485 28199 495 28227
rect 505 28227 519 28233
rect 544 28227 555 28265
rect 505 28199 525 28227
rect 544 28199 553 28227
rect 544 28179 548 28199
rect 579 28158 582 28248
rect 612 28230 624 28231
rect 599 28228 649 28230
rect 612 28227 624 28228
rect 610 28220 632 28227
rect 607 28219 632 28220
rect 586 28212 644 28219
rect 607 28211 644 28212
rect 607 28195 610 28211
rect 616 28195 644 28211
rect 607 28194 644 28195
rect 586 28187 644 28194
rect 607 28186 610 28187
rect 612 28179 632 28187
rect 612 28175 624 28179
rect 649 28178 651 28228
rect 544 28141 548 28149
rect 400 28109 408 28139
rect 420 28109 436 28139
rect 400 28105 436 28109
rect 400 28097 430 28105
rect 428 28081 430 28097
rect 476 28069 480 28137
rect 544 28107 552 28141
rect 578 28107 582 28141
rect 544 28099 548 28107
rect 544 28069 586 28070
rect 288 28029 292 28061
rect 296 28059 368 28067
rect 378 28059 450 28067
rect 544 28062 548 28069
rect 439 28031 444 28059
rect 120 28015 170 28017
rect 76 28011 130 28015
rect 110 28006 130 28011
rect 60 27981 67 27991
rect 76 27981 77 28001
rect 96 27972 99 28006
rect 109 27981 110 28001
rect 119 27981 126 27991
rect 76 27965 92 27971
rect 94 27965 110 27971
rect 170 27965 172 28015
rect 186 27949 190 27983
rect 216 27949 220 27983
rect 213 27917 224 27949
rect 282 27945 292 28029
rect 296 28023 368 28031
rect 378 28023 450 28031
rect 468 28028 473 28062
rect 428 27993 430 28009
rect 251 27917 292 27945
rect 318 27924 324 27993
rect 12 27912 62 27914
rect 28 27903 59 27911
rect 62 27903 64 27912
rect 251 27911 263 27917
rect 28 27895 64 27903
rect 127 27903 158 27911
rect 127 27896 182 27903
rect 127 27895 161 27896
rect 59 27879 64 27895
rect 158 27879 161 27895
rect 253 27883 263 27911
rect 273 27883 293 27917
rect 318 27914 335 27924
rect 303 27898 316 27908
rect 318 27898 324 27914
rect 346 27908 348 27993
rect 400 27985 430 27993
rect 476 27991 480 28059
rect 511 28028 582 28062
rect 544 28021 548 28028
rect 400 27981 436 27985
rect 400 27951 408 27981
rect 420 27951 436 27981
rect 544 27983 548 27991
rect 28 27871 64 27879
rect 127 27878 161 27879
rect 127 27871 182 27878
rect 62 27862 64 27871
rect 282 27825 292 27883
rect 295 27874 324 27898
rect 333 27898 353 27908
rect 428 27904 430 27951
rect 476 27911 480 27979
rect 544 27949 552 27983
rect 578 27949 582 27983
rect 544 27941 548 27949
rect 367 27898 380 27904
rect 333 27874 380 27898
rect 318 27861 324 27874
rect 346 27861 348 27874
rect 367 27870 380 27874
rect 396 27870 408 27904
rect 420 27870 436 27904
rect 544 27901 553 27929
rect 319 27850 346 27861
rect 120 27809 170 27811
rect 76 27803 92 27809
rect 94 27803 110 27809
rect 76 27793 99 27802
rect 60 27783 67 27793
rect 76 27773 77 27793
rect 96 27768 99 27793
rect 109 27773 110 27793
rect 119 27783 126 27793
rect 76 27759 110 27763
rect 170 27759 172 27809
rect 186 27791 190 27825
rect 216 27791 220 27825
rect 182 27753 224 27754
rect 186 27729 220 27746
rect 223 27729 257 27746
rect 182 27712 257 27729
rect 182 27711 224 27712
rect 160 27705 246 27711
rect 288 27705 292 27825
rect 296 27823 368 27831
rect 428 27823 430 27870
rect 476 27833 480 27901
rect 485 27857 495 27891
rect 505 27863 525 27891
rect 505 27857 519 27863
rect 544 27857 555 27901
rect 485 27833 492 27857
rect 579 27842 582 27932
rect 612 27914 624 27915
rect 599 27912 649 27914
rect 612 27911 624 27912
rect 610 27904 632 27911
rect 607 27903 632 27904
rect 586 27896 644 27903
rect 607 27895 644 27896
rect 607 27879 610 27895
rect 616 27879 644 27895
rect 607 27878 644 27879
rect 586 27871 644 27878
rect 607 27870 610 27871
rect 612 27863 632 27871
rect 612 27859 624 27863
rect 649 27862 651 27912
rect 544 27825 548 27833
rect 400 27793 408 27823
rect 420 27793 436 27823
rect 400 27789 436 27793
rect 400 27781 430 27789
rect 428 27765 430 27781
rect 476 27753 480 27821
rect 544 27791 552 27825
rect 578 27791 582 27825
rect 544 27783 548 27791
rect 295 27712 300 27746
rect 324 27712 329 27746
rect 378 27743 450 27751
rect 544 27748 548 27753
rect 544 27744 582 27748
rect 544 27729 552 27744
rect 578 27729 582 27744
rect 544 27711 586 27729
rect 522 27705 608 27711
rect 182 27689 224 27705
rect 544 27689 586 27705
rect 17 27675 67 27677
rect 119 27675 169 27677
rect 186 27675 220 27689
rect 548 27675 582 27689
rect 599 27675 649 27677
rect 42 27633 59 27667
rect 67 27625 69 27675
rect 160 27667 246 27675
rect 522 27667 608 27675
rect 76 27633 110 27667
rect 127 27633 144 27667
rect 152 27633 161 27667
rect 162 27665 195 27667
rect 224 27665 244 27667
rect 162 27633 244 27665
rect 524 27665 548 27667
rect 573 27665 582 27667
rect 586 27665 606 27667
rect 160 27625 246 27633
rect 186 27609 220 27625
rect 182 27595 224 27596
rect 160 27589 182 27595
rect 224 27589 246 27595
rect 186 27554 220 27588
rect 223 27554 257 27588
rect 120 27541 170 27543
rect 76 27537 130 27541
rect 110 27532 130 27537
rect 60 27507 67 27517
rect 76 27507 77 27527
rect 96 27498 99 27532
rect 109 27507 110 27527
rect 119 27507 126 27517
rect 76 27491 92 27497
rect 94 27491 110 27497
rect 170 27491 172 27541
rect 186 27475 190 27509
rect 216 27475 220 27509
rect 288 27475 292 27663
rect 476 27595 480 27663
rect 524 27633 606 27665
rect 607 27633 616 27667
rect 522 27625 608 27633
rect 649 27625 651 27675
rect 548 27609 582 27625
rect 522 27590 548 27595
rect 522 27589 582 27590
rect 586 27589 608 27595
rect 295 27554 300 27588
rect 324 27554 329 27588
rect 544 27586 582 27589
rect 378 27549 450 27557
rect 428 27519 430 27535
rect 400 27511 430 27519
rect 476 27517 480 27585
rect 544 27556 552 27586
rect 578 27556 582 27586
rect 544 27547 548 27556
rect 400 27507 436 27511
rect 400 27477 408 27507
rect 420 27477 436 27507
rect 544 27509 548 27517
rect 12 27438 62 27440
rect 28 27429 59 27437
rect 62 27429 64 27438
rect 28 27421 64 27429
rect 127 27429 158 27437
rect 127 27422 182 27429
rect 215 27427 224 27455
rect 127 27421 161 27422
rect 59 27405 64 27421
rect 158 27405 161 27421
rect 28 27397 64 27405
rect 127 27404 161 27405
rect 127 27397 182 27404
rect 62 27388 64 27397
rect 213 27389 224 27427
rect 282 27417 292 27475
rect 296 27469 368 27477
rect 319 27439 346 27450
rect 318 27426 324 27439
rect 346 27426 348 27439
rect 428 27430 430 27477
rect 443 27467 450 27469
rect 476 27437 480 27505
rect 544 27475 552 27509
rect 578 27475 582 27509
rect 481 27443 517 27471
rect 481 27437 495 27443
rect 367 27426 380 27430
rect 251 27383 263 27417
rect 273 27383 293 27417
rect 295 27402 324 27426
rect 303 27392 316 27402
rect 318 27386 324 27402
rect 333 27402 380 27426
rect 333 27392 353 27402
rect 367 27396 380 27402
rect 396 27396 408 27430
rect 420 27396 436 27430
rect 120 27335 170 27337
rect 76 27329 92 27335
rect 94 27329 110 27335
rect 76 27319 99 27328
rect 60 27309 67 27319
rect 76 27299 77 27319
rect 96 27294 99 27319
rect 109 27299 110 27319
rect 119 27309 126 27319
rect 76 27285 110 27289
rect 170 27285 172 27335
rect 186 27317 190 27351
rect 216 27317 220 27351
rect 186 27240 220 27274
rect 282 27271 292 27383
rect 318 27376 335 27386
rect 318 27307 324 27376
rect 346 27307 348 27392
rect 428 27349 430 27396
rect 476 27359 480 27427
rect 485 27409 495 27437
rect 505 27437 519 27443
rect 544 27437 555 27475
rect 505 27409 525 27437
rect 544 27409 553 27437
rect 544 27389 548 27409
rect 579 27368 582 27458
rect 612 27440 624 27441
rect 599 27438 649 27440
rect 612 27437 624 27438
rect 610 27430 632 27437
rect 607 27429 632 27430
rect 586 27422 644 27429
rect 607 27421 644 27422
rect 607 27405 610 27421
rect 616 27405 644 27421
rect 607 27404 644 27405
rect 586 27397 644 27404
rect 607 27396 610 27397
rect 612 27389 632 27397
rect 612 27385 624 27389
rect 649 27388 651 27438
rect 544 27351 548 27359
rect 400 27319 408 27349
rect 420 27319 436 27349
rect 400 27315 436 27319
rect 400 27307 430 27315
rect 428 27291 430 27307
rect 476 27279 480 27347
rect 544 27317 552 27351
rect 578 27317 582 27351
rect 544 27309 548 27317
rect 544 27279 586 27280
rect 288 27239 292 27271
rect 296 27269 368 27277
rect 378 27269 450 27277
rect 544 27272 548 27279
rect 439 27241 444 27269
rect 120 27225 170 27227
rect 76 27221 130 27225
rect 110 27216 130 27221
rect 60 27191 67 27201
rect 76 27191 77 27211
rect 96 27182 99 27216
rect 109 27191 110 27211
rect 119 27191 126 27201
rect 76 27175 92 27181
rect 94 27175 110 27181
rect 170 27175 172 27225
rect 186 27159 190 27193
rect 216 27159 220 27193
rect 213 27127 224 27159
rect 282 27155 292 27239
rect 296 27233 368 27241
rect 378 27233 450 27241
rect 468 27238 473 27272
rect 428 27203 430 27219
rect 251 27127 292 27155
rect 318 27134 324 27203
rect 12 27122 62 27124
rect 28 27113 59 27121
rect 62 27113 64 27122
rect 251 27121 263 27127
rect 28 27105 64 27113
rect 127 27113 158 27121
rect 127 27106 182 27113
rect 127 27105 161 27106
rect 59 27089 64 27105
rect 158 27089 161 27105
rect 253 27093 263 27121
rect 273 27093 293 27127
rect 318 27124 335 27134
rect 303 27108 316 27118
rect 318 27108 324 27124
rect 346 27118 348 27203
rect 400 27195 430 27203
rect 476 27201 480 27269
rect 511 27238 582 27272
rect 544 27231 548 27238
rect 400 27191 436 27195
rect 400 27161 408 27191
rect 420 27161 436 27191
rect 544 27193 548 27201
rect 28 27081 64 27089
rect 127 27088 161 27089
rect 127 27081 182 27088
rect 62 27072 64 27081
rect 282 27035 292 27093
rect 295 27084 324 27108
rect 333 27108 353 27118
rect 428 27114 430 27161
rect 476 27121 480 27189
rect 544 27159 552 27193
rect 578 27159 582 27193
rect 544 27151 548 27159
rect 367 27108 380 27114
rect 333 27084 380 27108
rect 318 27071 324 27084
rect 346 27071 348 27084
rect 367 27080 380 27084
rect 396 27080 408 27114
rect 420 27080 436 27114
rect 544 27111 553 27139
rect 319 27060 346 27071
rect 120 27019 170 27021
rect 76 27013 92 27019
rect 94 27013 110 27019
rect 76 27003 99 27012
rect 60 26993 67 27003
rect 76 26983 77 27003
rect 96 26978 99 27003
rect 109 26983 110 27003
rect 119 26993 126 27003
rect 76 26969 110 26973
rect 170 26969 172 27019
rect 186 27001 190 27035
rect 216 27001 220 27035
rect 182 26963 224 26964
rect 186 26939 220 26956
rect 223 26939 257 26956
rect 182 26922 257 26939
rect 182 26921 224 26922
rect 160 26915 246 26921
rect 288 26915 292 27035
rect 296 27033 368 27041
rect 428 27033 430 27080
rect 476 27043 480 27111
rect 485 27067 495 27101
rect 505 27073 525 27101
rect 505 27067 519 27073
rect 544 27067 555 27111
rect 485 27043 492 27067
rect 579 27052 582 27142
rect 612 27124 624 27125
rect 599 27122 649 27124
rect 612 27121 624 27122
rect 610 27114 632 27121
rect 607 27113 632 27114
rect 586 27106 644 27113
rect 607 27105 644 27106
rect 607 27089 610 27105
rect 616 27089 644 27105
rect 607 27088 644 27089
rect 586 27081 644 27088
rect 607 27080 610 27081
rect 612 27073 632 27081
rect 612 27069 624 27073
rect 649 27072 651 27122
rect 544 27035 548 27043
rect 400 27003 408 27033
rect 420 27003 436 27033
rect 400 26999 436 27003
rect 400 26991 430 26999
rect 428 26975 430 26991
rect 476 26963 480 27031
rect 544 27001 552 27035
rect 578 27001 582 27035
rect 544 26993 548 27001
rect 295 26922 300 26956
rect 324 26922 329 26956
rect 378 26953 450 26961
rect 544 26958 548 26963
rect 544 26954 582 26958
rect 544 26939 552 26954
rect 578 26939 582 26954
rect 544 26921 586 26939
rect 522 26915 608 26921
rect 182 26899 224 26915
rect 544 26899 586 26915
rect 17 26885 67 26887
rect 119 26885 169 26887
rect 186 26885 220 26899
rect 548 26885 582 26899
rect 599 26885 649 26887
rect 42 26843 59 26877
rect 67 26835 69 26885
rect 160 26877 246 26885
rect 522 26877 608 26885
rect 76 26843 110 26877
rect 127 26843 144 26877
rect 152 26843 161 26877
rect 162 26875 195 26877
rect 224 26875 244 26877
rect 162 26843 244 26875
rect 524 26875 548 26877
rect 573 26875 582 26877
rect 586 26875 606 26877
rect 160 26835 246 26843
rect 186 26819 220 26835
rect 182 26805 224 26806
rect 160 26799 182 26805
rect 224 26799 246 26805
rect 186 26764 220 26798
rect 223 26764 257 26798
rect 120 26751 170 26753
rect 76 26747 130 26751
rect 110 26742 130 26747
rect 60 26717 67 26727
rect 76 26717 77 26737
rect 96 26708 99 26742
rect 109 26717 110 26737
rect 119 26717 126 26727
rect 76 26701 92 26707
rect 94 26701 110 26707
rect 170 26701 172 26751
rect 186 26685 190 26719
rect 216 26685 220 26719
rect 288 26685 292 26873
rect 476 26805 480 26873
rect 524 26843 606 26875
rect 607 26843 616 26877
rect 522 26835 608 26843
rect 649 26835 651 26885
rect 548 26819 582 26835
rect 522 26800 548 26805
rect 522 26799 582 26800
rect 586 26799 608 26805
rect 295 26764 300 26798
rect 324 26764 329 26798
rect 544 26796 582 26799
rect 378 26759 450 26767
rect 428 26729 430 26745
rect 400 26721 430 26729
rect 476 26727 480 26795
rect 544 26766 552 26796
rect 578 26766 582 26796
rect 544 26757 548 26766
rect 400 26717 436 26721
rect 400 26687 408 26717
rect 420 26687 436 26717
rect 544 26719 548 26727
rect 12 26648 62 26650
rect 28 26639 59 26647
rect 62 26639 64 26648
rect 28 26631 64 26639
rect 127 26639 158 26647
rect 127 26632 182 26639
rect 215 26637 224 26665
rect 127 26631 161 26632
rect 59 26615 64 26631
rect 158 26615 161 26631
rect 28 26607 64 26615
rect 127 26614 161 26615
rect 127 26607 182 26614
rect 62 26598 64 26607
rect 213 26599 224 26637
rect 282 26627 292 26685
rect 296 26679 368 26687
rect 319 26649 346 26660
rect 318 26636 324 26649
rect 346 26636 348 26649
rect 428 26640 430 26687
rect 443 26677 450 26679
rect 476 26647 480 26715
rect 544 26685 552 26719
rect 578 26685 582 26719
rect 481 26653 517 26681
rect 481 26647 495 26653
rect 367 26636 380 26640
rect 251 26593 263 26627
rect 273 26593 293 26627
rect 295 26612 324 26636
rect 303 26602 316 26612
rect 318 26596 324 26612
rect 333 26612 380 26636
rect 333 26602 353 26612
rect 367 26606 380 26612
rect 396 26606 408 26640
rect 420 26606 436 26640
rect 120 26545 170 26547
rect 76 26539 92 26545
rect 94 26539 110 26545
rect 76 26529 99 26538
rect 60 26519 67 26529
rect 76 26509 77 26529
rect 96 26504 99 26529
rect 109 26509 110 26529
rect 119 26519 126 26529
rect 76 26495 110 26499
rect 170 26495 172 26545
rect 186 26527 190 26561
rect 216 26527 220 26561
rect 186 26450 220 26484
rect 282 26481 292 26593
rect 318 26586 335 26596
rect 318 26517 324 26586
rect 346 26517 348 26602
rect 428 26559 430 26606
rect 476 26569 480 26637
rect 485 26619 495 26647
rect 505 26647 519 26653
rect 544 26647 555 26685
rect 505 26619 525 26647
rect 544 26619 553 26647
rect 544 26599 548 26619
rect 579 26578 582 26668
rect 612 26650 624 26651
rect 599 26648 649 26650
rect 612 26647 624 26648
rect 610 26640 632 26647
rect 607 26639 632 26640
rect 586 26632 644 26639
rect 607 26631 644 26632
rect 607 26615 610 26631
rect 616 26615 644 26631
rect 607 26614 644 26615
rect 586 26607 644 26614
rect 607 26606 610 26607
rect 612 26599 632 26607
rect 612 26595 624 26599
rect 649 26598 651 26648
rect 544 26561 548 26569
rect 400 26529 408 26559
rect 420 26529 436 26559
rect 400 26525 436 26529
rect 400 26517 430 26525
rect 428 26501 430 26517
rect 476 26489 480 26557
rect 544 26527 552 26561
rect 578 26527 582 26561
rect 544 26519 548 26527
rect 544 26489 586 26490
rect 288 26449 292 26481
rect 296 26479 368 26487
rect 378 26479 450 26487
rect 544 26482 548 26489
rect 439 26451 444 26479
rect 120 26435 170 26437
rect 76 26431 130 26435
rect 110 26426 130 26431
rect 60 26401 67 26411
rect 76 26401 77 26421
rect 96 26392 99 26426
rect 109 26401 110 26421
rect 119 26401 126 26411
rect 76 26385 92 26391
rect 94 26385 110 26391
rect 170 26385 172 26435
rect 186 26369 190 26403
rect 216 26369 220 26403
rect 213 26337 224 26369
rect 282 26365 292 26449
rect 296 26443 368 26451
rect 378 26443 450 26451
rect 468 26448 473 26482
rect 428 26413 430 26429
rect 251 26337 292 26365
rect 318 26344 324 26413
rect 12 26332 62 26334
rect 28 26323 59 26331
rect 62 26323 64 26332
rect 251 26331 263 26337
rect 28 26315 64 26323
rect 127 26323 158 26331
rect 127 26316 182 26323
rect 127 26315 161 26316
rect 59 26299 64 26315
rect 158 26299 161 26315
rect 253 26303 263 26331
rect 273 26303 293 26337
rect 318 26334 335 26344
rect 303 26318 316 26328
rect 318 26318 324 26334
rect 346 26328 348 26413
rect 400 26405 430 26413
rect 476 26411 480 26479
rect 511 26448 582 26482
rect 544 26441 548 26448
rect 400 26401 436 26405
rect 400 26371 408 26401
rect 420 26371 436 26401
rect 544 26403 548 26411
rect 28 26291 64 26299
rect 127 26298 161 26299
rect 127 26291 182 26298
rect 62 26282 64 26291
rect 282 26245 292 26303
rect 295 26294 324 26318
rect 333 26318 353 26328
rect 428 26324 430 26371
rect 476 26331 480 26399
rect 544 26369 552 26403
rect 578 26369 582 26403
rect 544 26361 548 26369
rect 367 26318 380 26324
rect 333 26294 380 26318
rect 318 26281 324 26294
rect 346 26281 348 26294
rect 367 26290 380 26294
rect 396 26290 408 26324
rect 420 26290 436 26324
rect 544 26321 553 26349
rect 319 26270 346 26281
rect 120 26229 170 26231
rect 76 26223 92 26229
rect 94 26223 110 26229
rect 76 26213 99 26222
rect 60 26203 67 26213
rect 76 26193 77 26213
rect 96 26188 99 26213
rect 109 26193 110 26213
rect 119 26203 126 26213
rect 76 26179 110 26183
rect 170 26179 172 26229
rect 186 26211 190 26245
rect 216 26211 220 26245
rect 182 26173 224 26174
rect 186 26149 220 26166
rect 223 26149 257 26166
rect 182 26132 257 26149
rect 182 26131 224 26132
rect 160 26125 246 26131
rect 288 26125 292 26245
rect 296 26243 368 26251
rect 428 26243 430 26290
rect 476 26253 480 26321
rect 485 26277 495 26311
rect 505 26283 525 26311
rect 505 26277 519 26283
rect 544 26277 555 26321
rect 485 26253 492 26277
rect 579 26262 582 26352
rect 612 26334 624 26335
rect 599 26332 649 26334
rect 612 26331 624 26332
rect 610 26324 632 26331
rect 607 26323 632 26324
rect 586 26316 644 26323
rect 607 26315 644 26316
rect 607 26299 610 26315
rect 616 26299 644 26315
rect 607 26298 644 26299
rect 586 26291 644 26298
rect 607 26290 610 26291
rect 612 26283 632 26291
rect 612 26279 624 26283
rect 649 26282 651 26332
rect 544 26245 548 26253
rect 400 26213 408 26243
rect 420 26213 436 26243
rect 400 26209 436 26213
rect 400 26201 430 26209
rect 428 26185 430 26201
rect 476 26173 480 26241
rect 544 26211 552 26245
rect 578 26211 582 26245
rect 544 26203 548 26211
rect 295 26132 300 26166
rect 324 26132 329 26166
rect 378 26163 450 26171
rect 544 26168 548 26173
rect 544 26164 582 26168
rect 544 26149 552 26164
rect 578 26149 582 26164
rect 544 26131 586 26149
rect 522 26125 608 26131
rect 182 26109 224 26125
rect 544 26109 586 26125
rect 17 26095 67 26097
rect 119 26095 169 26097
rect 186 26095 220 26109
rect 548 26095 582 26109
rect 599 26095 649 26097
rect 42 26053 59 26087
rect 67 26045 69 26095
rect 160 26087 246 26095
rect 522 26087 608 26095
rect 76 26053 110 26087
rect 127 26053 144 26087
rect 152 26053 161 26087
rect 162 26085 195 26087
rect 224 26085 244 26087
rect 162 26053 244 26085
rect 524 26085 548 26087
rect 573 26085 582 26087
rect 586 26085 606 26087
rect 160 26045 246 26053
rect 186 26029 220 26045
rect 182 26015 224 26016
rect 160 26009 182 26015
rect 224 26009 246 26015
rect 186 25974 220 26008
rect 223 25974 257 26008
rect 120 25961 170 25963
rect 76 25957 130 25961
rect 110 25952 130 25957
rect 60 25927 67 25937
rect 76 25927 77 25947
rect 96 25918 99 25952
rect 109 25927 110 25947
rect 119 25927 126 25937
rect 76 25911 92 25917
rect 94 25911 110 25917
rect 170 25911 172 25961
rect 186 25895 190 25929
rect 216 25895 220 25929
rect 288 25895 292 26083
rect 476 26015 480 26083
rect 524 26053 606 26085
rect 607 26053 616 26087
rect 522 26045 608 26053
rect 649 26045 651 26095
rect 548 26029 582 26045
rect 522 26010 548 26015
rect 522 26009 582 26010
rect 586 26009 608 26015
rect 295 25974 300 26008
rect 324 25974 329 26008
rect 544 26006 582 26009
rect 378 25969 450 25977
rect 428 25939 430 25955
rect 400 25931 430 25939
rect 476 25937 480 26005
rect 544 25976 552 26006
rect 578 25976 582 26006
rect 544 25967 548 25976
rect 400 25927 436 25931
rect 400 25897 408 25927
rect 420 25897 436 25927
rect 544 25929 548 25937
rect 12 25858 62 25860
rect 28 25849 59 25857
rect 62 25849 64 25858
rect 28 25841 64 25849
rect 127 25849 158 25857
rect 127 25842 182 25849
rect 215 25847 224 25875
rect 127 25841 161 25842
rect 59 25825 64 25841
rect 158 25825 161 25841
rect 28 25817 64 25825
rect 127 25824 161 25825
rect 127 25817 182 25824
rect 62 25808 64 25817
rect 213 25809 224 25847
rect 282 25837 292 25895
rect 296 25889 368 25897
rect 319 25859 346 25870
rect 318 25846 324 25859
rect 346 25846 348 25859
rect 428 25850 430 25897
rect 443 25887 450 25889
rect 476 25857 480 25925
rect 544 25895 552 25929
rect 578 25895 582 25929
rect 481 25863 517 25891
rect 481 25857 495 25863
rect 367 25846 380 25850
rect 251 25803 263 25837
rect 273 25803 293 25837
rect 295 25822 324 25846
rect 303 25812 316 25822
rect 318 25806 324 25822
rect 333 25822 380 25846
rect 333 25812 353 25822
rect 367 25816 380 25822
rect 396 25816 408 25850
rect 420 25816 436 25850
rect 120 25755 170 25757
rect 76 25749 92 25755
rect 94 25749 110 25755
rect 76 25739 99 25748
rect 60 25729 67 25739
rect 76 25719 77 25739
rect 96 25714 99 25739
rect 109 25719 110 25739
rect 119 25729 126 25739
rect 76 25705 110 25709
rect 170 25705 172 25755
rect 186 25737 190 25771
rect 216 25737 220 25771
rect 186 25660 220 25694
rect 282 25691 292 25803
rect 318 25796 335 25806
rect 318 25727 324 25796
rect 346 25727 348 25812
rect 428 25769 430 25816
rect 476 25779 480 25847
rect 485 25829 495 25857
rect 505 25857 519 25863
rect 544 25857 555 25895
rect 505 25829 525 25857
rect 544 25829 553 25857
rect 544 25809 548 25829
rect 579 25788 582 25878
rect 612 25860 624 25861
rect 599 25858 649 25860
rect 612 25857 624 25858
rect 610 25850 632 25857
rect 607 25849 632 25850
rect 586 25842 644 25849
rect 607 25841 644 25842
rect 607 25825 610 25841
rect 616 25825 644 25841
rect 607 25824 644 25825
rect 586 25817 644 25824
rect 607 25816 610 25817
rect 612 25809 632 25817
rect 612 25805 624 25809
rect 649 25808 651 25858
rect 544 25771 548 25779
rect 400 25739 408 25769
rect 420 25739 436 25769
rect 400 25735 436 25739
rect 400 25727 430 25735
rect 428 25711 430 25727
rect 476 25699 480 25767
rect 544 25737 552 25771
rect 578 25737 582 25771
rect 544 25729 548 25737
rect 544 25699 586 25700
rect 288 25659 292 25691
rect 296 25689 368 25697
rect 378 25689 450 25697
rect 544 25692 548 25699
rect 439 25661 444 25689
rect 120 25645 170 25647
rect 76 25641 130 25645
rect 110 25636 130 25641
rect 60 25611 67 25621
rect 76 25611 77 25631
rect 96 25602 99 25636
rect 109 25611 110 25631
rect 119 25611 126 25621
rect 76 25595 92 25601
rect 94 25595 110 25601
rect 170 25595 172 25645
rect 186 25579 190 25613
rect 216 25579 220 25613
rect 213 25547 224 25579
rect 282 25575 292 25659
rect 296 25653 368 25661
rect 378 25653 450 25661
rect 468 25658 473 25692
rect 428 25623 430 25639
rect 251 25547 292 25575
rect 318 25554 324 25623
rect 12 25542 62 25544
rect 28 25533 59 25541
rect 62 25533 64 25542
rect 251 25541 263 25547
rect 28 25525 64 25533
rect 127 25533 158 25541
rect 127 25526 182 25533
rect 127 25525 161 25526
rect 59 25509 64 25525
rect 158 25509 161 25525
rect 253 25513 263 25541
rect 273 25513 293 25547
rect 318 25544 335 25554
rect 303 25528 316 25538
rect 318 25528 324 25544
rect 346 25538 348 25623
rect 400 25615 430 25623
rect 476 25621 480 25689
rect 511 25658 582 25692
rect 544 25651 548 25658
rect 400 25611 436 25615
rect 400 25581 408 25611
rect 420 25581 436 25611
rect 544 25613 548 25621
rect 28 25501 64 25509
rect 127 25508 161 25509
rect 127 25501 182 25508
rect 62 25492 64 25501
rect 282 25455 292 25513
rect 295 25504 324 25528
rect 333 25528 353 25538
rect 428 25534 430 25581
rect 476 25541 480 25609
rect 544 25579 552 25613
rect 578 25579 582 25613
rect 544 25571 548 25579
rect 367 25528 380 25534
rect 333 25504 380 25528
rect 318 25491 324 25504
rect 346 25491 348 25504
rect 367 25500 380 25504
rect 396 25500 408 25534
rect 420 25500 436 25534
rect 544 25531 553 25559
rect 319 25480 346 25491
rect 120 25439 170 25441
rect 76 25433 92 25439
rect 94 25433 110 25439
rect 76 25423 99 25432
rect 60 25413 67 25423
rect 76 25403 77 25423
rect 96 25398 99 25423
rect 109 25403 110 25423
rect 119 25413 126 25423
rect 76 25389 110 25393
rect 170 25389 172 25439
rect 186 25421 190 25455
rect 216 25421 220 25455
rect 182 25383 224 25384
rect 186 25359 220 25376
rect 223 25359 257 25376
rect 182 25342 257 25359
rect 182 25341 224 25342
rect 160 25335 246 25341
rect 288 25335 292 25455
rect 296 25453 368 25461
rect 428 25453 430 25500
rect 476 25463 480 25531
rect 485 25487 495 25521
rect 505 25493 525 25521
rect 505 25487 519 25493
rect 544 25487 555 25531
rect 485 25463 492 25487
rect 579 25472 582 25562
rect 612 25544 624 25545
rect 599 25542 649 25544
rect 612 25541 624 25542
rect 610 25534 632 25541
rect 607 25533 632 25534
rect 586 25526 644 25533
rect 607 25525 644 25526
rect 607 25509 610 25525
rect 616 25509 644 25525
rect 607 25508 644 25509
rect 586 25501 644 25508
rect 607 25500 610 25501
rect 612 25493 632 25501
rect 612 25489 624 25493
rect 649 25492 651 25542
rect 544 25455 548 25463
rect 400 25423 408 25453
rect 420 25423 436 25453
rect 400 25419 436 25423
rect 400 25411 430 25419
rect 428 25395 430 25411
rect 476 25383 480 25451
rect 544 25421 552 25455
rect 578 25421 582 25455
rect 544 25413 548 25421
rect 295 25342 300 25376
rect 324 25342 329 25376
rect 378 25373 450 25381
rect 544 25378 548 25383
rect 544 25374 582 25378
rect 544 25359 552 25374
rect 578 25359 582 25374
rect 544 25341 586 25359
rect 522 25335 608 25341
rect 182 25319 224 25335
rect 544 25319 586 25335
rect 17 25305 67 25307
rect 119 25305 169 25307
rect 186 25305 220 25319
rect 548 25305 582 25319
rect 599 25305 649 25307
rect 42 25263 59 25297
rect 67 25255 69 25305
rect 160 25297 246 25305
rect 522 25297 608 25305
rect 76 25263 110 25297
rect 127 25263 144 25297
rect 152 25263 161 25297
rect 162 25295 195 25297
rect 224 25295 244 25297
rect 162 25263 244 25295
rect 524 25295 548 25297
rect 573 25295 582 25297
rect 586 25295 606 25297
rect 160 25255 246 25263
rect 186 25239 220 25255
rect 182 25225 224 25226
rect 160 25219 182 25225
rect 224 25219 246 25225
rect 186 25184 220 25218
rect 223 25184 257 25218
rect 120 25171 170 25173
rect 76 25167 130 25171
rect 110 25162 130 25167
rect 60 25137 67 25147
rect 76 25137 77 25157
rect 96 25128 99 25162
rect 109 25137 110 25157
rect 119 25137 126 25147
rect 76 25121 92 25127
rect 94 25121 110 25127
rect 170 25121 172 25171
rect 186 25105 190 25139
rect 216 25105 220 25139
rect 288 25105 292 25293
rect 476 25225 480 25293
rect 524 25263 606 25295
rect 607 25263 616 25297
rect 522 25255 608 25263
rect 649 25255 651 25305
rect 548 25239 582 25255
rect 522 25220 548 25225
rect 522 25219 582 25220
rect 586 25219 608 25225
rect 295 25184 300 25218
rect 324 25184 329 25218
rect 544 25216 582 25219
rect 378 25179 450 25187
rect 428 25149 430 25165
rect 400 25141 430 25149
rect 476 25147 480 25215
rect 544 25186 552 25216
rect 578 25186 582 25216
rect 544 25177 548 25186
rect 400 25137 436 25141
rect 400 25107 408 25137
rect 420 25107 436 25137
rect 544 25139 548 25147
rect 12 25068 62 25070
rect 28 25059 59 25067
rect 62 25059 64 25068
rect 28 25051 64 25059
rect 127 25059 158 25067
rect 127 25052 182 25059
rect 215 25057 224 25085
rect 127 25051 161 25052
rect 59 25035 64 25051
rect 158 25035 161 25051
rect 28 25027 64 25035
rect 127 25034 161 25035
rect 127 25027 182 25034
rect 62 25018 64 25027
rect 213 25019 224 25057
rect 282 25047 292 25105
rect 296 25099 368 25107
rect 319 25069 346 25080
rect 318 25056 324 25069
rect 346 25056 348 25069
rect 428 25060 430 25107
rect 443 25097 450 25099
rect 476 25067 480 25135
rect 544 25105 552 25139
rect 578 25105 582 25139
rect 481 25073 517 25101
rect 481 25067 495 25073
rect 367 25056 380 25060
rect 251 25013 263 25047
rect 273 25013 293 25047
rect 295 25032 324 25056
rect 303 25022 316 25032
rect 318 25016 324 25032
rect 333 25032 380 25056
rect 333 25022 353 25032
rect 367 25026 380 25032
rect 396 25026 408 25060
rect 420 25026 436 25060
rect 120 24965 170 24967
rect 76 24959 92 24965
rect 94 24959 110 24965
rect 76 24949 99 24958
rect 60 24939 67 24949
rect 76 24929 77 24949
rect 96 24924 99 24949
rect 109 24929 110 24949
rect 119 24939 126 24949
rect 76 24915 110 24919
rect 170 24915 172 24965
rect 186 24947 190 24981
rect 216 24947 220 24981
rect 186 24870 220 24904
rect 282 24901 292 25013
rect 318 25006 335 25016
rect 318 24937 324 25006
rect 346 24937 348 25022
rect 428 24979 430 25026
rect 476 24989 480 25057
rect 485 25039 495 25067
rect 505 25067 519 25073
rect 544 25067 555 25105
rect 505 25039 525 25067
rect 544 25039 553 25067
rect 544 25019 548 25039
rect 579 24998 582 25088
rect 612 25070 624 25071
rect 599 25068 649 25070
rect 612 25067 624 25068
rect 610 25060 632 25067
rect 607 25059 632 25060
rect 586 25052 644 25059
rect 607 25051 644 25052
rect 607 25035 610 25051
rect 616 25035 644 25051
rect 607 25034 644 25035
rect 586 25027 644 25034
rect 607 25026 610 25027
rect 612 25019 632 25027
rect 612 25015 624 25019
rect 649 25018 651 25068
rect 544 24981 548 24989
rect 400 24949 408 24979
rect 420 24949 436 24979
rect 400 24945 436 24949
rect 400 24937 430 24945
rect 428 24921 430 24937
rect 476 24909 480 24977
rect 544 24947 552 24981
rect 578 24947 582 24981
rect 544 24939 548 24947
rect 544 24909 586 24910
rect 288 24869 292 24901
rect 296 24899 368 24907
rect 378 24899 450 24907
rect 544 24902 548 24909
rect 439 24871 444 24899
rect 120 24855 170 24857
rect 76 24851 130 24855
rect 110 24846 130 24851
rect 60 24821 67 24831
rect 76 24821 77 24841
rect 96 24812 99 24846
rect 109 24821 110 24841
rect 119 24821 126 24831
rect 76 24805 92 24811
rect 94 24805 110 24811
rect 170 24805 172 24855
rect 186 24789 190 24823
rect 216 24789 220 24823
rect 213 24757 224 24789
rect 282 24785 292 24869
rect 296 24863 368 24871
rect 378 24863 450 24871
rect 468 24868 473 24902
rect 428 24833 430 24849
rect 251 24757 292 24785
rect 318 24764 324 24833
rect 12 24752 62 24754
rect 28 24743 59 24751
rect 62 24743 64 24752
rect 251 24751 263 24757
rect 28 24735 64 24743
rect 127 24743 158 24751
rect 127 24736 182 24743
rect 127 24735 161 24736
rect 59 24719 64 24735
rect 158 24719 161 24735
rect 253 24723 263 24751
rect 273 24723 293 24757
rect 318 24754 335 24764
rect 303 24738 316 24748
rect 318 24738 324 24754
rect 346 24748 348 24833
rect 400 24825 430 24833
rect 476 24831 480 24899
rect 511 24868 582 24902
rect 544 24861 548 24868
rect 400 24821 436 24825
rect 400 24791 408 24821
rect 420 24791 436 24821
rect 544 24823 548 24831
rect 28 24711 64 24719
rect 127 24718 161 24719
rect 127 24711 182 24718
rect 62 24702 64 24711
rect 282 24665 292 24723
rect 295 24714 324 24738
rect 333 24738 353 24748
rect 428 24744 430 24791
rect 476 24751 480 24819
rect 544 24789 552 24823
rect 578 24789 582 24823
rect 544 24781 548 24789
rect 367 24738 380 24744
rect 333 24714 380 24738
rect 318 24701 324 24714
rect 346 24701 348 24714
rect 367 24710 380 24714
rect 396 24710 408 24744
rect 420 24710 436 24744
rect 544 24741 553 24769
rect 319 24690 346 24701
rect 120 24649 170 24651
rect 76 24643 92 24649
rect 94 24643 110 24649
rect 76 24633 99 24642
rect 60 24623 67 24633
rect 76 24613 77 24633
rect 96 24608 99 24633
rect 109 24613 110 24633
rect 119 24623 126 24633
rect 76 24599 110 24603
rect 170 24599 172 24649
rect 186 24631 190 24665
rect 216 24631 220 24665
rect 182 24593 224 24594
rect 186 24569 220 24586
rect 223 24569 257 24586
rect 182 24552 257 24569
rect 182 24551 224 24552
rect 160 24545 246 24551
rect 288 24545 292 24665
rect 296 24663 368 24671
rect 428 24663 430 24710
rect 476 24673 480 24741
rect 485 24697 495 24731
rect 505 24703 525 24731
rect 505 24697 519 24703
rect 544 24697 555 24741
rect 485 24673 492 24697
rect 579 24682 582 24772
rect 612 24754 624 24755
rect 599 24752 649 24754
rect 612 24751 624 24752
rect 610 24744 632 24751
rect 607 24743 632 24744
rect 586 24736 644 24743
rect 607 24735 644 24736
rect 607 24719 610 24735
rect 616 24719 644 24735
rect 607 24718 644 24719
rect 586 24711 644 24718
rect 607 24710 610 24711
rect 612 24703 632 24711
rect 612 24699 624 24703
rect 649 24702 651 24752
rect 544 24665 548 24673
rect 400 24633 408 24663
rect 420 24633 436 24663
rect 400 24629 436 24633
rect 400 24621 430 24629
rect 428 24605 430 24621
rect 476 24593 480 24661
rect 544 24631 552 24665
rect 578 24631 582 24665
rect 544 24623 548 24631
rect 295 24552 300 24586
rect 324 24552 329 24586
rect 378 24583 450 24591
rect 544 24588 548 24593
rect 544 24584 582 24588
rect 544 24569 552 24584
rect 578 24569 582 24584
rect 544 24551 586 24569
rect 522 24545 608 24551
rect 182 24529 224 24545
rect 544 24529 586 24545
rect 17 24515 67 24517
rect 119 24515 169 24517
rect 186 24515 220 24529
rect 548 24515 582 24529
rect 599 24515 649 24517
rect 42 24473 59 24507
rect 67 24465 69 24515
rect 160 24507 246 24515
rect 522 24507 608 24515
rect 76 24473 110 24507
rect 127 24473 144 24507
rect 152 24473 161 24507
rect 162 24505 195 24507
rect 224 24505 244 24507
rect 162 24473 244 24505
rect 524 24505 548 24507
rect 573 24505 582 24507
rect 586 24505 606 24507
rect 160 24465 246 24473
rect 186 24449 220 24465
rect 182 24435 224 24436
rect 160 24429 182 24435
rect 224 24429 246 24435
rect 186 24394 220 24428
rect 223 24394 257 24428
rect 120 24381 170 24383
rect 76 24377 130 24381
rect 110 24372 130 24377
rect 60 24347 67 24357
rect 76 24347 77 24367
rect 96 24338 99 24372
rect 109 24347 110 24367
rect 119 24347 126 24357
rect 76 24331 92 24337
rect 94 24331 110 24337
rect 170 24331 172 24381
rect 186 24315 190 24349
rect 216 24315 220 24349
rect 288 24315 292 24503
rect 476 24435 480 24503
rect 524 24473 606 24505
rect 607 24473 616 24507
rect 522 24465 608 24473
rect 649 24465 651 24515
rect 548 24449 582 24465
rect 522 24430 548 24435
rect 522 24429 582 24430
rect 586 24429 608 24435
rect 295 24394 300 24428
rect 324 24394 329 24428
rect 544 24426 582 24429
rect 378 24389 450 24397
rect 428 24359 430 24375
rect 400 24351 430 24359
rect 476 24357 480 24425
rect 544 24396 552 24426
rect 578 24396 582 24426
rect 544 24387 548 24396
rect 400 24347 436 24351
rect 400 24317 408 24347
rect 420 24317 436 24347
rect 544 24349 548 24357
rect 12 24278 62 24280
rect 28 24269 59 24277
rect 62 24269 64 24278
rect 28 24261 64 24269
rect 127 24269 158 24277
rect 127 24262 182 24269
rect 215 24267 224 24295
rect 127 24261 161 24262
rect 59 24245 64 24261
rect 158 24245 161 24261
rect 28 24237 64 24245
rect 127 24244 161 24245
rect 127 24237 182 24244
rect 62 24228 64 24237
rect 213 24229 224 24267
rect 282 24257 292 24315
rect 296 24309 368 24317
rect 319 24279 346 24290
rect 318 24266 324 24279
rect 346 24266 348 24279
rect 428 24270 430 24317
rect 443 24307 450 24309
rect 476 24277 480 24345
rect 544 24315 552 24349
rect 578 24315 582 24349
rect 481 24283 517 24311
rect 481 24277 495 24283
rect 367 24266 380 24270
rect 251 24223 263 24257
rect 273 24223 293 24257
rect 295 24242 324 24266
rect 303 24232 316 24242
rect 318 24226 324 24242
rect 333 24242 380 24266
rect 333 24232 353 24242
rect 367 24236 380 24242
rect 396 24236 408 24270
rect 420 24236 436 24270
rect 120 24175 170 24177
rect 76 24169 92 24175
rect 94 24169 110 24175
rect 76 24159 99 24168
rect 60 24149 67 24159
rect 76 24139 77 24159
rect 96 24134 99 24159
rect 109 24139 110 24159
rect 119 24149 126 24159
rect 76 24125 110 24129
rect 170 24125 172 24175
rect 186 24157 190 24191
rect 216 24157 220 24191
rect 186 24080 220 24114
rect 282 24111 292 24223
rect 318 24216 335 24226
rect 318 24147 324 24216
rect 346 24147 348 24232
rect 428 24189 430 24236
rect 476 24199 480 24267
rect 485 24249 495 24277
rect 505 24277 519 24283
rect 544 24277 555 24315
rect 505 24249 525 24277
rect 544 24249 553 24277
rect 544 24229 548 24249
rect 579 24208 582 24298
rect 612 24280 624 24281
rect 599 24278 649 24280
rect 612 24277 624 24278
rect 610 24270 632 24277
rect 607 24269 632 24270
rect 586 24262 644 24269
rect 607 24261 644 24262
rect 607 24245 610 24261
rect 616 24245 644 24261
rect 607 24244 644 24245
rect 586 24237 644 24244
rect 607 24236 610 24237
rect 612 24229 632 24237
rect 612 24225 624 24229
rect 649 24228 651 24278
rect 544 24191 548 24199
rect 400 24159 408 24189
rect 420 24159 436 24189
rect 400 24155 436 24159
rect 400 24147 430 24155
rect 428 24131 430 24147
rect 476 24119 480 24187
rect 544 24157 552 24191
rect 578 24157 582 24191
rect 544 24149 548 24157
rect 544 24119 586 24120
rect 288 24079 292 24111
rect 296 24109 368 24117
rect 378 24109 450 24117
rect 544 24112 548 24119
rect 439 24081 444 24109
rect 120 24065 170 24067
rect 76 24061 130 24065
rect 110 24056 130 24061
rect 60 24031 67 24041
rect 76 24031 77 24051
rect 96 24022 99 24056
rect 109 24031 110 24051
rect 119 24031 126 24041
rect 76 24015 92 24021
rect 94 24015 110 24021
rect 170 24015 172 24065
rect 186 23999 190 24033
rect 216 23999 220 24033
rect 213 23967 224 23999
rect 282 23995 292 24079
rect 296 24073 368 24081
rect 378 24073 450 24081
rect 468 24078 473 24112
rect 428 24043 430 24059
rect 251 23967 292 23995
rect 318 23974 324 24043
rect 12 23962 62 23964
rect 28 23953 59 23961
rect 62 23953 64 23962
rect 251 23961 263 23967
rect 28 23945 64 23953
rect 127 23953 158 23961
rect 127 23946 182 23953
rect 127 23945 161 23946
rect 59 23929 64 23945
rect 158 23929 161 23945
rect 253 23933 263 23961
rect 273 23933 293 23967
rect 318 23964 335 23974
rect 303 23948 316 23958
rect 318 23948 324 23964
rect 346 23958 348 24043
rect 400 24035 430 24043
rect 476 24041 480 24109
rect 511 24078 582 24112
rect 544 24071 548 24078
rect 400 24031 436 24035
rect 400 24001 408 24031
rect 420 24001 436 24031
rect 544 24033 548 24041
rect 28 23921 64 23929
rect 127 23928 161 23929
rect 127 23921 182 23928
rect 62 23912 64 23921
rect 282 23875 292 23933
rect 295 23924 324 23948
rect 333 23948 353 23958
rect 428 23954 430 24001
rect 476 23961 480 24029
rect 544 23999 552 24033
rect 578 23999 582 24033
rect 544 23991 548 23999
rect 367 23948 380 23954
rect 333 23924 380 23948
rect 318 23911 324 23924
rect 346 23911 348 23924
rect 367 23920 380 23924
rect 396 23920 408 23954
rect 420 23920 436 23954
rect 544 23951 553 23979
rect 319 23900 346 23911
rect 120 23859 170 23861
rect 76 23853 92 23859
rect 94 23853 110 23859
rect 76 23843 99 23852
rect 60 23833 67 23843
rect 76 23823 77 23843
rect 96 23818 99 23843
rect 109 23823 110 23843
rect 119 23833 126 23843
rect 76 23809 110 23813
rect 170 23809 172 23859
rect 186 23841 190 23875
rect 216 23841 220 23875
rect 182 23803 224 23804
rect 186 23779 220 23796
rect 223 23779 257 23796
rect 182 23762 257 23779
rect 182 23761 224 23762
rect 160 23755 246 23761
rect 288 23755 292 23875
rect 296 23873 368 23881
rect 428 23873 430 23920
rect 476 23883 480 23951
rect 485 23907 495 23941
rect 505 23913 525 23941
rect 505 23907 519 23913
rect 544 23907 555 23951
rect 485 23883 492 23907
rect 579 23892 582 23982
rect 612 23964 624 23965
rect 599 23962 649 23964
rect 612 23961 624 23962
rect 610 23954 632 23961
rect 607 23953 632 23954
rect 586 23946 644 23953
rect 607 23945 644 23946
rect 607 23929 610 23945
rect 616 23929 644 23945
rect 607 23928 644 23929
rect 586 23921 644 23928
rect 607 23920 610 23921
rect 612 23913 632 23921
rect 612 23909 624 23913
rect 649 23912 651 23962
rect 544 23875 548 23883
rect 400 23843 408 23873
rect 420 23843 436 23873
rect 400 23839 436 23843
rect 400 23831 430 23839
rect 428 23815 430 23831
rect 476 23803 480 23871
rect 544 23841 552 23875
rect 578 23841 582 23875
rect 544 23833 548 23841
rect 295 23762 300 23796
rect 324 23762 329 23796
rect 378 23793 450 23801
rect 544 23798 548 23803
rect 544 23794 582 23798
rect 544 23779 552 23794
rect 578 23779 582 23794
rect 544 23761 586 23779
rect 522 23755 608 23761
rect 182 23739 224 23755
rect 544 23739 586 23755
rect 17 23725 67 23727
rect 119 23725 169 23727
rect 186 23725 220 23739
rect 548 23725 582 23739
rect 599 23725 649 23727
rect 42 23683 59 23717
rect 67 23675 69 23725
rect 160 23717 246 23725
rect 522 23717 608 23725
rect 76 23683 110 23717
rect 127 23683 144 23717
rect 152 23683 161 23717
rect 162 23715 195 23717
rect 224 23715 244 23717
rect 162 23683 244 23715
rect 524 23715 548 23717
rect 573 23715 582 23717
rect 586 23715 606 23717
rect 160 23675 246 23683
rect 186 23659 220 23675
rect 182 23645 224 23646
rect 160 23639 182 23645
rect 224 23639 246 23645
rect 186 23604 220 23638
rect 223 23604 257 23638
rect 120 23591 170 23593
rect 76 23587 130 23591
rect 110 23582 130 23587
rect 60 23557 67 23567
rect 76 23557 77 23577
rect 96 23548 99 23582
rect 109 23557 110 23577
rect 119 23557 126 23567
rect 76 23541 92 23547
rect 94 23541 110 23547
rect 170 23541 172 23591
rect 186 23525 190 23559
rect 216 23525 220 23559
rect 288 23525 292 23713
rect 476 23645 480 23713
rect 524 23683 606 23715
rect 607 23683 616 23717
rect 522 23675 608 23683
rect 649 23675 651 23725
rect 548 23659 582 23675
rect 522 23640 548 23645
rect 522 23639 582 23640
rect 586 23639 608 23645
rect 295 23604 300 23638
rect 324 23604 329 23638
rect 544 23636 582 23639
rect 378 23599 450 23607
rect 428 23569 430 23585
rect 400 23561 430 23569
rect 476 23567 480 23635
rect 544 23606 552 23636
rect 578 23606 582 23636
rect 544 23597 548 23606
rect 400 23557 436 23561
rect 400 23527 408 23557
rect 420 23527 436 23557
rect 544 23559 548 23567
rect 12 23488 62 23490
rect 28 23479 59 23487
rect 62 23479 64 23488
rect 28 23471 64 23479
rect 127 23479 158 23487
rect 127 23472 182 23479
rect 215 23477 224 23505
rect 127 23471 161 23472
rect 59 23455 64 23471
rect 158 23455 161 23471
rect 28 23447 64 23455
rect 127 23454 161 23455
rect 127 23447 182 23454
rect 62 23438 64 23447
rect 213 23439 224 23477
rect 282 23467 292 23525
rect 296 23519 368 23527
rect 319 23489 346 23500
rect 318 23476 324 23489
rect 346 23476 348 23489
rect 428 23480 430 23527
rect 443 23517 450 23519
rect 476 23487 480 23555
rect 544 23525 552 23559
rect 578 23525 582 23559
rect 481 23493 517 23521
rect 481 23487 495 23493
rect 367 23476 380 23480
rect 251 23433 263 23467
rect 273 23433 293 23467
rect 295 23452 324 23476
rect 303 23442 316 23452
rect 318 23436 324 23452
rect 333 23452 380 23476
rect 333 23442 353 23452
rect 367 23446 380 23452
rect 396 23446 408 23480
rect 420 23446 436 23480
rect 120 23385 170 23387
rect 76 23379 92 23385
rect 94 23379 110 23385
rect 76 23369 99 23378
rect 60 23359 67 23369
rect 76 23349 77 23369
rect 96 23344 99 23369
rect 109 23349 110 23369
rect 119 23359 126 23369
rect 76 23335 110 23339
rect 170 23335 172 23385
rect 186 23367 190 23401
rect 216 23367 220 23401
rect 186 23290 220 23324
rect 282 23321 292 23433
rect 318 23426 335 23436
rect 318 23357 324 23426
rect 346 23357 348 23442
rect 428 23399 430 23446
rect 476 23409 480 23477
rect 485 23459 495 23487
rect 505 23487 519 23493
rect 544 23487 555 23525
rect 505 23459 525 23487
rect 544 23459 553 23487
rect 544 23439 548 23459
rect 579 23418 582 23508
rect 612 23490 624 23491
rect 599 23488 649 23490
rect 612 23487 624 23488
rect 610 23480 632 23487
rect 607 23479 632 23480
rect 586 23472 644 23479
rect 607 23471 644 23472
rect 607 23455 610 23471
rect 616 23455 644 23471
rect 607 23454 644 23455
rect 586 23447 644 23454
rect 607 23446 610 23447
rect 612 23439 632 23447
rect 612 23435 624 23439
rect 649 23438 651 23488
rect 544 23401 548 23409
rect 400 23369 408 23399
rect 420 23369 436 23399
rect 400 23365 436 23369
rect 400 23357 430 23365
rect 428 23341 430 23357
rect 476 23329 480 23397
rect 544 23367 552 23401
rect 578 23367 582 23401
rect 544 23359 548 23367
rect 544 23329 586 23330
rect 288 23289 292 23321
rect 296 23319 368 23327
rect 378 23319 450 23327
rect 544 23322 548 23329
rect 439 23291 444 23319
rect 120 23275 170 23277
rect 76 23271 130 23275
rect 110 23266 130 23271
rect 60 23241 67 23251
rect 76 23241 77 23261
rect 96 23232 99 23266
rect 109 23241 110 23261
rect 119 23241 126 23251
rect 76 23225 92 23231
rect 94 23225 110 23231
rect 170 23225 172 23275
rect 186 23209 190 23243
rect 216 23209 220 23243
rect 213 23177 224 23209
rect 282 23205 292 23289
rect 296 23283 368 23291
rect 378 23283 450 23291
rect 468 23288 473 23322
rect 428 23253 430 23269
rect 251 23177 292 23205
rect 318 23184 324 23253
rect 12 23172 62 23174
rect 28 23163 59 23171
rect 62 23163 64 23172
rect 251 23171 263 23177
rect 28 23155 64 23163
rect 127 23163 158 23171
rect 127 23156 182 23163
rect 127 23155 161 23156
rect 59 23139 64 23155
rect 158 23139 161 23155
rect 253 23143 263 23171
rect 273 23143 293 23177
rect 318 23174 335 23184
rect 303 23158 316 23168
rect 318 23158 324 23174
rect 346 23168 348 23253
rect 400 23245 430 23253
rect 476 23251 480 23319
rect 511 23288 582 23322
rect 544 23281 548 23288
rect 400 23241 436 23245
rect 400 23211 408 23241
rect 420 23211 436 23241
rect 544 23243 548 23251
rect 28 23131 64 23139
rect 127 23138 161 23139
rect 127 23131 182 23138
rect 62 23122 64 23131
rect 282 23085 292 23143
rect 295 23134 324 23158
rect 333 23158 353 23168
rect 428 23164 430 23211
rect 476 23171 480 23239
rect 544 23209 552 23243
rect 578 23209 582 23243
rect 544 23201 548 23209
rect 367 23158 380 23164
rect 333 23134 380 23158
rect 318 23121 324 23134
rect 346 23121 348 23134
rect 367 23130 380 23134
rect 396 23130 408 23164
rect 420 23130 436 23164
rect 544 23161 553 23189
rect 319 23110 346 23121
rect 120 23069 170 23071
rect 76 23063 92 23069
rect 94 23063 110 23069
rect 76 23053 99 23062
rect 60 23043 67 23053
rect 76 23033 77 23053
rect 96 23028 99 23053
rect 109 23033 110 23053
rect 119 23043 126 23053
rect 76 23019 110 23023
rect 170 23019 172 23069
rect 186 23051 190 23085
rect 216 23051 220 23085
rect 182 23013 224 23014
rect 186 22989 220 23006
rect 223 22989 257 23006
rect 182 22972 257 22989
rect 182 22971 224 22972
rect 160 22965 246 22971
rect 288 22965 292 23085
rect 296 23083 368 23091
rect 428 23083 430 23130
rect 476 23093 480 23161
rect 485 23117 495 23151
rect 505 23123 525 23151
rect 505 23117 519 23123
rect 544 23117 555 23161
rect 485 23093 492 23117
rect 579 23102 582 23192
rect 612 23174 624 23175
rect 599 23172 649 23174
rect 612 23171 624 23172
rect 610 23164 632 23171
rect 607 23163 632 23164
rect 586 23156 644 23163
rect 607 23155 644 23156
rect 607 23139 610 23155
rect 616 23139 644 23155
rect 607 23138 644 23139
rect 586 23131 644 23138
rect 607 23130 610 23131
rect 612 23123 632 23131
rect 612 23119 624 23123
rect 649 23122 651 23172
rect 544 23085 548 23093
rect 400 23053 408 23083
rect 420 23053 436 23083
rect 400 23049 436 23053
rect 400 23041 430 23049
rect 428 23025 430 23041
rect 476 23013 480 23081
rect 544 23051 552 23085
rect 578 23051 582 23085
rect 544 23043 548 23051
rect 295 22972 300 23006
rect 324 22972 329 23006
rect 378 23003 450 23011
rect 544 23008 548 23013
rect 544 23004 582 23008
rect 544 22989 552 23004
rect 578 22989 582 23004
rect 544 22971 586 22989
rect 522 22965 608 22971
rect 182 22949 224 22965
rect 544 22949 586 22965
rect 17 22935 67 22937
rect 119 22935 169 22937
rect 186 22935 220 22949
rect 548 22935 582 22949
rect 599 22935 649 22937
rect 42 22893 59 22927
rect 67 22885 69 22935
rect 160 22927 246 22935
rect 522 22927 608 22935
rect 76 22893 110 22927
rect 127 22893 144 22927
rect 152 22893 161 22927
rect 162 22925 195 22927
rect 224 22925 244 22927
rect 162 22893 244 22925
rect 524 22925 548 22927
rect 573 22925 582 22927
rect 586 22925 606 22927
rect 160 22885 246 22893
rect 186 22869 220 22885
rect 182 22855 224 22856
rect 160 22849 182 22855
rect 224 22849 246 22855
rect 186 22814 220 22848
rect 223 22814 257 22848
rect 120 22801 170 22803
rect 76 22797 130 22801
rect 110 22792 130 22797
rect 60 22767 67 22777
rect 76 22767 77 22787
rect 96 22758 99 22792
rect 109 22767 110 22787
rect 119 22767 126 22777
rect 76 22751 92 22757
rect 94 22751 110 22757
rect 170 22751 172 22801
rect 186 22735 190 22769
rect 216 22735 220 22769
rect 288 22735 292 22923
rect 476 22855 480 22923
rect 524 22893 606 22925
rect 607 22893 616 22927
rect 522 22885 608 22893
rect 649 22885 651 22935
rect 548 22869 582 22885
rect 522 22850 548 22855
rect 522 22849 582 22850
rect 586 22849 608 22855
rect 295 22814 300 22848
rect 324 22814 329 22848
rect 544 22846 582 22849
rect 378 22809 450 22817
rect 428 22779 430 22795
rect 400 22771 430 22779
rect 476 22777 480 22845
rect 544 22816 552 22846
rect 578 22816 582 22846
rect 544 22807 548 22816
rect 400 22767 436 22771
rect 400 22737 408 22767
rect 420 22737 436 22767
rect 544 22769 548 22777
rect 12 22698 62 22700
rect 28 22689 59 22697
rect 62 22689 64 22698
rect 28 22681 64 22689
rect 127 22689 158 22697
rect 127 22682 182 22689
rect 215 22687 224 22715
rect 127 22681 161 22682
rect 59 22665 64 22681
rect 158 22665 161 22681
rect 28 22657 64 22665
rect 127 22664 161 22665
rect 127 22657 182 22664
rect 62 22648 64 22657
rect 213 22649 224 22687
rect 282 22677 292 22735
rect 296 22729 368 22737
rect 319 22699 346 22710
rect 318 22686 324 22699
rect 346 22686 348 22699
rect 428 22690 430 22737
rect 443 22727 450 22729
rect 476 22697 480 22765
rect 544 22735 552 22769
rect 578 22735 582 22769
rect 481 22703 517 22731
rect 481 22697 495 22703
rect 367 22686 380 22690
rect 251 22643 263 22677
rect 273 22643 293 22677
rect 295 22662 324 22686
rect 303 22652 316 22662
rect 318 22646 324 22662
rect 333 22662 380 22686
rect 333 22652 353 22662
rect 367 22656 380 22662
rect 396 22656 408 22690
rect 420 22656 436 22690
rect 120 22595 170 22597
rect 76 22589 92 22595
rect 94 22589 110 22595
rect 76 22579 99 22588
rect 60 22569 67 22579
rect 76 22559 77 22579
rect 96 22554 99 22579
rect 109 22559 110 22579
rect 119 22569 126 22579
rect 76 22545 110 22549
rect 170 22545 172 22595
rect 186 22577 190 22611
rect 216 22577 220 22611
rect 186 22500 220 22534
rect 282 22531 292 22643
rect 318 22636 335 22646
rect 318 22567 324 22636
rect 346 22567 348 22652
rect 428 22609 430 22656
rect 476 22619 480 22687
rect 485 22669 495 22697
rect 505 22697 519 22703
rect 544 22697 555 22735
rect 505 22669 525 22697
rect 544 22669 553 22697
rect 544 22649 548 22669
rect 579 22628 582 22718
rect 612 22700 624 22701
rect 599 22698 649 22700
rect 612 22697 624 22698
rect 610 22690 632 22697
rect 607 22689 632 22690
rect 586 22682 644 22689
rect 607 22681 644 22682
rect 607 22665 610 22681
rect 616 22665 644 22681
rect 607 22664 644 22665
rect 586 22657 644 22664
rect 607 22656 610 22657
rect 612 22649 632 22657
rect 612 22645 624 22649
rect 649 22648 651 22698
rect 544 22611 548 22619
rect 400 22579 408 22609
rect 420 22579 436 22609
rect 400 22575 436 22579
rect 400 22567 430 22575
rect 428 22551 430 22567
rect 476 22539 480 22607
rect 544 22577 552 22611
rect 578 22577 582 22611
rect 544 22569 548 22577
rect 544 22539 586 22540
rect 288 22499 292 22531
rect 296 22529 368 22537
rect 378 22529 450 22537
rect 544 22532 548 22539
rect 439 22501 444 22529
rect 120 22485 170 22487
rect 76 22481 130 22485
rect 110 22476 130 22481
rect 60 22451 67 22461
rect 76 22451 77 22471
rect 96 22442 99 22476
rect 109 22451 110 22471
rect 119 22451 126 22461
rect 76 22435 92 22441
rect 94 22435 110 22441
rect 170 22435 172 22485
rect 186 22419 190 22453
rect 216 22419 220 22453
rect 213 22387 224 22419
rect 282 22415 292 22499
rect 296 22493 368 22501
rect 378 22493 450 22501
rect 468 22498 473 22532
rect 428 22463 430 22479
rect 251 22387 292 22415
rect 318 22394 324 22463
rect 12 22382 62 22384
rect 28 22373 59 22381
rect 62 22373 64 22382
rect 251 22381 263 22387
rect 28 22365 64 22373
rect 127 22373 158 22381
rect 127 22366 182 22373
rect 127 22365 161 22366
rect 59 22349 64 22365
rect 158 22349 161 22365
rect 253 22353 263 22381
rect 273 22353 293 22387
rect 318 22384 335 22394
rect 303 22368 316 22378
rect 318 22368 324 22384
rect 346 22378 348 22463
rect 400 22455 430 22463
rect 476 22461 480 22529
rect 511 22498 582 22532
rect 544 22491 548 22498
rect 400 22451 436 22455
rect 400 22421 408 22451
rect 420 22421 436 22451
rect 544 22453 548 22461
rect 28 22341 64 22349
rect 127 22348 161 22349
rect 127 22341 182 22348
rect 62 22332 64 22341
rect 282 22295 292 22353
rect 295 22344 324 22368
rect 333 22368 353 22378
rect 428 22374 430 22421
rect 476 22381 480 22449
rect 544 22419 552 22453
rect 578 22419 582 22453
rect 544 22411 548 22419
rect 367 22368 380 22374
rect 333 22344 380 22368
rect 318 22331 324 22344
rect 346 22331 348 22344
rect 367 22340 380 22344
rect 396 22340 408 22374
rect 420 22340 436 22374
rect 544 22371 553 22399
rect 319 22320 346 22331
rect 120 22279 170 22281
rect 76 22273 92 22279
rect 94 22273 110 22279
rect 76 22263 99 22272
rect 60 22253 67 22263
rect 76 22243 77 22263
rect 96 22238 99 22263
rect 109 22243 110 22263
rect 119 22253 126 22263
rect 76 22229 110 22233
rect 170 22229 172 22279
rect 186 22261 190 22295
rect 216 22261 220 22295
rect 182 22223 224 22224
rect 186 22199 220 22216
rect 223 22199 257 22216
rect 182 22182 257 22199
rect 182 22181 224 22182
rect 160 22175 246 22181
rect 288 22175 292 22295
rect 296 22293 368 22301
rect 428 22293 430 22340
rect 476 22303 480 22371
rect 485 22327 495 22361
rect 505 22333 525 22361
rect 505 22327 519 22333
rect 544 22327 555 22371
rect 485 22303 492 22327
rect 579 22312 582 22402
rect 612 22384 624 22385
rect 599 22382 649 22384
rect 612 22381 624 22382
rect 610 22374 632 22381
rect 607 22373 632 22374
rect 586 22366 644 22373
rect 607 22365 644 22366
rect 607 22349 610 22365
rect 616 22349 644 22365
rect 607 22348 644 22349
rect 586 22341 644 22348
rect 607 22340 610 22341
rect 612 22333 632 22341
rect 612 22329 624 22333
rect 649 22332 651 22382
rect 544 22295 548 22303
rect 400 22263 408 22293
rect 420 22263 436 22293
rect 400 22259 436 22263
rect 400 22251 430 22259
rect 428 22235 430 22251
rect 476 22223 480 22291
rect 544 22261 552 22295
rect 578 22261 582 22295
rect 544 22253 548 22261
rect 295 22182 300 22216
rect 324 22182 329 22216
rect 378 22213 450 22221
rect 544 22218 548 22223
rect 544 22214 582 22218
rect 544 22199 552 22214
rect 578 22199 582 22214
rect 544 22181 586 22199
rect 522 22175 608 22181
rect 182 22159 224 22175
rect 544 22159 586 22175
rect 17 22145 67 22147
rect 119 22145 169 22147
rect 186 22145 220 22159
rect 548 22145 582 22159
rect 599 22145 649 22147
rect 42 22103 59 22137
rect 67 22095 69 22145
rect 160 22137 246 22145
rect 522 22137 608 22145
rect 76 22103 110 22137
rect 127 22103 144 22137
rect 152 22103 161 22137
rect 162 22135 195 22137
rect 224 22135 244 22137
rect 162 22103 244 22135
rect 524 22135 548 22137
rect 573 22135 582 22137
rect 586 22135 606 22137
rect 160 22095 246 22103
rect 186 22079 220 22095
rect 182 22065 224 22066
rect 160 22059 182 22065
rect 224 22059 246 22065
rect 186 22024 220 22058
rect 223 22024 257 22058
rect 120 22011 170 22013
rect 76 22007 130 22011
rect 110 22002 130 22007
rect 60 21977 67 21987
rect 76 21977 77 21997
rect 96 21968 99 22002
rect 109 21977 110 21997
rect 119 21977 126 21987
rect 76 21961 92 21967
rect 94 21961 110 21967
rect 170 21961 172 22011
rect 186 21945 190 21979
rect 216 21945 220 21979
rect 288 21945 292 22133
rect 476 22065 480 22133
rect 524 22103 606 22135
rect 607 22103 616 22137
rect 522 22095 608 22103
rect 649 22095 651 22145
rect 548 22079 582 22095
rect 522 22060 548 22065
rect 522 22059 582 22060
rect 586 22059 608 22065
rect 295 22024 300 22058
rect 324 22024 329 22058
rect 544 22056 582 22059
rect 378 22019 450 22027
rect 428 21989 430 22005
rect 400 21981 430 21989
rect 476 21987 480 22055
rect 544 22026 552 22056
rect 578 22026 582 22056
rect 544 22017 548 22026
rect 400 21977 436 21981
rect 400 21947 408 21977
rect 420 21947 436 21977
rect 544 21979 548 21987
rect 12 21908 62 21910
rect 28 21899 59 21907
rect 62 21899 64 21908
rect 28 21891 64 21899
rect 127 21899 158 21907
rect 127 21892 182 21899
rect 215 21897 224 21925
rect 127 21891 161 21892
rect 59 21875 64 21891
rect 158 21875 161 21891
rect 28 21867 64 21875
rect 127 21874 161 21875
rect 127 21867 182 21874
rect 62 21858 64 21867
rect 213 21859 224 21897
rect 282 21887 292 21945
rect 296 21939 368 21947
rect 319 21909 346 21920
rect 318 21896 324 21909
rect 346 21896 348 21909
rect 428 21900 430 21947
rect 443 21937 450 21939
rect 476 21907 480 21975
rect 544 21945 552 21979
rect 578 21945 582 21979
rect 481 21913 517 21941
rect 481 21907 495 21913
rect 367 21896 380 21900
rect 251 21853 263 21887
rect 273 21853 293 21887
rect 295 21872 324 21896
rect 303 21862 316 21872
rect 318 21856 324 21872
rect 333 21872 380 21896
rect 333 21862 353 21872
rect 367 21866 380 21872
rect 396 21866 408 21900
rect 420 21866 436 21900
rect 120 21805 170 21807
rect 76 21799 92 21805
rect 94 21799 110 21805
rect 76 21789 99 21798
rect 60 21779 67 21789
rect 76 21769 77 21789
rect 96 21764 99 21789
rect 109 21769 110 21789
rect 119 21779 126 21789
rect 76 21755 110 21759
rect 170 21755 172 21805
rect 186 21787 190 21821
rect 216 21787 220 21821
rect 186 21710 220 21744
rect 282 21741 292 21853
rect 318 21846 335 21856
rect 318 21777 324 21846
rect 346 21777 348 21862
rect 428 21819 430 21866
rect 476 21829 480 21897
rect 485 21879 495 21907
rect 505 21907 519 21913
rect 544 21907 555 21945
rect 505 21879 525 21907
rect 544 21879 553 21907
rect 544 21859 548 21879
rect 579 21838 582 21928
rect 612 21910 624 21911
rect 599 21908 649 21910
rect 612 21907 624 21908
rect 610 21900 632 21907
rect 607 21899 632 21900
rect 586 21892 644 21899
rect 607 21891 644 21892
rect 607 21875 610 21891
rect 616 21875 644 21891
rect 607 21874 644 21875
rect 586 21867 644 21874
rect 607 21866 610 21867
rect 612 21859 632 21867
rect 612 21855 624 21859
rect 649 21858 651 21908
rect 544 21821 548 21829
rect 400 21789 408 21819
rect 420 21789 436 21819
rect 400 21785 436 21789
rect 400 21777 430 21785
rect 428 21761 430 21777
rect 476 21749 480 21817
rect 544 21787 552 21821
rect 578 21787 582 21821
rect 544 21779 548 21787
rect 544 21749 586 21750
rect 288 21709 292 21741
rect 296 21739 368 21747
rect 378 21739 450 21747
rect 544 21742 548 21749
rect 439 21711 444 21739
rect 120 21695 170 21697
rect 76 21691 130 21695
rect 110 21686 130 21691
rect 60 21661 67 21671
rect 76 21661 77 21681
rect 96 21652 99 21686
rect 109 21661 110 21681
rect 119 21661 126 21671
rect 76 21645 92 21651
rect 94 21645 110 21651
rect 170 21645 172 21695
rect 186 21629 190 21663
rect 216 21629 220 21663
rect 213 21597 224 21629
rect 282 21625 292 21709
rect 296 21703 368 21711
rect 378 21703 450 21711
rect 468 21708 473 21742
rect 428 21673 430 21689
rect 251 21597 292 21625
rect 318 21604 324 21673
rect 12 21592 62 21594
rect 28 21583 59 21591
rect 62 21583 64 21592
rect 251 21591 263 21597
rect 28 21575 64 21583
rect 127 21583 158 21591
rect 127 21576 182 21583
rect 127 21575 161 21576
rect 59 21559 64 21575
rect 158 21559 161 21575
rect 253 21563 263 21591
rect 273 21563 293 21597
rect 318 21594 335 21604
rect 303 21578 316 21588
rect 318 21578 324 21594
rect 346 21588 348 21673
rect 400 21665 430 21673
rect 476 21671 480 21739
rect 511 21708 582 21742
rect 544 21701 548 21708
rect 400 21661 436 21665
rect 400 21631 408 21661
rect 420 21631 436 21661
rect 544 21663 548 21671
rect 28 21551 64 21559
rect 127 21558 161 21559
rect 127 21551 182 21558
rect 62 21542 64 21551
rect 282 21505 292 21563
rect 295 21554 324 21578
rect 333 21578 353 21588
rect 428 21584 430 21631
rect 476 21591 480 21659
rect 544 21629 552 21663
rect 578 21629 582 21663
rect 544 21621 548 21629
rect 367 21578 380 21584
rect 333 21554 380 21578
rect 318 21541 324 21554
rect 346 21541 348 21554
rect 367 21550 380 21554
rect 396 21550 408 21584
rect 420 21550 436 21584
rect 544 21581 553 21609
rect 319 21530 346 21541
rect 120 21489 170 21491
rect 76 21483 92 21489
rect 94 21483 110 21489
rect 76 21473 99 21482
rect 60 21463 67 21473
rect 76 21453 77 21473
rect 96 21448 99 21473
rect 109 21453 110 21473
rect 119 21463 126 21473
rect 76 21439 110 21443
rect 170 21439 172 21489
rect 186 21471 190 21505
rect 216 21471 220 21505
rect 182 21433 224 21434
rect 186 21409 220 21426
rect 223 21409 257 21426
rect 182 21392 257 21409
rect 182 21391 224 21392
rect 160 21385 246 21391
rect 288 21385 292 21505
rect 296 21503 368 21511
rect 428 21503 430 21550
rect 476 21513 480 21581
rect 485 21537 495 21571
rect 505 21543 525 21571
rect 505 21537 519 21543
rect 544 21537 555 21581
rect 485 21513 492 21537
rect 579 21522 582 21612
rect 612 21594 624 21595
rect 599 21592 649 21594
rect 612 21591 624 21592
rect 610 21584 632 21591
rect 607 21583 632 21584
rect 586 21576 644 21583
rect 607 21575 644 21576
rect 607 21559 610 21575
rect 616 21559 644 21575
rect 607 21558 644 21559
rect 586 21551 644 21558
rect 607 21550 610 21551
rect 612 21543 632 21551
rect 612 21539 624 21543
rect 649 21542 651 21592
rect 544 21505 548 21513
rect 400 21473 408 21503
rect 420 21473 436 21503
rect 400 21469 436 21473
rect 400 21461 430 21469
rect 428 21445 430 21461
rect 476 21433 480 21501
rect 544 21471 552 21505
rect 578 21471 582 21505
rect 544 21463 548 21471
rect 295 21392 300 21426
rect 324 21392 329 21426
rect 378 21423 450 21431
rect 544 21428 548 21433
rect 544 21424 582 21428
rect 544 21409 552 21424
rect 578 21409 582 21424
rect 544 21391 586 21409
rect 522 21385 608 21391
rect 182 21369 224 21385
rect 544 21369 586 21385
rect 17 21355 67 21357
rect 119 21355 169 21357
rect 186 21355 220 21369
rect 548 21355 582 21369
rect 599 21355 649 21357
rect 42 21313 59 21347
rect 67 21305 69 21355
rect 160 21347 246 21355
rect 522 21347 608 21355
rect 76 21313 110 21347
rect 127 21313 144 21347
rect 152 21313 161 21347
rect 162 21345 195 21347
rect 224 21345 244 21347
rect 162 21313 244 21345
rect 524 21345 548 21347
rect 573 21345 582 21347
rect 586 21345 606 21347
rect 160 21305 246 21313
rect 186 21289 220 21305
rect 182 21275 224 21276
rect 160 21269 182 21275
rect 224 21269 246 21275
rect 186 21234 220 21268
rect 223 21234 257 21268
rect 120 21221 170 21223
rect 76 21217 130 21221
rect 110 21212 130 21217
rect 60 21187 67 21197
rect 76 21187 77 21207
rect 96 21178 99 21212
rect 109 21187 110 21207
rect 119 21187 126 21197
rect 76 21171 92 21177
rect 94 21171 110 21177
rect 170 21171 172 21221
rect 186 21155 190 21189
rect 216 21155 220 21189
rect 288 21155 292 21343
rect 476 21275 480 21343
rect 524 21313 606 21345
rect 607 21313 616 21347
rect 522 21305 608 21313
rect 649 21305 651 21355
rect 548 21289 582 21305
rect 522 21270 548 21275
rect 522 21269 582 21270
rect 586 21269 608 21275
rect 295 21234 300 21268
rect 324 21234 329 21268
rect 544 21266 582 21269
rect 378 21229 450 21237
rect 428 21199 430 21215
rect 400 21191 430 21199
rect 476 21197 480 21265
rect 544 21236 552 21266
rect 578 21236 582 21266
rect 544 21227 548 21236
rect 400 21187 436 21191
rect 400 21157 408 21187
rect 420 21157 436 21187
rect 544 21189 548 21197
rect 12 21118 62 21120
rect 28 21109 59 21117
rect 62 21109 64 21118
rect 28 21101 64 21109
rect 127 21109 158 21117
rect 127 21102 182 21109
rect 215 21107 224 21135
rect 127 21101 161 21102
rect 59 21085 64 21101
rect 158 21085 161 21101
rect 28 21077 64 21085
rect 127 21084 161 21085
rect 127 21077 182 21084
rect 62 21068 64 21077
rect 213 21069 224 21107
rect 282 21097 292 21155
rect 296 21149 368 21157
rect 319 21119 346 21130
rect 318 21106 324 21119
rect 346 21106 348 21119
rect 428 21110 430 21157
rect 443 21147 450 21149
rect 476 21117 480 21185
rect 544 21155 552 21189
rect 578 21155 582 21189
rect 481 21123 517 21151
rect 481 21117 495 21123
rect 367 21106 380 21110
rect 251 21063 263 21097
rect 273 21063 293 21097
rect 295 21082 324 21106
rect 303 21072 316 21082
rect 318 21066 324 21082
rect 333 21082 380 21106
rect 333 21072 353 21082
rect 367 21076 380 21082
rect 396 21076 408 21110
rect 420 21076 436 21110
rect 120 21015 170 21017
rect 76 21009 92 21015
rect 94 21009 110 21015
rect 76 20999 99 21008
rect 60 20989 67 20999
rect 76 20979 77 20999
rect 96 20974 99 20999
rect 109 20979 110 20999
rect 119 20989 126 20999
rect 76 20965 110 20969
rect 170 20965 172 21015
rect 186 20997 190 21031
rect 216 20997 220 21031
rect 186 20920 220 20954
rect 282 20951 292 21063
rect 318 21056 335 21066
rect 318 20987 324 21056
rect 346 20987 348 21072
rect 428 21029 430 21076
rect 476 21039 480 21107
rect 485 21089 495 21117
rect 505 21117 519 21123
rect 544 21117 555 21155
rect 505 21089 525 21117
rect 544 21089 553 21117
rect 544 21069 548 21089
rect 579 21048 582 21138
rect 612 21120 624 21121
rect 599 21118 649 21120
rect 612 21117 624 21118
rect 610 21110 632 21117
rect 607 21109 632 21110
rect 586 21102 644 21109
rect 607 21101 644 21102
rect 607 21085 610 21101
rect 616 21085 644 21101
rect 607 21084 644 21085
rect 586 21077 644 21084
rect 607 21076 610 21077
rect 612 21069 632 21077
rect 612 21065 624 21069
rect 649 21068 651 21118
rect 544 21031 548 21039
rect 400 20999 408 21029
rect 420 20999 436 21029
rect 400 20995 436 20999
rect 400 20987 430 20995
rect 428 20971 430 20987
rect 476 20959 480 21027
rect 544 20997 552 21031
rect 578 20997 582 21031
rect 544 20989 548 20997
rect 544 20959 586 20960
rect 288 20919 292 20951
rect 296 20949 368 20957
rect 378 20949 450 20957
rect 544 20952 548 20959
rect 439 20921 444 20949
rect 120 20905 170 20907
rect 76 20901 130 20905
rect 110 20896 130 20901
rect 60 20871 67 20881
rect 76 20871 77 20891
rect 96 20862 99 20896
rect 109 20871 110 20891
rect 119 20871 126 20881
rect 76 20855 92 20861
rect 94 20855 110 20861
rect 170 20855 172 20905
rect 186 20839 190 20873
rect 216 20839 220 20873
rect 213 20807 224 20839
rect 282 20835 292 20919
rect 296 20913 368 20921
rect 378 20913 450 20921
rect 468 20918 473 20952
rect 428 20883 430 20899
rect 251 20807 292 20835
rect 318 20814 324 20883
rect 12 20802 62 20804
rect 28 20793 59 20801
rect 62 20793 64 20802
rect 251 20801 263 20807
rect 28 20785 64 20793
rect 127 20793 158 20801
rect 127 20786 182 20793
rect 127 20785 161 20786
rect 59 20769 64 20785
rect 158 20769 161 20785
rect 253 20773 263 20801
rect 273 20773 293 20807
rect 318 20804 335 20814
rect 303 20788 316 20798
rect 318 20788 324 20804
rect 346 20798 348 20883
rect 400 20875 430 20883
rect 476 20881 480 20949
rect 511 20918 582 20952
rect 544 20911 548 20918
rect 400 20871 436 20875
rect 400 20841 408 20871
rect 420 20841 436 20871
rect 544 20873 548 20881
rect 28 20761 64 20769
rect 127 20768 161 20769
rect 127 20761 182 20768
rect 62 20752 64 20761
rect 282 20715 292 20773
rect 295 20764 324 20788
rect 333 20788 353 20798
rect 428 20794 430 20841
rect 476 20801 480 20869
rect 544 20839 552 20873
rect 578 20839 582 20873
rect 544 20831 548 20839
rect 367 20788 380 20794
rect 333 20764 380 20788
rect 318 20751 324 20764
rect 346 20751 348 20764
rect 367 20760 380 20764
rect 396 20760 408 20794
rect 420 20760 436 20794
rect 544 20791 553 20819
rect 319 20740 346 20751
rect 120 20699 170 20701
rect 76 20693 92 20699
rect 94 20693 110 20699
rect 76 20683 99 20692
rect 60 20673 67 20683
rect 76 20663 77 20683
rect 96 20658 99 20683
rect 109 20663 110 20683
rect 119 20673 126 20683
rect 76 20649 110 20653
rect 170 20649 172 20699
rect 186 20681 190 20715
rect 216 20681 220 20715
rect 182 20643 224 20644
rect 186 20619 220 20636
rect 223 20619 257 20636
rect 182 20602 257 20619
rect 182 20601 224 20602
rect 160 20595 246 20601
rect 288 20595 292 20715
rect 296 20713 368 20721
rect 428 20713 430 20760
rect 476 20723 480 20791
rect 485 20747 495 20781
rect 505 20753 525 20781
rect 505 20747 519 20753
rect 544 20747 555 20791
rect 485 20723 492 20747
rect 579 20732 582 20822
rect 612 20804 624 20805
rect 599 20802 649 20804
rect 612 20801 624 20802
rect 610 20794 632 20801
rect 607 20793 632 20794
rect 586 20786 644 20793
rect 607 20785 644 20786
rect 607 20769 610 20785
rect 616 20769 644 20785
rect 607 20768 644 20769
rect 586 20761 644 20768
rect 607 20760 610 20761
rect 612 20753 632 20761
rect 612 20749 624 20753
rect 649 20752 651 20802
rect 544 20715 548 20723
rect 400 20683 408 20713
rect 420 20683 436 20713
rect 400 20679 436 20683
rect 400 20671 430 20679
rect 428 20655 430 20671
rect 476 20643 480 20711
rect 544 20681 552 20715
rect 578 20681 582 20715
rect 544 20673 548 20681
rect 295 20602 300 20636
rect 324 20602 329 20636
rect 378 20633 450 20641
rect 544 20638 548 20643
rect 544 20634 582 20638
rect 544 20619 552 20634
rect 578 20619 582 20634
rect 544 20601 586 20619
rect 522 20595 608 20601
rect 182 20579 224 20595
rect 544 20579 586 20595
rect 17 20565 67 20567
rect 119 20565 169 20567
rect 186 20565 220 20579
rect 548 20565 582 20579
rect 599 20565 649 20567
rect 42 20523 59 20557
rect 67 20515 69 20565
rect 160 20557 246 20565
rect 522 20557 608 20565
rect 76 20523 110 20557
rect 127 20523 144 20557
rect 152 20523 161 20557
rect 162 20555 195 20557
rect 224 20555 244 20557
rect 162 20523 244 20555
rect 524 20555 548 20557
rect 573 20555 582 20557
rect 586 20555 606 20557
rect 160 20515 246 20523
rect 186 20499 220 20515
rect 182 20485 224 20486
rect 160 20479 182 20485
rect 224 20479 246 20485
rect 186 20444 220 20478
rect 223 20444 257 20478
rect 120 20431 170 20433
rect 76 20427 130 20431
rect 110 20422 130 20427
rect 60 20397 67 20407
rect 76 20397 77 20417
rect 96 20388 99 20422
rect 109 20397 110 20417
rect 119 20397 126 20407
rect 76 20381 92 20387
rect 94 20381 110 20387
rect 170 20381 172 20431
rect 186 20365 190 20399
rect 216 20365 220 20399
rect 288 20365 292 20553
rect 476 20485 480 20553
rect 524 20523 606 20555
rect 607 20523 616 20557
rect 522 20515 608 20523
rect 649 20515 651 20565
rect 548 20499 582 20515
rect 522 20480 548 20485
rect 522 20479 582 20480
rect 586 20479 608 20485
rect 295 20444 300 20478
rect 324 20444 329 20478
rect 544 20476 582 20479
rect 378 20439 450 20447
rect 428 20409 430 20425
rect 400 20401 430 20409
rect 476 20407 480 20475
rect 544 20446 552 20476
rect 578 20446 582 20476
rect 544 20437 548 20446
rect 400 20397 436 20401
rect 400 20367 408 20397
rect 420 20367 436 20397
rect 544 20399 548 20407
rect 12 20328 62 20330
rect 28 20319 59 20327
rect 62 20319 64 20328
rect 28 20311 64 20319
rect 127 20319 158 20327
rect 127 20312 182 20319
rect 215 20317 224 20345
rect 127 20311 161 20312
rect 59 20295 64 20311
rect 158 20295 161 20311
rect 28 20287 64 20295
rect 127 20294 161 20295
rect 127 20287 182 20294
rect 62 20278 64 20287
rect 213 20279 224 20317
rect 282 20307 292 20365
rect 296 20359 368 20367
rect 319 20329 346 20340
rect 318 20316 324 20329
rect 346 20316 348 20329
rect 428 20320 430 20367
rect 443 20357 450 20359
rect 476 20327 480 20395
rect 544 20365 552 20399
rect 578 20365 582 20399
rect 481 20333 517 20361
rect 481 20327 495 20333
rect 367 20316 380 20320
rect 251 20273 263 20307
rect 273 20273 293 20307
rect 295 20292 324 20316
rect 303 20282 316 20292
rect 318 20276 324 20292
rect 333 20292 380 20316
rect 333 20282 353 20292
rect 367 20286 380 20292
rect 396 20286 408 20320
rect 420 20286 436 20320
rect 120 20225 170 20227
rect 76 20219 92 20225
rect 94 20219 110 20225
rect 76 20209 99 20218
rect 60 20199 67 20209
rect 76 20189 77 20209
rect 96 20184 99 20209
rect 109 20189 110 20209
rect 119 20199 126 20209
rect 76 20175 110 20179
rect 170 20175 172 20225
rect 186 20207 190 20241
rect 216 20207 220 20241
rect 186 20130 220 20164
rect 282 20161 292 20273
rect 318 20266 335 20276
rect 318 20197 324 20266
rect 346 20197 348 20282
rect 428 20239 430 20286
rect 476 20249 480 20317
rect 485 20299 495 20327
rect 505 20327 519 20333
rect 544 20327 555 20365
rect 505 20299 525 20327
rect 544 20299 553 20327
rect 544 20279 548 20299
rect 579 20258 582 20348
rect 612 20330 624 20331
rect 599 20328 649 20330
rect 612 20327 624 20328
rect 610 20320 632 20327
rect 607 20319 632 20320
rect 586 20312 644 20319
rect 607 20311 644 20312
rect 607 20295 610 20311
rect 616 20295 644 20311
rect 607 20294 644 20295
rect 586 20287 644 20294
rect 607 20286 610 20287
rect 612 20279 632 20287
rect 612 20275 624 20279
rect 649 20278 651 20328
rect 544 20241 548 20249
rect 400 20209 408 20239
rect 420 20209 436 20239
rect 400 20205 436 20209
rect 400 20197 430 20205
rect 428 20181 430 20197
rect 476 20169 480 20237
rect 544 20207 552 20241
rect 578 20207 582 20241
rect 544 20199 548 20207
rect 544 20169 586 20170
rect 288 20129 292 20161
rect 296 20159 368 20167
rect 378 20159 450 20167
rect 544 20162 548 20169
rect 439 20131 444 20159
rect 120 20115 170 20117
rect 76 20111 130 20115
rect 110 20106 130 20111
rect 60 20081 67 20091
rect 76 20081 77 20101
rect 96 20072 99 20106
rect 109 20081 110 20101
rect 119 20081 126 20091
rect 76 20065 92 20071
rect 94 20065 110 20071
rect 170 20065 172 20115
rect 186 20049 190 20083
rect 216 20049 220 20083
rect 213 20017 224 20049
rect 282 20045 292 20129
rect 296 20123 368 20131
rect 378 20123 450 20131
rect 468 20128 473 20162
rect 428 20093 430 20109
rect 251 20017 292 20045
rect 318 20024 324 20093
rect 12 20012 62 20014
rect 28 20003 59 20011
rect 62 20003 64 20012
rect 251 20011 263 20017
rect 28 19995 64 20003
rect 127 20003 158 20011
rect 127 19996 182 20003
rect 127 19995 161 19996
rect 59 19979 64 19995
rect 158 19979 161 19995
rect 253 19983 263 20011
rect 273 19983 293 20017
rect 318 20014 335 20024
rect 303 19998 316 20008
rect 318 19998 324 20014
rect 346 20008 348 20093
rect 400 20085 430 20093
rect 476 20091 480 20159
rect 511 20128 582 20162
rect 544 20121 548 20128
rect 400 20081 436 20085
rect 400 20051 408 20081
rect 420 20051 436 20081
rect 544 20083 548 20091
rect 28 19971 64 19979
rect 127 19978 161 19979
rect 127 19971 182 19978
rect 62 19962 64 19971
rect 282 19925 292 19983
rect 295 19974 324 19998
rect 333 19998 353 20008
rect 428 20004 430 20051
rect 476 20011 480 20079
rect 544 20049 552 20083
rect 578 20049 582 20083
rect 544 20041 548 20049
rect 367 19998 380 20004
rect 333 19974 380 19998
rect 318 19961 324 19974
rect 346 19961 348 19974
rect 367 19970 380 19974
rect 396 19970 408 20004
rect 420 19970 436 20004
rect 544 20001 553 20029
rect 319 19950 346 19961
rect 120 19909 170 19911
rect 76 19903 92 19909
rect 94 19903 110 19909
rect 76 19893 99 19902
rect 60 19883 67 19893
rect 76 19873 77 19893
rect 96 19868 99 19893
rect 109 19873 110 19893
rect 119 19883 126 19893
rect 76 19859 110 19863
rect 170 19859 172 19909
rect 186 19891 190 19925
rect 216 19891 220 19925
rect 182 19853 224 19854
rect 186 19829 220 19846
rect 223 19829 257 19846
rect 182 19812 257 19829
rect 182 19811 224 19812
rect 160 19805 246 19811
rect 288 19805 292 19925
rect 296 19923 368 19931
rect 428 19923 430 19970
rect 476 19933 480 20001
rect 485 19957 495 19991
rect 505 19963 525 19991
rect 505 19957 519 19963
rect 544 19957 555 20001
rect 485 19933 492 19957
rect 579 19942 582 20032
rect 612 20014 624 20015
rect 599 20012 649 20014
rect 612 20011 624 20012
rect 610 20004 632 20011
rect 607 20003 632 20004
rect 586 19996 644 20003
rect 607 19995 644 19996
rect 607 19979 610 19995
rect 616 19979 644 19995
rect 607 19978 644 19979
rect 586 19971 644 19978
rect 607 19970 610 19971
rect 612 19963 632 19971
rect 612 19959 624 19963
rect 649 19962 651 20012
rect 544 19925 548 19933
rect 400 19893 408 19923
rect 420 19893 436 19923
rect 400 19889 436 19893
rect 400 19881 430 19889
rect 428 19865 430 19881
rect 476 19853 480 19921
rect 544 19891 552 19925
rect 578 19891 582 19925
rect 544 19883 548 19891
rect 295 19812 300 19846
rect 324 19812 329 19846
rect 378 19843 450 19851
rect 544 19848 548 19853
rect 544 19844 582 19848
rect 544 19829 552 19844
rect 578 19829 582 19844
rect 544 19811 586 19829
rect 522 19805 608 19811
rect 182 19789 224 19805
rect 544 19789 586 19805
rect 17 19775 67 19777
rect 119 19775 169 19777
rect 186 19775 220 19789
rect 548 19775 582 19789
rect 599 19775 649 19777
rect 42 19733 59 19767
rect 67 19725 69 19775
rect 160 19767 246 19775
rect 522 19767 608 19775
rect 76 19733 110 19767
rect 127 19733 144 19767
rect 152 19733 161 19767
rect 162 19765 195 19767
rect 224 19765 244 19767
rect 162 19733 244 19765
rect 524 19765 548 19767
rect 573 19765 582 19767
rect 586 19765 606 19767
rect 160 19725 246 19733
rect 186 19709 220 19725
rect 182 19695 224 19696
rect 160 19689 182 19695
rect 224 19689 246 19695
rect 186 19654 220 19688
rect 223 19654 257 19688
rect 120 19641 170 19643
rect 76 19637 130 19641
rect 110 19632 130 19637
rect 60 19607 67 19617
rect 76 19607 77 19627
rect 96 19598 99 19632
rect 109 19607 110 19627
rect 119 19607 126 19617
rect 76 19591 92 19597
rect 94 19591 110 19597
rect 170 19591 172 19641
rect 186 19575 190 19609
rect 216 19575 220 19609
rect 288 19575 292 19763
rect 476 19695 480 19763
rect 524 19733 606 19765
rect 607 19733 616 19767
rect 522 19725 608 19733
rect 649 19725 651 19775
rect 548 19709 582 19725
rect 522 19690 548 19695
rect 522 19689 582 19690
rect 586 19689 608 19695
rect 295 19654 300 19688
rect 324 19654 329 19688
rect 544 19686 582 19689
rect 378 19649 450 19657
rect 428 19619 430 19635
rect 400 19611 430 19619
rect 476 19617 480 19685
rect 544 19656 552 19686
rect 578 19656 582 19686
rect 544 19647 548 19656
rect 400 19607 436 19611
rect 400 19577 408 19607
rect 420 19577 436 19607
rect 544 19609 548 19617
rect 12 19538 62 19540
rect 28 19529 59 19537
rect 62 19529 64 19538
rect 28 19521 64 19529
rect 127 19529 158 19537
rect 127 19522 182 19529
rect 215 19527 224 19555
rect 127 19521 161 19522
rect 59 19505 64 19521
rect 158 19505 161 19521
rect 28 19497 64 19505
rect 127 19504 161 19505
rect 127 19497 182 19504
rect 62 19488 64 19497
rect 213 19489 224 19527
rect 282 19517 292 19575
rect 296 19569 368 19577
rect 319 19539 346 19550
rect 318 19526 324 19539
rect 346 19526 348 19539
rect 428 19530 430 19577
rect 443 19567 450 19569
rect 476 19537 480 19605
rect 544 19575 552 19609
rect 578 19575 582 19609
rect 481 19543 517 19571
rect 481 19537 495 19543
rect 367 19526 380 19530
rect 251 19483 263 19517
rect 273 19483 293 19517
rect 295 19502 324 19526
rect 303 19492 316 19502
rect 318 19486 324 19502
rect 333 19502 380 19526
rect 333 19492 353 19502
rect 367 19496 380 19502
rect 396 19496 408 19530
rect 420 19496 436 19530
rect 120 19435 170 19437
rect 76 19429 92 19435
rect 94 19429 110 19435
rect 76 19419 99 19428
rect 60 19409 67 19419
rect 76 19399 77 19419
rect 96 19394 99 19419
rect 109 19399 110 19419
rect 119 19409 126 19419
rect 76 19385 110 19389
rect 170 19385 172 19435
rect 186 19417 190 19451
rect 216 19417 220 19451
rect 186 19340 220 19374
rect 282 19371 292 19483
rect 318 19476 335 19486
rect 318 19407 324 19476
rect 346 19407 348 19492
rect 428 19449 430 19496
rect 476 19459 480 19527
rect 485 19509 495 19537
rect 505 19537 519 19543
rect 544 19537 555 19575
rect 505 19509 525 19537
rect 544 19509 553 19537
rect 544 19489 548 19509
rect 579 19468 582 19558
rect 612 19540 624 19541
rect 599 19538 649 19540
rect 612 19537 624 19538
rect 610 19530 632 19537
rect 607 19529 632 19530
rect 586 19522 644 19529
rect 607 19521 644 19522
rect 607 19505 610 19521
rect 616 19505 644 19521
rect 607 19504 644 19505
rect 586 19497 644 19504
rect 607 19496 610 19497
rect 612 19489 632 19497
rect 612 19485 624 19489
rect 649 19488 651 19538
rect 544 19451 548 19459
rect 400 19419 408 19449
rect 420 19419 436 19449
rect 400 19415 436 19419
rect 400 19407 430 19415
rect 428 19391 430 19407
rect 476 19379 480 19447
rect 544 19417 552 19451
rect 578 19417 582 19451
rect 544 19409 548 19417
rect 544 19379 586 19380
rect 288 19339 292 19371
rect 296 19369 368 19377
rect 378 19369 450 19377
rect 544 19372 548 19379
rect 439 19341 444 19369
rect 120 19325 170 19327
rect 76 19321 130 19325
rect 110 19316 130 19321
rect 60 19291 67 19301
rect 76 19291 77 19311
rect 96 19282 99 19316
rect 109 19291 110 19311
rect 119 19291 126 19301
rect 76 19275 92 19281
rect 94 19275 110 19281
rect 170 19275 172 19325
rect 186 19259 190 19293
rect 216 19259 220 19293
rect 213 19227 224 19259
rect 282 19255 292 19339
rect 296 19333 368 19341
rect 378 19333 450 19341
rect 468 19338 473 19372
rect 428 19303 430 19319
rect 251 19227 292 19255
rect 318 19234 324 19303
rect 12 19222 62 19224
rect 28 19213 59 19221
rect 62 19213 64 19222
rect 251 19221 263 19227
rect 28 19205 64 19213
rect 127 19213 158 19221
rect 127 19206 182 19213
rect 127 19205 161 19206
rect 59 19189 64 19205
rect 158 19189 161 19205
rect 253 19193 263 19221
rect 273 19193 293 19227
rect 318 19224 335 19234
rect 303 19208 316 19218
rect 318 19208 324 19224
rect 346 19218 348 19303
rect 400 19295 430 19303
rect 476 19301 480 19369
rect 511 19338 582 19372
rect 544 19331 548 19338
rect 400 19291 436 19295
rect 400 19261 408 19291
rect 420 19261 436 19291
rect 544 19293 548 19301
rect 28 19181 64 19189
rect 127 19188 161 19189
rect 127 19181 182 19188
rect 62 19172 64 19181
rect 282 19135 292 19193
rect 295 19184 324 19208
rect 333 19208 353 19218
rect 428 19214 430 19261
rect 476 19221 480 19289
rect 544 19259 552 19293
rect 578 19259 582 19293
rect 544 19251 548 19259
rect 367 19208 380 19214
rect 333 19184 380 19208
rect 318 19171 324 19184
rect 346 19171 348 19184
rect 367 19180 380 19184
rect 396 19180 408 19214
rect 420 19180 436 19214
rect 544 19211 553 19239
rect 319 19160 346 19171
rect 120 19119 170 19121
rect 76 19113 92 19119
rect 94 19113 110 19119
rect 76 19103 99 19112
rect 60 19093 67 19103
rect 76 19083 77 19103
rect 96 19078 99 19103
rect 109 19083 110 19103
rect 119 19093 126 19103
rect 76 19069 110 19073
rect 170 19069 172 19119
rect 186 19101 190 19135
rect 216 19101 220 19135
rect 182 19063 224 19064
rect 186 19039 220 19056
rect 223 19039 257 19056
rect 182 19022 257 19039
rect 182 19021 224 19022
rect 160 19015 246 19021
rect 288 19015 292 19135
rect 296 19133 368 19141
rect 428 19133 430 19180
rect 476 19143 480 19211
rect 485 19167 495 19201
rect 505 19173 525 19201
rect 505 19167 519 19173
rect 544 19167 555 19211
rect 485 19143 492 19167
rect 579 19152 582 19242
rect 612 19224 624 19225
rect 599 19222 649 19224
rect 612 19221 624 19222
rect 610 19214 632 19221
rect 607 19213 632 19214
rect 586 19206 644 19213
rect 607 19205 644 19206
rect 607 19189 610 19205
rect 616 19189 644 19205
rect 607 19188 644 19189
rect 586 19181 644 19188
rect 607 19180 610 19181
rect 612 19173 632 19181
rect 612 19169 624 19173
rect 649 19172 651 19222
rect 544 19135 548 19143
rect 400 19103 408 19133
rect 420 19103 436 19133
rect 400 19099 436 19103
rect 400 19091 430 19099
rect 428 19075 430 19091
rect 476 19063 480 19131
rect 544 19101 552 19135
rect 578 19101 582 19135
rect 544 19093 548 19101
rect 295 19022 300 19056
rect 324 19022 329 19056
rect 378 19053 450 19061
rect 544 19058 548 19063
rect 544 19054 582 19058
rect 544 19039 552 19054
rect 578 19039 582 19054
rect 544 19021 586 19039
rect 522 19015 608 19021
rect 182 18999 224 19015
rect 544 18999 586 19015
rect 17 18985 67 18987
rect 119 18985 169 18987
rect 186 18985 220 18999
rect 548 18985 582 18999
rect 599 18985 649 18987
rect 42 18943 59 18977
rect 67 18935 69 18985
rect 160 18977 246 18985
rect 522 18977 608 18985
rect 76 18943 110 18977
rect 127 18943 144 18977
rect 152 18943 161 18977
rect 162 18975 195 18977
rect 224 18975 244 18977
rect 162 18943 244 18975
rect 524 18975 548 18977
rect 573 18975 582 18977
rect 586 18975 606 18977
rect 160 18935 246 18943
rect 186 18919 220 18935
rect 182 18905 224 18906
rect 160 18899 182 18905
rect 224 18899 246 18905
rect 186 18864 220 18898
rect 223 18864 257 18898
rect 120 18851 170 18853
rect 76 18847 130 18851
rect 110 18842 130 18847
rect 60 18817 67 18827
rect 76 18817 77 18837
rect 96 18808 99 18842
rect 109 18817 110 18837
rect 119 18817 126 18827
rect 76 18801 92 18807
rect 94 18801 110 18807
rect 170 18801 172 18851
rect 186 18785 190 18819
rect 216 18785 220 18819
rect 288 18785 292 18973
rect 476 18905 480 18973
rect 524 18943 606 18975
rect 607 18943 616 18977
rect 522 18935 608 18943
rect 649 18935 651 18985
rect 548 18919 582 18935
rect 522 18900 548 18905
rect 522 18899 582 18900
rect 586 18899 608 18905
rect 295 18864 300 18898
rect 324 18864 329 18898
rect 544 18896 582 18899
rect 378 18859 450 18867
rect 428 18829 430 18845
rect 400 18821 430 18829
rect 476 18827 480 18895
rect 544 18866 552 18896
rect 578 18866 582 18896
rect 544 18857 548 18866
rect 400 18817 436 18821
rect 400 18787 408 18817
rect 420 18787 436 18817
rect 544 18819 548 18827
rect 12 18748 62 18750
rect 28 18739 59 18747
rect 62 18739 64 18748
rect 28 18731 64 18739
rect 127 18739 158 18747
rect 127 18732 182 18739
rect 215 18737 224 18765
rect 127 18731 161 18732
rect 59 18715 64 18731
rect 158 18715 161 18731
rect 28 18707 64 18715
rect 127 18714 161 18715
rect 127 18707 182 18714
rect 62 18698 64 18707
rect 213 18699 224 18737
rect 282 18727 292 18785
rect 296 18779 368 18787
rect 319 18749 346 18760
rect 318 18736 324 18749
rect 346 18736 348 18749
rect 428 18740 430 18787
rect 443 18777 450 18779
rect 476 18747 480 18815
rect 544 18785 552 18819
rect 578 18785 582 18819
rect 481 18753 517 18781
rect 481 18747 495 18753
rect 367 18736 380 18740
rect 251 18693 263 18727
rect 273 18693 293 18727
rect 295 18712 324 18736
rect 303 18702 316 18712
rect 318 18696 324 18712
rect 333 18712 380 18736
rect 333 18702 353 18712
rect 367 18706 380 18712
rect 396 18706 408 18740
rect 420 18706 436 18740
rect 120 18645 170 18647
rect 76 18639 92 18645
rect 94 18639 110 18645
rect 76 18629 99 18638
rect 60 18619 67 18629
rect 76 18609 77 18629
rect 96 18604 99 18629
rect 109 18609 110 18629
rect 119 18619 126 18629
rect 76 18595 110 18599
rect 170 18595 172 18645
rect 186 18627 190 18661
rect 216 18627 220 18661
rect 186 18550 220 18584
rect 282 18581 292 18693
rect 318 18686 335 18696
rect 318 18617 324 18686
rect 346 18617 348 18702
rect 428 18659 430 18706
rect 476 18669 480 18737
rect 485 18719 495 18747
rect 505 18747 519 18753
rect 544 18747 555 18785
rect 505 18719 525 18747
rect 544 18719 553 18747
rect 544 18699 548 18719
rect 579 18678 582 18768
rect 612 18750 624 18751
rect 599 18748 649 18750
rect 612 18747 624 18748
rect 610 18740 632 18747
rect 607 18739 632 18740
rect 586 18732 644 18739
rect 607 18731 644 18732
rect 607 18715 610 18731
rect 616 18715 644 18731
rect 607 18714 644 18715
rect 586 18707 644 18714
rect 607 18706 610 18707
rect 612 18699 632 18707
rect 612 18695 624 18699
rect 649 18698 651 18748
rect 544 18661 548 18669
rect 400 18629 408 18659
rect 420 18629 436 18659
rect 400 18625 436 18629
rect 400 18617 430 18625
rect 428 18601 430 18617
rect 476 18589 480 18657
rect 544 18627 552 18661
rect 578 18627 582 18661
rect 544 18619 548 18627
rect 544 18589 586 18590
rect 288 18549 292 18581
rect 296 18579 368 18587
rect 378 18579 450 18587
rect 544 18582 548 18589
rect 439 18551 444 18579
rect 120 18535 170 18537
rect 76 18531 130 18535
rect 110 18526 130 18531
rect 60 18501 67 18511
rect 76 18501 77 18521
rect 96 18492 99 18526
rect 109 18501 110 18521
rect 119 18501 126 18511
rect 76 18485 92 18491
rect 94 18485 110 18491
rect 170 18485 172 18535
rect 186 18469 190 18503
rect 216 18469 220 18503
rect 213 18437 224 18469
rect 282 18465 292 18549
rect 296 18543 368 18551
rect 378 18543 450 18551
rect 468 18548 473 18582
rect 428 18513 430 18529
rect 251 18437 292 18465
rect 318 18444 324 18513
rect 12 18432 62 18434
rect 28 18423 59 18431
rect 62 18423 64 18432
rect 251 18431 263 18437
rect 28 18415 64 18423
rect 127 18423 158 18431
rect 127 18416 182 18423
rect 127 18415 161 18416
rect 59 18399 64 18415
rect 158 18399 161 18415
rect 253 18403 263 18431
rect 273 18403 293 18437
rect 318 18434 335 18444
rect 303 18418 316 18428
rect 318 18418 324 18434
rect 346 18428 348 18513
rect 400 18505 430 18513
rect 476 18511 480 18579
rect 511 18548 582 18582
rect 544 18541 548 18548
rect 400 18501 436 18505
rect 400 18471 408 18501
rect 420 18471 436 18501
rect 544 18503 548 18511
rect 28 18391 64 18399
rect 127 18398 161 18399
rect 127 18391 182 18398
rect 62 18382 64 18391
rect 282 18345 292 18403
rect 295 18394 324 18418
rect 333 18418 353 18428
rect 428 18424 430 18471
rect 476 18431 480 18499
rect 544 18469 552 18503
rect 578 18469 582 18503
rect 544 18461 548 18469
rect 367 18418 380 18424
rect 333 18394 380 18418
rect 318 18381 324 18394
rect 346 18381 348 18394
rect 367 18390 380 18394
rect 396 18390 408 18424
rect 420 18390 436 18424
rect 544 18421 553 18449
rect 319 18370 346 18381
rect 120 18329 170 18331
rect 76 18323 92 18329
rect 94 18323 110 18329
rect 76 18313 99 18322
rect 60 18303 67 18313
rect 76 18293 77 18313
rect 96 18288 99 18313
rect 109 18293 110 18313
rect 119 18303 126 18313
rect 76 18279 110 18283
rect 170 18279 172 18329
rect 186 18311 190 18345
rect 216 18311 220 18345
rect 182 18273 224 18274
rect 186 18249 220 18266
rect 223 18249 257 18266
rect 182 18232 257 18249
rect 182 18231 224 18232
rect 160 18225 246 18231
rect 288 18225 292 18345
rect 296 18343 368 18351
rect 428 18343 430 18390
rect 476 18353 480 18421
rect 485 18377 495 18411
rect 505 18383 525 18411
rect 505 18377 519 18383
rect 544 18377 555 18421
rect 485 18353 492 18377
rect 579 18362 582 18452
rect 612 18434 624 18435
rect 599 18432 649 18434
rect 612 18431 624 18432
rect 610 18424 632 18431
rect 607 18423 632 18424
rect 586 18416 644 18423
rect 607 18415 644 18416
rect 607 18399 610 18415
rect 616 18399 644 18415
rect 607 18398 644 18399
rect 586 18391 644 18398
rect 607 18390 610 18391
rect 612 18383 632 18391
rect 612 18379 624 18383
rect 649 18382 651 18432
rect 544 18345 548 18353
rect 400 18313 408 18343
rect 420 18313 436 18343
rect 400 18309 436 18313
rect 400 18301 430 18309
rect 428 18285 430 18301
rect 476 18273 480 18341
rect 544 18311 552 18345
rect 578 18311 582 18345
rect 544 18303 548 18311
rect 295 18232 300 18266
rect 324 18232 329 18266
rect 378 18263 450 18271
rect 544 18268 548 18273
rect 544 18264 582 18268
rect 544 18249 552 18264
rect 578 18249 582 18264
rect 544 18231 586 18249
rect 522 18225 608 18231
rect 182 18209 224 18225
rect 544 18209 586 18225
rect 17 18195 67 18197
rect 119 18195 169 18197
rect 186 18195 220 18209
rect 548 18195 582 18209
rect 599 18195 649 18197
rect 42 18153 59 18187
rect 67 18145 69 18195
rect 160 18187 246 18195
rect 522 18187 608 18195
rect 76 18153 110 18187
rect 127 18153 144 18187
rect 152 18153 161 18187
rect 162 18185 195 18187
rect 224 18185 244 18187
rect 162 18153 244 18185
rect 524 18185 548 18187
rect 573 18185 582 18187
rect 586 18185 606 18187
rect 160 18145 246 18153
rect 186 18129 220 18145
rect 182 18115 224 18116
rect 160 18109 182 18115
rect 224 18109 246 18115
rect 186 18074 220 18108
rect 223 18074 257 18108
rect 120 18061 170 18063
rect 76 18057 130 18061
rect 110 18052 130 18057
rect 60 18027 67 18037
rect 76 18027 77 18047
rect 96 18018 99 18052
rect 109 18027 110 18047
rect 119 18027 126 18037
rect 76 18011 92 18017
rect 94 18011 110 18017
rect 170 18011 172 18061
rect 186 17995 190 18029
rect 216 17995 220 18029
rect 288 17995 292 18183
rect 476 18115 480 18183
rect 524 18153 606 18185
rect 607 18153 616 18187
rect 522 18145 608 18153
rect 649 18145 651 18195
rect 548 18129 582 18145
rect 522 18110 548 18115
rect 522 18109 582 18110
rect 586 18109 608 18115
rect 295 18074 300 18108
rect 324 18074 329 18108
rect 544 18106 582 18109
rect 378 18069 450 18077
rect 428 18039 430 18055
rect 400 18031 430 18039
rect 476 18037 480 18105
rect 544 18076 552 18106
rect 578 18076 582 18106
rect 544 18067 548 18076
rect 400 18027 436 18031
rect 400 17997 408 18027
rect 420 17997 436 18027
rect 544 18029 548 18037
rect 12 17958 62 17960
rect 28 17949 59 17957
rect 62 17949 64 17958
rect 28 17941 64 17949
rect 127 17949 158 17957
rect 127 17942 182 17949
rect 215 17947 224 17975
rect 127 17941 161 17942
rect 59 17925 64 17941
rect 158 17925 161 17941
rect 28 17917 64 17925
rect 127 17924 161 17925
rect 127 17917 182 17924
rect 62 17908 64 17917
rect 213 17909 224 17947
rect 282 17937 292 17995
rect 296 17989 368 17997
rect 319 17959 346 17970
rect 318 17946 324 17959
rect 346 17946 348 17959
rect 428 17950 430 17997
rect 443 17987 450 17989
rect 476 17957 480 18025
rect 544 17995 552 18029
rect 578 17995 582 18029
rect 481 17963 517 17991
rect 481 17957 495 17963
rect 367 17946 380 17950
rect 251 17903 263 17937
rect 273 17903 293 17937
rect 295 17922 324 17946
rect 303 17912 316 17922
rect 318 17906 324 17922
rect 333 17922 380 17946
rect 333 17912 353 17922
rect 367 17916 380 17922
rect 396 17916 408 17950
rect 420 17916 436 17950
rect 120 17855 170 17857
rect 76 17849 92 17855
rect 94 17849 110 17855
rect 76 17839 99 17848
rect 60 17829 67 17839
rect 76 17819 77 17839
rect 96 17814 99 17839
rect 109 17819 110 17839
rect 119 17829 126 17839
rect 76 17805 110 17809
rect 170 17805 172 17855
rect 186 17837 190 17871
rect 216 17837 220 17871
rect 186 17760 220 17794
rect 282 17791 292 17903
rect 318 17896 335 17906
rect 318 17827 324 17896
rect 346 17827 348 17912
rect 428 17869 430 17916
rect 476 17879 480 17947
rect 485 17929 495 17957
rect 505 17957 519 17963
rect 544 17957 555 17995
rect 505 17929 525 17957
rect 544 17929 553 17957
rect 544 17909 548 17929
rect 579 17888 582 17978
rect 612 17960 624 17961
rect 599 17958 649 17960
rect 612 17957 624 17958
rect 610 17950 632 17957
rect 607 17949 632 17950
rect 586 17942 644 17949
rect 607 17941 644 17942
rect 607 17925 610 17941
rect 616 17925 644 17941
rect 607 17924 644 17925
rect 586 17917 644 17924
rect 607 17916 610 17917
rect 612 17909 632 17917
rect 612 17905 624 17909
rect 649 17908 651 17958
rect 544 17871 548 17879
rect 400 17839 408 17869
rect 420 17839 436 17869
rect 400 17835 436 17839
rect 400 17827 430 17835
rect 428 17811 430 17827
rect 476 17799 480 17867
rect 544 17837 552 17871
rect 578 17837 582 17871
rect 544 17829 548 17837
rect 544 17799 586 17800
rect 288 17759 292 17791
rect 296 17789 368 17797
rect 378 17789 450 17797
rect 544 17792 548 17799
rect 439 17761 444 17789
rect 120 17745 170 17747
rect 76 17741 130 17745
rect 110 17736 130 17741
rect 60 17711 67 17721
rect 76 17711 77 17731
rect 96 17702 99 17736
rect 109 17711 110 17731
rect 119 17711 126 17721
rect 76 17695 92 17701
rect 94 17695 110 17701
rect 170 17695 172 17745
rect 186 17679 190 17713
rect 216 17679 220 17713
rect 213 17647 224 17679
rect 282 17675 292 17759
rect 296 17753 368 17761
rect 378 17753 450 17761
rect 468 17758 473 17792
rect 428 17723 430 17739
rect 251 17647 292 17675
rect 318 17654 324 17723
rect 12 17642 62 17644
rect 28 17633 59 17641
rect 62 17633 64 17642
rect 251 17641 263 17647
rect 28 17625 64 17633
rect 127 17633 158 17641
rect 127 17626 182 17633
rect 127 17625 161 17626
rect 59 17609 64 17625
rect 158 17609 161 17625
rect 253 17613 263 17641
rect 273 17613 293 17647
rect 318 17644 335 17654
rect 303 17628 316 17638
rect 318 17628 324 17644
rect 346 17638 348 17723
rect 400 17715 430 17723
rect 476 17721 480 17789
rect 511 17758 582 17792
rect 544 17751 548 17758
rect 400 17711 436 17715
rect 400 17681 408 17711
rect 420 17681 436 17711
rect 544 17713 548 17721
rect 28 17601 64 17609
rect 127 17608 161 17609
rect 127 17601 182 17608
rect 62 17592 64 17601
rect 282 17555 292 17613
rect 295 17604 324 17628
rect 333 17628 353 17638
rect 428 17634 430 17681
rect 476 17641 480 17709
rect 544 17679 552 17713
rect 578 17679 582 17713
rect 544 17671 548 17679
rect 367 17628 380 17634
rect 333 17604 380 17628
rect 318 17591 324 17604
rect 346 17591 348 17604
rect 367 17600 380 17604
rect 396 17600 408 17634
rect 420 17600 436 17634
rect 544 17631 553 17659
rect 319 17580 346 17591
rect 120 17539 170 17541
rect 76 17533 92 17539
rect 94 17533 110 17539
rect 76 17523 99 17532
rect 60 17513 67 17523
rect 76 17503 77 17523
rect 96 17498 99 17523
rect 109 17503 110 17523
rect 119 17513 126 17523
rect 76 17489 110 17493
rect 170 17489 172 17539
rect 186 17521 190 17555
rect 216 17521 220 17555
rect 182 17483 224 17484
rect 186 17459 220 17476
rect 223 17459 257 17476
rect 182 17442 257 17459
rect 182 17441 224 17442
rect 160 17435 246 17441
rect 288 17435 292 17555
rect 296 17553 368 17561
rect 428 17553 430 17600
rect 476 17563 480 17631
rect 485 17587 495 17621
rect 505 17593 525 17621
rect 505 17587 519 17593
rect 544 17587 555 17631
rect 485 17563 492 17587
rect 579 17572 582 17662
rect 612 17644 624 17645
rect 599 17642 649 17644
rect 612 17641 624 17642
rect 610 17634 632 17641
rect 607 17633 632 17634
rect 586 17626 644 17633
rect 607 17625 644 17626
rect 607 17609 610 17625
rect 616 17609 644 17625
rect 607 17608 644 17609
rect 586 17601 644 17608
rect 607 17600 610 17601
rect 612 17593 632 17601
rect 612 17589 624 17593
rect 649 17592 651 17642
rect 544 17555 548 17563
rect 400 17523 408 17553
rect 420 17523 436 17553
rect 400 17519 436 17523
rect 400 17511 430 17519
rect 428 17495 430 17511
rect 476 17483 480 17551
rect 544 17521 552 17555
rect 578 17521 582 17555
rect 544 17513 548 17521
rect 295 17442 300 17476
rect 324 17442 329 17476
rect 378 17473 450 17481
rect 544 17478 548 17483
rect 544 17474 582 17478
rect 544 17459 552 17474
rect 578 17459 582 17474
rect 544 17441 586 17459
rect 522 17435 608 17441
rect 182 17419 224 17435
rect 544 17419 586 17435
rect 17 17405 67 17407
rect 119 17405 169 17407
rect 186 17405 220 17419
rect 548 17405 582 17419
rect 599 17405 649 17407
rect 42 17363 59 17397
rect 67 17355 69 17405
rect 160 17397 246 17405
rect 522 17397 608 17405
rect 76 17363 110 17397
rect 127 17363 144 17397
rect 152 17363 161 17397
rect 162 17395 195 17397
rect 224 17395 244 17397
rect 162 17363 244 17395
rect 524 17395 548 17397
rect 573 17395 582 17397
rect 586 17395 606 17397
rect 160 17355 246 17363
rect 186 17339 220 17355
rect 182 17325 224 17326
rect 160 17319 182 17325
rect 224 17319 246 17325
rect 186 17284 220 17318
rect 223 17284 257 17318
rect 120 17271 170 17273
rect 76 17267 130 17271
rect 110 17262 130 17267
rect 60 17237 67 17247
rect 76 17237 77 17257
rect 96 17228 99 17262
rect 109 17237 110 17257
rect 119 17237 126 17247
rect 76 17221 92 17227
rect 94 17221 110 17227
rect 170 17221 172 17271
rect 186 17205 190 17239
rect 216 17205 220 17239
rect 288 17205 292 17393
rect 476 17325 480 17393
rect 524 17363 606 17395
rect 607 17363 616 17397
rect 522 17355 608 17363
rect 649 17355 651 17405
rect 548 17339 582 17355
rect 522 17320 548 17325
rect 522 17319 582 17320
rect 586 17319 608 17325
rect 295 17284 300 17318
rect 324 17284 329 17318
rect 544 17316 582 17319
rect 378 17279 450 17287
rect 428 17249 430 17265
rect 400 17241 430 17249
rect 476 17247 480 17315
rect 544 17286 552 17316
rect 578 17286 582 17316
rect 544 17277 548 17286
rect 400 17237 436 17241
rect 400 17207 408 17237
rect 420 17207 436 17237
rect 544 17239 548 17247
rect 12 17168 62 17170
rect 28 17159 59 17167
rect 62 17159 64 17168
rect 28 17151 64 17159
rect 127 17159 158 17167
rect 127 17152 182 17159
rect 215 17157 224 17185
rect 127 17151 161 17152
rect 59 17135 64 17151
rect 158 17135 161 17151
rect 28 17127 64 17135
rect 127 17134 161 17135
rect 127 17127 182 17134
rect 62 17118 64 17127
rect 213 17119 224 17157
rect 282 17147 292 17205
rect 296 17199 368 17207
rect 319 17169 346 17180
rect 318 17156 324 17169
rect 346 17156 348 17169
rect 428 17160 430 17207
rect 443 17197 450 17199
rect 476 17167 480 17235
rect 544 17205 552 17239
rect 578 17205 582 17239
rect 481 17173 517 17201
rect 481 17167 495 17173
rect 367 17156 380 17160
rect 251 17113 263 17147
rect 273 17113 293 17147
rect 295 17132 324 17156
rect 303 17122 316 17132
rect 318 17116 324 17132
rect 333 17132 380 17156
rect 333 17122 353 17132
rect 367 17126 380 17132
rect 396 17126 408 17160
rect 420 17126 436 17160
rect 120 17065 170 17067
rect 76 17059 92 17065
rect 94 17059 110 17065
rect 76 17049 99 17058
rect 60 17039 67 17049
rect 76 17029 77 17049
rect 96 17024 99 17049
rect 109 17029 110 17049
rect 119 17039 126 17049
rect 76 17015 110 17019
rect 170 17015 172 17065
rect 186 17047 190 17081
rect 216 17047 220 17081
rect 186 16970 220 17004
rect 282 17001 292 17113
rect 318 17106 335 17116
rect 318 17037 324 17106
rect 346 17037 348 17122
rect 428 17079 430 17126
rect 476 17089 480 17157
rect 485 17139 495 17167
rect 505 17167 519 17173
rect 544 17167 555 17205
rect 505 17139 525 17167
rect 544 17139 553 17167
rect 544 17119 548 17139
rect 579 17098 582 17188
rect 612 17170 624 17171
rect 599 17168 649 17170
rect 612 17167 624 17168
rect 610 17160 632 17167
rect 607 17159 632 17160
rect 586 17152 644 17159
rect 607 17151 644 17152
rect 607 17135 610 17151
rect 616 17135 644 17151
rect 607 17134 644 17135
rect 586 17127 644 17134
rect 607 17126 610 17127
rect 612 17119 632 17127
rect 612 17115 624 17119
rect 649 17118 651 17168
rect 544 17081 548 17089
rect 400 17049 408 17079
rect 420 17049 436 17079
rect 400 17045 436 17049
rect 400 17037 430 17045
rect 428 17021 430 17037
rect 476 17009 480 17077
rect 544 17047 552 17081
rect 578 17047 582 17081
rect 544 17039 548 17047
rect 544 17009 586 17010
rect 288 16969 292 17001
rect 296 16999 368 17007
rect 378 16999 450 17007
rect 544 17002 548 17009
rect 439 16971 444 16999
rect 120 16955 170 16957
rect 76 16951 130 16955
rect 110 16946 130 16951
rect 60 16921 67 16931
rect 76 16921 77 16941
rect 96 16912 99 16946
rect 109 16921 110 16941
rect 119 16921 126 16931
rect 76 16905 92 16911
rect 94 16905 110 16911
rect 170 16905 172 16955
rect 186 16889 190 16923
rect 216 16889 220 16923
rect 213 16857 224 16889
rect 282 16885 292 16969
rect 296 16963 368 16971
rect 378 16963 450 16971
rect 468 16968 473 17002
rect 428 16933 430 16949
rect 251 16857 292 16885
rect 318 16864 324 16933
rect 12 16852 62 16854
rect 28 16843 59 16851
rect 62 16843 64 16852
rect 251 16851 263 16857
rect 28 16835 64 16843
rect 127 16843 158 16851
rect 127 16836 182 16843
rect 127 16835 161 16836
rect 59 16819 64 16835
rect 158 16819 161 16835
rect 253 16823 263 16851
rect 273 16823 293 16857
rect 318 16854 335 16864
rect 303 16838 316 16848
rect 318 16838 324 16854
rect 346 16848 348 16933
rect 400 16925 430 16933
rect 476 16931 480 16999
rect 511 16968 582 17002
rect 544 16961 548 16968
rect 400 16921 436 16925
rect 400 16891 408 16921
rect 420 16891 436 16921
rect 544 16923 548 16931
rect 28 16811 64 16819
rect 127 16818 161 16819
rect 127 16811 182 16818
rect 62 16802 64 16811
rect 282 16765 292 16823
rect 295 16814 324 16838
rect 333 16838 353 16848
rect 428 16844 430 16891
rect 476 16851 480 16919
rect 544 16889 552 16923
rect 578 16889 582 16923
rect 544 16881 548 16889
rect 367 16838 380 16844
rect 333 16814 380 16838
rect 318 16801 324 16814
rect 346 16801 348 16814
rect 367 16810 380 16814
rect 396 16810 408 16844
rect 420 16810 436 16844
rect 544 16841 553 16869
rect 319 16790 346 16801
rect 120 16749 170 16751
rect 76 16743 92 16749
rect 94 16743 110 16749
rect 76 16733 99 16742
rect 60 16723 67 16733
rect 76 16713 77 16733
rect 96 16708 99 16733
rect 109 16713 110 16733
rect 119 16723 126 16733
rect 76 16699 110 16703
rect 170 16699 172 16749
rect 186 16731 190 16765
rect 216 16731 220 16765
rect 182 16693 224 16694
rect 186 16669 220 16686
rect 223 16669 257 16686
rect 182 16652 257 16669
rect 182 16651 224 16652
rect 160 16645 246 16651
rect 288 16645 292 16765
rect 296 16763 368 16771
rect 428 16763 430 16810
rect 476 16773 480 16841
rect 485 16797 495 16831
rect 505 16803 525 16831
rect 505 16797 519 16803
rect 544 16797 555 16841
rect 485 16773 492 16797
rect 579 16782 582 16872
rect 612 16854 624 16855
rect 599 16852 649 16854
rect 612 16851 624 16852
rect 610 16844 632 16851
rect 607 16843 632 16844
rect 586 16836 644 16843
rect 607 16835 644 16836
rect 607 16819 610 16835
rect 616 16819 644 16835
rect 607 16818 644 16819
rect 586 16811 644 16818
rect 607 16810 610 16811
rect 612 16803 632 16811
rect 612 16799 624 16803
rect 649 16802 651 16852
rect 544 16765 548 16773
rect 400 16733 408 16763
rect 420 16733 436 16763
rect 400 16729 436 16733
rect 400 16721 430 16729
rect 428 16705 430 16721
rect 476 16693 480 16761
rect 544 16731 552 16765
rect 578 16731 582 16765
rect 544 16723 548 16731
rect 295 16652 300 16686
rect 324 16652 329 16686
rect 378 16683 450 16691
rect 544 16688 548 16693
rect 544 16684 582 16688
rect 544 16669 552 16684
rect 578 16669 582 16684
rect 544 16651 586 16669
rect 522 16645 608 16651
rect 182 16629 224 16645
rect 544 16629 586 16645
rect 17 16615 67 16617
rect 119 16615 169 16617
rect 186 16615 220 16629
rect 548 16615 582 16629
rect 599 16615 649 16617
rect 42 16573 59 16607
rect 67 16565 69 16615
rect 160 16607 246 16615
rect 522 16607 608 16615
rect 76 16573 110 16607
rect 127 16573 144 16607
rect 152 16573 161 16607
rect 162 16605 195 16607
rect 224 16605 244 16607
rect 162 16573 244 16605
rect 524 16605 548 16607
rect 573 16605 582 16607
rect 586 16605 606 16607
rect 160 16565 246 16573
rect 186 16549 220 16565
rect 182 16535 224 16536
rect 160 16529 182 16535
rect 224 16529 246 16535
rect 186 16494 220 16528
rect 223 16494 257 16528
rect 120 16481 170 16483
rect 76 16477 130 16481
rect 110 16472 130 16477
rect 60 16447 67 16457
rect 76 16447 77 16467
rect 96 16438 99 16472
rect 109 16447 110 16467
rect 119 16447 126 16457
rect 76 16431 92 16437
rect 94 16431 110 16437
rect 170 16431 172 16481
rect 186 16415 190 16449
rect 216 16415 220 16449
rect 288 16415 292 16603
rect 476 16535 480 16603
rect 524 16573 606 16605
rect 607 16573 616 16607
rect 522 16565 608 16573
rect 649 16565 651 16615
rect 548 16549 582 16565
rect 522 16530 548 16535
rect 522 16529 582 16530
rect 586 16529 608 16535
rect 295 16494 300 16528
rect 324 16494 329 16528
rect 544 16526 582 16529
rect 378 16489 450 16497
rect 428 16459 430 16475
rect 400 16451 430 16459
rect 476 16457 480 16525
rect 544 16496 552 16526
rect 578 16496 582 16526
rect 544 16487 548 16496
rect 400 16447 436 16451
rect 400 16417 408 16447
rect 420 16417 436 16447
rect 544 16449 548 16457
rect 12 16378 62 16380
rect 28 16369 59 16377
rect 62 16369 64 16378
rect 28 16361 64 16369
rect 127 16369 158 16377
rect 127 16362 182 16369
rect 215 16367 224 16395
rect 127 16361 161 16362
rect 59 16345 64 16361
rect 158 16345 161 16361
rect 28 16337 64 16345
rect 127 16344 161 16345
rect 127 16337 182 16344
rect 62 16328 64 16337
rect 213 16329 224 16367
rect 282 16357 292 16415
rect 296 16409 368 16417
rect 319 16379 346 16390
rect 318 16366 324 16379
rect 346 16366 348 16379
rect 428 16370 430 16417
rect 443 16407 450 16409
rect 476 16377 480 16445
rect 544 16415 552 16449
rect 578 16415 582 16449
rect 481 16383 517 16411
rect 481 16377 495 16383
rect 367 16366 380 16370
rect 251 16323 263 16357
rect 273 16323 293 16357
rect 295 16342 324 16366
rect 303 16332 316 16342
rect 318 16326 324 16342
rect 333 16342 380 16366
rect 333 16332 353 16342
rect 367 16336 380 16342
rect 396 16336 408 16370
rect 420 16336 436 16370
rect 120 16275 170 16277
rect 76 16269 92 16275
rect 94 16269 110 16275
rect 76 16259 99 16268
rect 60 16249 67 16259
rect 76 16239 77 16259
rect 96 16234 99 16259
rect 109 16239 110 16259
rect 119 16249 126 16259
rect 76 16225 110 16229
rect 170 16225 172 16275
rect 186 16257 190 16291
rect 216 16257 220 16291
rect 186 16180 220 16214
rect 282 16211 292 16323
rect 318 16316 335 16326
rect 318 16247 324 16316
rect 346 16247 348 16332
rect 428 16289 430 16336
rect 476 16299 480 16367
rect 485 16349 495 16377
rect 505 16377 519 16383
rect 544 16377 555 16415
rect 505 16349 525 16377
rect 544 16349 553 16377
rect 544 16329 548 16349
rect 579 16308 582 16398
rect 612 16380 624 16381
rect 599 16378 649 16380
rect 612 16377 624 16378
rect 610 16370 632 16377
rect 607 16369 632 16370
rect 586 16362 644 16369
rect 607 16361 644 16362
rect 607 16345 610 16361
rect 616 16345 644 16361
rect 607 16344 644 16345
rect 586 16337 644 16344
rect 607 16336 610 16337
rect 612 16329 632 16337
rect 612 16325 624 16329
rect 649 16328 651 16378
rect 544 16291 548 16299
rect 400 16259 408 16289
rect 420 16259 436 16289
rect 400 16255 436 16259
rect 400 16247 430 16255
rect 428 16231 430 16247
rect 476 16219 480 16287
rect 544 16257 552 16291
rect 578 16257 582 16291
rect 544 16249 548 16257
rect 544 16219 586 16220
rect 288 16179 292 16211
rect 296 16209 368 16217
rect 378 16209 450 16217
rect 544 16212 548 16219
rect 439 16181 444 16209
rect 120 16165 170 16167
rect 76 16161 130 16165
rect 110 16156 130 16161
rect 60 16131 67 16141
rect 76 16131 77 16151
rect 96 16122 99 16156
rect 109 16131 110 16151
rect 119 16131 126 16141
rect 76 16115 92 16121
rect 94 16115 110 16121
rect 170 16115 172 16165
rect 186 16099 190 16133
rect 216 16099 220 16133
rect 213 16067 224 16099
rect 282 16095 292 16179
rect 296 16173 368 16181
rect 378 16173 450 16181
rect 468 16178 473 16212
rect 428 16143 430 16159
rect 251 16067 292 16095
rect 318 16074 324 16143
rect 12 16062 62 16064
rect 28 16053 59 16061
rect 62 16053 64 16062
rect 251 16061 263 16067
rect 28 16045 64 16053
rect 127 16053 158 16061
rect 127 16046 182 16053
rect 127 16045 161 16046
rect 59 16029 64 16045
rect 158 16029 161 16045
rect 253 16033 263 16061
rect 273 16033 293 16067
rect 318 16064 335 16074
rect 303 16048 316 16058
rect 318 16048 324 16064
rect 346 16058 348 16143
rect 400 16135 430 16143
rect 476 16141 480 16209
rect 511 16178 582 16212
rect 544 16171 548 16178
rect 400 16131 436 16135
rect 400 16101 408 16131
rect 420 16101 436 16131
rect 544 16133 548 16141
rect 28 16021 64 16029
rect 127 16028 161 16029
rect 127 16021 182 16028
rect 62 16012 64 16021
rect 282 15975 292 16033
rect 295 16024 324 16048
rect 333 16048 353 16058
rect 428 16054 430 16101
rect 476 16061 480 16129
rect 544 16099 552 16133
rect 578 16099 582 16133
rect 544 16091 548 16099
rect 367 16048 380 16054
rect 333 16024 380 16048
rect 318 16011 324 16024
rect 346 16011 348 16024
rect 367 16020 380 16024
rect 396 16020 408 16054
rect 420 16020 436 16054
rect 544 16051 553 16079
rect 319 16000 346 16011
rect 120 15959 170 15961
rect 76 15953 92 15959
rect 94 15953 110 15959
rect 76 15943 99 15952
rect 60 15933 67 15943
rect 76 15923 77 15943
rect 96 15918 99 15943
rect 109 15923 110 15943
rect 119 15933 126 15943
rect 76 15909 110 15913
rect 170 15909 172 15959
rect 186 15941 190 15975
rect 216 15941 220 15975
rect 182 15903 224 15904
rect 186 15879 220 15896
rect 223 15879 257 15896
rect 182 15862 257 15879
rect 182 15861 224 15862
rect 160 15855 246 15861
rect 288 15855 292 15975
rect 296 15973 368 15981
rect 428 15973 430 16020
rect 476 15983 480 16051
rect 485 16007 495 16041
rect 505 16013 525 16041
rect 505 16007 519 16013
rect 544 16007 555 16051
rect 485 15983 492 16007
rect 579 15992 582 16082
rect 612 16064 624 16065
rect 599 16062 649 16064
rect 612 16061 624 16062
rect 610 16054 632 16061
rect 607 16053 632 16054
rect 586 16046 644 16053
rect 607 16045 644 16046
rect 607 16029 610 16045
rect 616 16029 644 16045
rect 607 16028 644 16029
rect 586 16021 644 16028
rect 607 16020 610 16021
rect 612 16013 632 16021
rect 612 16009 624 16013
rect 649 16012 651 16062
rect 544 15975 548 15983
rect 400 15943 408 15973
rect 420 15943 436 15973
rect 400 15939 436 15943
rect 400 15931 430 15939
rect 428 15915 430 15931
rect 476 15903 480 15971
rect 544 15941 552 15975
rect 578 15941 582 15975
rect 544 15933 548 15941
rect 295 15862 300 15896
rect 324 15862 329 15896
rect 378 15893 450 15901
rect 544 15898 548 15903
rect 544 15894 582 15898
rect 544 15879 552 15894
rect 578 15879 582 15894
rect 544 15861 586 15879
rect 522 15855 608 15861
rect 182 15839 224 15855
rect 544 15839 586 15855
rect 17 15825 67 15827
rect 119 15825 169 15827
rect 186 15825 220 15839
rect 548 15825 582 15839
rect 599 15825 649 15827
rect 42 15783 59 15817
rect 67 15775 69 15825
rect 160 15817 246 15825
rect 522 15817 608 15825
rect 76 15783 110 15817
rect 127 15783 144 15817
rect 152 15783 161 15817
rect 162 15815 195 15817
rect 224 15815 244 15817
rect 162 15783 244 15815
rect 524 15815 548 15817
rect 573 15815 582 15817
rect 586 15815 606 15817
rect 160 15775 246 15783
rect 186 15759 220 15775
rect 182 15745 224 15746
rect 160 15739 182 15745
rect 224 15739 246 15745
rect 186 15704 220 15738
rect 223 15704 257 15738
rect 120 15691 170 15693
rect 76 15687 130 15691
rect 110 15682 130 15687
rect 60 15657 67 15667
rect 76 15657 77 15677
rect 96 15648 99 15682
rect 109 15657 110 15677
rect 119 15657 126 15667
rect 76 15641 92 15647
rect 94 15641 110 15647
rect 170 15641 172 15691
rect 186 15625 190 15659
rect 216 15625 220 15659
rect 288 15625 292 15813
rect 476 15745 480 15813
rect 524 15783 606 15815
rect 607 15783 616 15817
rect 522 15775 608 15783
rect 649 15775 651 15825
rect 548 15759 582 15775
rect 522 15740 548 15745
rect 522 15739 582 15740
rect 586 15739 608 15745
rect 295 15704 300 15738
rect 324 15704 329 15738
rect 544 15736 582 15739
rect 378 15699 450 15707
rect 428 15669 430 15685
rect 400 15661 430 15669
rect 476 15667 480 15735
rect 544 15706 552 15736
rect 578 15706 582 15736
rect 544 15697 548 15706
rect 400 15657 436 15661
rect 400 15627 408 15657
rect 420 15627 436 15657
rect 544 15659 548 15667
rect 12 15588 62 15590
rect 28 15579 59 15587
rect 62 15579 64 15588
rect 28 15571 64 15579
rect 127 15579 158 15587
rect 127 15572 182 15579
rect 215 15577 224 15605
rect 127 15571 161 15572
rect 59 15555 64 15571
rect 158 15555 161 15571
rect 28 15547 64 15555
rect 127 15554 161 15555
rect 127 15547 182 15554
rect 62 15538 64 15547
rect 213 15539 224 15577
rect 282 15567 292 15625
rect 296 15619 368 15627
rect 319 15589 346 15600
rect 318 15576 324 15589
rect 346 15576 348 15589
rect 428 15580 430 15627
rect 443 15617 450 15619
rect 476 15587 480 15655
rect 544 15625 552 15659
rect 578 15625 582 15659
rect 481 15593 517 15621
rect 481 15587 495 15593
rect 367 15576 380 15580
rect 251 15533 263 15567
rect 273 15533 293 15567
rect 295 15552 324 15576
rect 303 15542 316 15552
rect 318 15536 324 15552
rect 333 15552 380 15576
rect 333 15542 353 15552
rect 367 15546 380 15552
rect 396 15546 408 15580
rect 420 15546 436 15580
rect 120 15485 170 15487
rect 76 15479 92 15485
rect 94 15479 110 15485
rect 76 15469 99 15478
rect 60 15459 67 15469
rect 76 15449 77 15469
rect 96 15444 99 15469
rect 109 15449 110 15469
rect 119 15459 126 15469
rect 76 15435 110 15439
rect 170 15435 172 15485
rect 186 15467 190 15501
rect 216 15467 220 15501
rect 186 15390 220 15424
rect 282 15421 292 15533
rect 318 15526 335 15536
rect 318 15457 324 15526
rect 346 15457 348 15542
rect 428 15499 430 15546
rect 476 15509 480 15577
rect 485 15559 495 15587
rect 505 15587 519 15593
rect 544 15587 555 15625
rect 505 15559 525 15587
rect 544 15559 553 15587
rect 544 15539 548 15559
rect 579 15518 582 15608
rect 612 15590 624 15591
rect 599 15588 649 15590
rect 612 15587 624 15588
rect 610 15580 632 15587
rect 607 15579 632 15580
rect 586 15572 644 15579
rect 607 15571 644 15572
rect 607 15555 610 15571
rect 616 15555 644 15571
rect 607 15554 644 15555
rect 586 15547 644 15554
rect 607 15546 610 15547
rect 612 15539 632 15547
rect 612 15535 624 15539
rect 649 15538 651 15588
rect 544 15501 548 15509
rect 400 15469 408 15499
rect 420 15469 436 15499
rect 400 15465 436 15469
rect 400 15457 430 15465
rect 428 15441 430 15457
rect 476 15429 480 15497
rect 544 15467 552 15501
rect 578 15467 582 15501
rect 544 15459 548 15467
rect 544 15429 586 15430
rect 288 15389 292 15421
rect 296 15419 368 15427
rect 378 15419 450 15427
rect 544 15422 548 15429
rect 439 15391 444 15419
rect 120 15375 170 15377
rect 76 15371 130 15375
rect 110 15366 130 15371
rect 60 15341 67 15351
rect 76 15341 77 15361
rect 96 15332 99 15366
rect 109 15341 110 15361
rect 119 15341 126 15351
rect 76 15325 92 15331
rect 94 15325 110 15331
rect 170 15325 172 15375
rect 186 15309 190 15343
rect 216 15309 220 15343
rect 213 15277 224 15309
rect 282 15305 292 15389
rect 296 15383 368 15391
rect 378 15383 450 15391
rect 468 15388 473 15422
rect 428 15353 430 15369
rect 251 15277 292 15305
rect 318 15284 324 15353
rect 12 15272 62 15274
rect 28 15263 59 15271
rect 62 15263 64 15272
rect 251 15271 263 15277
rect 28 15255 64 15263
rect 127 15263 158 15271
rect 127 15256 182 15263
rect 127 15255 161 15256
rect 59 15239 64 15255
rect 158 15239 161 15255
rect 253 15243 263 15271
rect 273 15243 293 15277
rect 318 15274 335 15284
rect 303 15258 316 15268
rect 318 15258 324 15274
rect 346 15268 348 15353
rect 400 15345 430 15353
rect 476 15351 480 15419
rect 511 15388 582 15422
rect 544 15381 548 15388
rect 400 15341 436 15345
rect 400 15311 408 15341
rect 420 15311 436 15341
rect 544 15343 548 15351
rect 28 15231 64 15239
rect 127 15238 161 15239
rect 127 15231 182 15238
rect 62 15222 64 15231
rect 282 15185 292 15243
rect 295 15234 324 15258
rect 333 15258 353 15268
rect 428 15264 430 15311
rect 476 15271 480 15339
rect 544 15309 552 15343
rect 578 15309 582 15343
rect 544 15301 548 15309
rect 367 15258 380 15264
rect 333 15234 380 15258
rect 318 15221 324 15234
rect 346 15221 348 15234
rect 367 15230 380 15234
rect 396 15230 408 15264
rect 420 15230 436 15264
rect 544 15261 553 15289
rect 319 15210 346 15221
rect 120 15169 170 15171
rect 76 15163 92 15169
rect 94 15163 110 15169
rect 76 15153 99 15162
rect 60 15143 67 15153
rect 76 15133 77 15153
rect 96 15128 99 15153
rect 109 15133 110 15153
rect 119 15143 126 15153
rect 76 15119 110 15123
rect 170 15119 172 15169
rect 186 15151 190 15185
rect 216 15151 220 15185
rect 182 15113 224 15114
rect 186 15089 220 15106
rect 223 15089 257 15106
rect 182 15072 257 15089
rect 182 15071 224 15072
rect 160 15065 246 15071
rect 288 15065 292 15185
rect 296 15183 368 15191
rect 428 15183 430 15230
rect 476 15193 480 15261
rect 485 15217 495 15251
rect 505 15223 525 15251
rect 505 15217 519 15223
rect 544 15217 555 15261
rect 485 15193 492 15217
rect 579 15202 582 15292
rect 612 15274 624 15275
rect 599 15272 649 15274
rect 612 15271 624 15272
rect 610 15264 632 15271
rect 607 15263 632 15264
rect 586 15256 644 15263
rect 607 15255 644 15256
rect 607 15239 610 15255
rect 616 15239 644 15255
rect 607 15238 644 15239
rect 586 15231 644 15238
rect 607 15230 610 15231
rect 612 15223 632 15231
rect 612 15219 624 15223
rect 649 15222 651 15272
rect 544 15185 548 15193
rect 400 15153 408 15183
rect 420 15153 436 15183
rect 400 15149 436 15153
rect 400 15141 430 15149
rect 428 15125 430 15141
rect 476 15113 480 15181
rect 544 15151 552 15185
rect 578 15151 582 15185
rect 544 15143 548 15151
rect 295 15072 300 15106
rect 324 15072 329 15106
rect 378 15103 450 15111
rect 544 15108 548 15113
rect 544 15104 582 15108
rect 544 15089 552 15104
rect 578 15089 582 15104
rect 544 15071 586 15089
rect 522 15065 608 15071
rect 182 15049 224 15065
rect 544 15049 586 15065
rect 17 15035 67 15037
rect 119 15035 169 15037
rect 186 15035 220 15049
rect 548 15035 582 15049
rect 599 15035 649 15037
rect 42 14993 59 15027
rect 67 14985 69 15035
rect 160 15027 246 15035
rect 522 15027 608 15035
rect 76 14993 110 15027
rect 127 14993 144 15027
rect 152 14993 161 15027
rect 162 15025 195 15027
rect 224 15025 244 15027
rect 162 14993 244 15025
rect 524 15025 548 15027
rect 573 15025 582 15027
rect 586 15025 606 15027
rect 160 14985 246 14993
rect 186 14969 220 14985
rect 182 14955 224 14956
rect 160 14949 182 14955
rect 224 14949 246 14955
rect 186 14914 220 14948
rect 223 14914 257 14948
rect 120 14901 170 14903
rect 76 14897 130 14901
rect 110 14892 130 14897
rect 60 14867 67 14877
rect 76 14867 77 14887
rect 96 14858 99 14892
rect 109 14867 110 14887
rect 119 14867 126 14877
rect 76 14851 92 14857
rect 94 14851 110 14857
rect 170 14851 172 14901
rect 186 14835 190 14869
rect 216 14835 220 14869
rect 288 14835 292 15023
rect 476 14955 480 15023
rect 524 14993 606 15025
rect 607 14993 616 15027
rect 522 14985 608 14993
rect 649 14985 651 15035
rect 548 14969 582 14985
rect 522 14950 548 14955
rect 522 14949 582 14950
rect 586 14949 608 14955
rect 295 14914 300 14948
rect 324 14914 329 14948
rect 544 14946 582 14949
rect 378 14909 450 14917
rect 428 14879 430 14895
rect 400 14871 430 14879
rect 476 14877 480 14945
rect 544 14916 552 14946
rect 578 14916 582 14946
rect 544 14907 548 14916
rect 400 14867 436 14871
rect 400 14837 408 14867
rect 420 14837 436 14867
rect 544 14869 548 14877
rect 12 14798 62 14800
rect 28 14789 59 14797
rect 62 14789 64 14798
rect 28 14781 64 14789
rect 127 14789 158 14797
rect 127 14782 182 14789
rect 215 14787 224 14815
rect 127 14781 161 14782
rect 59 14765 64 14781
rect 158 14765 161 14781
rect 28 14757 64 14765
rect 127 14764 161 14765
rect 127 14757 182 14764
rect 62 14748 64 14757
rect 213 14749 224 14787
rect 282 14777 292 14835
rect 296 14829 368 14837
rect 319 14799 346 14810
rect 318 14786 324 14799
rect 346 14786 348 14799
rect 428 14790 430 14837
rect 443 14827 450 14829
rect 476 14797 480 14865
rect 544 14835 552 14869
rect 578 14835 582 14869
rect 481 14803 517 14831
rect 481 14797 495 14803
rect 367 14786 380 14790
rect 251 14743 263 14777
rect 273 14743 293 14777
rect 295 14762 324 14786
rect 303 14752 316 14762
rect 318 14746 324 14762
rect 333 14762 380 14786
rect 333 14752 353 14762
rect 367 14756 380 14762
rect 396 14756 408 14790
rect 420 14756 436 14790
rect 120 14695 170 14697
rect 76 14689 92 14695
rect 94 14689 110 14695
rect 76 14679 99 14688
rect 60 14669 67 14679
rect 76 14659 77 14679
rect 96 14654 99 14679
rect 109 14659 110 14679
rect 119 14669 126 14679
rect 76 14645 110 14649
rect 170 14645 172 14695
rect 186 14677 190 14711
rect 216 14677 220 14711
rect 186 14600 220 14634
rect 282 14631 292 14743
rect 318 14736 335 14746
rect 318 14667 324 14736
rect 346 14667 348 14752
rect 428 14709 430 14756
rect 476 14719 480 14787
rect 485 14769 495 14797
rect 505 14797 519 14803
rect 544 14797 555 14835
rect 505 14769 525 14797
rect 544 14769 553 14797
rect 544 14749 548 14769
rect 579 14728 582 14818
rect 612 14800 624 14801
rect 599 14798 649 14800
rect 612 14797 624 14798
rect 610 14790 632 14797
rect 607 14789 632 14790
rect 586 14782 644 14789
rect 607 14781 644 14782
rect 607 14765 610 14781
rect 616 14765 644 14781
rect 607 14764 644 14765
rect 586 14757 644 14764
rect 607 14756 610 14757
rect 612 14749 632 14757
rect 612 14745 624 14749
rect 649 14748 651 14798
rect 544 14711 548 14719
rect 400 14679 408 14709
rect 420 14679 436 14709
rect 400 14675 436 14679
rect 400 14667 430 14675
rect 428 14651 430 14667
rect 476 14639 480 14707
rect 544 14677 552 14711
rect 578 14677 582 14711
rect 544 14669 548 14677
rect 544 14639 586 14640
rect 288 14599 292 14631
rect 296 14629 368 14637
rect 378 14629 450 14637
rect 544 14632 548 14639
rect 439 14601 444 14629
rect 120 14585 170 14587
rect 76 14581 130 14585
rect 110 14576 130 14581
rect 60 14551 67 14561
rect 76 14551 77 14571
rect 96 14542 99 14576
rect 109 14551 110 14571
rect 119 14551 126 14561
rect 76 14535 92 14541
rect 94 14535 110 14541
rect 170 14535 172 14585
rect 186 14519 190 14553
rect 216 14519 220 14553
rect 213 14487 224 14519
rect 282 14515 292 14599
rect 296 14593 368 14601
rect 378 14593 450 14601
rect 468 14598 473 14632
rect 428 14563 430 14579
rect 251 14487 292 14515
rect 318 14494 324 14563
rect 12 14482 62 14484
rect 28 14473 59 14481
rect 62 14473 64 14482
rect 251 14481 263 14487
rect 28 14465 64 14473
rect 127 14473 158 14481
rect 127 14466 182 14473
rect 127 14465 161 14466
rect 59 14449 64 14465
rect 158 14449 161 14465
rect 253 14453 263 14481
rect 273 14453 293 14487
rect 318 14484 335 14494
rect 303 14468 316 14478
rect 318 14468 324 14484
rect 346 14478 348 14563
rect 400 14555 430 14563
rect 476 14561 480 14629
rect 511 14598 582 14632
rect 544 14591 548 14598
rect 400 14551 436 14555
rect 400 14521 408 14551
rect 420 14521 436 14551
rect 544 14553 548 14561
rect 28 14441 64 14449
rect 127 14448 161 14449
rect 127 14441 182 14448
rect 62 14432 64 14441
rect 282 14395 292 14453
rect 295 14444 324 14468
rect 333 14468 353 14478
rect 428 14474 430 14521
rect 476 14481 480 14549
rect 544 14519 552 14553
rect 578 14519 582 14553
rect 544 14511 548 14519
rect 367 14468 380 14474
rect 333 14444 380 14468
rect 318 14431 324 14444
rect 346 14431 348 14444
rect 367 14440 380 14444
rect 396 14440 408 14474
rect 420 14440 436 14474
rect 544 14471 553 14499
rect 319 14420 346 14431
rect 120 14379 170 14381
rect 76 14373 92 14379
rect 94 14373 110 14379
rect 76 14363 99 14372
rect 60 14353 67 14363
rect 76 14343 77 14363
rect 96 14338 99 14363
rect 109 14343 110 14363
rect 119 14353 126 14363
rect 76 14329 110 14333
rect 170 14329 172 14379
rect 186 14361 190 14395
rect 216 14361 220 14395
rect 182 14323 224 14324
rect 186 14299 220 14316
rect 223 14299 257 14316
rect 182 14282 257 14299
rect 182 14281 224 14282
rect 160 14275 246 14281
rect 288 14275 292 14395
rect 296 14393 368 14401
rect 428 14393 430 14440
rect 476 14403 480 14471
rect 485 14427 495 14461
rect 505 14433 525 14461
rect 505 14427 519 14433
rect 544 14427 555 14471
rect 485 14403 492 14427
rect 579 14412 582 14502
rect 612 14484 624 14485
rect 599 14482 649 14484
rect 612 14481 624 14482
rect 610 14474 632 14481
rect 607 14473 632 14474
rect 586 14466 644 14473
rect 607 14465 644 14466
rect 607 14449 610 14465
rect 616 14449 644 14465
rect 607 14448 644 14449
rect 586 14441 644 14448
rect 607 14440 610 14441
rect 612 14433 632 14441
rect 612 14429 624 14433
rect 649 14432 651 14482
rect 544 14395 548 14403
rect 400 14363 408 14393
rect 420 14363 436 14393
rect 400 14359 436 14363
rect 400 14351 430 14359
rect 428 14335 430 14351
rect 476 14323 480 14391
rect 544 14361 552 14395
rect 578 14361 582 14395
rect 544 14353 548 14361
rect 295 14282 300 14316
rect 324 14282 329 14316
rect 378 14313 450 14321
rect 544 14318 548 14323
rect 544 14314 582 14318
rect 544 14299 552 14314
rect 578 14299 582 14314
rect 544 14281 586 14299
rect 522 14275 608 14281
rect 182 14259 224 14275
rect 544 14259 586 14275
rect 17 14245 67 14247
rect 119 14245 169 14247
rect 186 14245 220 14259
rect 548 14245 582 14259
rect 599 14245 649 14247
rect 42 14203 59 14237
rect 67 14195 69 14245
rect 160 14237 246 14245
rect 522 14237 608 14245
rect 76 14203 110 14237
rect 127 14203 144 14237
rect 152 14203 161 14237
rect 162 14235 195 14237
rect 224 14235 244 14237
rect 162 14203 244 14235
rect 524 14235 548 14237
rect 573 14235 582 14237
rect 586 14235 606 14237
rect 160 14195 246 14203
rect 186 14179 220 14195
rect 182 14165 224 14166
rect 160 14159 182 14165
rect 224 14159 246 14165
rect 186 14124 220 14158
rect 223 14124 257 14158
rect 120 14111 170 14113
rect 76 14107 130 14111
rect 110 14102 130 14107
rect 60 14077 67 14087
rect 76 14077 77 14097
rect 96 14068 99 14102
rect 109 14077 110 14097
rect 119 14077 126 14087
rect 76 14061 92 14067
rect 94 14061 110 14067
rect 170 14061 172 14111
rect 186 14045 190 14079
rect 216 14045 220 14079
rect 288 14045 292 14233
rect 476 14165 480 14233
rect 524 14203 606 14235
rect 607 14203 616 14237
rect 522 14195 608 14203
rect 649 14195 651 14245
rect 548 14179 582 14195
rect 522 14160 548 14165
rect 522 14159 582 14160
rect 586 14159 608 14165
rect 295 14124 300 14158
rect 324 14124 329 14158
rect 544 14156 582 14159
rect 378 14119 450 14127
rect 428 14089 430 14105
rect 400 14081 430 14089
rect 476 14087 480 14155
rect 544 14126 552 14156
rect 578 14126 582 14156
rect 544 14117 548 14126
rect 400 14077 436 14081
rect 400 14047 408 14077
rect 420 14047 436 14077
rect 544 14079 548 14087
rect 12 14008 62 14010
rect 28 13999 59 14007
rect 62 13999 64 14008
rect 28 13991 64 13999
rect 127 13999 158 14007
rect 127 13992 182 13999
rect 215 13997 224 14025
rect 127 13991 161 13992
rect 59 13975 64 13991
rect 158 13975 161 13991
rect 28 13967 64 13975
rect 127 13974 161 13975
rect 127 13967 182 13974
rect 62 13958 64 13967
rect 213 13959 224 13997
rect 282 13987 292 14045
rect 296 14039 368 14047
rect 319 14009 346 14020
rect 318 13996 324 14009
rect 346 13996 348 14009
rect 428 14000 430 14047
rect 443 14037 450 14039
rect 476 14007 480 14075
rect 544 14045 552 14079
rect 578 14045 582 14079
rect 481 14013 517 14041
rect 481 14007 495 14013
rect 367 13996 380 14000
rect 251 13953 263 13987
rect 273 13953 293 13987
rect 295 13972 324 13996
rect 303 13962 316 13972
rect 318 13956 324 13972
rect 333 13972 380 13996
rect 333 13962 353 13972
rect 367 13966 380 13972
rect 396 13966 408 14000
rect 420 13966 436 14000
rect 120 13905 170 13907
rect 76 13899 92 13905
rect 94 13899 110 13905
rect 76 13889 99 13898
rect 60 13879 67 13889
rect 76 13869 77 13889
rect 96 13864 99 13889
rect 109 13869 110 13889
rect 119 13879 126 13889
rect 76 13855 110 13859
rect 170 13855 172 13905
rect 186 13887 190 13921
rect 216 13887 220 13921
rect 186 13810 220 13844
rect 282 13841 292 13953
rect 318 13946 335 13956
rect 318 13877 324 13946
rect 346 13877 348 13962
rect 428 13919 430 13966
rect 476 13929 480 13997
rect 485 13979 495 14007
rect 505 14007 519 14013
rect 544 14007 555 14045
rect 505 13979 525 14007
rect 544 13979 553 14007
rect 544 13959 548 13979
rect 579 13938 582 14028
rect 612 14010 624 14011
rect 599 14008 649 14010
rect 612 14007 624 14008
rect 610 14000 632 14007
rect 607 13999 632 14000
rect 586 13992 644 13999
rect 607 13991 644 13992
rect 607 13975 610 13991
rect 616 13975 644 13991
rect 607 13974 644 13975
rect 586 13967 644 13974
rect 607 13966 610 13967
rect 612 13959 632 13967
rect 612 13955 624 13959
rect 649 13958 651 14008
rect 544 13921 548 13929
rect 400 13889 408 13919
rect 420 13889 436 13919
rect 400 13885 436 13889
rect 400 13877 430 13885
rect 428 13861 430 13877
rect 476 13849 480 13917
rect 544 13887 552 13921
rect 578 13887 582 13921
rect 544 13879 548 13887
rect 544 13849 586 13850
rect 288 13809 292 13841
rect 296 13839 368 13847
rect 378 13839 450 13847
rect 544 13842 548 13849
rect 439 13811 444 13839
rect 120 13795 170 13797
rect 76 13791 130 13795
rect 110 13786 130 13791
rect 60 13761 67 13771
rect 76 13761 77 13781
rect 96 13752 99 13786
rect 109 13761 110 13781
rect 119 13761 126 13771
rect 76 13745 92 13751
rect 94 13745 110 13751
rect 170 13745 172 13795
rect 186 13729 190 13763
rect 216 13729 220 13763
rect 213 13697 224 13729
rect 282 13725 292 13809
rect 296 13803 368 13811
rect 378 13803 450 13811
rect 468 13808 473 13842
rect 428 13773 430 13789
rect 251 13697 292 13725
rect 318 13704 324 13773
rect 12 13692 62 13694
rect 28 13683 59 13691
rect 62 13683 64 13692
rect 251 13691 263 13697
rect 28 13675 64 13683
rect 127 13683 158 13691
rect 127 13676 182 13683
rect 127 13675 161 13676
rect 59 13659 64 13675
rect 158 13659 161 13675
rect 253 13663 263 13691
rect 273 13663 293 13697
rect 318 13694 335 13704
rect 303 13678 316 13688
rect 318 13678 324 13694
rect 346 13688 348 13773
rect 400 13765 430 13773
rect 476 13771 480 13839
rect 511 13808 582 13842
rect 544 13801 548 13808
rect 400 13761 436 13765
rect 400 13731 408 13761
rect 420 13731 436 13761
rect 544 13763 548 13771
rect 28 13651 64 13659
rect 127 13658 161 13659
rect 127 13651 182 13658
rect 62 13642 64 13651
rect 282 13605 292 13663
rect 295 13654 324 13678
rect 333 13678 353 13688
rect 428 13684 430 13731
rect 476 13691 480 13759
rect 544 13729 552 13763
rect 578 13729 582 13763
rect 544 13721 548 13729
rect 367 13678 380 13684
rect 333 13654 380 13678
rect 318 13641 324 13654
rect 346 13641 348 13654
rect 367 13650 380 13654
rect 396 13650 408 13684
rect 420 13650 436 13684
rect 544 13681 553 13709
rect 319 13630 346 13641
rect 120 13589 170 13591
rect 76 13583 92 13589
rect 94 13583 110 13589
rect 76 13573 99 13582
rect 60 13563 67 13573
rect 76 13553 77 13573
rect 96 13548 99 13573
rect 109 13553 110 13573
rect 119 13563 126 13573
rect 76 13539 110 13543
rect 170 13539 172 13589
rect 186 13571 190 13605
rect 216 13571 220 13605
rect 182 13533 224 13534
rect 186 13509 220 13526
rect 223 13509 257 13526
rect 182 13492 257 13509
rect 182 13491 224 13492
rect 160 13485 246 13491
rect 288 13485 292 13605
rect 296 13603 368 13611
rect 428 13603 430 13650
rect 476 13613 480 13681
rect 485 13637 495 13671
rect 505 13643 525 13671
rect 505 13637 519 13643
rect 544 13637 555 13681
rect 485 13613 492 13637
rect 579 13622 582 13712
rect 612 13694 624 13695
rect 599 13692 649 13694
rect 612 13691 624 13692
rect 610 13684 632 13691
rect 607 13683 632 13684
rect 586 13676 644 13683
rect 607 13675 644 13676
rect 607 13659 610 13675
rect 616 13659 644 13675
rect 607 13658 644 13659
rect 586 13651 644 13658
rect 607 13650 610 13651
rect 612 13643 632 13651
rect 612 13639 624 13643
rect 649 13642 651 13692
rect 544 13605 548 13613
rect 400 13573 408 13603
rect 420 13573 436 13603
rect 400 13569 436 13573
rect 400 13561 430 13569
rect 428 13545 430 13561
rect 476 13533 480 13601
rect 544 13571 552 13605
rect 578 13571 582 13605
rect 544 13563 548 13571
rect 295 13492 300 13526
rect 324 13492 329 13526
rect 378 13523 450 13531
rect 544 13528 548 13533
rect 544 13524 582 13528
rect 544 13509 552 13524
rect 578 13509 582 13524
rect 544 13491 586 13509
rect 522 13485 608 13491
rect 182 13469 224 13485
rect 544 13469 586 13485
rect 17 13455 67 13457
rect 119 13455 169 13457
rect 186 13455 220 13469
rect 548 13455 582 13469
rect 599 13455 649 13457
rect 42 13413 59 13447
rect 67 13405 69 13455
rect 160 13447 246 13455
rect 522 13447 608 13455
rect 76 13413 110 13447
rect 127 13413 144 13447
rect 152 13413 161 13447
rect 162 13445 195 13447
rect 224 13445 244 13447
rect 162 13413 244 13445
rect 524 13445 548 13447
rect 573 13445 582 13447
rect 586 13445 606 13447
rect 160 13405 246 13413
rect 186 13389 220 13405
rect 182 13375 224 13376
rect 160 13369 182 13375
rect 224 13369 246 13375
rect 186 13334 220 13368
rect 223 13334 257 13368
rect 120 13321 170 13323
rect 76 13317 130 13321
rect 110 13312 130 13317
rect 60 13287 67 13297
rect 76 13287 77 13307
rect 96 13278 99 13312
rect 109 13287 110 13307
rect 119 13287 126 13297
rect 76 13271 92 13277
rect 94 13271 110 13277
rect 170 13271 172 13321
rect 186 13255 190 13289
rect 216 13255 220 13289
rect 288 13255 292 13443
rect 476 13375 480 13443
rect 524 13413 606 13445
rect 607 13413 616 13447
rect 522 13405 608 13413
rect 649 13405 651 13455
rect 548 13389 582 13405
rect 522 13370 548 13375
rect 522 13369 582 13370
rect 586 13369 608 13375
rect 295 13334 300 13368
rect 324 13334 329 13368
rect 544 13366 582 13369
rect 378 13329 450 13337
rect 428 13299 430 13315
rect 400 13291 430 13299
rect 476 13297 480 13365
rect 544 13336 552 13366
rect 578 13336 582 13366
rect 544 13327 548 13336
rect 400 13287 436 13291
rect 400 13257 408 13287
rect 420 13257 436 13287
rect 544 13289 548 13297
rect 12 13218 62 13220
rect 28 13209 59 13217
rect 62 13209 64 13218
rect 28 13201 64 13209
rect 127 13209 158 13217
rect 127 13202 182 13209
rect 215 13207 224 13235
rect 127 13201 161 13202
rect 59 13185 64 13201
rect 158 13185 161 13201
rect 28 13177 64 13185
rect 127 13184 161 13185
rect 127 13177 182 13184
rect 62 13168 64 13177
rect 213 13169 224 13207
rect 282 13197 292 13255
rect 296 13249 368 13257
rect 319 13219 346 13230
rect 318 13206 324 13219
rect 346 13206 348 13219
rect 428 13210 430 13257
rect 443 13247 450 13249
rect 476 13217 480 13285
rect 544 13255 552 13289
rect 578 13255 582 13289
rect 481 13223 517 13251
rect 481 13217 495 13223
rect 367 13206 380 13210
rect 251 13163 263 13197
rect 273 13163 293 13197
rect 295 13182 324 13206
rect 303 13172 316 13182
rect 318 13166 324 13182
rect 333 13182 380 13206
rect 333 13172 353 13182
rect 367 13176 380 13182
rect 396 13176 408 13210
rect 420 13176 436 13210
rect 120 13115 170 13117
rect 76 13109 92 13115
rect 94 13109 110 13115
rect 76 13099 99 13108
rect 60 13089 67 13099
rect 76 13079 77 13099
rect 96 13074 99 13099
rect 109 13079 110 13099
rect 119 13089 126 13099
rect 76 13065 110 13069
rect 170 13065 172 13115
rect 186 13097 190 13131
rect 216 13097 220 13131
rect 186 13020 220 13054
rect 282 13051 292 13163
rect 318 13156 335 13166
rect 318 13087 324 13156
rect 346 13087 348 13172
rect 428 13129 430 13176
rect 476 13139 480 13207
rect 485 13189 495 13217
rect 505 13217 519 13223
rect 544 13217 555 13255
rect 505 13189 525 13217
rect 544 13189 553 13217
rect 544 13169 548 13189
rect 579 13148 582 13238
rect 612 13220 624 13221
rect 599 13218 649 13220
rect 612 13217 624 13218
rect 610 13210 632 13217
rect 607 13209 632 13210
rect 586 13202 644 13209
rect 607 13201 644 13202
rect 607 13185 610 13201
rect 616 13185 644 13201
rect 607 13184 644 13185
rect 586 13177 644 13184
rect 607 13176 610 13177
rect 612 13169 632 13177
rect 612 13165 624 13169
rect 649 13168 651 13218
rect 544 13131 548 13139
rect 400 13099 408 13129
rect 420 13099 436 13129
rect 400 13095 436 13099
rect 400 13087 430 13095
rect 428 13071 430 13087
rect 476 13059 480 13127
rect 544 13097 552 13131
rect 578 13097 582 13131
rect 544 13089 548 13097
rect 544 13059 586 13060
rect 288 13019 292 13051
rect 296 13049 368 13057
rect 378 13049 450 13057
rect 544 13052 548 13059
rect 439 13021 444 13049
rect 120 13005 170 13007
rect 76 13001 130 13005
rect 110 12996 130 13001
rect 60 12971 67 12981
rect 76 12971 77 12991
rect 96 12962 99 12996
rect 109 12971 110 12991
rect 119 12971 126 12981
rect 76 12955 92 12961
rect 94 12955 110 12961
rect 170 12955 172 13005
rect 186 12939 190 12973
rect 216 12939 220 12973
rect 213 12907 224 12939
rect 282 12935 292 13019
rect 296 13013 368 13021
rect 378 13013 450 13021
rect 468 13018 473 13052
rect 428 12983 430 12999
rect 251 12907 292 12935
rect 318 12914 324 12983
rect 12 12902 62 12904
rect 28 12893 59 12901
rect 62 12893 64 12902
rect 251 12901 263 12907
rect 28 12885 64 12893
rect 127 12893 158 12901
rect 127 12886 182 12893
rect 127 12885 161 12886
rect 59 12869 64 12885
rect 158 12869 161 12885
rect 253 12873 263 12901
rect 273 12873 293 12907
rect 318 12904 335 12914
rect 303 12888 316 12898
rect 318 12888 324 12904
rect 346 12898 348 12983
rect 400 12975 430 12983
rect 476 12981 480 13049
rect 511 13018 582 13052
rect 544 13011 548 13018
rect 400 12971 436 12975
rect 400 12941 408 12971
rect 420 12941 436 12971
rect 544 12973 548 12981
rect 28 12861 64 12869
rect 127 12868 161 12869
rect 127 12861 182 12868
rect 62 12852 64 12861
rect 282 12815 292 12873
rect 295 12864 324 12888
rect 333 12888 353 12898
rect 428 12894 430 12941
rect 476 12901 480 12969
rect 544 12939 552 12973
rect 578 12939 582 12973
rect 544 12931 548 12939
rect 367 12888 380 12894
rect 333 12864 380 12888
rect 318 12851 324 12864
rect 346 12851 348 12864
rect 367 12860 380 12864
rect 396 12860 408 12894
rect 420 12860 436 12894
rect 544 12891 553 12919
rect 319 12840 346 12851
rect 120 12799 170 12801
rect 76 12793 92 12799
rect 94 12793 110 12799
rect 76 12783 99 12792
rect 60 12773 67 12783
rect 76 12763 77 12783
rect 96 12758 99 12783
rect 109 12763 110 12783
rect 119 12773 126 12783
rect 76 12749 110 12753
rect 170 12749 172 12799
rect 186 12781 190 12815
rect 216 12781 220 12815
rect 182 12743 224 12744
rect 186 12719 220 12736
rect 223 12719 257 12736
rect 182 12702 257 12719
rect 182 12701 224 12702
rect 160 12695 246 12701
rect 288 12695 292 12815
rect 296 12813 368 12821
rect 428 12813 430 12860
rect 476 12823 480 12891
rect 485 12847 495 12881
rect 505 12853 525 12881
rect 505 12847 519 12853
rect 544 12847 555 12891
rect 485 12823 492 12847
rect 579 12832 582 12922
rect 612 12904 624 12905
rect 599 12902 649 12904
rect 612 12901 624 12902
rect 610 12894 632 12901
rect 607 12893 632 12894
rect 586 12886 644 12893
rect 607 12885 644 12886
rect 607 12869 610 12885
rect 616 12869 644 12885
rect 607 12868 644 12869
rect 586 12861 644 12868
rect 607 12860 610 12861
rect 612 12853 632 12861
rect 612 12849 624 12853
rect 649 12852 651 12902
rect 544 12815 548 12823
rect 400 12783 408 12813
rect 420 12783 436 12813
rect 400 12779 436 12783
rect 400 12771 430 12779
rect 428 12755 430 12771
rect 476 12743 480 12811
rect 544 12781 552 12815
rect 578 12781 582 12815
rect 544 12773 548 12781
rect 295 12702 300 12736
rect 324 12702 329 12736
rect 378 12733 450 12741
rect 544 12738 548 12743
rect 544 12734 582 12738
rect 544 12719 552 12734
rect 578 12719 582 12734
rect 544 12701 586 12719
rect 522 12695 608 12701
rect 182 12679 224 12695
rect 544 12679 586 12695
rect 17 12665 67 12667
rect 119 12665 169 12667
rect 186 12665 220 12679
rect 548 12665 582 12679
rect 599 12665 649 12667
rect 42 12623 59 12657
rect 67 12615 69 12665
rect 160 12657 246 12665
rect 522 12657 608 12665
rect 76 12623 110 12657
rect 127 12623 144 12657
rect 152 12623 161 12657
rect 162 12655 195 12657
rect 224 12655 244 12657
rect 162 12623 244 12655
rect 524 12655 548 12657
rect 573 12655 582 12657
rect 586 12655 606 12657
rect 160 12615 246 12623
rect 186 12599 220 12615
rect 182 12585 224 12586
rect 160 12579 182 12585
rect 224 12579 246 12585
rect 186 12544 220 12578
rect 223 12544 257 12578
rect 120 12531 170 12533
rect 76 12527 130 12531
rect 110 12522 130 12527
rect 60 12497 67 12507
rect 76 12497 77 12517
rect 96 12488 99 12522
rect 109 12497 110 12517
rect 119 12497 126 12507
rect 76 12481 92 12487
rect 94 12481 110 12487
rect 170 12481 172 12531
rect 186 12465 190 12499
rect 216 12465 220 12499
rect 288 12465 292 12653
rect 476 12585 480 12653
rect 524 12623 606 12655
rect 607 12623 616 12657
rect 522 12615 608 12623
rect 649 12615 651 12665
rect 548 12599 582 12615
rect 522 12580 548 12585
rect 522 12579 582 12580
rect 586 12579 608 12585
rect 295 12544 300 12578
rect 324 12544 329 12578
rect 544 12576 582 12579
rect 378 12539 450 12547
rect 428 12509 430 12525
rect 400 12501 430 12509
rect 476 12507 480 12575
rect 544 12546 552 12576
rect 578 12546 582 12576
rect 544 12537 548 12546
rect 400 12497 436 12501
rect 400 12467 408 12497
rect 420 12467 436 12497
rect 544 12499 548 12507
rect 12 12428 62 12430
rect 28 12419 59 12427
rect 62 12419 64 12428
rect 28 12411 64 12419
rect 127 12419 158 12427
rect 127 12412 182 12419
rect 215 12417 224 12445
rect 127 12411 161 12412
rect 59 12395 64 12411
rect 158 12395 161 12411
rect 28 12387 64 12395
rect 127 12394 161 12395
rect 127 12387 182 12394
rect 62 12378 64 12387
rect 213 12379 224 12417
rect 282 12407 292 12465
rect 296 12459 368 12467
rect 319 12429 346 12440
rect 318 12416 324 12429
rect 346 12416 348 12429
rect 428 12420 430 12467
rect 443 12457 450 12459
rect 476 12427 480 12495
rect 544 12465 552 12499
rect 578 12465 582 12499
rect 481 12433 517 12461
rect 481 12427 495 12433
rect 367 12416 380 12420
rect 251 12373 263 12407
rect 273 12373 293 12407
rect 295 12392 324 12416
rect 303 12382 316 12392
rect 318 12376 324 12392
rect 333 12392 380 12416
rect 333 12382 353 12392
rect 367 12386 380 12392
rect 396 12386 408 12420
rect 420 12386 436 12420
rect 120 12325 170 12327
rect 76 12319 92 12325
rect 94 12319 110 12325
rect 76 12309 99 12318
rect 60 12299 67 12309
rect 76 12289 77 12309
rect 96 12284 99 12309
rect 109 12289 110 12309
rect 119 12299 126 12309
rect 76 12275 110 12279
rect 170 12275 172 12325
rect 186 12307 190 12341
rect 216 12307 220 12341
rect 186 12230 220 12264
rect 282 12261 292 12373
rect 318 12366 335 12376
rect 318 12297 324 12366
rect 346 12297 348 12382
rect 428 12339 430 12386
rect 476 12349 480 12417
rect 485 12399 495 12427
rect 505 12427 519 12433
rect 544 12427 555 12465
rect 505 12399 525 12427
rect 544 12399 553 12427
rect 544 12379 548 12399
rect 579 12358 582 12448
rect 612 12430 624 12431
rect 599 12428 649 12430
rect 612 12427 624 12428
rect 610 12420 632 12427
rect 607 12419 632 12420
rect 586 12412 644 12419
rect 607 12411 644 12412
rect 607 12395 610 12411
rect 616 12395 644 12411
rect 607 12394 644 12395
rect 586 12387 644 12394
rect 607 12386 610 12387
rect 612 12379 632 12387
rect 612 12375 624 12379
rect 649 12378 651 12428
rect 544 12341 548 12349
rect 400 12309 408 12339
rect 420 12309 436 12339
rect 400 12305 436 12309
rect 400 12297 430 12305
rect 428 12281 430 12297
rect 476 12269 480 12337
rect 544 12307 552 12341
rect 578 12307 582 12341
rect 544 12299 548 12307
rect 544 12269 586 12270
rect 288 12229 292 12261
rect 296 12259 368 12267
rect 378 12259 450 12267
rect 544 12262 548 12269
rect 439 12231 444 12259
rect 120 12215 170 12217
rect 76 12211 130 12215
rect 110 12206 130 12211
rect 60 12181 67 12191
rect 76 12181 77 12201
rect 96 12172 99 12206
rect 109 12181 110 12201
rect 119 12181 126 12191
rect 76 12165 92 12171
rect 94 12165 110 12171
rect 170 12165 172 12215
rect 186 12149 190 12183
rect 216 12149 220 12183
rect 213 12117 224 12149
rect 282 12145 292 12229
rect 296 12223 368 12231
rect 378 12223 450 12231
rect 468 12228 473 12262
rect 428 12193 430 12209
rect 251 12117 292 12145
rect 318 12124 324 12193
rect 12 12112 62 12114
rect 28 12103 59 12111
rect 62 12103 64 12112
rect 251 12111 263 12117
rect 28 12095 64 12103
rect 127 12103 158 12111
rect 127 12096 182 12103
rect 127 12095 161 12096
rect 59 12079 64 12095
rect 158 12079 161 12095
rect 253 12083 263 12111
rect 273 12083 293 12117
rect 318 12114 335 12124
rect 303 12098 316 12108
rect 318 12098 324 12114
rect 346 12108 348 12193
rect 400 12185 430 12193
rect 476 12191 480 12259
rect 511 12228 582 12262
rect 544 12221 548 12228
rect 400 12181 436 12185
rect 400 12151 408 12181
rect 420 12151 436 12181
rect 544 12183 548 12191
rect 28 12071 64 12079
rect 127 12078 161 12079
rect 127 12071 182 12078
rect 62 12062 64 12071
rect 282 12025 292 12083
rect 295 12074 324 12098
rect 333 12098 353 12108
rect 428 12104 430 12151
rect 476 12111 480 12179
rect 544 12149 552 12183
rect 578 12149 582 12183
rect 544 12141 548 12149
rect 367 12098 380 12104
rect 333 12074 380 12098
rect 318 12061 324 12074
rect 346 12061 348 12074
rect 367 12070 380 12074
rect 396 12070 408 12104
rect 420 12070 436 12104
rect 544 12101 553 12129
rect 319 12050 346 12061
rect 120 12009 170 12011
rect 76 12003 92 12009
rect 94 12003 110 12009
rect 76 11993 99 12002
rect 60 11983 67 11993
rect 76 11973 77 11993
rect 96 11968 99 11993
rect 109 11973 110 11993
rect 119 11983 126 11993
rect 76 11959 110 11963
rect 170 11959 172 12009
rect 186 11991 190 12025
rect 216 11991 220 12025
rect 182 11953 224 11954
rect 186 11929 220 11946
rect 223 11929 257 11946
rect 182 11912 257 11929
rect 182 11911 224 11912
rect 160 11905 246 11911
rect 288 11905 292 12025
rect 296 12023 368 12031
rect 428 12023 430 12070
rect 476 12033 480 12101
rect 485 12057 495 12091
rect 505 12063 525 12091
rect 505 12057 519 12063
rect 544 12057 555 12101
rect 485 12033 492 12057
rect 579 12042 582 12132
rect 612 12114 624 12115
rect 599 12112 649 12114
rect 612 12111 624 12112
rect 610 12104 632 12111
rect 607 12103 632 12104
rect 586 12096 644 12103
rect 607 12095 644 12096
rect 607 12079 610 12095
rect 616 12079 644 12095
rect 607 12078 644 12079
rect 586 12071 644 12078
rect 607 12070 610 12071
rect 612 12063 632 12071
rect 612 12059 624 12063
rect 649 12062 651 12112
rect 544 12025 548 12033
rect 400 11993 408 12023
rect 420 11993 436 12023
rect 400 11989 436 11993
rect 400 11981 430 11989
rect 428 11965 430 11981
rect 476 11953 480 12021
rect 544 11991 552 12025
rect 578 11991 582 12025
rect 544 11983 548 11991
rect 295 11912 300 11946
rect 324 11912 329 11946
rect 378 11943 450 11951
rect 544 11948 548 11953
rect 544 11944 582 11948
rect 544 11929 552 11944
rect 578 11929 582 11944
rect 544 11911 586 11929
rect 522 11905 608 11911
rect 182 11889 224 11905
rect 544 11889 586 11905
rect 17 11875 67 11877
rect 119 11875 169 11877
rect 186 11875 220 11889
rect 548 11875 582 11889
rect 599 11875 649 11877
rect 42 11833 59 11867
rect 67 11825 69 11875
rect 160 11867 246 11875
rect 522 11867 608 11875
rect 76 11833 110 11867
rect 127 11833 144 11867
rect 152 11833 161 11867
rect 162 11865 195 11867
rect 224 11865 244 11867
rect 162 11833 244 11865
rect 524 11865 548 11867
rect 573 11865 582 11867
rect 586 11865 606 11867
rect 160 11825 246 11833
rect 186 11809 220 11825
rect 182 11795 224 11796
rect 160 11789 182 11795
rect 224 11789 246 11795
rect 186 11754 220 11788
rect 223 11754 257 11788
rect 120 11741 170 11743
rect 76 11737 130 11741
rect 110 11732 130 11737
rect 60 11707 67 11717
rect 76 11707 77 11727
rect 96 11698 99 11732
rect 109 11707 110 11727
rect 119 11707 126 11717
rect 76 11691 92 11697
rect 94 11691 110 11697
rect 170 11691 172 11741
rect 186 11675 190 11709
rect 216 11675 220 11709
rect 288 11675 292 11863
rect 476 11795 480 11863
rect 524 11833 606 11865
rect 607 11833 616 11867
rect 522 11825 608 11833
rect 649 11825 651 11875
rect 548 11809 582 11825
rect 522 11790 548 11795
rect 522 11789 582 11790
rect 586 11789 608 11795
rect 295 11754 300 11788
rect 324 11754 329 11788
rect 544 11786 582 11789
rect 378 11749 450 11757
rect 428 11719 430 11735
rect 400 11711 430 11719
rect 476 11717 480 11785
rect 544 11756 552 11786
rect 578 11756 582 11786
rect 544 11747 548 11756
rect 400 11707 436 11711
rect 400 11677 408 11707
rect 420 11677 436 11707
rect 544 11709 548 11717
rect 12 11638 62 11640
rect 28 11629 59 11637
rect 62 11629 64 11638
rect 28 11621 64 11629
rect 127 11629 158 11637
rect 127 11622 182 11629
rect 215 11627 224 11655
rect 127 11621 161 11622
rect 59 11605 64 11621
rect 158 11605 161 11621
rect 28 11597 64 11605
rect 127 11604 161 11605
rect 127 11597 182 11604
rect 62 11588 64 11597
rect 213 11589 224 11627
rect 282 11617 292 11675
rect 296 11669 368 11677
rect 319 11639 346 11650
rect 318 11626 324 11639
rect 346 11626 348 11639
rect 428 11630 430 11677
rect 443 11667 450 11669
rect 476 11637 480 11705
rect 544 11675 552 11709
rect 578 11675 582 11709
rect 481 11643 517 11671
rect 481 11637 495 11643
rect 367 11626 380 11630
rect 251 11583 263 11617
rect 273 11583 293 11617
rect 295 11602 324 11626
rect 303 11592 316 11602
rect 318 11586 324 11602
rect 333 11602 380 11626
rect 333 11592 353 11602
rect 367 11596 380 11602
rect 396 11596 408 11630
rect 420 11596 436 11630
rect 120 11535 170 11537
rect 76 11529 92 11535
rect 94 11529 110 11535
rect 76 11519 99 11528
rect 60 11509 67 11519
rect 76 11499 77 11519
rect 96 11494 99 11519
rect 109 11499 110 11519
rect 119 11509 126 11519
rect 76 11485 110 11489
rect 170 11485 172 11535
rect 186 11517 190 11551
rect 216 11517 220 11551
rect 186 11440 220 11474
rect 282 11471 292 11583
rect 318 11576 335 11586
rect 318 11507 324 11576
rect 346 11507 348 11592
rect 428 11549 430 11596
rect 476 11559 480 11627
rect 485 11609 495 11637
rect 505 11637 519 11643
rect 544 11637 555 11675
rect 505 11609 525 11637
rect 544 11609 553 11637
rect 544 11589 548 11609
rect 579 11568 582 11658
rect 612 11640 624 11641
rect 599 11638 649 11640
rect 612 11637 624 11638
rect 610 11630 632 11637
rect 607 11629 632 11630
rect 586 11622 644 11629
rect 607 11621 644 11622
rect 607 11605 610 11621
rect 616 11605 644 11621
rect 607 11604 644 11605
rect 586 11597 644 11604
rect 607 11596 610 11597
rect 612 11589 632 11597
rect 612 11585 624 11589
rect 649 11588 651 11638
rect 544 11551 548 11559
rect 400 11519 408 11549
rect 420 11519 436 11549
rect 400 11515 436 11519
rect 400 11507 430 11515
rect 428 11491 430 11507
rect 476 11479 480 11547
rect 544 11517 552 11551
rect 578 11517 582 11551
rect 544 11509 548 11517
rect 544 11479 586 11480
rect 288 11439 292 11471
rect 296 11469 368 11477
rect 378 11469 450 11477
rect 544 11472 548 11479
rect 439 11441 444 11469
rect 120 11425 170 11427
rect 76 11421 130 11425
rect 110 11416 130 11421
rect 60 11391 67 11401
rect 76 11391 77 11411
rect 96 11382 99 11416
rect 109 11391 110 11411
rect 119 11391 126 11401
rect 76 11375 92 11381
rect 94 11375 110 11381
rect 170 11375 172 11425
rect 186 11359 190 11393
rect 216 11359 220 11393
rect 213 11327 224 11359
rect 282 11355 292 11439
rect 296 11433 368 11441
rect 378 11433 450 11441
rect 468 11438 473 11472
rect 428 11403 430 11419
rect 251 11327 292 11355
rect 318 11334 324 11403
rect 12 11322 62 11324
rect 28 11313 59 11321
rect 62 11313 64 11322
rect 251 11321 263 11327
rect 28 11305 64 11313
rect 127 11313 158 11321
rect 127 11306 182 11313
rect 127 11305 161 11306
rect 59 11289 64 11305
rect 158 11289 161 11305
rect 253 11293 263 11321
rect 273 11293 293 11327
rect 318 11324 335 11334
rect 303 11308 316 11318
rect 318 11308 324 11324
rect 346 11318 348 11403
rect 400 11395 430 11403
rect 476 11401 480 11469
rect 511 11438 582 11472
rect 544 11431 548 11438
rect 400 11391 436 11395
rect 400 11361 408 11391
rect 420 11361 436 11391
rect 544 11393 548 11401
rect 28 11281 64 11289
rect 127 11288 161 11289
rect 127 11281 182 11288
rect 62 11272 64 11281
rect 282 11235 292 11293
rect 295 11284 324 11308
rect 333 11308 353 11318
rect 428 11314 430 11361
rect 476 11321 480 11389
rect 544 11359 552 11393
rect 578 11359 582 11393
rect 544 11351 548 11359
rect 367 11308 380 11314
rect 333 11284 380 11308
rect 318 11271 324 11284
rect 346 11271 348 11284
rect 367 11280 380 11284
rect 396 11280 408 11314
rect 420 11280 436 11314
rect 544 11311 553 11339
rect 319 11260 346 11271
rect 120 11219 170 11221
rect 76 11213 92 11219
rect 94 11213 110 11219
rect 76 11203 99 11212
rect 60 11193 67 11203
rect 76 11183 77 11203
rect 96 11178 99 11203
rect 109 11183 110 11203
rect 119 11193 126 11203
rect 76 11169 110 11173
rect 170 11169 172 11219
rect 186 11201 190 11235
rect 216 11201 220 11235
rect 182 11163 224 11164
rect 186 11139 220 11156
rect 223 11139 257 11156
rect 182 11122 257 11139
rect 182 11121 224 11122
rect 160 11115 246 11121
rect 288 11115 292 11235
rect 296 11233 368 11241
rect 428 11233 430 11280
rect 476 11243 480 11311
rect 485 11267 495 11301
rect 505 11273 525 11301
rect 505 11267 519 11273
rect 544 11267 555 11311
rect 485 11243 492 11267
rect 579 11252 582 11342
rect 612 11324 624 11325
rect 599 11322 649 11324
rect 612 11321 624 11322
rect 610 11314 632 11321
rect 607 11313 632 11314
rect 586 11306 644 11313
rect 607 11305 644 11306
rect 607 11289 610 11305
rect 616 11289 644 11305
rect 607 11288 644 11289
rect 586 11281 644 11288
rect 607 11280 610 11281
rect 612 11273 632 11281
rect 612 11269 624 11273
rect 649 11272 651 11322
rect 544 11235 548 11243
rect 400 11203 408 11233
rect 420 11203 436 11233
rect 400 11199 436 11203
rect 400 11191 430 11199
rect 428 11175 430 11191
rect 476 11163 480 11231
rect 544 11201 552 11235
rect 578 11201 582 11235
rect 544 11193 548 11201
rect 295 11122 300 11156
rect 324 11122 329 11156
rect 378 11153 450 11161
rect 544 11158 548 11163
rect 544 11154 582 11158
rect 544 11139 552 11154
rect 578 11139 582 11154
rect 544 11121 586 11139
rect 522 11115 608 11121
rect 182 11099 224 11115
rect 544 11099 586 11115
rect 17 11085 67 11087
rect 119 11085 169 11087
rect 186 11085 220 11099
rect 548 11085 582 11099
rect 599 11085 649 11087
rect 42 11043 59 11077
rect 67 11035 69 11085
rect 160 11077 246 11085
rect 522 11077 608 11085
rect 76 11043 110 11077
rect 127 11043 144 11077
rect 152 11043 161 11077
rect 162 11075 195 11077
rect 224 11075 244 11077
rect 162 11043 244 11075
rect 524 11075 548 11077
rect 573 11075 582 11077
rect 586 11075 606 11077
rect 160 11035 246 11043
rect 186 11019 220 11035
rect 182 11005 224 11006
rect 160 10999 182 11005
rect 224 10999 246 11005
rect 186 10964 220 10998
rect 223 10964 257 10998
rect 120 10951 170 10953
rect 76 10947 130 10951
rect 110 10942 130 10947
rect 60 10917 67 10927
rect 76 10917 77 10937
rect 96 10908 99 10942
rect 109 10917 110 10937
rect 119 10917 126 10927
rect 76 10901 92 10907
rect 94 10901 110 10907
rect 170 10901 172 10951
rect 186 10885 190 10919
rect 216 10885 220 10919
rect 288 10885 292 11073
rect 476 11005 480 11073
rect 524 11043 606 11075
rect 607 11043 616 11077
rect 522 11035 608 11043
rect 649 11035 651 11085
rect 548 11019 582 11035
rect 522 11000 548 11005
rect 522 10999 582 11000
rect 586 10999 608 11005
rect 295 10964 300 10998
rect 324 10964 329 10998
rect 544 10996 582 10999
rect 378 10959 450 10967
rect 428 10929 430 10945
rect 400 10921 430 10929
rect 476 10927 480 10995
rect 544 10966 552 10996
rect 578 10966 582 10996
rect 544 10957 548 10966
rect 400 10917 436 10921
rect 400 10887 408 10917
rect 420 10887 436 10917
rect 544 10919 548 10927
rect 12 10848 62 10850
rect 28 10839 59 10847
rect 62 10839 64 10848
rect 28 10831 64 10839
rect 127 10839 158 10847
rect 127 10832 182 10839
rect 215 10837 224 10865
rect 127 10831 161 10832
rect 59 10815 64 10831
rect 158 10815 161 10831
rect 28 10807 64 10815
rect 127 10814 161 10815
rect 127 10807 182 10814
rect 62 10798 64 10807
rect 213 10799 224 10837
rect 282 10827 292 10885
rect 296 10879 368 10887
rect 319 10849 346 10860
rect 318 10836 324 10849
rect 346 10836 348 10849
rect 428 10840 430 10887
rect 443 10877 450 10879
rect 476 10847 480 10915
rect 544 10885 552 10919
rect 578 10885 582 10919
rect 481 10853 517 10881
rect 481 10847 495 10853
rect 367 10836 380 10840
rect 251 10793 263 10827
rect 273 10793 293 10827
rect 295 10812 324 10836
rect 303 10802 316 10812
rect 318 10796 324 10812
rect 333 10812 380 10836
rect 333 10802 353 10812
rect 367 10806 380 10812
rect 396 10806 408 10840
rect 420 10806 436 10840
rect 120 10745 170 10747
rect 76 10739 92 10745
rect 94 10739 110 10745
rect 76 10729 99 10738
rect 60 10719 67 10729
rect 76 10709 77 10729
rect 96 10704 99 10729
rect 109 10709 110 10729
rect 119 10719 126 10729
rect 76 10695 110 10699
rect 170 10695 172 10745
rect 186 10727 190 10761
rect 216 10727 220 10761
rect 186 10650 220 10684
rect 282 10681 292 10793
rect 318 10786 335 10796
rect 318 10717 324 10786
rect 346 10717 348 10802
rect 428 10759 430 10806
rect 476 10769 480 10837
rect 485 10819 495 10847
rect 505 10847 519 10853
rect 544 10847 555 10885
rect 505 10819 525 10847
rect 544 10819 553 10847
rect 544 10799 548 10819
rect 579 10778 582 10868
rect 612 10850 624 10851
rect 599 10848 649 10850
rect 612 10847 624 10848
rect 610 10840 632 10847
rect 607 10839 632 10840
rect 586 10832 644 10839
rect 607 10831 644 10832
rect 607 10815 610 10831
rect 616 10815 644 10831
rect 607 10814 644 10815
rect 586 10807 644 10814
rect 607 10806 610 10807
rect 612 10799 632 10807
rect 612 10795 624 10799
rect 649 10798 651 10848
rect 544 10761 548 10769
rect 400 10729 408 10759
rect 420 10729 436 10759
rect 400 10725 436 10729
rect 400 10717 430 10725
rect 428 10701 430 10717
rect 476 10689 480 10757
rect 544 10727 552 10761
rect 578 10727 582 10761
rect 544 10719 548 10727
rect 544 10689 586 10690
rect 288 10649 292 10681
rect 296 10679 368 10687
rect 378 10679 450 10687
rect 544 10682 548 10689
rect 439 10651 444 10679
rect 120 10635 170 10637
rect 76 10631 130 10635
rect 110 10626 130 10631
rect 60 10601 67 10611
rect 76 10601 77 10621
rect 96 10592 99 10626
rect 109 10601 110 10621
rect 119 10601 126 10611
rect 76 10585 92 10591
rect 94 10585 110 10591
rect 170 10585 172 10635
rect 186 10569 190 10603
rect 216 10569 220 10603
rect 213 10537 224 10569
rect 282 10565 292 10649
rect 296 10643 368 10651
rect 378 10643 450 10651
rect 468 10648 473 10682
rect 428 10613 430 10629
rect 251 10537 292 10565
rect 318 10544 324 10613
rect 12 10532 62 10534
rect 28 10523 59 10531
rect 62 10523 64 10532
rect 251 10531 263 10537
rect 28 10515 64 10523
rect 127 10523 158 10531
rect 127 10516 182 10523
rect 127 10515 161 10516
rect 59 10499 64 10515
rect 158 10499 161 10515
rect 253 10503 263 10531
rect 273 10503 293 10537
rect 318 10534 335 10544
rect 303 10518 316 10528
rect 318 10518 324 10534
rect 346 10528 348 10613
rect 400 10605 430 10613
rect 476 10611 480 10679
rect 511 10648 582 10682
rect 544 10641 548 10648
rect 400 10601 436 10605
rect 400 10571 408 10601
rect 420 10571 436 10601
rect 544 10603 548 10611
rect 28 10491 64 10499
rect 127 10498 161 10499
rect 127 10491 182 10498
rect 62 10482 64 10491
rect 282 10445 292 10503
rect 295 10494 324 10518
rect 333 10518 353 10528
rect 428 10524 430 10571
rect 476 10531 480 10599
rect 544 10569 552 10603
rect 578 10569 582 10603
rect 544 10561 548 10569
rect 367 10518 380 10524
rect 333 10494 380 10518
rect 318 10481 324 10494
rect 346 10481 348 10494
rect 367 10490 380 10494
rect 396 10490 408 10524
rect 420 10490 436 10524
rect 544 10521 553 10549
rect 319 10470 346 10481
rect 120 10429 170 10431
rect 76 10423 92 10429
rect 94 10423 110 10429
rect 76 10413 99 10422
rect 60 10403 67 10413
rect 76 10393 77 10413
rect 96 10388 99 10413
rect 109 10393 110 10413
rect 119 10403 126 10413
rect 76 10379 110 10383
rect 170 10379 172 10429
rect 186 10411 190 10445
rect 216 10411 220 10445
rect 182 10373 224 10374
rect 186 10349 220 10366
rect 223 10349 257 10366
rect 182 10332 257 10349
rect 182 10331 224 10332
rect 160 10325 246 10331
rect 288 10325 292 10445
rect 296 10443 368 10451
rect 428 10443 430 10490
rect 476 10453 480 10521
rect 485 10477 495 10511
rect 505 10483 525 10511
rect 505 10477 519 10483
rect 544 10477 555 10521
rect 485 10453 492 10477
rect 579 10462 582 10552
rect 612 10534 624 10535
rect 599 10532 649 10534
rect 612 10531 624 10532
rect 610 10524 632 10531
rect 607 10523 632 10524
rect 586 10516 644 10523
rect 607 10515 644 10516
rect 607 10499 610 10515
rect 616 10499 644 10515
rect 607 10498 644 10499
rect 586 10491 644 10498
rect 607 10490 610 10491
rect 612 10483 632 10491
rect 612 10479 624 10483
rect 649 10482 651 10532
rect 544 10445 548 10453
rect 400 10413 408 10443
rect 420 10413 436 10443
rect 400 10409 436 10413
rect 400 10401 430 10409
rect 428 10385 430 10401
rect 476 10373 480 10441
rect 544 10411 552 10445
rect 578 10411 582 10445
rect 544 10403 548 10411
rect 295 10332 300 10366
rect 324 10332 329 10366
rect 378 10363 450 10371
rect 544 10368 548 10373
rect 544 10364 582 10368
rect 544 10349 552 10364
rect 578 10349 582 10364
rect 544 10331 586 10349
rect 522 10325 608 10331
rect 182 10309 224 10325
rect 544 10309 586 10325
rect 17 10295 67 10297
rect 119 10295 169 10297
rect 186 10295 220 10309
rect 548 10295 582 10309
rect 599 10295 649 10297
rect 42 10253 59 10287
rect 67 10245 69 10295
rect 160 10287 246 10295
rect 522 10287 608 10295
rect 76 10253 110 10287
rect 127 10253 144 10287
rect 152 10253 161 10287
rect 162 10285 195 10287
rect 224 10285 244 10287
rect 162 10253 244 10285
rect 524 10285 548 10287
rect 573 10285 582 10287
rect 586 10285 606 10287
rect 160 10245 246 10253
rect 186 10229 220 10245
rect 182 10215 224 10216
rect 160 10209 182 10215
rect 224 10209 246 10215
rect 186 10174 220 10208
rect 223 10174 257 10208
rect 120 10161 170 10163
rect 76 10157 130 10161
rect 110 10152 130 10157
rect 60 10127 67 10137
rect 76 10127 77 10147
rect 96 10118 99 10152
rect 109 10127 110 10147
rect 119 10127 126 10137
rect 76 10111 92 10117
rect 94 10111 110 10117
rect 170 10111 172 10161
rect 186 10095 190 10129
rect 216 10095 220 10129
rect 288 10095 292 10283
rect 476 10215 480 10283
rect 524 10253 606 10285
rect 607 10253 616 10287
rect 522 10245 608 10253
rect 649 10245 651 10295
rect 548 10229 582 10245
rect 522 10210 548 10215
rect 522 10209 582 10210
rect 586 10209 608 10215
rect 295 10174 300 10208
rect 324 10174 329 10208
rect 544 10206 582 10209
rect 378 10169 450 10177
rect 428 10139 430 10155
rect 400 10131 430 10139
rect 476 10137 480 10205
rect 544 10176 552 10206
rect 578 10176 582 10206
rect 544 10167 548 10176
rect 400 10127 436 10131
rect 400 10097 408 10127
rect 420 10097 436 10127
rect 544 10129 548 10137
rect 12 10058 62 10060
rect 28 10049 59 10057
rect 62 10049 64 10058
rect 28 10041 64 10049
rect 127 10049 158 10057
rect 127 10042 182 10049
rect 215 10047 224 10075
rect 127 10041 161 10042
rect 59 10025 64 10041
rect 158 10025 161 10041
rect 28 10017 64 10025
rect 127 10024 161 10025
rect 127 10017 182 10024
rect 62 10008 64 10017
rect 213 10009 224 10047
rect 282 10037 292 10095
rect 296 10089 368 10097
rect 319 10059 346 10070
rect 318 10046 324 10059
rect 346 10046 348 10059
rect 428 10050 430 10097
rect 443 10087 450 10089
rect 476 10057 480 10125
rect 544 10095 552 10129
rect 578 10095 582 10129
rect 481 10063 517 10091
rect 481 10057 495 10063
rect 367 10046 380 10050
rect 251 10003 263 10037
rect 273 10003 293 10037
rect 295 10022 324 10046
rect 303 10012 316 10022
rect 318 10006 324 10022
rect 333 10022 380 10046
rect 333 10012 353 10022
rect 367 10016 380 10022
rect 396 10016 408 10050
rect 420 10016 436 10050
rect 120 9955 170 9957
rect 76 9949 92 9955
rect 94 9949 110 9955
rect 76 9939 99 9948
rect 60 9929 67 9939
rect 76 9919 77 9939
rect 96 9914 99 9939
rect 109 9919 110 9939
rect 119 9929 126 9939
rect 76 9905 110 9909
rect 170 9905 172 9955
rect 186 9937 190 9971
rect 216 9937 220 9971
rect 186 9860 220 9894
rect 282 9891 292 10003
rect 318 9996 335 10006
rect 318 9927 324 9996
rect 346 9927 348 10012
rect 428 9969 430 10016
rect 476 9979 480 10047
rect 485 10029 495 10057
rect 505 10057 519 10063
rect 544 10057 555 10095
rect 505 10029 525 10057
rect 544 10029 553 10057
rect 544 10009 548 10029
rect 579 9988 582 10078
rect 612 10060 624 10061
rect 599 10058 649 10060
rect 612 10057 624 10058
rect 610 10050 632 10057
rect 607 10049 632 10050
rect 586 10042 644 10049
rect 607 10041 644 10042
rect 607 10025 610 10041
rect 616 10025 644 10041
rect 607 10024 644 10025
rect 586 10017 644 10024
rect 607 10016 610 10017
rect 612 10009 632 10017
rect 612 10005 624 10009
rect 649 10008 651 10058
rect 544 9971 548 9979
rect 400 9939 408 9969
rect 420 9939 436 9969
rect 400 9935 436 9939
rect 400 9927 430 9935
rect 428 9911 430 9927
rect 476 9899 480 9967
rect 544 9937 552 9971
rect 578 9937 582 9971
rect 544 9929 548 9937
rect 544 9899 586 9900
rect 288 9859 292 9891
rect 296 9889 368 9897
rect 378 9889 450 9897
rect 544 9892 548 9899
rect 439 9861 444 9889
rect 120 9845 170 9847
rect 76 9841 130 9845
rect 110 9836 130 9841
rect 60 9811 67 9821
rect 76 9811 77 9831
rect 96 9802 99 9836
rect 109 9811 110 9831
rect 119 9811 126 9821
rect 76 9795 92 9801
rect 94 9795 110 9801
rect 170 9795 172 9845
rect 186 9779 190 9813
rect 216 9779 220 9813
rect 213 9747 224 9779
rect 282 9775 292 9859
rect 296 9853 368 9861
rect 378 9853 450 9861
rect 468 9858 473 9892
rect 428 9823 430 9839
rect 251 9747 292 9775
rect 318 9754 324 9823
rect 12 9742 62 9744
rect 28 9733 59 9741
rect 62 9733 64 9742
rect 251 9741 263 9747
rect 28 9725 64 9733
rect 127 9733 158 9741
rect 127 9726 182 9733
rect 127 9725 161 9726
rect 59 9709 64 9725
rect 158 9709 161 9725
rect 253 9713 263 9741
rect 273 9713 293 9747
rect 318 9744 335 9754
rect 303 9728 316 9738
rect 318 9728 324 9744
rect 346 9738 348 9823
rect 400 9815 430 9823
rect 476 9821 480 9889
rect 511 9858 582 9892
rect 544 9851 548 9858
rect 400 9811 436 9815
rect 400 9781 408 9811
rect 420 9781 436 9811
rect 544 9813 548 9821
rect 28 9701 64 9709
rect 127 9708 161 9709
rect 127 9701 182 9708
rect 62 9692 64 9701
rect 282 9655 292 9713
rect 295 9704 324 9728
rect 333 9728 353 9738
rect 428 9734 430 9781
rect 476 9741 480 9809
rect 544 9779 552 9813
rect 578 9779 582 9813
rect 544 9771 548 9779
rect 367 9728 380 9734
rect 333 9704 380 9728
rect 318 9691 324 9704
rect 346 9691 348 9704
rect 367 9700 380 9704
rect 396 9700 408 9734
rect 420 9700 436 9734
rect 544 9731 553 9759
rect 319 9680 346 9691
rect 120 9639 170 9641
rect 76 9633 92 9639
rect 94 9633 110 9639
rect 76 9623 99 9632
rect 60 9613 67 9623
rect 76 9603 77 9623
rect 96 9598 99 9623
rect 109 9603 110 9623
rect 119 9613 126 9623
rect 76 9589 110 9593
rect 170 9589 172 9639
rect 186 9621 190 9655
rect 216 9621 220 9655
rect 182 9583 224 9584
rect 186 9559 220 9576
rect 223 9559 257 9576
rect 182 9542 257 9559
rect 182 9541 224 9542
rect 160 9535 246 9541
rect 288 9535 292 9655
rect 296 9653 368 9661
rect 428 9653 430 9700
rect 476 9663 480 9731
rect 485 9687 495 9721
rect 505 9693 525 9721
rect 505 9687 519 9693
rect 544 9687 555 9731
rect 485 9663 492 9687
rect 579 9672 582 9762
rect 612 9744 624 9745
rect 599 9742 649 9744
rect 612 9741 624 9742
rect 610 9734 632 9741
rect 607 9733 632 9734
rect 586 9726 644 9733
rect 607 9725 644 9726
rect 607 9709 610 9725
rect 616 9709 644 9725
rect 607 9708 644 9709
rect 586 9701 644 9708
rect 607 9700 610 9701
rect 612 9693 632 9701
rect 612 9689 624 9693
rect 649 9692 651 9742
rect 544 9655 548 9663
rect 400 9623 408 9653
rect 420 9623 436 9653
rect 400 9619 436 9623
rect 400 9611 430 9619
rect 428 9595 430 9611
rect 476 9583 480 9651
rect 544 9621 552 9655
rect 578 9621 582 9655
rect 544 9613 548 9621
rect 295 9542 300 9576
rect 324 9542 329 9576
rect 378 9573 450 9581
rect 544 9578 548 9583
rect 544 9574 582 9578
rect 544 9559 552 9574
rect 578 9559 582 9574
rect 544 9541 586 9559
rect 522 9535 608 9541
rect 182 9519 224 9535
rect 544 9519 586 9535
rect 17 9505 67 9507
rect 119 9505 169 9507
rect 186 9505 220 9519
rect 548 9505 582 9519
rect 599 9505 649 9507
rect 42 9463 59 9497
rect 67 9455 69 9505
rect 160 9497 246 9505
rect 522 9497 608 9505
rect 76 9463 110 9497
rect 127 9463 144 9497
rect 152 9463 161 9497
rect 162 9495 195 9497
rect 224 9495 244 9497
rect 162 9463 244 9495
rect 524 9495 548 9497
rect 573 9495 582 9497
rect 586 9495 606 9497
rect 160 9455 246 9463
rect 186 9439 220 9455
rect 182 9425 224 9426
rect 160 9419 182 9425
rect 224 9419 246 9425
rect 186 9384 220 9418
rect 223 9384 257 9418
rect 120 9371 170 9373
rect 76 9367 130 9371
rect 110 9362 130 9367
rect 60 9337 67 9347
rect 76 9337 77 9357
rect 96 9328 99 9362
rect 109 9337 110 9357
rect 119 9337 126 9347
rect 76 9321 92 9327
rect 94 9321 110 9327
rect 170 9321 172 9371
rect 186 9305 190 9339
rect 216 9305 220 9339
rect 288 9305 292 9493
rect 476 9425 480 9493
rect 524 9463 606 9495
rect 607 9463 616 9497
rect 522 9455 608 9463
rect 649 9455 651 9505
rect 548 9439 582 9455
rect 522 9420 548 9425
rect 522 9419 582 9420
rect 586 9419 608 9425
rect 295 9384 300 9418
rect 324 9384 329 9418
rect 544 9416 582 9419
rect 378 9379 450 9387
rect 428 9349 430 9365
rect 400 9341 430 9349
rect 476 9347 480 9415
rect 544 9386 552 9416
rect 578 9386 582 9416
rect 544 9377 548 9386
rect 400 9337 436 9341
rect 400 9307 408 9337
rect 420 9307 436 9337
rect 544 9339 548 9347
rect 12 9268 62 9270
rect 28 9259 59 9267
rect 62 9259 64 9268
rect 28 9251 64 9259
rect 127 9259 158 9267
rect 127 9252 182 9259
rect 215 9257 224 9285
rect 127 9251 161 9252
rect 59 9235 64 9251
rect 158 9235 161 9251
rect 28 9227 64 9235
rect 127 9234 161 9235
rect 127 9227 182 9234
rect 62 9218 64 9227
rect 213 9219 224 9257
rect 282 9247 292 9305
rect 296 9299 368 9307
rect 319 9269 346 9280
rect 318 9256 324 9269
rect 346 9256 348 9269
rect 428 9260 430 9307
rect 443 9297 450 9299
rect 476 9267 480 9335
rect 544 9305 552 9339
rect 578 9305 582 9339
rect 481 9273 517 9301
rect 481 9267 495 9273
rect 367 9256 380 9260
rect 251 9213 263 9247
rect 273 9213 293 9247
rect 295 9232 324 9256
rect 303 9222 316 9232
rect 318 9216 324 9232
rect 333 9232 380 9256
rect 333 9222 353 9232
rect 367 9226 380 9232
rect 396 9226 408 9260
rect 420 9226 436 9260
rect 120 9165 170 9167
rect 76 9159 92 9165
rect 94 9159 110 9165
rect 76 9149 99 9158
rect 60 9139 67 9149
rect 76 9129 77 9149
rect 96 9124 99 9149
rect 109 9129 110 9149
rect 119 9139 126 9149
rect 76 9115 110 9119
rect 170 9115 172 9165
rect 186 9147 190 9181
rect 216 9147 220 9181
rect 186 9070 220 9104
rect 282 9101 292 9213
rect 318 9206 335 9216
rect 318 9137 324 9206
rect 346 9137 348 9222
rect 428 9179 430 9226
rect 476 9189 480 9257
rect 485 9239 495 9267
rect 505 9267 519 9273
rect 544 9267 555 9305
rect 505 9239 525 9267
rect 544 9239 553 9267
rect 544 9219 548 9239
rect 579 9198 582 9288
rect 612 9270 624 9271
rect 599 9268 649 9270
rect 612 9267 624 9268
rect 610 9260 632 9267
rect 607 9259 632 9260
rect 586 9252 644 9259
rect 607 9251 644 9252
rect 607 9235 610 9251
rect 616 9235 644 9251
rect 607 9234 644 9235
rect 586 9227 644 9234
rect 607 9226 610 9227
rect 612 9219 632 9227
rect 612 9215 624 9219
rect 649 9218 651 9268
rect 544 9181 548 9189
rect 400 9149 408 9179
rect 420 9149 436 9179
rect 400 9145 436 9149
rect 400 9137 430 9145
rect 428 9121 430 9137
rect 476 9109 480 9177
rect 544 9147 552 9181
rect 578 9147 582 9181
rect 544 9139 548 9147
rect 544 9109 586 9110
rect 288 9069 292 9101
rect 296 9099 368 9107
rect 378 9099 450 9107
rect 544 9102 548 9109
rect 439 9071 444 9099
rect 120 9055 170 9057
rect 76 9051 130 9055
rect 110 9046 130 9051
rect 60 9021 67 9031
rect 76 9021 77 9041
rect 96 9012 99 9046
rect 109 9021 110 9041
rect 119 9021 126 9031
rect 76 9005 92 9011
rect 94 9005 110 9011
rect 170 9005 172 9055
rect 186 8989 190 9023
rect 216 8989 220 9023
rect 213 8957 224 8989
rect 282 8985 292 9069
rect 296 9063 368 9071
rect 378 9063 450 9071
rect 468 9068 473 9102
rect 428 9033 430 9049
rect 251 8957 292 8985
rect 318 8964 324 9033
rect 12 8952 62 8954
rect 28 8943 59 8951
rect 62 8943 64 8952
rect 251 8951 263 8957
rect 28 8935 64 8943
rect 127 8943 158 8951
rect 127 8936 182 8943
rect 127 8935 161 8936
rect 59 8919 64 8935
rect 158 8919 161 8935
rect 253 8923 263 8951
rect 273 8923 293 8957
rect 318 8954 335 8964
rect 303 8938 316 8948
rect 318 8938 324 8954
rect 346 8948 348 9033
rect 400 9025 430 9033
rect 476 9031 480 9099
rect 511 9068 582 9102
rect 544 9061 548 9068
rect 400 9021 436 9025
rect 400 8991 408 9021
rect 420 8991 436 9021
rect 544 9023 548 9031
rect 28 8911 64 8919
rect 127 8918 161 8919
rect 127 8911 182 8918
rect 62 8902 64 8911
rect 282 8865 292 8923
rect 295 8914 324 8938
rect 333 8938 353 8948
rect 428 8944 430 8991
rect 476 8951 480 9019
rect 544 8989 552 9023
rect 578 8989 582 9023
rect 544 8981 548 8989
rect 367 8938 380 8944
rect 333 8914 380 8938
rect 318 8901 324 8914
rect 346 8901 348 8914
rect 367 8910 380 8914
rect 396 8910 408 8944
rect 420 8910 436 8944
rect 544 8941 553 8969
rect 319 8890 346 8901
rect 120 8849 170 8851
rect 76 8843 92 8849
rect 94 8843 110 8849
rect 76 8833 99 8842
rect 60 8823 67 8833
rect 76 8813 77 8833
rect 96 8808 99 8833
rect 109 8813 110 8833
rect 119 8823 126 8833
rect 76 8799 110 8803
rect 170 8799 172 8849
rect 186 8831 190 8865
rect 216 8831 220 8865
rect 182 8793 224 8794
rect 186 8769 220 8786
rect 223 8769 257 8786
rect 182 8752 257 8769
rect 182 8751 224 8752
rect 160 8745 246 8751
rect 288 8745 292 8865
rect 296 8863 368 8871
rect 428 8863 430 8910
rect 476 8873 480 8941
rect 485 8897 495 8931
rect 505 8903 525 8931
rect 505 8897 519 8903
rect 544 8897 555 8941
rect 485 8873 492 8897
rect 579 8882 582 8972
rect 612 8954 624 8955
rect 599 8952 649 8954
rect 612 8951 624 8952
rect 610 8944 632 8951
rect 607 8943 632 8944
rect 586 8936 644 8943
rect 607 8935 644 8936
rect 607 8919 610 8935
rect 616 8919 644 8935
rect 607 8918 644 8919
rect 586 8911 644 8918
rect 607 8910 610 8911
rect 612 8903 632 8911
rect 612 8899 624 8903
rect 649 8902 651 8952
rect 544 8865 548 8873
rect 400 8833 408 8863
rect 420 8833 436 8863
rect 400 8829 436 8833
rect 400 8821 430 8829
rect 428 8805 430 8821
rect 476 8793 480 8861
rect 544 8831 552 8865
rect 578 8831 582 8865
rect 544 8823 548 8831
rect 295 8752 300 8786
rect 324 8752 329 8786
rect 378 8783 450 8791
rect 544 8788 548 8793
rect 544 8784 582 8788
rect 544 8769 552 8784
rect 578 8769 582 8784
rect 544 8751 586 8769
rect 522 8745 608 8751
rect 182 8729 224 8745
rect 544 8729 586 8745
rect 17 8715 67 8717
rect 119 8715 169 8717
rect 186 8715 220 8729
rect 548 8715 582 8729
rect 599 8715 649 8717
rect 42 8673 59 8707
rect 67 8665 69 8715
rect 160 8707 246 8715
rect 522 8707 608 8715
rect 76 8673 110 8707
rect 127 8673 144 8707
rect 152 8673 161 8707
rect 162 8705 195 8707
rect 224 8705 244 8707
rect 162 8673 244 8705
rect 524 8705 548 8707
rect 573 8705 582 8707
rect 586 8705 606 8707
rect 160 8665 246 8673
rect 186 8649 220 8665
rect 182 8635 224 8636
rect 160 8629 182 8635
rect 224 8629 246 8635
rect 186 8594 220 8628
rect 223 8594 257 8628
rect 120 8581 170 8583
rect 76 8577 130 8581
rect 110 8572 130 8577
rect 60 8547 67 8557
rect 76 8547 77 8567
rect 96 8538 99 8572
rect 109 8547 110 8567
rect 119 8547 126 8557
rect 76 8531 92 8537
rect 94 8531 110 8537
rect 170 8531 172 8581
rect 186 8515 190 8549
rect 216 8515 220 8549
rect 288 8515 292 8703
rect 476 8635 480 8703
rect 524 8673 606 8705
rect 607 8673 616 8707
rect 522 8665 608 8673
rect 649 8665 651 8715
rect 548 8649 582 8665
rect 522 8630 548 8635
rect 522 8629 582 8630
rect 586 8629 608 8635
rect 295 8594 300 8628
rect 324 8594 329 8628
rect 544 8626 582 8629
rect 378 8589 450 8597
rect 428 8559 430 8575
rect 400 8551 430 8559
rect 476 8557 480 8625
rect 544 8596 552 8626
rect 578 8596 582 8626
rect 544 8587 548 8596
rect 400 8547 436 8551
rect 400 8517 408 8547
rect 420 8517 436 8547
rect 544 8549 548 8557
rect 12 8478 62 8480
rect 28 8469 59 8477
rect 62 8469 64 8478
rect 28 8461 64 8469
rect 127 8469 158 8477
rect 127 8462 182 8469
rect 215 8467 224 8495
rect 127 8461 161 8462
rect 59 8445 64 8461
rect 158 8445 161 8461
rect 28 8437 64 8445
rect 127 8444 161 8445
rect 127 8437 182 8444
rect 62 8428 64 8437
rect 213 8429 224 8467
rect 282 8457 292 8515
rect 296 8509 368 8517
rect 319 8479 346 8490
rect 318 8466 324 8479
rect 346 8466 348 8479
rect 428 8470 430 8517
rect 443 8507 450 8509
rect 476 8477 480 8545
rect 544 8515 552 8549
rect 578 8515 582 8549
rect 481 8483 517 8511
rect 481 8477 495 8483
rect 367 8466 380 8470
rect 251 8423 263 8457
rect 273 8423 293 8457
rect 295 8442 324 8466
rect 303 8432 316 8442
rect 318 8426 324 8442
rect 333 8442 380 8466
rect 333 8432 353 8442
rect 367 8436 380 8442
rect 396 8436 408 8470
rect 420 8436 436 8470
rect 120 8375 170 8377
rect 76 8369 92 8375
rect 94 8369 110 8375
rect 76 8359 99 8368
rect 60 8349 67 8359
rect 76 8339 77 8359
rect 96 8334 99 8359
rect 109 8339 110 8359
rect 119 8349 126 8359
rect 76 8325 110 8329
rect 170 8325 172 8375
rect 186 8357 190 8391
rect 216 8357 220 8391
rect 186 8280 220 8314
rect 282 8311 292 8423
rect 318 8416 335 8426
rect 318 8347 324 8416
rect 346 8347 348 8432
rect 428 8389 430 8436
rect 476 8399 480 8467
rect 485 8449 495 8477
rect 505 8477 519 8483
rect 544 8477 555 8515
rect 505 8449 525 8477
rect 544 8449 553 8477
rect 544 8429 548 8449
rect 579 8408 582 8498
rect 612 8480 624 8481
rect 599 8478 649 8480
rect 612 8477 624 8478
rect 610 8470 632 8477
rect 607 8469 632 8470
rect 586 8462 644 8469
rect 607 8461 644 8462
rect 607 8445 610 8461
rect 616 8445 644 8461
rect 607 8444 644 8445
rect 586 8437 644 8444
rect 607 8436 610 8437
rect 612 8429 632 8437
rect 612 8425 624 8429
rect 649 8428 651 8478
rect 544 8391 548 8399
rect 400 8359 408 8389
rect 420 8359 436 8389
rect 400 8355 436 8359
rect 400 8347 430 8355
rect 428 8331 430 8347
rect 476 8319 480 8387
rect 544 8357 552 8391
rect 578 8357 582 8391
rect 544 8349 548 8357
rect 544 8319 586 8320
rect 288 8279 292 8311
rect 296 8309 368 8317
rect 378 8309 450 8317
rect 544 8312 548 8319
rect 439 8281 444 8309
rect 120 8265 170 8267
rect 76 8261 130 8265
rect 110 8256 130 8261
rect 60 8231 67 8241
rect 76 8231 77 8251
rect 96 8222 99 8256
rect 109 8231 110 8251
rect 119 8231 126 8241
rect 76 8215 92 8221
rect 94 8215 110 8221
rect 170 8215 172 8265
rect 186 8199 190 8233
rect 216 8199 220 8233
rect 213 8167 224 8199
rect 282 8195 292 8279
rect 296 8273 368 8281
rect 378 8273 450 8281
rect 468 8278 473 8312
rect 428 8243 430 8259
rect 251 8167 292 8195
rect 318 8174 324 8243
rect 12 8162 62 8164
rect 28 8153 59 8161
rect 62 8153 64 8162
rect 251 8161 263 8167
rect 28 8145 64 8153
rect 127 8153 158 8161
rect 127 8146 182 8153
rect 127 8145 161 8146
rect 59 8129 64 8145
rect 158 8129 161 8145
rect 253 8133 263 8161
rect 273 8133 293 8167
rect 318 8164 335 8174
rect 303 8148 316 8158
rect 318 8148 324 8164
rect 346 8158 348 8243
rect 400 8235 430 8243
rect 476 8241 480 8309
rect 511 8278 582 8312
rect 544 8271 548 8278
rect 400 8231 436 8235
rect 400 8201 408 8231
rect 420 8201 436 8231
rect 544 8233 548 8241
rect 28 8121 64 8129
rect 127 8128 161 8129
rect 127 8121 182 8128
rect 62 8112 64 8121
rect 282 8075 292 8133
rect 295 8124 324 8148
rect 333 8148 353 8158
rect 428 8154 430 8201
rect 476 8161 480 8229
rect 544 8199 552 8233
rect 578 8199 582 8233
rect 544 8191 548 8199
rect 367 8148 380 8154
rect 333 8124 380 8148
rect 318 8111 324 8124
rect 346 8111 348 8124
rect 367 8120 380 8124
rect 396 8120 408 8154
rect 420 8120 436 8154
rect 544 8151 553 8179
rect 319 8100 346 8111
rect 120 8059 170 8061
rect 76 8053 92 8059
rect 94 8053 110 8059
rect 76 8043 99 8052
rect 60 8033 67 8043
rect 76 8023 77 8043
rect 96 8018 99 8043
rect 109 8023 110 8043
rect 119 8033 126 8043
rect 76 8009 110 8013
rect 170 8009 172 8059
rect 186 8041 190 8075
rect 216 8041 220 8075
rect 182 8003 224 8004
rect 186 7979 220 7996
rect 223 7979 257 7996
rect 182 7962 257 7979
rect 182 7961 224 7962
rect 160 7955 246 7961
rect 288 7955 292 8075
rect 296 8073 368 8081
rect 428 8073 430 8120
rect 476 8083 480 8151
rect 485 8107 495 8141
rect 505 8113 525 8141
rect 505 8107 519 8113
rect 544 8107 555 8151
rect 485 8083 492 8107
rect 579 8092 582 8182
rect 612 8164 624 8165
rect 599 8162 649 8164
rect 612 8161 624 8162
rect 610 8154 632 8161
rect 607 8153 632 8154
rect 586 8146 644 8153
rect 607 8145 644 8146
rect 607 8129 610 8145
rect 616 8129 644 8145
rect 607 8128 644 8129
rect 586 8121 644 8128
rect 607 8120 610 8121
rect 612 8113 632 8121
rect 612 8109 624 8113
rect 649 8112 651 8162
rect 544 8075 548 8083
rect 400 8043 408 8073
rect 420 8043 436 8073
rect 400 8039 436 8043
rect 400 8031 430 8039
rect 428 8015 430 8031
rect 476 8003 480 8071
rect 544 8041 552 8075
rect 578 8041 582 8075
rect 544 8033 548 8041
rect 295 7962 300 7996
rect 324 7962 329 7996
rect 378 7993 450 8001
rect 544 7998 548 8003
rect 544 7994 582 7998
rect 544 7979 552 7994
rect 578 7979 582 7994
rect 544 7961 586 7979
rect 522 7955 608 7961
rect 182 7939 224 7955
rect 544 7939 586 7955
rect 17 7925 67 7927
rect 119 7925 169 7927
rect 186 7925 220 7939
rect 548 7925 582 7939
rect 599 7925 649 7927
rect 42 7883 59 7917
rect 67 7875 69 7925
rect 160 7917 246 7925
rect 522 7917 608 7925
rect 76 7883 110 7917
rect 127 7883 144 7917
rect 152 7883 161 7917
rect 162 7915 195 7917
rect 224 7915 244 7917
rect 162 7883 244 7915
rect 524 7915 548 7917
rect 573 7915 582 7917
rect 586 7915 606 7917
rect 160 7875 246 7883
rect 186 7859 220 7875
rect 182 7845 224 7846
rect 160 7839 182 7845
rect 224 7839 246 7845
rect 186 7804 220 7838
rect 223 7804 257 7838
rect 120 7791 170 7793
rect 76 7787 130 7791
rect 110 7782 130 7787
rect 60 7757 67 7767
rect 76 7757 77 7777
rect 96 7748 99 7782
rect 109 7757 110 7777
rect 119 7757 126 7767
rect 76 7741 92 7747
rect 94 7741 110 7747
rect 170 7741 172 7791
rect 186 7725 190 7759
rect 216 7725 220 7759
rect 288 7725 292 7913
rect 476 7845 480 7913
rect 524 7883 606 7915
rect 607 7883 616 7917
rect 522 7875 608 7883
rect 649 7875 651 7925
rect 548 7859 582 7875
rect 522 7840 548 7845
rect 522 7839 582 7840
rect 586 7839 608 7845
rect 295 7804 300 7838
rect 324 7804 329 7838
rect 544 7836 582 7839
rect 378 7799 450 7807
rect 428 7769 430 7785
rect 400 7761 430 7769
rect 476 7767 480 7835
rect 544 7806 552 7836
rect 578 7806 582 7836
rect 544 7797 548 7806
rect 400 7757 436 7761
rect 400 7727 408 7757
rect 420 7727 436 7757
rect 544 7759 548 7767
rect 12 7688 62 7690
rect 28 7679 59 7687
rect 62 7679 64 7688
rect 28 7671 64 7679
rect 127 7679 158 7687
rect 127 7672 182 7679
rect 215 7677 224 7705
rect 127 7671 161 7672
rect 59 7655 64 7671
rect 158 7655 161 7671
rect 28 7647 64 7655
rect 127 7654 161 7655
rect 127 7647 182 7654
rect 62 7638 64 7647
rect 213 7639 224 7677
rect 282 7667 292 7725
rect 296 7719 368 7727
rect 319 7689 346 7700
rect 318 7676 324 7689
rect 346 7676 348 7689
rect 428 7680 430 7727
rect 443 7717 450 7719
rect 476 7687 480 7755
rect 544 7725 552 7759
rect 578 7725 582 7759
rect 481 7693 517 7721
rect 481 7687 495 7693
rect 367 7676 380 7680
rect 251 7633 263 7667
rect 273 7633 293 7667
rect 295 7652 324 7676
rect 303 7642 316 7652
rect 318 7636 324 7652
rect 333 7652 380 7676
rect 333 7642 353 7652
rect 367 7646 380 7652
rect 396 7646 408 7680
rect 420 7646 436 7680
rect 120 7585 170 7587
rect 76 7579 92 7585
rect 94 7579 110 7585
rect 76 7569 99 7578
rect 60 7559 67 7569
rect 76 7549 77 7569
rect 96 7544 99 7569
rect 109 7549 110 7569
rect 119 7559 126 7569
rect 76 7535 110 7539
rect 170 7535 172 7585
rect 186 7567 190 7601
rect 216 7567 220 7601
rect 186 7490 220 7524
rect 282 7521 292 7633
rect 318 7626 335 7636
rect 318 7557 324 7626
rect 346 7557 348 7642
rect 428 7599 430 7646
rect 476 7609 480 7677
rect 485 7659 495 7687
rect 505 7687 519 7693
rect 544 7687 555 7725
rect 505 7659 525 7687
rect 544 7659 553 7687
rect 544 7639 548 7659
rect 579 7618 582 7708
rect 612 7690 624 7691
rect 599 7688 649 7690
rect 612 7687 624 7688
rect 610 7680 632 7687
rect 607 7679 632 7680
rect 586 7672 644 7679
rect 607 7671 644 7672
rect 607 7655 610 7671
rect 616 7655 644 7671
rect 607 7654 644 7655
rect 586 7647 644 7654
rect 607 7646 610 7647
rect 612 7639 632 7647
rect 612 7635 624 7639
rect 649 7638 651 7688
rect 544 7601 548 7609
rect 400 7569 408 7599
rect 420 7569 436 7599
rect 400 7565 436 7569
rect 400 7557 430 7565
rect 428 7541 430 7557
rect 476 7529 480 7597
rect 544 7567 552 7601
rect 578 7567 582 7601
rect 544 7559 548 7567
rect 544 7529 586 7530
rect 288 7489 292 7521
rect 296 7519 368 7527
rect 378 7519 450 7527
rect 544 7522 548 7529
rect 439 7491 444 7519
rect 120 7475 170 7477
rect 76 7471 130 7475
rect 110 7466 130 7471
rect 60 7441 67 7451
rect 76 7441 77 7461
rect 96 7432 99 7466
rect 109 7441 110 7461
rect 119 7441 126 7451
rect 76 7425 92 7431
rect 94 7425 110 7431
rect 170 7425 172 7475
rect 186 7409 190 7443
rect 216 7409 220 7443
rect 213 7377 224 7409
rect 282 7405 292 7489
rect 296 7483 368 7491
rect 378 7483 450 7491
rect 468 7488 473 7522
rect 428 7453 430 7469
rect 251 7377 292 7405
rect 318 7384 324 7453
rect 12 7372 62 7374
rect 28 7363 59 7371
rect 62 7363 64 7372
rect 251 7371 263 7377
rect 28 7355 64 7363
rect 127 7363 158 7371
rect 127 7356 182 7363
rect 127 7355 161 7356
rect 59 7339 64 7355
rect 158 7339 161 7355
rect 253 7343 263 7371
rect 273 7343 293 7377
rect 318 7374 335 7384
rect 303 7358 316 7368
rect 318 7358 324 7374
rect 346 7368 348 7453
rect 400 7445 430 7453
rect 476 7451 480 7519
rect 511 7488 582 7522
rect 544 7481 548 7488
rect 400 7441 436 7445
rect 400 7411 408 7441
rect 420 7411 436 7441
rect 544 7443 548 7451
rect 28 7331 64 7339
rect 127 7338 161 7339
rect 127 7331 182 7338
rect 62 7322 64 7331
rect 282 7285 292 7343
rect 295 7334 324 7358
rect 333 7358 353 7368
rect 428 7364 430 7411
rect 476 7371 480 7439
rect 544 7409 552 7443
rect 578 7409 582 7443
rect 544 7401 548 7409
rect 367 7358 380 7364
rect 333 7334 380 7358
rect 318 7321 324 7334
rect 346 7321 348 7334
rect 367 7330 380 7334
rect 396 7330 408 7364
rect 420 7330 436 7364
rect 544 7361 553 7389
rect 319 7310 346 7321
rect 120 7269 170 7271
rect 76 7263 92 7269
rect 94 7263 110 7269
rect 76 7253 99 7262
rect 60 7243 67 7253
rect 76 7233 77 7253
rect 96 7228 99 7253
rect 109 7233 110 7253
rect 119 7243 126 7253
rect 76 7219 110 7223
rect 170 7219 172 7269
rect 186 7251 190 7285
rect 216 7251 220 7285
rect 182 7213 224 7214
rect 186 7189 220 7206
rect 223 7189 257 7206
rect 182 7172 257 7189
rect 182 7171 224 7172
rect 160 7165 246 7171
rect 288 7165 292 7285
rect 296 7283 368 7291
rect 428 7283 430 7330
rect 476 7293 480 7361
rect 485 7317 495 7351
rect 505 7323 525 7351
rect 505 7317 519 7323
rect 544 7317 555 7361
rect 485 7293 492 7317
rect 579 7302 582 7392
rect 612 7374 624 7375
rect 599 7372 649 7374
rect 612 7371 624 7372
rect 610 7364 632 7371
rect 607 7363 632 7364
rect 586 7356 644 7363
rect 607 7355 644 7356
rect 607 7339 610 7355
rect 616 7339 644 7355
rect 607 7338 644 7339
rect 586 7331 644 7338
rect 607 7330 610 7331
rect 612 7323 632 7331
rect 612 7319 624 7323
rect 649 7322 651 7372
rect 544 7285 548 7293
rect 400 7253 408 7283
rect 420 7253 436 7283
rect 400 7249 436 7253
rect 400 7241 430 7249
rect 428 7225 430 7241
rect 476 7213 480 7281
rect 544 7251 552 7285
rect 578 7251 582 7285
rect 544 7243 548 7251
rect 295 7172 300 7206
rect 324 7172 329 7206
rect 378 7203 450 7211
rect 544 7208 548 7213
rect 544 7204 582 7208
rect 544 7189 552 7204
rect 578 7189 582 7204
rect 544 7171 586 7189
rect 522 7165 608 7171
rect 182 7149 224 7165
rect 544 7149 586 7165
rect 17 7135 67 7137
rect 119 7135 169 7137
rect 186 7135 220 7149
rect 548 7135 582 7149
rect 599 7135 649 7137
rect 42 7093 59 7127
rect 67 7085 69 7135
rect 160 7127 246 7135
rect 522 7127 608 7135
rect 76 7093 110 7127
rect 127 7093 144 7127
rect 152 7093 161 7127
rect 162 7125 195 7127
rect 224 7125 244 7127
rect 162 7093 244 7125
rect 524 7125 548 7127
rect 573 7125 582 7127
rect 586 7125 606 7127
rect 160 7085 246 7093
rect 186 7069 220 7085
rect 182 7055 224 7056
rect 160 7049 182 7055
rect 224 7049 246 7055
rect 186 7014 220 7048
rect 223 7014 257 7048
rect 120 7001 170 7003
rect 76 6997 130 7001
rect 110 6992 130 6997
rect 60 6967 67 6977
rect 76 6967 77 6987
rect 96 6958 99 6992
rect 109 6967 110 6987
rect 119 6967 126 6977
rect 76 6951 92 6957
rect 94 6951 110 6957
rect 170 6951 172 7001
rect 186 6935 190 6969
rect 216 6935 220 6969
rect 288 6935 292 7123
rect 476 7055 480 7123
rect 524 7093 606 7125
rect 607 7093 616 7127
rect 522 7085 608 7093
rect 649 7085 651 7135
rect 548 7069 582 7085
rect 522 7050 548 7055
rect 522 7049 582 7050
rect 586 7049 608 7055
rect 295 7014 300 7048
rect 324 7014 329 7048
rect 544 7046 582 7049
rect 378 7009 450 7017
rect 428 6979 430 6995
rect 400 6971 430 6979
rect 476 6977 480 7045
rect 544 7016 552 7046
rect 578 7016 582 7046
rect 544 7007 548 7016
rect 400 6967 436 6971
rect 400 6937 408 6967
rect 420 6937 436 6967
rect 544 6969 548 6977
rect 12 6898 62 6900
rect 28 6889 59 6897
rect 62 6889 64 6898
rect 28 6881 64 6889
rect 127 6889 158 6897
rect 127 6882 182 6889
rect 215 6887 224 6915
rect 127 6881 161 6882
rect 59 6865 64 6881
rect 158 6865 161 6881
rect 28 6857 64 6865
rect 127 6864 161 6865
rect 127 6857 182 6864
rect 62 6848 64 6857
rect 213 6849 224 6887
rect 282 6877 292 6935
rect 296 6929 368 6937
rect 319 6899 346 6910
rect 318 6886 324 6899
rect 346 6886 348 6899
rect 428 6890 430 6937
rect 443 6927 450 6929
rect 476 6897 480 6965
rect 544 6935 552 6969
rect 578 6935 582 6969
rect 481 6903 517 6931
rect 481 6897 495 6903
rect 367 6886 380 6890
rect 251 6843 263 6877
rect 273 6843 293 6877
rect 295 6862 324 6886
rect 303 6852 316 6862
rect 318 6846 324 6862
rect 333 6862 380 6886
rect 333 6852 353 6862
rect 367 6856 380 6862
rect 396 6856 408 6890
rect 420 6856 436 6890
rect 120 6795 170 6797
rect 76 6789 92 6795
rect 94 6789 110 6795
rect 76 6779 99 6788
rect 60 6769 67 6779
rect 76 6759 77 6779
rect 96 6754 99 6779
rect 109 6759 110 6779
rect 119 6769 126 6779
rect 76 6745 110 6749
rect 170 6745 172 6795
rect 186 6777 190 6811
rect 216 6777 220 6811
rect 186 6700 220 6734
rect 282 6731 292 6843
rect 318 6836 335 6846
rect 318 6767 324 6836
rect 346 6767 348 6852
rect 428 6809 430 6856
rect 476 6819 480 6887
rect 485 6869 495 6897
rect 505 6897 519 6903
rect 544 6897 555 6935
rect 505 6869 525 6897
rect 544 6869 553 6897
rect 544 6849 548 6869
rect 579 6828 582 6918
rect 612 6900 624 6901
rect 599 6898 649 6900
rect 612 6897 624 6898
rect 610 6890 632 6897
rect 607 6889 632 6890
rect 586 6882 644 6889
rect 607 6881 644 6882
rect 607 6865 610 6881
rect 616 6865 644 6881
rect 607 6864 644 6865
rect 586 6857 644 6864
rect 607 6856 610 6857
rect 612 6849 632 6857
rect 612 6845 624 6849
rect 649 6848 651 6898
rect 544 6811 548 6819
rect 400 6779 408 6809
rect 420 6779 436 6809
rect 400 6775 436 6779
rect 400 6767 430 6775
rect 428 6751 430 6767
rect 476 6739 480 6807
rect 544 6777 552 6811
rect 578 6777 582 6811
rect 544 6769 548 6777
rect 544 6739 586 6740
rect 288 6699 292 6731
rect 296 6729 368 6737
rect 378 6729 450 6737
rect 544 6732 548 6739
rect 439 6701 444 6729
rect 120 6685 170 6687
rect 76 6681 130 6685
rect 110 6676 130 6681
rect 60 6651 67 6661
rect 76 6651 77 6671
rect 96 6642 99 6676
rect 109 6651 110 6671
rect 119 6651 126 6661
rect 76 6635 92 6641
rect 94 6635 110 6641
rect 170 6635 172 6685
rect 186 6619 190 6653
rect 216 6619 220 6653
rect 213 6587 224 6619
rect 282 6615 292 6699
rect 296 6693 368 6701
rect 378 6693 450 6701
rect 468 6698 473 6732
rect 428 6663 430 6679
rect 251 6587 292 6615
rect 318 6594 324 6663
rect 12 6582 62 6584
rect 28 6573 59 6581
rect 62 6573 64 6582
rect 251 6581 263 6587
rect 28 6565 64 6573
rect 127 6573 158 6581
rect 127 6566 182 6573
rect 127 6565 161 6566
rect 59 6549 64 6565
rect 158 6549 161 6565
rect 253 6553 263 6581
rect 273 6553 293 6587
rect 318 6584 335 6594
rect 303 6568 316 6578
rect 318 6568 324 6584
rect 346 6578 348 6663
rect 400 6655 430 6663
rect 476 6661 480 6729
rect 511 6698 582 6732
rect 544 6691 548 6698
rect 400 6651 436 6655
rect 400 6621 408 6651
rect 420 6621 436 6651
rect 544 6653 548 6661
rect 28 6541 64 6549
rect 127 6548 161 6549
rect 127 6541 182 6548
rect 62 6532 64 6541
rect 282 6495 292 6553
rect 295 6544 324 6568
rect 333 6568 353 6578
rect 428 6574 430 6621
rect 476 6581 480 6649
rect 544 6619 552 6653
rect 578 6619 582 6653
rect 544 6611 548 6619
rect 367 6568 380 6574
rect 333 6544 380 6568
rect 318 6531 324 6544
rect 346 6531 348 6544
rect 367 6540 380 6544
rect 396 6540 408 6574
rect 420 6540 436 6574
rect 544 6571 553 6599
rect 319 6520 346 6531
rect 120 6479 170 6481
rect 76 6473 92 6479
rect 94 6473 110 6479
rect 76 6463 99 6472
rect 60 6453 67 6463
rect 76 6443 77 6463
rect 96 6438 99 6463
rect 109 6443 110 6463
rect 119 6453 126 6463
rect 76 6429 110 6433
rect 170 6429 172 6479
rect 186 6461 190 6495
rect 216 6461 220 6495
rect 182 6423 224 6424
rect 186 6399 220 6416
rect 223 6399 257 6416
rect 182 6382 257 6399
rect 182 6381 224 6382
rect 160 6375 246 6381
rect 288 6375 292 6495
rect 296 6493 368 6501
rect 428 6493 430 6540
rect 476 6503 480 6571
rect 485 6527 495 6561
rect 505 6533 525 6561
rect 505 6527 519 6533
rect 544 6527 555 6571
rect 485 6503 492 6527
rect 579 6512 582 6602
rect 612 6584 624 6585
rect 599 6582 649 6584
rect 612 6581 624 6582
rect 610 6574 632 6581
rect 607 6573 632 6574
rect 586 6566 644 6573
rect 607 6565 644 6566
rect 607 6549 610 6565
rect 616 6549 644 6565
rect 607 6548 644 6549
rect 586 6541 644 6548
rect 607 6540 610 6541
rect 612 6533 632 6541
rect 612 6529 624 6533
rect 649 6532 651 6582
rect 544 6495 548 6503
rect 400 6463 408 6493
rect 420 6463 436 6493
rect 400 6459 436 6463
rect 400 6451 430 6459
rect 428 6435 430 6451
rect 476 6423 480 6491
rect 544 6461 552 6495
rect 578 6461 582 6495
rect 544 6453 548 6461
rect 295 6382 300 6416
rect 324 6382 329 6416
rect 378 6413 450 6421
rect 544 6418 548 6423
rect 544 6414 582 6418
rect 544 6399 552 6414
rect 578 6399 582 6414
rect 544 6381 586 6399
rect 522 6375 608 6381
rect 182 6359 224 6375
rect 544 6359 586 6375
rect 17 6345 67 6347
rect 119 6345 169 6347
rect 186 6345 220 6359
rect 548 6345 582 6359
rect 599 6345 649 6347
rect 42 6303 59 6337
rect 67 6295 69 6345
rect 160 6337 246 6345
rect 522 6337 608 6345
rect 76 6303 110 6337
rect 127 6303 144 6337
rect 152 6303 161 6337
rect 162 6335 195 6337
rect 224 6335 244 6337
rect 162 6303 244 6335
rect 524 6335 548 6337
rect 573 6335 582 6337
rect 586 6335 606 6337
rect 160 6295 246 6303
rect 186 6279 220 6295
rect 182 6265 224 6266
rect 160 6259 182 6265
rect 224 6259 246 6265
rect 186 6224 220 6258
rect 223 6224 257 6258
rect 120 6211 170 6213
rect 76 6207 130 6211
rect 110 6202 130 6207
rect 60 6177 67 6187
rect 76 6177 77 6197
rect 96 6168 99 6202
rect 109 6177 110 6197
rect 119 6177 126 6187
rect 76 6161 92 6167
rect 94 6161 110 6167
rect 170 6161 172 6211
rect 186 6145 190 6179
rect 216 6145 220 6179
rect 288 6145 292 6333
rect 476 6265 480 6333
rect 524 6303 606 6335
rect 607 6303 616 6337
rect 522 6295 608 6303
rect 649 6295 651 6345
rect 548 6279 582 6295
rect 522 6260 548 6265
rect 522 6259 582 6260
rect 586 6259 608 6265
rect 295 6224 300 6258
rect 324 6224 329 6258
rect 544 6256 582 6259
rect 378 6219 450 6227
rect 428 6189 430 6205
rect 400 6181 430 6189
rect 476 6187 480 6255
rect 544 6226 552 6256
rect 578 6226 582 6256
rect 544 6217 548 6226
rect 400 6177 436 6181
rect 400 6147 408 6177
rect 420 6147 436 6177
rect 544 6179 548 6187
rect 12 6108 62 6110
rect 28 6099 59 6107
rect 62 6099 64 6108
rect 28 6091 64 6099
rect 127 6099 158 6107
rect 127 6092 182 6099
rect 215 6097 224 6125
rect 127 6091 161 6092
rect 59 6075 64 6091
rect 158 6075 161 6091
rect 28 6067 64 6075
rect 127 6074 161 6075
rect 127 6067 182 6074
rect 62 6058 64 6067
rect 213 6059 224 6097
rect 282 6087 292 6145
rect 296 6139 368 6147
rect 319 6109 346 6120
rect 318 6096 324 6109
rect 346 6096 348 6109
rect 428 6100 430 6147
rect 443 6137 450 6139
rect 476 6107 480 6175
rect 544 6145 552 6179
rect 578 6145 582 6179
rect 481 6113 517 6141
rect 481 6107 495 6113
rect 367 6096 380 6100
rect 251 6053 263 6087
rect 273 6053 293 6087
rect 295 6072 324 6096
rect 303 6062 316 6072
rect 318 6056 324 6072
rect 333 6072 380 6096
rect 333 6062 353 6072
rect 367 6066 380 6072
rect 396 6066 408 6100
rect 420 6066 436 6100
rect 120 6005 170 6007
rect 76 5999 92 6005
rect 94 5999 110 6005
rect 76 5989 99 5998
rect 60 5979 67 5989
rect 76 5969 77 5989
rect 96 5964 99 5989
rect 109 5969 110 5989
rect 119 5979 126 5989
rect 76 5955 110 5959
rect 170 5955 172 6005
rect 186 5987 190 6021
rect 216 5987 220 6021
rect 186 5910 220 5944
rect 282 5941 292 6053
rect 318 6046 335 6056
rect 318 5977 324 6046
rect 346 5977 348 6062
rect 428 6019 430 6066
rect 476 6029 480 6097
rect 485 6079 495 6107
rect 505 6107 519 6113
rect 544 6107 555 6145
rect 505 6079 525 6107
rect 544 6079 553 6107
rect 544 6059 548 6079
rect 579 6038 582 6128
rect 612 6110 624 6111
rect 599 6108 649 6110
rect 612 6107 624 6108
rect 610 6100 632 6107
rect 607 6099 632 6100
rect 586 6092 644 6099
rect 607 6091 644 6092
rect 607 6075 610 6091
rect 616 6075 644 6091
rect 607 6074 644 6075
rect 586 6067 644 6074
rect 607 6066 610 6067
rect 612 6059 632 6067
rect 612 6055 624 6059
rect 649 6058 651 6108
rect 544 6021 548 6029
rect 400 5989 408 6019
rect 420 5989 436 6019
rect 400 5985 436 5989
rect 400 5977 430 5985
rect 428 5961 430 5977
rect 476 5949 480 6017
rect 544 5987 552 6021
rect 578 5987 582 6021
rect 544 5979 548 5987
rect 544 5949 586 5950
rect 288 5909 292 5941
rect 296 5939 368 5947
rect 378 5939 450 5947
rect 544 5942 548 5949
rect 439 5911 444 5939
rect 120 5895 170 5897
rect 76 5891 130 5895
rect 110 5886 130 5891
rect 60 5861 67 5871
rect 76 5861 77 5881
rect 96 5852 99 5886
rect 109 5861 110 5881
rect 119 5861 126 5871
rect 76 5845 92 5851
rect 94 5845 110 5851
rect 170 5845 172 5895
rect 186 5829 190 5863
rect 216 5829 220 5863
rect 213 5797 224 5829
rect 282 5825 292 5909
rect 296 5903 368 5911
rect 378 5903 450 5911
rect 468 5908 473 5942
rect 428 5873 430 5889
rect 251 5797 292 5825
rect 318 5804 324 5873
rect 12 5792 62 5794
rect 28 5783 59 5791
rect 62 5783 64 5792
rect 251 5791 263 5797
rect 28 5775 64 5783
rect 127 5783 158 5791
rect 127 5776 182 5783
rect 127 5775 161 5776
rect 59 5759 64 5775
rect 158 5759 161 5775
rect 253 5763 263 5791
rect 273 5763 293 5797
rect 318 5794 335 5804
rect 303 5778 316 5788
rect 318 5778 324 5794
rect 346 5788 348 5873
rect 400 5865 430 5873
rect 476 5871 480 5939
rect 511 5908 582 5942
rect 544 5901 548 5908
rect 400 5861 436 5865
rect 400 5831 408 5861
rect 420 5831 436 5861
rect 544 5863 548 5871
rect 28 5751 64 5759
rect 127 5758 161 5759
rect 127 5751 182 5758
rect 62 5742 64 5751
rect 282 5705 292 5763
rect 295 5754 324 5778
rect 333 5778 353 5788
rect 428 5784 430 5831
rect 476 5791 480 5859
rect 544 5829 552 5863
rect 578 5829 582 5863
rect 544 5821 548 5829
rect 367 5778 380 5784
rect 333 5754 380 5778
rect 318 5741 324 5754
rect 346 5741 348 5754
rect 367 5750 380 5754
rect 396 5750 408 5784
rect 420 5750 436 5784
rect 544 5781 553 5809
rect 319 5730 346 5741
rect 120 5689 170 5691
rect 76 5683 92 5689
rect 94 5683 110 5689
rect 76 5673 99 5682
rect 60 5663 67 5673
rect 76 5653 77 5673
rect 96 5648 99 5673
rect 109 5653 110 5673
rect 119 5663 126 5673
rect 76 5639 110 5643
rect 170 5639 172 5689
rect 186 5671 190 5705
rect 216 5671 220 5705
rect 182 5633 224 5634
rect 186 5609 220 5626
rect 223 5609 257 5626
rect 182 5592 257 5609
rect 182 5591 224 5592
rect 160 5585 246 5591
rect 288 5585 292 5705
rect 296 5703 368 5711
rect 428 5703 430 5750
rect 476 5713 480 5781
rect 485 5737 495 5771
rect 505 5743 525 5771
rect 505 5737 519 5743
rect 544 5737 555 5781
rect 485 5713 492 5737
rect 579 5722 582 5812
rect 612 5794 624 5795
rect 599 5792 649 5794
rect 612 5791 624 5792
rect 610 5784 632 5791
rect 607 5783 632 5784
rect 586 5776 644 5783
rect 607 5775 644 5776
rect 607 5759 610 5775
rect 616 5759 644 5775
rect 607 5758 644 5759
rect 586 5751 644 5758
rect 607 5750 610 5751
rect 612 5743 632 5751
rect 612 5739 624 5743
rect 649 5742 651 5792
rect 544 5705 548 5713
rect 400 5673 408 5703
rect 420 5673 436 5703
rect 400 5669 436 5673
rect 400 5661 430 5669
rect 428 5645 430 5661
rect 476 5633 480 5701
rect 544 5671 552 5705
rect 578 5671 582 5705
rect 544 5663 548 5671
rect 295 5592 300 5626
rect 324 5592 329 5626
rect 378 5623 450 5631
rect 544 5628 548 5633
rect 544 5624 582 5628
rect 544 5609 552 5624
rect 578 5609 582 5624
rect 544 5591 586 5609
rect 522 5585 608 5591
rect 182 5569 224 5585
rect 544 5569 586 5585
rect 17 5555 67 5557
rect 119 5555 169 5557
rect 186 5555 220 5569
rect 548 5555 582 5569
rect 599 5555 649 5557
rect 42 5513 59 5547
rect 67 5505 69 5555
rect 160 5547 246 5555
rect 522 5547 608 5555
rect 76 5513 110 5547
rect 127 5513 144 5547
rect 152 5513 161 5547
rect 162 5545 195 5547
rect 224 5545 244 5547
rect 162 5513 244 5545
rect 524 5545 548 5547
rect 573 5545 582 5547
rect 586 5545 606 5547
rect 160 5505 246 5513
rect 186 5489 220 5505
rect 182 5475 224 5476
rect 160 5469 182 5475
rect 224 5469 246 5475
rect 186 5434 220 5468
rect 223 5434 257 5468
rect 120 5421 170 5423
rect 76 5417 130 5421
rect 110 5412 130 5417
rect 60 5387 67 5397
rect 76 5387 77 5407
rect 96 5378 99 5412
rect 109 5387 110 5407
rect 119 5387 126 5397
rect 76 5371 92 5377
rect 94 5371 110 5377
rect 170 5371 172 5421
rect 186 5355 190 5389
rect 216 5355 220 5389
rect 288 5355 292 5543
rect 476 5475 480 5543
rect 524 5513 606 5545
rect 607 5513 616 5547
rect 522 5505 608 5513
rect 649 5505 651 5555
rect 548 5489 582 5505
rect 522 5470 548 5475
rect 522 5469 582 5470
rect 586 5469 608 5475
rect 295 5434 300 5468
rect 324 5434 329 5468
rect 544 5466 582 5469
rect 378 5429 450 5437
rect 428 5399 430 5415
rect 400 5391 430 5399
rect 476 5397 480 5465
rect 544 5436 552 5466
rect 578 5436 582 5466
rect 544 5427 548 5436
rect 400 5387 436 5391
rect 400 5357 408 5387
rect 420 5357 436 5387
rect 544 5389 548 5397
rect 12 5318 62 5320
rect 28 5309 59 5317
rect 62 5309 64 5318
rect 28 5301 64 5309
rect 127 5309 158 5317
rect 127 5302 182 5309
rect 215 5307 224 5335
rect 127 5301 161 5302
rect 59 5285 64 5301
rect 158 5285 161 5301
rect 28 5277 64 5285
rect 127 5284 161 5285
rect 127 5277 182 5284
rect 62 5268 64 5277
rect 213 5269 224 5307
rect 282 5297 292 5355
rect 296 5349 368 5357
rect 319 5319 346 5330
rect 318 5306 324 5319
rect 346 5306 348 5319
rect 428 5310 430 5357
rect 443 5347 450 5349
rect 476 5317 480 5385
rect 544 5355 552 5389
rect 578 5355 582 5389
rect 481 5323 517 5351
rect 481 5317 495 5323
rect 367 5306 380 5310
rect 251 5263 263 5297
rect 273 5263 293 5297
rect 295 5282 324 5306
rect 303 5272 316 5282
rect 318 5266 324 5282
rect 333 5282 380 5306
rect 333 5272 353 5282
rect 367 5276 380 5282
rect 396 5276 408 5310
rect 420 5276 436 5310
rect 120 5215 170 5217
rect 76 5209 92 5215
rect 94 5209 110 5215
rect 76 5199 99 5208
rect 60 5189 67 5199
rect 76 5179 77 5199
rect 96 5174 99 5199
rect 109 5179 110 5199
rect 119 5189 126 5199
rect 76 5165 110 5169
rect 170 5165 172 5215
rect 186 5197 190 5231
rect 216 5197 220 5231
rect 186 5120 220 5154
rect 282 5151 292 5263
rect 318 5256 335 5266
rect 318 5187 324 5256
rect 346 5187 348 5272
rect 428 5229 430 5276
rect 476 5239 480 5307
rect 485 5289 495 5317
rect 505 5317 519 5323
rect 544 5317 555 5355
rect 505 5289 525 5317
rect 544 5289 553 5317
rect 544 5269 548 5289
rect 579 5248 582 5338
rect 612 5320 624 5321
rect 599 5318 649 5320
rect 612 5317 624 5318
rect 610 5310 632 5317
rect 607 5309 632 5310
rect 586 5302 644 5309
rect 607 5301 644 5302
rect 607 5285 610 5301
rect 616 5285 644 5301
rect 607 5284 644 5285
rect 586 5277 644 5284
rect 607 5276 610 5277
rect 612 5269 632 5277
rect 612 5265 624 5269
rect 649 5268 651 5318
rect 544 5231 548 5239
rect 400 5199 408 5229
rect 420 5199 436 5229
rect 400 5195 436 5199
rect 400 5187 430 5195
rect 428 5171 430 5187
rect 476 5159 480 5227
rect 544 5197 552 5231
rect 578 5197 582 5231
rect 544 5189 548 5197
rect 544 5159 586 5160
rect 288 5119 292 5151
rect 296 5149 368 5157
rect 378 5149 450 5157
rect 544 5152 548 5159
rect 439 5121 444 5149
rect 120 5105 170 5107
rect 76 5101 130 5105
rect 110 5096 130 5101
rect 60 5071 67 5081
rect 76 5071 77 5091
rect 96 5062 99 5096
rect 109 5071 110 5091
rect 119 5071 126 5081
rect 76 5055 92 5061
rect 94 5055 110 5061
rect 170 5055 172 5105
rect 186 5039 190 5073
rect 216 5039 220 5073
rect 213 5007 224 5039
rect 282 5035 292 5119
rect 296 5113 368 5121
rect 378 5113 450 5121
rect 468 5118 473 5152
rect 428 5083 430 5099
rect 251 5007 292 5035
rect 318 5014 324 5083
rect 12 5002 62 5004
rect 28 4993 59 5001
rect 62 4993 64 5002
rect 251 5001 263 5007
rect 28 4985 64 4993
rect 127 4993 158 5001
rect 127 4986 182 4993
rect 127 4985 161 4986
rect 59 4969 64 4985
rect 158 4969 161 4985
rect 253 4973 263 5001
rect 273 4973 293 5007
rect 318 5004 335 5014
rect 303 4988 316 4998
rect 318 4988 324 5004
rect 346 4998 348 5083
rect 400 5075 430 5083
rect 476 5081 480 5149
rect 511 5118 582 5152
rect 544 5111 548 5118
rect 400 5071 436 5075
rect 400 5041 408 5071
rect 420 5041 436 5071
rect 544 5073 548 5081
rect 28 4961 64 4969
rect 127 4968 161 4969
rect 127 4961 182 4968
rect 62 4952 64 4961
rect 282 4915 292 4973
rect 295 4964 324 4988
rect 333 4988 353 4998
rect 428 4994 430 5041
rect 476 5001 480 5069
rect 544 5039 552 5073
rect 578 5039 582 5073
rect 544 5031 548 5039
rect 367 4988 380 4994
rect 333 4964 380 4988
rect 318 4951 324 4964
rect 346 4951 348 4964
rect 367 4960 380 4964
rect 396 4960 408 4994
rect 420 4960 436 4994
rect 544 4991 553 5019
rect 319 4940 346 4951
rect 120 4899 170 4901
rect 76 4893 92 4899
rect 94 4893 110 4899
rect 76 4883 99 4892
rect 60 4873 67 4883
rect 76 4863 77 4883
rect 96 4858 99 4883
rect 109 4863 110 4883
rect 119 4873 126 4883
rect 76 4849 110 4853
rect 170 4849 172 4899
rect 186 4881 190 4915
rect 216 4881 220 4915
rect 182 4843 224 4844
rect 186 4819 220 4836
rect 223 4819 257 4836
rect 182 4802 257 4819
rect 182 4801 224 4802
rect 160 4795 246 4801
rect 288 4795 292 4915
rect 296 4913 368 4921
rect 428 4913 430 4960
rect 476 4923 480 4991
rect 485 4947 495 4981
rect 505 4953 525 4981
rect 505 4947 519 4953
rect 544 4947 555 4991
rect 485 4923 492 4947
rect 579 4932 582 5022
rect 612 5004 624 5005
rect 599 5002 649 5004
rect 612 5001 624 5002
rect 610 4994 632 5001
rect 607 4993 632 4994
rect 586 4986 644 4993
rect 607 4985 644 4986
rect 607 4969 610 4985
rect 616 4969 644 4985
rect 607 4968 644 4969
rect 586 4961 644 4968
rect 607 4960 610 4961
rect 612 4953 632 4961
rect 612 4949 624 4953
rect 649 4952 651 5002
rect 544 4915 548 4923
rect 400 4883 408 4913
rect 420 4883 436 4913
rect 400 4879 436 4883
rect 400 4871 430 4879
rect 428 4855 430 4871
rect 476 4843 480 4911
rect 544 4881 552 4915
rect 578 4881 582 4915
rect 544 4873 548 4881
rect 295 4802 300 4836
rect 324 4802 329 4836
rect 378 4833 450 4841
rect 544 4838 548 4843
rect 544 4834 582 4838
rect 544 4819 552 4834
rect 578 4819 582 4834
rect 544 4801 586 4819
rect 522 4795 608 4801
rect 182 4779 224 4795
rect 544 4779 586 4795
rect 17 4765 67 4767
rect 119 4765 169 4767
rect 186 4765 220 4779
rect 548 4765 582 4779
rect 599 4765 649 4767
rect 42 4723 59 4757
rect 67 4715 69 4765
rect 160 4757 246 4765
rect 522 4757 608 4765
rect 76 4723 110 4757
rect 127 4723 144 4757
rect 152 4723 161 4757
rect 162 4755 195 4757
rect 224 4755 244 4757
rect 162 4723 244 4755
rect 524 4755 548 4757
rect 573 4755 582 4757
rect 586 4755 606 4757
rect 160 4715 246 4723
rect 186 4699 220 4715
rect 182 4685 224 4686
rect 160 4679 182 4685
rect 224 4679 246 4685
rect 186 4644 220 4678
rect 223 4644 257 4678
rect 120 4631 170 4633
rect 76 4627 130 4631
rect 110 4622 130 4627
rect 60 4597 67 4607
rect 76 4597 77 4617
rect 96 4588 99 4622
rect 109 4597 110 4617
rect 119 4597 126 4607
rect 76 4581 92 4587
rect 94 4581 110 4587
rect 170 4581 172 4631
rect 186 4565 190 4599
rect 216 4565 220 4599
rect 288 4565 292 4753
rect 476 4685 480 4753
rect 524 4723 606 4755
rect 607 4723 616 4757
rect 522 4715 608 4723
rect 649 4715 651 4765
rect 548 4699 582 4715
rect 522 4680 548 4685
rect 522 4679 582 4680
rect 586 4679 608 4685
rect 295 4644 300 4678
rect 324 4644 329 4678
rect 544 4676 582 4679
rect 378 4639 450 4647
rect 428 4609 430 4625
rect 400 4601 430 4609
rect 476 4607 480 4675
rect 544 4646 552 4676
rect 578 4646 582 4676
rect 544 4637 548 4646
rect 400 4597 436 4601
rect 400 4567 408 4597
rect 420 4567 436 4597
rect 544 4599 548 4607
rect 12 4528 62 4530
rect 28 4519 59 4527
rect 62 4519 64 4528
rect 28 4511 64 4519
rect 127 4519 158 4527
rect 127 4512 182 4519
rect 215 4517 224 4545
rect 127 4511 161 4512
rect 59 4495 64 4511
rect 158 4495 161 4511
rect 28 4487 64 4495
rect 127 4494 161 4495
rect 127 4487 182 4494
rect 62 4478 64 4487
rect 213 4479 224 4517
rect 282 4507 292 4565
rect 296 4559 368 4567
rect 319 4529 346 4540
rect 318 4516 324 4529
rect 346 4516 348 4529
rect 428 4520 430 4567
rect 443 4557 450 4559
rect 476 4527 480 4595
rect 544 4565 552 4599
rect 578 4565 582 4599
rect 481 4533 517 4561
rect 481 4527 495 4533
rect 367 4516 380 4520
rect 251 4473 263 4507
rect 273 4473 293 4507
rect 295 4492 324 4516
rect 303 4482 316 4492
rect 318 4476 324 4492
rect 333 4492 380 4516
rect 333 4482 353 4492
rect 367 4486 380 4492
rect 396 4486 408 4520
rect 420 4486 436 4520
rect 120 4425 170 4427
rect 76 4419 92 4425
rect 94 4419 110 4425
rect 76 4409 99 4418
rect 60 4399 67 4409
rect 76 4389 77 4409
rect 96 4384 99 4409
rect 109 4389 110 4409
rect 119 4399 126 4409
rect 76 4375 110 4379
rect 170 4375 172 4425
rect 186 4407 190 4441
rect 216 4407 220 4441
rect 186 4330 220 4364
rect 282 4361 292 4473
rect 318 4466 335 4476
rect 318 4397 324 4466
rect 346 4397 348 4482
rect 428 4439 430 4486
rect 476 4449 480 4517
rect 485 4499 495 4527
rect 505 4527 519 4533
rect 544 4527 555 4565
rect 505 4499 525 4527
rect 544 4499 553 4527
rect 544 4479 548 4499
rect 579 4458 582 4548
rect 612 4530 624 4531
rect 599 4528 649 4530
rect 612 4527 624 4528
rect 610 4520 632 4527
rect 607 4519 632 4520
rect 586 4512 644 4519
rect 607 4511 644 4512
rect 607 4495 610 4511
rect 616 4495 644 4511
rect 607 4494 644 4495
rect 586 4487 644 4494
rect 607 4486 610 4487
rect 612 4479 632 4487
rect 612 4475 624 4479
rect 649 4478 651 4528
rect 544 4441 548 4449
rect 400 4409 408 4439
rect 420 4409 436 4439
rect 400 4405 436 4409
rect 400 4397 430 4405
rect 428 4381 430 4397
rect 476 4369 480 4437
rect 544 4407 552 4441
rect 578 4407 582 4441
rect 544 4399 548 4407
rect 544 4369 586 4370
rect 288 4329 292 4361
rect 296 4359 368 4367
rect 378 4359 450 4367
rect 544 4362 548 4369
rect 439 4331 444 4359
rect 120 4315 170 4317
rect 76 4311 130 4315
rect 110 4306 130 4311
rect 60 4281 67 4291
rect 76 4281 77 4301
rect 96 4272 99 4306
rect 109 4281 110 4301
rect 119 4281 126 4291
rect 76 4265 92 4271
rect 94 4265 110 4271
rect 170 4265 172 4315
rect 186 4249 190 4283
rect 216 4249 220 4283
rect 213 4217 224 4249
rect 282 4245 292 4329
rect 296 4323 368 4331
rect 378 4323 450 4331
rect 468 4328 473 4362
rect 428 4293 430 4309
rect 251 4217 292 4245
rect 318 4224 324 4293
rect 12 4212 62 4214
rect 28 4203 59 4211
rect 62 4203 64 4212
rect 251 4211 263 4217
rect 28 4195 64 4203
rect 127 4203 158 4211
rect 127 4196 182 4203
rect 127 4195 161 4196
rect 59 4179 64 4195
rect 158 4179 161 4195
rect 253 4183 263 4211
rect 273 4183 293 4217
rect 318 4214 335 4224
rect 303 4198 316 4208
rect 318 4198 324 4214
rect 346 4208 348 4293
rect 400 4285 430 4293
rect 476 4291 480 4359
rect 511 4328 582 4362
rect 544 4321 548 4328
rect 400 4281 436 4285
rect 400 4251 408 4281
rect 420 4251 436 4281
rect 544 4283 548 4291
rect 28 4171 64 4179
rect 127 4178 161 4179
rect 127 4171 182 4178
rect 62 4162 64 4171
rect 282 4125 292 4183
rect 295 4174 324 4198
rect 333 4198 353 4208
rect 428 4204 430 4251
rect 476 4211 480 4279
rect 544 4249 552 4283
rect 578 4249 582 4283
rect 544 4241 548 4249
rect 367 4198 380 4204
rect 333 4174 380 4198
rect 318 4161 324 4174
rect 346 4161 348 4174
rect 367 4170 380 4174
rect 396 4170 408 4204
rect 420 4170 436 4204
rect 544 4201 553 4229
rect 319 4150 346 4161
rect 120 4109 170 4111
rect 76 4103 92 4109
rect 94 4103 110 4109
rect 76 4093 99 4102
rect 60 4083 67 4093
rect 76 4073 77 4093
rect 96 4068 99 4093
rect 109 4073 110 4093
rect 119 4083 126 4093
rect 76 4059 110 4063
rect 170 4059 172 4109
rect 186 4091 190 4125
rect 216 4091 220 4125
rect 182 4053 224 4054
rect 186 4029 220 4046
rect 223 4029 257 4046
rect 182 4012 257 4029
rect 182 4011 224 4012
rect 160 4005 246 4011
rect 288 4005 292 4125
rect 296 4123 368 4131
rect 428 4123 430 4170
rect 476 4133 480 4201
rect 485 4157 495 4191
rect 505 4163 525 4191
rect 505 4157 519 4163
rect 544 4157 555 4201
rect 485 4133 492 4157
rect 579 4142 582 4232
rect 612 4214 624 4215
rect 599 4212 649 4214
rect 612 4211 624 4212
rect 610 4204 632 4211
rect 607 4203 632 4204
rect 586 4196 644 4203
rect 607 4195 644 4196
rect 607 4179 610 4195
rect 616 4179 644 4195
rect 607 4178 644 4179
rect 586 4171 644 4178
rect 607 4170 610 4171
rect 612 4163 632 4171
rect 612 4159 624 4163
rect 649 4162 651 4212
rect 544 4125 548 4133
rect 400 4093 408 4123
rect 420 4093 436 4123
rect 400 4089 436 4093
rect 400 4081 430 4089
rect 428 4065 430 4081
rect 476 4053 480 4121
rect 544 4091 552 4125
rect 578 4091 582 4125
rect 544 4083 548 4091
rect 295 4012 300 4046
rect 324 4012 329 4046
rect 378 4043 450 4051
rect 544 4048 548 4053
rect 544 4044 582 4048
rect 544 4029 552 4044
rect 578 4029 582 4044
rect 544 4011 586 4029
rect 522 4005 608 4011
rect 182 3989 224 4005
rect 544 3989 586 4005
rect 17 3975 67 3977
rect 119 3975 169 3977
rect 186 3975 220 3989
rect 548 3975 582 3989
rect 599 3975 649 3977
rect 42 3933 59 3967
rect 67 3925 69 3975
rect 160 3967 246 3975
rect 522 3967 608 3975
rect 76 3933 110 3967
rect 127 3933 144 3967
rect 152 3933 161 3967
rect 162 3965 195 3967
rect 224 3965 244 3967
rect 162 3933 244 3965
rect 524 3965 548 3967
rect 573 3965 582 3967
rect 586 3965 606 3967
rect 160 3925 246 3933
rect 186 3909 220 3925
rect 182 3895 224 3896
rect 160 3889 182 3895
rect 224 3889 246 3895
rect 186 3854 220 3888
rect 223 3854 257 3888
rect 120 3841 170 3843
rect 76 3837 130 3841
rect 110 3832 130 3837
rect 60 3807 67 3817
rect 76 3807 77 3827
rect 96 3798 99 3832
rect 109 3807 110 3827
rect 119 3807 126 3817
rect 76 3791 92 3797
rect 94 3791 110 3797
rect 170 3791 172 3841
rect 186 3775 190 3809
rect 216 3775 220 3809
rect 288 3775 292 3963
rect 476 3895 480 3963
rect 524 3933 606 3965
rect 607 3933 616 3967
rect 522 3925 608 3933
rect 649 3925 651 3975
rect 548 3909 582 3925
rect 522 3890 548 3895
rect 522 3889 582 3890
rect 586 3889 608 3895
rect 295 3854 300 3888
rect 324 3854 329 3888
rect 544 3886 582 3889
rect 378 3849 450 3857
rect 428 3819 430 3835
rect 400 3811 430 3819
rect 476 3817 480 3885
rect 544 3856 552 3886
rect 578 3856 582 3886
rect 544 3847 548 3856
rect 400 3807 436 3811
rect 400 3777 408 3807
rect 420 3777 436 3807
rect 544 3809 548 3817
rect 12 3738 62 3740
rect 28 3729 59 3737
rect 62 3729 64 3738
rect 28 3721 64 3729
rect 127 3729 158 3737
rect 127 3722 182 3729
rect 215 3727 224 3755
rect 127 3721 161 3722
rect 59 3705 64 3721
rect 158 3705 161 3721
rect 28 3697 64 3705
rect 127 3704 161 3705
rect 127 3697 182 3704
rect 62 3688 64 3697
rect 213 3689 224 3727
rect 282 3717 292 3775
rect 296 3769 368 3777
rect 319 3739 346 3750
rect 318 3726 324 3739
rect 346 3726 348 3739
rect 428 3730 430 3777
rect 443 3767 450 3769
rect 476 3737 480 3805
rect 544 3775 552 3809
rect 578 3775 582 3809
rect 481 3743 517 3771
rect 481 3737 495 3743
rect 367 3726 380 3730
rect 251 3683 263 3717
rect 273 3683 293 3717
rect 295 3702 324 3726
rect 303 3692 316 3702
rect 318 3686 324 3702
rect 333 3702 380 3726
rect 333 3692 353 3702
rect 367 3696 380 3702
rect 396 3696 408 3730
rect 420 3696 436 3730
rect 120 3635 170 3637
rect 76 3629 92 3635
rect 94 3629 110 3635
rect 76 3619 99 3628
rect 60 3609 67 3619
rect 76 3599 77 3619
rect 96 3594 99 3619
rect 109 3599 110 3619
rect 119 3609 126 3619
rect 76 3585 110 3589
rect 170 3585 172 3635
rect 186 3617 190 3651
rect 216 3617 220 3651
rect 186 3540 220 3574
rect 282 3571 292 3683
rect 318 3676 335 3686
rect 318 3607 324 3676
rect 346 3607 348 3692
rect 428 3649 430 3696
rect 476 3659 480 3727
rect 485 3709 495 3737
rect 505 3737 519 3743
rect 544 3737 555 3775
rect 505 3709 525 3737
rect 544 3709 553 3737
rect 544 3689 548 3709
rect 579 3668 582 3758
rect 612 3740 624 3741
rect 599 3738 649 3740
rect 612 3737 624 3738
rect 610 3730 632 3737
rect 607 3729 632 3730
rect 586 3722 644 3729
rect 607 3721 644 3722
rect 607 3705 610 3721
rect 616 3705 644 3721
rect 607 3704 644 3705
rect 586 3697 644 3704
rect 607 3696 610 3697
rect 612 3689 632 3697
rect 612 3685 624 3689
rect 649 3688 651 3738
rect 544 3651 548 3659
rect 400 3619 408 3649
rect 420 3619 436 3649
rect 400 3615 436 3619
rect 400 3607 430 3615
rect 428 3591 430 3607
rect 476 3579 480 3647
rect 544 3617 552 3651
rect 578 3617 582 3651
rect 544 3609 548 3617
rect 544 3579 586 3580
rect 288 3539 292 3571
rect 296 3569 368 3577
rect 378 3569 450 3577
rect 544 3572 548 3579
rect 439 3541 444 3569
rect 120 3525 170 3527
rect 76 3521 130 3525
rect 110 3516 130 3521
rect 60 3491 67 3501
rect 76 3491 77 3511
rect 96 3482 99 3516
rect 109 3491 110 3511
rect 119 3491 126 3501
rect 76 3475 92 3481
rect 94 3475 110 3481
rect 170 3475 172 3525
rect 186 3459 190 3493
rect 216 3459 220 3493
rect 213 3427 224 3459
rect 282 3455 292 3539
rect 296 3533 368 3541
rect 378 3533 450 3541
rect 468 3538 473 3572
rect 428 3503 430 3519
rect 251 3427 292 3455
rect 318 3434 324 3503
rect 12 3422 62 3424
rect 28 3413 59 3421
rect 62 3413 64 3422
rect 251 3421 263 3427
rect 28 3405 64 3413
rect 127 3413 158 3421
rect 127 3406 182 3413
rect 127 3405 161 3406
rect 59 3389 64 3405
rect 158 3389 161 3405
rect 253 3393 263 3421
rect 273 3393 293 3427
rect 318 3424 335 3434
rect 303 3408 316 3418
rect 318 3408 324 3424
rect 346 3418 348 3503
rect 400 3495 430 3503
rect 476 3501 480 3569
rect 511 3538 582 3572
rect 544 3531 548 3538
rect 400 3491 436 3495
rect 400 3461 408 3491
rect 420 3461 436 3491
rect 544 3493 548 3501
rect 28 3381 64 3389
rect 127 3388 161 3389
rect 127 3381 182 3388
rect 62 3372 64 3381
rect 282 3335 292 3393
rect 295 3384 324 3408
rect 333 3408 353 3418
rect 428 3414 430 3461
rect 476 3421 480 3489
rect 544 3459 552 3493
rect 578 3459 582 3493
rect 544 3451 548 3459
rect 367 3408 380 3414
rect 333 3384 380 3408
rect 318 3371 324 3384
rect 346 3371 348 3384
rect 367 3380 380 3384
rect 396 3380 408 3414
rect 420 3380 436 3414
rect 544 3411 553 3439
rect 319 3360 346 3371
rect 120 3319 170 3321
rect 76 3313 92 3319
rect 94 3313 110 3319
rect 76 3303 99 3312
rect 60 3293 67 3303
rect 76 3283 77 3303
rect 96 3278 99 3303
rect 109 3283 110 3303
rect 119 3293 126 3303
rect 76 3269 110 3273
rect 170 3269 172 3319
rect 186 3301 190 3335
rect 216 3301 220 3335
rect 182 3263 224 3264
rect 186 3239 220 3256
rect 223 3239 257 3256
rect 182 3222 257 3239
rect 182 3221 224 3222
rect 160 3215 246 3221
rect 288 3215 292 3335
rect 296 3333 368 3341
rect 428 3333 430 3380
rect 476 3343 480 3411
rect 485 3367 495 3401
rect 505 3373 525 3401
rect 505 3367 519 3373
rect 544 3367 555 3411
rect 485 3343 492 3367
rect 579 3352 582 3442
rect 612 3424 624 3425
rect 599 3422 649 3424
rect 612 3421 624 3422
rect 610 3414 632 3421
rect 607 3413 632 3414
rect 586 3406 644 3413
rect 607 3405 644 3406
rect 607 3389 610 3405
rect 616 3389 644 3405
rect 607 3388 644 3389
rect 586 3381 644 3388
rect 607 3380 610 3381
rect 612 3373 632 3381
rect 612 3369 624 3373
rect 649 3372 651 3422
rect 544 3335 548 3343
rect 400 3303 408 3333
rect 420 3303 436 3333
rect 400 3299 436 3303
rect 400 3291 430 3299
rect 428 3275 430 3291
rect 476 3263 480 3331
rect 544 3301 552 3335
rect 578 3301 582 3335
rect 544 3293 548 3301
rect 295 3222 300 3256
rect 324 3222 329 3256
rect 378 3253 450 3261
rect 544 3258 548 3263
rect 544 3254 582 3258
rect 544 3239 552 3254
rect 578 3239 582 3254
rect 544 3221 586 3239
rect 522 3215 608 3221
rect 182 3199 224 3215
rect 544 3199 586 3215
rect 17 3185 67 3187
rect 119 3185 169 3187
rect 186 3185 220 3199
rect 548 3185 582 3199
rect 599 3185 649 3187
rect 42 3143 59 3177
rect 67 3135 69 3185
rect 160 3177 246 3185
rect 522 3177 608 3185
rect 76 3143 110 3177
rect 127 3143 144 3177
rect 152 3143 161 3177
rect 162 3175 195 3177
rect 224 3175 244 3177
rect 162 3143 244 3175
rect 524 3175 548 3177
rect 573 3175 582 3177
rect 586 3175 606 3177
rect 160 3135 246 3143
rect 186 3119 220 3135
rect 182 3105 224 3106
rect 160 3099 182 3105
rect 224 3099 246 3105
rect 186 3064 220 3098
rect 223 3064 257 3098
rect 120 3051 170 3053
rect 76 3047 130 3051
rect 110 3042 130 3047
rect 60 3017 67 3027
rect 76 3017 77 3037
rect 96 3008 99 3042
rect 109 3017 110 3037
rect 119 3017 126 3027
rect 76 3001 92 3007
rect 94 3001 110 3007
rect 170 3001 172 3051
rect 186 2985 190 3019
rect 216 2985 220 3019
rect 288 2985 292 3173
rect 476 3105 480 3173
rect 524 3143 606 3175
rect 607 3143 616 3177
rect 522 3135 608 3143
rect 649 3135 651 3185
rect 548 3119 582 3135
rect 522 3100 548 3105
rect 522 3099 582 3100
rect 586 3099 608 3105
rect 295 3064 300 3098
rect 324 3064 329 3098
rect 544 3096 582 3099
rect 378 3059 450 3067
rect 428 3029 430 3045
rect 400 3021 430 3029
rect 476 3027 480 3095
rect 544 3066 552 3096
rect 578 3066 582 3096
rect 544 3057 548 3066
rect 400 3017 436 3021
rect 400 2987 408 3017
rect 420 2987 436 3017
rect 544 3019 548 3027
rect 12 2948 62 2950
rect 28 2939 59 2947
rect 62 2939 64 2948
rect 28 2931 64 2939
rect 127 2939 158 2947
rect 127 2932 182 2939
rect 215 2937 224 2965
rect 127 2931 161 2932
rect 59 2915 64 2931
rect 158 2915 161 2931
rect 28 2907 64 2915
rect 127 2914 161 2915
rect 127 2907 182 2914
rect 62 2898 64 2907
rect 213 2899 224 2937
rect 282 2927 292 2985
rect 296 2979 368 2987
rect 319 2949 346 2960
rect 318 2936 324 2949
rect 346 2936 348 2949
rect 428 2940 430 2987
rect 443 2977 450 2979
rect 476 2947 480 3015
rect 544 2985 552 3019
rect 578 2985 582 3019
rect 481 2953 517 2981
rect 481 2947 495 2953
rect 367 2936 380 2940
rect 251 2893 263 2927
rect 273 2893 293 2927
rect 295 2912 324 2936
rect 303 2902 316 2912
rect 318 2896 324 2912
rect 333 2912 380 2936
rect 333 2902 353 2912
rect 367 2906 380 2912
rect 396 2906 408 2940
rect 420 2906 436 2940
rect 120 2845 170 2847
rect 76 2839 92 2845
rect 94 2839 110 2845
rect 76 2829 99 2838
rect 60 2819 67 2829
rect 76 2809 77 2829
rect 96 2804 99 2829
rect 109 2809 110 2829
rect 119 2819 126 2829
rect 76 2795 110 2799
rect 170 2795 172 2845
rect 186 2827 190 2861
rect 216 2827 220 2861
rect 186 2750 220 2784
rect 282 2781 292 2893
rect 318 2886 335 2896
rect 318 2817 324 2886
rect 346 2817 348 2902
rect 428 2859 430 2906
rect 476 2869 480 2937
rect 485 2919 495 2947
rect 505 2947 519 2953
rect 544 2947 555 2985
rect 505 2919 525 2947
rect 544 2919 553 2947
rect 544 2899 548 2919
rect 579 2878 582 2968
rect 612 2950 624 2951
rect 599 2948 649 2950
rect 612 2947 624 2948
rect 610 2940 632 2947
rect 607 2939 632 2940
rect 586 2932 644 2939
rect 607 2931 644 2932
rect 607 2915 610 2931
rect 616 2915 644 2931
rect 607 2914 644 2915
rect 586 2907 644 2914
rect 607 2906 610 2907
rect 612 2899 632 2907
rect 612 2895 624 2899
rect 649 2898 651 2948
rect 544 2861 548 2869
rect 400 2829 408 2859
rect 420 2829 436 2859
rect 400 2825 436 2829
rect 400 2817 430 2825
rect 428 2801 430 2817
rect 476 2789 480 2857
rect 544 2827 552 2861
rect 578 2827 582 2861
rect 544 2819 548 2827
rect 544 2789 586 2790
rect 288 2749 292 2781
rect 296 2779 368 2787
rect 378 2779 450 2787
rect 544 2782 548 2789
rect 439 2751 444 2779
rect 120 2735 170 2737
rect 76 2731 130 2735
rect 110 2726 130 2731
rect 60 2701 67 2711
rect 76 2701 77 2721
rect 96 2692 99 2726
rect 109 2701 110 2721
rect 119 2701 126 2711
rect 76 2685 92 2691
rect 94 2685 110 2691
rect 170 2685 172 2735
rect 186 2669 190 2703
rect 216 2669 220 2703
rect 213 2637 224 2669
rect 282 2665 292 2749
rect 296 2743 368 2751
rect 378 2743 450 2751
rect 468 2748 473 2782
rect 428 2713 430 2729
rect 251 2637 292 2665
rect 318 2644 324 2713
rect 12 2632 62 2634
rect 28 2623 59 2631
rect 62 2623 64 2632
rect 251 2631 263 2637
rect 28 2615 64 2623
rect 127 2623 158 2631
rect 127 2616 182 2623
rect 127 2615 161 2616
rect 59 2599 64 2615
rect 158 2599 161 2615
rect 253 2603 263 2631
rect 273 2603 293 2637
rect 318 2634 335 2644
rect 303 2618 316 2628
rect 318 2618 324 2634
rect 346 2628 348 2713
rect 400 2705 430 2713
rect 476 2711 480 2779
rect 511 2748 582 2782
rect 544 2741 548 2748
rect 400 2701 436 2705
rect 400 2671 408 2701
rect 420 2671 436 2701
rect 544 2703 548 2711
rect 28 2591 64 2599
rect 127 2598 161 2599
rect 127 2591 182 2598
rect 62 2582 64 2591
rect 282 2545 292 2603
rect 295 2594 324 2618
rect 333 2618 353 2628
rect 428 2624 430 2671
rect 476 2631 480 2699
rect 544 2669 552 2703
rect 578 2669 582 2703
rect 544 2661 548 2669
rect 367 2618 380 2624
rect 333 2594 380 2618
rect 318 2581 324 2594
rect 346 2581 348 2594
rect 367 2590 380 2594
rect 396 2590 408 2624
rect 420 2590 436 2624
rect 544 2621 553 2649
rect 319 2570 346 2581
rect 120 2529 170 2531
rect 76 2523 92 2529
rect 94 2523 110 2529
rect 76 2513 99 2522
rect 60 2503 67 2513
rect 76 2493 77 2513
rect 96 2488 99 2513
rect 109 2493 110 2513
rect 119 2503 126 2513
rect 76 2479 110 2483
rect 170 2479 172 2529
rect 186 2511 190 2545
rect 216 2511 220 2545
rect 182 2473 224 2474
rect 186 2449 220 2466
rect 223 2449 257 2466
rect 182 2432 257 2449
rect 182 2431 224 2432
rect 160 2425 246 2431
rect 288 2425 292 2545
rect 296 2543 368 2551
rect 428 2543 430 2590
rect 476 2553 480 2621
rect 485 2577 495 2611
rect 505 2583 525 2611
rect 505 2577 519 2583
rect 544 2577 555 2621
rect 485 2553 492 2577
rect 579 2562 582 2652
rect 612 2634 624 2635
rect 599 2632 649 2634
rect 612 2631 624 2632
rect 610 2624 632 2631
rect 607 2623 632 2624
rect 586 2616 644 2623
rect 607 2615 644 2616
rect 607 2599 610 2615
rect 616 2599 644 2615
rect 607 2598 644 2599
rect 586 2591 644 2598
rect 607 2590 610 2591
rect 612 2583 632 2591
rect 612 2579 624 2583
rect 649 2582 651 2632
rect 544 2545 548 2553
rect 400 2513 408 2543
rect 420 2513 436 2543
rect 400 2509 436 2513
rect 400 2501 430 2509
rect 428 2485 430 2501
rect 476 2473 480 2541
rect 544 2511 552 2545
rect 578 2511 582 2545
rect 544 2503 548 2511
rect 295 2432 300 2466
rect 324 2432 329 2466
rect 378 2463 450 2471
rect 544 2468 548 2473
rect 544 2464 582 2468
rect 544 2449 552 2464
rect 578 2449 582 2464
rect 544 2431 586 2449
rect 522 2425 608 2431
rect 182 2409 224 2425
rect 544 2409 586 2425
rect 17 2395 67 2397
rect 119 2395 169 2397
rect 186 2395 220 2409
rect 548 2395 582 2409
rect 599 2395 649 2397
rect 42 2353 59 2387
rect 67 2345 69 2395
rect 160 2387 246 2395
rect 522 2387 608 2395
rect 76 2353 110 2387
rect 127 2353 144 2387
rect 152 2353 161 2387
rect 162 2385 195 2387
rect 224 2385 244 2387
rect 162 2353 244 2385
rect 524 2385 548 2387
rect 573 2385 582 2387
rect 586 2385 606 2387
rect 160 2345 246 2353
rect 186 2329 220 2345
rect 182 2315 224 2316
rect 160 2309 182 2315
rect 224 2309 246 2315
rect 186 2274 220 2308
rect 223 2274 257 2308
rect 120 2261 170 2263
rect 76 2257 130 2261
rect 110 2252 130 2257
rect 60 2227 67 2237
rect 76 2227 77 2247
rect 96 2218 99 2252
rect 109 2227 110 2247
rect 119 2227 126 2237
rect 76 2211 92 2217
rect 94 2211 110 2217
rect 170 2211 172 2261
rect 186 2195 190 2229
rect 216 2195 220 2229
rect 288 2195 292 2383
rect 476 2315 480 2383
rect 524 2353 606 2385
rect 607 2353 616 2387
rect 522 2345 608 2353
rect 649 2345 651 2395
rect 548 2329 582 2345
rect 522 2310 548 2315
rect 522 2309 582 2310
rect 586 2309 608 2315
rect 295 2274 300 2308
rect 324 2274 329 2308
rect 544 2306 582 2309
rect 378 2269 450 2277
rect 428 2239 430 2255
rect 400 2231 430 2239
rect 476 2237 480 2305
rect 544 2276 552 2306
rect 578 2276 582 2306
rect 544 2267 548 2276
rect 400 2227 436 2231
rect 400 2197 408 2227
rect 420 2197 436 2227
rect 544 2229 548 2237
rect 12 2158 62 2160
rect 28 2149 59 2157
rect 62 2149 64 2158
rect 28 2141 64 2149
rect 127 2149 158 2157
rect 127 2142 182 2149
rect 215 2147 224 2175
rect 127 2141 161 2142
rect 59 2125 64 2141
rect 158 2125 161 2141
rect 28 2117 64 2125
rect 127 2124 161 2125
rect 127 2117 182 2124
rect 62 2108 64 2117
rect 213 2109 224 2147
rect 282 2137 292 2195
rect 296 2189 368 2197
rect 319 2159 346 2170
rect 318 2146 324 2159
rect 346 2146 348 2159
rect 428 2150 430 2197
rect 443 2187 450 2189
rect 476 2157 480 2225
rect 544 2195 552 2229
rect 578 2195 582 2229
rect 481 2163 517 2191
rect 481 2157 495 2163
rect 367 2146 380 2150
rect 251 2103 263 2137
rect 273 2103 293 2137
rect 295 2122 324 2146
rect 303 2112 316 2122
rect 318 2106 324 2122
rect 333 2122 380 2146
rect 333 2112 353 2122
rect 367 2116 380 2122
rect 396 2116 408 2150
rect 420 2116 436 2150
rect 120 2055 170 2057
rect 76 2049 92 2055
rect 94 2049 110 2055
rect 76 2039 99 2048
rect 60 2029 67 2039
rect 76 2019 77 2039
rect 96 2014 99 2039
rect 109 2019 110 2039
rect 119 2029 126 2039
rect 76 2005 110 2009
rect 170 2005 172 2055
rect 186 2037 190 2071
rect 216 2037 220 2071
rect 186 1960 220 1994
rect 282 1991 292 2103
rect 318 2096 335 2106
rect 318 2027 324 2096
rect 346 2027 348 2112
rect 428 2069 430 2116
rect 476 2079 480 2147
rect 485 2129 495 2157
rect 505 2157 519 2163
rect 544 2157 555 2195
rect 505 2129 525 2157
rect 544 2129 553 2157
rect 544 2109 548 2129
rect 579 2088 582 2178
rect 612 2160 624 2161
rect 599 2158 649 2160
rect 612 2157 624 2158
rect 610 2150 632 2157
rect 607 2149 632 2150
rect 586 2142 644 2149
rect 607 2141 644 2142
rect 607 2125 610 2141
rect 616 2125 644 2141
rect 607 2124 644 2125
rect 586 2117 644 2124
rect 607 2116 610 2117
rect 612 2109 632 2117
rect 612 2105 624 2109
rect 649 2108 651 2158
rect 544 2071 548 2079
rect 400 2039 408 2069
rect 420 2039 436 2069
rect 400 2035 436 2039
rect 400 2027 430 2035
rect 428 2011 430 2027
rect 476 1999 480 2067
rect 544 2037 552 2071
rect 578 2037 582 2071
rect 544 2029 548 2037
rect 544 1999 586 2000
rect 288 1959 292 1991
rect 296 1989 368 1997
rect 378 1989 450 1997
rect 544 1992 548 1999
rect 439 1961 444 1989
rect 120 1945 170 1947
rect 76 1941 130 1945
rect 110 1936 130 1941
rect 60 1911 67 1921
rect 76 1911 77 1931
rect 96 1902 99 1936
rect 109 1911 110 1931
rect 119 1911 126 1921
rect 76 1895 92 1901
rect 94 1895 110 1901
rect 170 1895 172 1945
rect 186 1879 190 1913
rect 216 1879 220 1913
rect 213 1847 224 1879
rect 282 1875 292 1959
rect 296 1953 368 1961
rect 378 1953 450 1961
rect 468 1958 473 1992
rect 428 1923 430 1939
rect 251 1847 292 1875
rect 318 1854 324 1923
rect 12 1842 62 1844
rect 28 1833 59 1841
rect 62 1833 64 1842
rect 251 1841 263 1847
rect 28 1825 64 1833
rect 127 1833 158 1841
rect 127 1826 182 1833
rect 127 1825 161 1826
rect 59 1809 64 1825
rect 158 1809 161 1825
rect 253 1813 263 1841
rect 273 1813 293 1847
rect 318 1844 335 1854
rect 303 1828 316 1838
rect 318 1828 324 1844
rect 346 1838 348 1923
rect 400 1915 430 1923
rect 476 1921 480 1989
rect 511 1958 582 1992
rect 544 1951 548 1958
rect 400 1911 436 1915
rect 400 1881 408 1911
rect 420 1881 436 1911
rect 544 1913 548 1921
rect 28 1801 64 1809
rect 127 1808 161 1809
rect 127 1801 182 1808
rect 62 1792 64 1801
rect 282 1755 292 1813
rect 295 1804 324 1828
rect 333 1828 353 1838
rect 428 1834 430 1881
rect 476 1841 480 1909
rect 544 1879 552 1913
rect 578 1879 582 1913
rect 544 1871 548 1879
rect 367 1828 380 1834
rect 333 1804 380 1828
rect 318 1791 324 1804
rect 346 1791 348 1804
rect 367 1800 380 1804
rect 396 1800 408 1834
rect 420 1800 436 1834
rect 544 1831 553 1859
rect 319 1780 346 1791
rect 120 1739 170 1741
rect 76 1733 92 1739
rect 94 1733 110 1739
rect 76 1723 99 1732
rect 60 1713 67 1723
rect 76 1703 77 1723
rect 96 1698 99 1723
rect 109 1703 110 1723
rect 119 1713 126 1723
rect 76 1689 110 1693
rect 170 1689 172 1739
rect 186 1721 190 1755
rect 216 1721 220 1755
rect 182 1683 224 1684
rect 186 1659 220 1676
rect 223 1659 257 1676
rect 182 1642 257 1659
rect 182 1641 224 1642
rect 160 1635 246 1641
rect 288 1635 292 1755
rect 296 1753 368 1761
rect 428 1753 430 1800
rect 476 1763 480 1831
rect 485 1787 495 1821
rect 505 1793 525 1821
rect 505 1787 519 1793
rect 544 1787 555 1831
rect 485 1763 492 1787
rect 579 1772 582 1862
rect 612 1844 624 1845
rect 599 1842 649 1844
rect 612 1841 624 1842
rect 610 1834 632 1841
rect 607 1833 632 1834
rect 586 1826 644 1833
rect 607 1825 644 1826
rect 607 1809 610 1825
rect 616 1809 644 1825
rect 607 1808 644 1809
rect 586 1801 644 1808
rect 607 1800 610 1801
rect 612 1793 632 1801
rect 612 1789 624 1793
rect 649 1792 651 1842
rect 544 1755 548 1763
rect 400 1723 408 1753
rect 420 1723 436 1753
rect 400 1719 436 1723
rect 400 1711 430 1719
rect 428 1695 430 1711
rect 476 1683 480 1751
rect 544 1721 552 1755
rect 578 1721 582 1755
rect 544 1713 548 1721
rect 295 1642 300 1676
rect 324 1642 329 1676
rect 378 1673 450 1681
rect 544 1678 548 1683
rect 544 1674 582 1678
rect 544 1659 552 1674
rect 578 1659 582 1674
rect 544 1641 586 1659
rect 522 1635 608 1641
rect 182 1619 224 1635
rect 544 1619 586 1635
rect 17 1605 67 1607
rect 119 1605 169 1607
rect 186 1605 220 1619
rect 548 1605 582 1619
rect 599 1605 649 1607
rect 42 1563 59 1597
rect 67 1555 69 1605
rect 160 1597 246 1605
rect 522 1597 608 1605
rect 76 1563 110 1597
rect 127 1563 144 1597
rect 152 1563 161 1597
rect 162 1595 195 1597
rect 224 1595 244 1597
rect 162 1563 244 1595
rect 524 1595 548 1597
rect 573 1595 582 1597
rect 586 1595 606 1597
rect 160 1555 246 1563
rect 186 1539 220 1555
rect 182 1525 224 1526
rect 160 1519 182 1525
rect 224 1519 246 1525
rect 186 1484 220 1518
rect 223 1484 257 1518
rect 120 1471 170 1473
rect 76 1467 130 1471
rect 110 1462 130 1467
rect 60 1437 67 1447
rect 76 1437 77 1457
rect 96 1428 99 1462
rect 109 1437 110 1457
rect 119 1437 126 1447
rect 76 1421 92 1427
rect 94 1421 110 1427
rect 170 1421 172 1471
rect 186 1405 190 1439
rect 216 1405 220 1439
rect 288 1405 292 1593
rect 476 1525 480 1593
rect 524 1563 606 1595
rect 607 1563 616 1597
rect 522 1555 608 1563
rect 649 1555 651 1605
rect 548 1539 582 1555
rect 522 1520 548 1525
rect 522 1519 582 1520
rect 586 1519 608 1525
rect 295 1484 300 1518
rect 324 1484 329 1518
rect 544 1516 582 1519
rect 378 1479 450 1487
rect 428 1449 430 1465
rect 400 1441 430 1449
rect 476 1447 480 1515
rect 544 1486 552 1516
rect 578 1486 582 1516
rect 544 1477 548 1486
rect 400 1437 436 1441
rect 400 1407 408 1437
rect 420 1407 436 1437
rect 544 1439 548 1447
rect 12 1368 62 1370
rect 28 1359 59 1367
rect 62 1359 64 1368
rect 28 1351 64 1359
rect 127 1359 158 1367
rect 127 1352 182 1359
rect 215 1357 224 1385
rect 127 1351 161 1352
rect 59 1335 64 1351
rect 158 1335 161 1351
rect 28 1327 64 1335
rect 127 1334 161 1335
rect 127 1327 182 1334
rect 62 1318 64 1327
rect 213 1319 224 1357
rect 282 1347 292 1405
rect 296 1399 368 1407
rect 319 1369 346 1380
rect 318 1356 324 1369
rect 346 1356 348 1369
rect 428 1360 430 1407
rect 443 1397 450 1399
rect 476 1367 480 1435
rect 544 1405 552 1439
rect 578 1405 582 1439
rect 481 1373 517 1401
rect 481 1367 495 1373
rect 367 1356 380 1360
rect 251 1313 263 1347
rect 273 1313 293 1347
rect 295 1332 324 1356
rect 303 1322 316 1332
rect 318 1316 324 1332
rect 333 1332 380 1356
rect 333 1322 353 1332
rect 367 1326 380 1332
rect 396 1326 408 1360
rect 420 1326 436 1360
rect 120 1265 170 1267
rect 76 1259 92 1265
rect 94 1259 110 1265
rect 76 1249 99 1258
rect 60 1239 67 1249
rect 76 1229 77 1249
rect 96 1224 99 1249
rect 109 1229 110 1249
rect 119 1239 126 1249
rect 76 1215 110 1219
rect 170 1215 172 1265
rect 186 1247 190 1281
rect 216 1247 220 1281
rect 186 1170 220 1204
rect 282 1201 292 1313
rect 318 1306 335 1316
rect 318 1237 324 1306
rect 346 1237 348 1322
rect 428 1279 430 1326
rect 476 1289 480 1357
rect 485 1339 495 1367
rect 505 1367 519 1373
rect 544 1367 555 1405
rect 505 1339 525 1367
rect 544 1339 553 1367
rect 544 1319 548 1339
rect 579 1298 582 1388
rect 612 1370 624 1371
rect 599 1368 649 1370
rect 612 1367 624 1368
rect 610 1360 632 1367
rect 607 1359 632 1360
rect 586 1352 644 1359
rect 607 1351 644 1352
rect 607 1335 610 1351
rect 616 1335 644 1351
rect 607 1334 644 1335
rect 586 1327 644 1334
rect 607 1326 610 1327
rect 612 1319 632 1327
rect 612 1315 624 1319
rect 649 1318 651 1368
rect 544 1281 548 1289
rect 400 1249 408 1279
rect 420 1249 436 1279
rect 400 1245 436 1249
rect 400 1237 430 1245
rect 428 1221 430 1237
rect 476 1209 480 1277
rect 544 1247 552 1281
rect 578 1247 582 1281
rect 544 1239 548 1247
rect 544 1209 586 1210
rect 288 1169 292 1201
rect 296 1199 368 1207
rect 378 1199 450 1207
rect 544 1202 548 1209
rect 439 1171 444 1199
rect 120 1155 170 1157
rect 76 1151 130 1155
rect 110 1146 130 1151
rect 60 1121 67 1131
rect 76 1121 77 1141
rect 96 1112 99 1146
rect 109 1121 110 1141
rect 119 1121 126 1131
rect 76 1105 92 1111
rect 94 1105 110 1111
rect 170 1105 172 1155
rect 186 1089 190 1123
rect 216 1089 220 1123
rect 213 1057 224 1089
rect 282 1085 292 1169
rect 296 1163 368 1171
rect 378 1163 450 1171
rect 468 1168 473 1202
rect 428 1133 430 1149
rect 251 1057 292 1085
rect 318 1064 324 1133
rect 12 1052 62 1054
rect 28 1043 59 1051
rect 62 1043 64 1052
rect 251 1051 263 1057
rect 28 1035 64 1043
rect 127 1043 158 1051
rect 127 1036 182 1043
rect 127 1035 161 1036
rect 59 1019 64 1035
rect 158 1019 161 1035
rect 253 1023 263 1051
rect 273 1023 293 1057
rect 318 1054 335 1064
rect 303 1038 316 1048
rect 318 1038 324 1054
rect 346 1048 348 1133
rect 400 1125 430 1133
rect 476 1131 480 1199
rect 511 1168 582 1202
rect 544 1161 548 1168
rect 400 1121 436 1125
rect 400 1091 408 1121
rect 420 1091 436 1121
rect 544 1123 548 1131
rect 28 1011 64 1019
rect 127 1018 161 1019
rect 127 1011 182 1018
rect 62 1002 64 1011
rect 282 965 292 1023
rect 295 1014 324 1038
rect 333 1038 353 1048
rect 428 1044 430 1091
rect 476 1051 480 1119
rect 544 1089 552 1123
rect 578 1089 582 1123
rect 544 1081 548 1089
rect 367 1038 380 1044
rect 333 1014 380 1038
rect 318 1001 324 1014
rect 346 1001 348 1014
rect 367 1010 380 1014
rect 396 1010 408 1044
rect 420 1010 436 1044
rect 544 1041 553 1069
rect 319 990 346 1001
rect 120 949 170 951
rect 76 943 92 949
rect 94 943 110 949
rect 76 933 99 942
rect 60 923 67 933
rect 76 913 77 933
rect 96 908 99 933
rect 109 913 110 933
rect 119 923 126 933
rect 76 899 110 903
rect 170 899 172 949
rect 186 931 190 965
rect 216 931 220 965
rect 182 893 224 894
rect 186 869 220 886
rect 223 869 257 886
rect 182 852 257 869
rect 182 851 224 852
rect 160 845 246 851
rect 288 845 292 965
rect 296 963 368 971
rect 428 963 430 1010
rect 476 973 480 1041
rect 485 997 495 1031
rect 505 1003 525 1031
rect 505 997 519 1003
rect 544 997 555 1041
rect 485 973 492 997
rect 579 982 582 1072
rect 612 1054 624 1055
rect 599 1052 649 1054
rect 612 1051 624 1052
rect 610 1044 632 1051
rect 607 1043 632 1044
rect 586 1036 644 1043
rect 607 1035 644 1036
rect 607 1019 610 1035
rect 616 1019 644 1035
rect 607 1018 644 1019
rect 586 1011 644 1018
rect 607 1010 610 1011
rect 612 1003 632 1011
rect 612 999 624 1003
rect 649 1002 651 1052
rect 544 965 548 973
rect 400 933 408 963
rect 420 933 436 963
rect 400 929 436 933
rect 400 921 430 929
rect 428 905 430 921
rect 476 893 480 961
rect 544 931 552 965
rect 578 931 582 965
rect 544 923 548 931
rect 295 852 300 886
rect 324 852 329 886
rect 378 883 450 891
rect 544 888 548 893
rect 544 884 582 888
rect 544 869 552 884
rect 578 869 582 884
rect 544 851 586 869
rect 522 845 608 851
rect 182 829 224 845
rect 544 829 586 845
rect 17 815 67 817
rect 119 815 169 817
rect 186 815 220 829
rect 548 815 582 829
rect 599 815 649 817
rect 42 773 59 807
rect 67 765 69 815
rect 160 807 246 815
rect 522 807 608 815
rect 76 773 110 807
rect 127 773 144 807
rect 152 773 161 807
rect 162 805 195 807
rect 224 805 244 807
rect 162 773 244 805
rect 524 805 548 807
rect 573 805 582 807
rect 586 805 606 807
rect 160 765 246 773
rect 186 749 220 765
rect 182 735 224 736
rect 160 729 182 735
rect 224 729 246 735
rect 186 694 220 728
rect 223 694 257 728
rect 120 681 170 683
rect 76 677 130 681
rect 110 672 130 677
rect 60 647 67 657
rect 76 647 77 667
rect 96 638 99 672
rect 109 647 110 667
rect 119 647 126 657
rect 76 631 92 637
rect 94 631 110 637
rect 170 631 172 681
rect 186 615 190 649
rect 216 615 220 649
rect 288 615 292 803
rect 476 735 480 803
rect 524 773 606 805
rect 607 773 616 807
rect 522 765 608 773
rect 649 765 651 815
rect 548 749 582 765
rect 522 730 548 735
rect 522 729 582 730
rect 586 729 608 735
rect 295 694 300 728
rect 324 694 329 728
rect 544 726 582 729
rect 378 689 450 697
rect 428 659 430 675
rect 400 651 430 659
rect 476 657 480 725
rect 544 696 552 726
rect 578 696 582 726
rect 544 687 548 696
rect 400 647 436 651
rect 400 617 408 647
rect 420 617 436 647
rect 544 649 548 657
rect 12 578 62 580
rect 28 569 59 577
rect 62 569 64 578
rect 28 561 64 569
rect 127 569 158 577
rect 127 562 182 569
rect 215 567 224 595
rect 127 561 161 562
rect 59 545 64 561
rect 158 545 161 561
rect 28 537 64 545
rect 127 544 161 545
rect 127 537 182 544
rect 62 528 64 537
rect 213 529 224 567
rect 282 557 292 615
rect 296 609 368 617
rect 319 579 346 590
rect 318 566 324 579
rect 346 566 348 579
rect 428 570 430 617
rect 443 607 450 609
rect 476 577 480 645
rect 544 615 552 649
rect 578 615 582 649
rect 481 583 517 611
rect 481 577 495 583
rect 367 566 380 570
rect 251 523 263 557
rect 273 523 293 557
rect 295 542 324 566
rect 303 532 316 542
rect 318 526 324 542
rect 333 542 380 566
rect 333 532 353 542
rect 367 536 380 542
rect 396 536 408 570
rect 420 536 436 570
rect 120 475 170 477
rect 76 469 92 475
rect 94 469 110 475
rect 76 459 99 468
rect 60 449 67 459
rect 76 439 77 459
rect 96 434 99 459
rect 109 439 110 459
rect 119 449 126 459
rect 76 425 110 429
rect 170 425 172 475
rect 186 457 190 491
rect 216 457 220 491
rect 186 411 220 429
rect 282 411 292 523
rect 318 516 335 526
rect 318 447 324 516
rect 346 447 348 532
rect 428 489 430 536
rect 476 499 480 567
rect 485 549 495 577
rect 505 577 519 583
rect 544 577 555 615
rect 505 549 525 577
rect 544 549 553 577
rect 544 529 548 549
rect 579 508 582 598
rect 612 580 624 581
rect 599 578 649 580
rect 612 577 624 578
rect 610 570 632 577
rect 607 569 632 570
rect 586 562 644 569
rect 607 561 644 562
rect 607 545 610 561
rect 616 545 644 561
rect 607 544 644 545
rect 586 537 644 544
rect 607 536 610 537
rect 612 529 632 537
rect 612 525 624 529
rect 649 528 651 578
rect 544 491 548 499
rect 400 459 408 489
rect 420 459 436 489
rect 400 455 436 459
rect 400 447 430 455
rect 428 431 430 447
rect 476 419 480 487
rect 544 457 552 491
rect 578 457 582 491
rect 544 449 548 457
rect 548 420 582 429
rect 544 419 586 420
rect 170 410 236 411
rect 186 403 190 410
rect 216 403 220 410
rect 186 395 220 403
rect 288 395 292 411
rect 296 409 368 417
rect 378 409 450 417
rect 544 412 582 419
rect 182 369 224 395
rect 439 378 444 409
rect 468 378 473 412
rect 511 395 582 412
rect 511 378 586 395
rect 544 369 586 378
<< metal1 >>
rect 222 0 258 102700
rect 294 0 330 102700
rect 366 101989 402 102330
rect 366 101199 402 101831
rect 366 100409 402 101041
rect 366 99619 402 100251
rect 366 98829 402 99461
rect 366 98039 402 98671
rect 366 97249 402 97881
rect 366 96459 402 97091
rect 366 95669 402 96301
rect 366 94879 402 95511
rect 366 94089 402 94721
rect 366 93299 402 93931
rect 366 92509 402 93141
rect 366 91719 402 92351
rect 366 90929 402 91561
rect 366 90139 402 90771
rect 366 89349 402 89981
rect 366 88559 402 89191
rect 366 87769 402 88401
rect 366 86979 402 87611
rect 366 86189 402 86821
rect 366 85399 402 86031
rect 366 84609 402 85241
rect 366 83819 402 84451
rect 366 83029 402 83661
rect 366 82239 402 82871
rect 366 81449 402 82081
rect 366 80659 402 81291
rect 366 79869 402 80501
rect 366 79079 402 79711
rect 366 78289 402 78921
rect 366 77499 402 78131
rect 366 76709 402 77341
rect 366 75919 402 76551
rect 366 75129 402 75761
rect 366 74339 402 74971
rect 366 73549 402 74181
rect 366 72759 402 73391
rect 366 71969 402 72601
rect 366 71179 402 71811
rect 366 70389 402 71021
rect 366 69599 402 70231
rect 366 68809 402 69441
rect 366 68019 402 68651
rect 366 67229 402 67861
rect 366 66439 402 67071
rect 366 65649 402 66281
rect 366 64859 402 65491
rect 366 64069 402 64701
rect 366 63279 402 63911
rect 366 62489 402 63121
rect 366 61699 402 62331
rect 366 60909 402 61541
rect 366 60119 402 60751
rect 366 59329 402 59961
rect 366 58539 402 59171
rect 366 57749 402 58381
rect 366 56959 402 57591
rect 366 56169 402 56801
rect 366 55379 402 56011
rect 366 54589 402 55221
rect 366 53799 402 54431
rect 366 53009 402 53641
rect 366 52219 402 52851
rect 366 51429 402 52061
rect 366 50639 402 51271
rect 366 49849 402 50481
rect 366 49059 402 49691
rect 366 48269 402 48901
rect 366 47479 402 48111
rect 366 46689 402 47321
rect 366 45899 402 46531
rect 366 45109 402 45741
rect 366 44319 402 44951
rect 366 43529 402 44161
rect 366 42739 402 43371
rect 366 41949 402 42581
rect 366 41159 402 41791
rect 366 40369 402 41001
rect 366 39579 402 40211
rect 366 38789 402 39421
rect 366 37999 402 38631
rect 366 37209 402 37841
rect 366 36419 402 37051
rect 366 35629 402 36261
rect 366 34839 402 35471
rect 366 34049 402 34681
rect 366 33259 402 33891
rect 366 32469 402 33101
rect 366 31679 402 32311
rect 366 30889 402 31521
rect 366 30099 402 30731
rect 366 29309 402 29941
rect 366 28519 402 29151
rect 366 27729 402 28361
rect 366 26939 402 27571
rect 366 26149 402 26781
rect 366 25359 402 25991
rect 366 24569 402 25201
rect 366 23779 402 24411
rect 366 22989 402 23621
rect 366 22199 402 22831
rect 366 21409 402 22041
rect 366 20619 402 21251
rect 366 19829 402 20461
rect 366 19039 402 19671
rect 366 18249 402 18881
rect 366 17459 402 18091
rect 366 16669 402 17301
rect 366 15879 402 16511
rect 366 15089 402 15721
rect 366 14299 402 14931
rect 366 13509 402 14141
rect 366 12719 402 13351
rect 366 11929 402 12561
rect 366 11139 402 11771
rect 366 10349 402 10981
rect 366 9559 402 10191
rect 366 8769 402 9401
rect 366 7979 402 8611
rect 366 7189 402 7821
rect 366 6399 402 7031
rect 366 5609 402 6241
rect 366 4819 402 5451
rect 366 4029 402 4661
rect 366 3239 402 3871
rect 366 2449 402 3081
rect 366 1659 402 2291
rect 366 869 402 1501
rect 366 370 402 711
rect 438 0 474 102700
rect 510 0 546 102700
<< metal2 >>
rect 0 102233 624 102281
rect 330 102109 438 102185
rect 0 102013 624 102061
rect 330 101855 438 101965
rect 0 101759 624 101807
rect 330 101635 438 101711
rect 0 101539 624 101587
rect 0 101443 624 101491
rect 330 101319 438 101395
rect 0 101223 624 101271
rect 330 101065 438 101175
rect 0 100969 624 101017
rect 330 100845 438 100921
rect 0 100749 624 100797
rect 0 100653 624 100701
rect 330 100529 438 100605
rect 0 100433 624 100481
rect 330 100275 438 100385
rect 0 100179 624 100227
rect 330 100055 438 100131
rect 0 99959 624 100007
rect 0 99863 624 99911
rect 330 99739 438 99815
rect 0 99643 624 99691
rect 330 99485 438 99595
rect 0 99389 624 99437
rect 330 99265 438 99341
rect 0 99169 624 99217
rect 0 99073 624 99121
rect 330 98949 438 99025
rect 0 98853 624 98901
rect 330 98695 438 98805
rect 0 98599 624 98647
rect 330 98475 438 98551
rect 0 98379 624 98427
rect 0 98283 624 98331
rect 330 98159 438 98235
rect 0 98063 624 98111
rect 330 97905 438 98015
rect 0 97809 624 97857
rect 330 97685 438 97761
rect 0 97589 624 97637
rect 0 97493 624 97541
rect 330 97369 438 97445
rect 0 97273 624 97321
rect 330 97115 438 97225
rect 0 97019 624 97067
rect 330 96895 438 96971
rect 0 96799 624 96847
rect 0 96703 624 96751
rect 330 96579 438 96655
rect 0 96483 624 96531
rect 330 96325 438 96435
rect 0 96229 624 96277
rect 330 96105 438 96181
rect 0 96009 624 96057
rect 0 95913 624 95961
rect 330 95789 438 95865
rect 0 95693 624 95741
rect 330 95535 438 95645
rect 0 95439 624 95487
rect 330 95315 438 95391
rect 0 95219 624 95267
rect 0 95123 624 95171
rect 330 94999 438 95075
rect 0 94903 624 94951
rect 330 94745 438 94855
rect 0 94649 624 94697
rect 330 94525 438 94601
rect 0 94429 624 94477
rect 0 94333 624 94381
rect 330 94209 438 94285
rect 0 94113 624 94161
rect 330 93955 438 94065
rect 0 93859 624 93907
rect 330 93735 438 93811
rect 0 93639 624 93687
rect 0 93543 624 93591
rect 330 93419 438 93495
rect 0 93323 624 93371
rect 330 93165 438 93275
rect 0 93069 624 93117
rect 330 92945 438 93021
rect 0 92849 624 92897
rect 0 92753 624 92801
rect 330 92629 438 92705
rect 0 92533 624 92581
rect 330 92375 438 92485
rect 0 92279 624 92327
rect 330 92155 438 92231
rect 0 92059 624 92107
rect 0 91963 624 92011
rect 330 91839 438 91915
rect 0 91743 624 91791
rect 330 91585 438 91695
rect 0 91489 624 91537
rect 330 91365 438 91441
rect 0 91269 624 91317
rect 0 91173 624 91221
rect 330 91049 438 91125
rect 0 90953 624 91001
rect 330 90795 438 90905
rect 0 90699 624 90747
rect 330 90575 438 90651
rect 0 90479 624 90527
rect 0 90383 624 90431
rect 330 90259 438 90335
rect 0 90163 624 90211
rect 330 90005 438 90115
rect 0 89909 624 89957
rect 330 89785 438 89861
rect 0 89689 624 89737
rect 0 89593 624 89641
rect 330 89469 438 89545
rect 0 89373 624 89421
rect 330 89215 438 89325
rect 0 89119 624 89167
rect 330 88995 438 89071
rect 0 88899 624 88947
rect 0 88803 624 88851
rect 330 88679 438 88755
rect 0 88583 624 88631
rect 330 88425 438 88535
rect 0 88329 624 88377
rect 330 88205 438 88281
rect 0 88109 624 88157
rect 0 88013 624 88061
rect 330 87889 438 87965
rect 0 87793 624 87841
rect 330 87635 438 87745
rect 0 87539 624 87587
rect 330 87415 438 87491
rect 0 87319 624 87367
rect 0 87223 624 87271
rect 330 87099 438 87175
rect 0 87003 624 87051
rect 330 86845 438 86955
rect 0 86749 624 86797
rect 330 86625 438 86701
rect 0 86529 624 86577
rect 0 86433 624 86481
rect 330 86309 438 86385
rect 0 86213 624 86261
rect 330 86055 438 86165
rect 0 85959 624 86007
rect 330 85835 438 85911
rect 0 85739 624 85787
rect 0 85643 624 85691
rect 330 85519 438 85595
rect 0 85423 624 85471
rect 330 85265 438 85375
rect 0 85169 624 85217
rect 330 85045 438 85121
rect 0 84949 624 84997
rect 0 84853 624 84901
rect 330 84729 438 84805
rect 0 84633 624 84681
rect 330 84475 438 84585
rect 0 84379 624 84427
rect 330 84255 438 84331
rect 0 84159 624 84207
rect 0 84063 624 84111
rect 330 83939 438 84015
rect 0 83843 624 83891
rect 330 83685 438 83795
rect 0 83589 624 83637
rect 330 83465 438 83541
rect 0 83369 624 83417
rect 0 83273 624 83321
rect 330 83149 438 83225
rect 0 83053 624 83101
rect 330 82895 438 83005
rect 0 82799 624 82847
rect 330 82675 438 82751
rect 0 82579 624 82627
rect 0 82483 624 82531
rect 330 82359 438 82435
rect 0 82263 624 82311
rect 330 82105 438 82215
rect 0 82009 624 82057
rect 330 81885 438 81961
rect 0 81789 624 81837
rect 0 81693 624 81741
rect 330 81569 438 81645
rect 0 81473 624 81521
rect 330 81315 438 81425
rect 0 81219 624 81267
rect 330 81095 438 81171
rect 0 80999 624 81047
rect 0 80903 624 80951
rect 330 80779 438 80855
rect 0 80683 624 80731
rect 330 80525 438 80635
rect 0 80429 624 80477
rect 330 80305 438 80381
rect 0 80209 624 80257
rect 0 80113 624 80161
rect 330 79989 438 80065
rect 0 79893 624 79941
rect 330 79735 438 79845
rect 0 79639 624 79687
rect 330 79515 438 79591
rect 0 79419 624 79467
rect 0 79323 624 79371
rect 330 79199 438 79275
rect 0 79103 624 79151
rect 330 78945 438 79055
rect 0 78849 624 78897
rect 330 78725 438 78801
rect 0 78629 624 78677
rect 0 78533 624 78581
rect 330 78409 438 78485
rect 0 78313 624 78361
rect 330 78155 438 78265
rect 0 78059 624 78107
rect 330 77935 438 78011
rect 0 77839 624 77887
rect 0 77743 624 77791
rect 330 77619 438 77695
rect 0 77523 624 77571
rect 330 77365 438 77475
rect 0 77269 624 77317
rect 330 77145 438 77221
rect 0 77049 624 77097
rect 0 76953 624 77001
rect 330 76829 438 76905
rect 0 76733 624 76781
rect 330 76575 438 76685
rect 0 76479 624 76527
rect 330 76355 438 76431
rect 0 76259 624 76307
rect 0 76163 624 76211
rect 330 76039 438 76115
rect 0 75943 624 75991
rect 330 75785 438 75895
rect 0 75689 624 75737
rect 330 75565 438 75641
rect 0 75469 624 75517
rect 0 75373 624 75421
rect 330 75249 438 75325
rect 0 75153 624 75201
rect 330 74995 438 75105
rect 0 74899 624 74947
rect 330 74775 438 74851
rect 0 74679 624 74727
rect 0 74583 624 74631
rect 330 74459 438 74535
rect 0 74363 624 74411
rect 330 74205 438 74315
rect 0 74109 624 74157
rect 330 73985 438 74061
rect 0 73889 624 73937
rect 0 73793 624 73841
rect 330 73669 438 73745
rect 0 73573 624 73621
rect 330 73415 438 73525
rect 0 73319 624 73367
rect 330 73195 438 73271
rect 0 73099 624 73147
rect 0 73003 624 73051
rect 330 72879 438 72955
rect 0 72783 624 72831
rect 330 72625 438 72735
rect 0 72529 624 72577
rect 330 72405 438 72481
rect 0 72309 624 72357
rect 0 72213 624 72261
rect 330 72089 438 72165
rect 0 71993 624 72041
rect 330 71835 438 71945
rect 0 71739 624 71787
rect 330 71615 438 71691
rect 0 71519 624 71567
rect 0 71423 624 71471
rect 330 71299 438 71375
rect 0 71203 624 71251
rect 330 71045 438 71155
rect 0 70949 624 70997
rect 330 70825 438 70901
rect 0 70729 624 70777
rect 0 70633 624 70681
rect 330 70509 438 70585
rect 0 70413 624 70461
rect 330 70255 438 70365
rect 0 70159 624 70207
rect 330 70035 438 70111
rect 0 69939 624 69987
rect 0 69843 624 69891
rect 330 69719 438 69795
rect 0 69623 624 69671
rect 330 69465 438 69575
rect 0 69369 624 69417
rect 330 69245 438 69321
rect 0 69149 624 69197
rect 0 69053 624 69101
rect 330 68929 438 69005
rect 0 68833 624 68881
rect 330 68675 438 68785
rect 0 68579 624 68627
rect 330 68455 438 68531
rect 0 68359 624 68407
rect 0 68263 624 68311
rect 330 68139 438 68215
rect 0 68043 624 68091
rect 330 67885 438 67995
rect 0 67789 624 67837
rect 330 67665 438 67741
rect 0 67569 624 67617
rect 0 67473 624 67521
rect 330 67349 438 67425
rect 0 67253 624 67301
rect 330 67095 438 67205
rect 0 66999 624 67047
rect 330 66875 438 66951
rect 0 66779 624 66827
rect 0 66683 624 66731
rect 330 66559 438 66635
rect 0 66463 624 66511
rect 330 66305 438 66415
rect 0 66209 624 66257
rect 330 66085 438 66161
rect 0 65989 624 66037
rect 0 65893 624 65941
rect 330 65769 438 65845
rect 0 65673 624 65721
rect 330 65515 438 65625
rect 0 65419 624 65467
rect 330 65295 438 65371
rect 0 65199 624 65247
rect 0 65103 624 65151
rect 330 64979 438 65055
rect 0 64883 624 64931
rect 330 64725 438 64835
rect 0 64629 624 64677
rect 330 64505 438 64581
rect 0 64409 624 64457
rect 0 64313 624 64361
rect 330 64189 438 64265
rect 0 64093 624 64141
rect 330 63935 438 64045
rect 0 63839 624 63887
rect 330 63715 438 63791
rect 0 63619 624 63667
rect 0 63523 624 63571
rect 330 63399 438 63475
rect 0 63303 624 63351
rect 330 63145 438 63255
rect 0 63049 624 63097
rect 330 62925 438 63001
rect 0 62829 624 62877
rect 0 62733 624 62781
rect 330 62609 438 62685
rect 0 62513 624 62561
rect 330 62355 438 62465
rect 0 62259 624 62307
rect 330 62135 438 62211
rect 0 62039 624 62087
rect 0 61943 624 61991
rect 330 61819 438 61895
rect 0 61723 624 61771
rect 330 61565 438 61675
rect 0 61469 624 61517
rect 330 61345 438 61421
rect 0 61249 624 61297
rect 0 61153 624 61201
rect 330 61029 438 61105
rect 0 60933 624 60981
rect 330 60775 438 60885
rect 0 60679 624 60727
rect 330 60555 438 60631
rect 0 60459 624 60507
rect 0 60363 624 60411
rect 330 60239 438 60315
rect 0 60143 624 60191
rect 330 59985 438 60095
rect 0 59889 624 59937
rect 330 59765 438 59841
rect 0 59669 624 59717
rect 0 59573 624 59621
rect 330 59449 438 59525
rect 0 59353 624 59401
rect 330 59195 438 59305
rect 0 59099 624 59147
rect 330 58975 438 59051
rect 0 58879 624 58927
rect 0 58783 624 58831
rect 330 58659 438 58735
rect 0 58563 624 58611
rect 330 58405 438 58515
rect 0 58309 624 58357
rect 330 58185 438 58261
rect 0 58089 624 58137
rect 0 57993 624 58041
rect 330 57869 438 57945
rect 0 57773 624 57821
rect 330 57615 438 57725
rect 0 57519 624 57567
rect 330 57395 438 57471
rect 0 57299 624 57347
rect 0 57203 624 57251
rect 330 57079 438 57155
rect 0 56983 624 57031
rect 330 56825 438 56935
rect 0 56729 624 56777
rect 330 56605 438 56681
rect 0 56509 624 56557
rect 0 56413 624 56461
rect 330 56289 438 56365
rect 0 56193 624 56241
rect 330 56035 438 56145
rect 0 55939 624 55987
rect 330 55815 438 55891
rect 0 55719 624 55767
rect 0 55623 624 55671
rect 330 55499 438 55575
rect 0 55403 624 55451
rect 330 55245 438 55355
rect 0 55149 624 55197
rect 330 55025 438 55101
rect 0 54929 624 54977
rect 0 54833 624 54881
rect 330 54709 438 54785
rect 0 54613 624 54661
rect 330 54455 438 54565
rect 0 54359 624 54407
rect 330 54235 438 54311
rect 0 54139 624 54187
rect 0 54043 624 54091
rect 330 53919 438 53995
rect 0 53823 624 53871
rect 330 53665 438 53775
rect 0 53569 624 53617
rect 330 53445 438 53521
rect 0 53349 624 53397
rect 0 53253 624 53301
rect 330 53129 438 53205
rect 0 53033 624 53081
rect 330 52875 438 52985
rect 0 52779 624 52827
rect 330 52655 438 52731
rect 0 52559 624 52607
rect 0 52463 624 52511
rect 330 52339 438 52415
rect 0 52243 624 52291
rect 330 52085 438 52195
rect 0 51989 624 52037
rect 330 51865 438 51941
rect 0 51769 624 51817
rect 0 51673 624 51721
rect 330 51549 438 51625
rect 0 51453 624 51501
rect 330 51295 438 51405
rect 0 51199 624 51247
rect 330 51075 438 51151
rect 0 50979 624 51027
rect 0 50883 624 50931
rect 330 50759 438 50835
rect 0 50663 624 50711
rect 330 50505 438 50615
rect 0 50409 624 50457
rect 330 50285 438 50361
rect 0 50189 624 50237
rect 0 50093 624 50141
rect 330 49969 438 50045
rect 0 49873 624 49921
rect 330 49715 438 49825
rect 0 49619 624 49667
rect 330 49495 438 49571
rect 0 49399 624 49447
rect 0 49303 624 49351
rect 330 49179 438 49255
rect 0 49083 624 49131
rect 330 48925 438 49035
rect 0 48829 624 48877
rect 330 48705 438 48781
rect 0 48609 624 48657
rect 0 48513 624 48561
rect 330 48389 438 48465
rect 0 48293 624 48341
rect 330 48135 438 48245
rect 0 48039 624 48087
rect 330 47915 438 47991
rect 0 47819 624 47867
rect 0 47723 624 47771
rect 330 47599 438 47675
rect 0 47503 624 47551
rect 330 47345 438 47455
rect 0 47249 624 47297
rect 330 47125 438 47201
rect 0 47029 624 47077
rect 0 46933 624 46981
rect 330 46809 438 46885
rect 0 46713 624 46761
rect 330 46555 438 46665
rect 0 46459 624 46507
rect 330 46335 438 46411
rect 0 46239 624 46287
rect 0 46143 624 46191
rect 330 46019 438 46095
rect 0 45923 624 45971
rect 330 45765 438 45875
rect 0 45669 624 45717
rect 330 45545 438 45621
rect 0 45449 624 45497
rect 0 45353 624 45401
rect 330 45229 438 45305
rect 0 45133 624 45181
rect 330 44975 438 45085
rect 0 44879 624 44927
rect 330 44755 438 44831
rect 0 44659 624 44707
rect 0 44563 624 44611
rect 330 44439 438 44515
rect 0 44343 624 44391
rect 330 44185 438 44295
rect 0 44089 624 44137
rect 330 43965 438 44041
rect 0 43869 624 43917
rect 0 43773 624 43821
rect 330 43649 438 43725
rect 0 43553 624 43601
rect 330 43395 438 43505
rect 0 43299 624 43347
rect 330 43175 438 43251
rect 0 43079 624 43127
rect 0 42983 624 43031
rect 330 42859 438 42935
rect 0 42763 624 42811
rect 330 42605 438 42715
rect 0 42509 624 42557
rect 330 42385 438 42461
rect 0 42289 624 42337
rect 0 42193 624 42241
rect 330 42069 438 42145
rect 0 41973 624 42021
rect 330 41815 438 41925
rect 0 41719 624 41767
rect 330 41595 438 41671
rect 0 41499 624 41547
rect 0 41403 624 41451
rect 330 41279 438 41355
rect 0 41183 624 41231
rect 330 41025 438 41135
rect 0 40929 624 40977
rect 330 40805 438 40881
rect 0 40709 624 40757
rect 0 40613 624 40661
rect 330 40489 438 40565
rect 0 40393 624 40441
rect 330 40235 438 40345
rect 0 40139 624 40187
rect 330 40015 438 40091
rect 0 39919 624 39967
rect 0 39823 624 39871
rect 330 39699 438 39775
rect 0 39603 624 39651
rect 330 39445 438 39555
rect 0 39349 624 39397
rect 330 39225 438 39301
rect 0 39129 624 39177
rect 0 39033 624 39081
rect 330 38909 438 38985
rect 0 38813 624 38861
rect 330 38655 438 38765
rect 0 38559 624 38607
rect 330 38435 438 38511
rect 0 38339 624 38387
rect 0 38243 624 38291
rect 330 38119 438 38195
rect 0 38023 624 38071
rect 330 37865 438 37975
rect 0 37769 624 37817
rect 330 37645 438 37721
rect 0 37549 624 37597
rect 0 37453 624 37501
rect 330 37329 438 37405
rect 0 37233 624 37281
rect 330 37075 438 37185
rect 0 36979 624 37027
rect 330 36855 438 36931
rect 0 36759 624 36807
rect 0 36663 624 36711
rect 330 36539 438 36615
rect 0 36443 624 36491
rect 330 36285 438 36395
rect 0 36189 624 36237
rect 330 36065 438 36141
rect 0 35969 624 36017
rect 0 35873 624 35921
rect 330 35749 438 35825
rect 0 35653 624 35701
rect 330 35495 438 35605
rect 0 35399 624 35447
rect 330 35275 438 35351
rect 0 35179 624 35227
rect 0 35083 624 35131
rect 330 34959 438 35035
rect 0 34863 624 34911
rect 330 34705 438 34815
rect 0 34609 624 34657
rect 330 34485 438 34561
rect 0 34389 624 34437
rect 0 34293 624 34341
rect 330 34169 438 34245
rect 0 34073 624 34121
rect 330 33915 438 34025
rect 0 33819 624 33867
rect 330 33695 438 33771
rect 0 33599 624 33647
rect 0 33503 624 33551
rect 330 33379 438 33455
rect 0 33283 624 33331
rect 330 33125 438 33235
rect 0 33029 624 33077
rect 330 32905 438 32981
rect 0 32809 624 32857
rect 0 32713 624 32761
rect 330 32589 438 32665
rect 0 32493 624 32541
rect 330 32335 438 32445
rect 0 32239 624 32287
rect 330 32115 438 32191
rect 0 32019 624 32067
rect 0 31923 624 31971
rect 330 31799 438 31875
rect 0 31703 624 31751
rect 330 31545 438 31655
rect 0 31449 624 31497
rect 330 31325 438 31401
rect 0 31229 624 31277
rect 0 31133 624 31181
rect 330 31009 438 31085
rect 0 30913 624 30961
rect 330 30755 438 30865
rect 0 30659 624 30707
rect 330 30535 438 30611
rect 0 30439 624 30487
rect 0 30343 624 30391
rect 330 30219 438 30295
rect 0 30123 624 30171
rect 330 29965 438 30075
rect 0 29869 624 29917
rect 330 29745 438 29821
rect 0 29649 624 29697
rect 0 29553 624 29601
rect 330 29429 438 29505
rect 0 29333 624 29381
rect 330 29175 438 29285
rect 0 29079 624 29127
rect 330 28955 438 29031
rect 0 28859 624 28907
rect 0 28763 624 28811
rect 330 28639 438 28715
rect 0 28543 624 28591
rect 330 28385 438 28495
rect 0 28289 624 28337
rect 330 28165 438 28241
rect 0 28069 624 28117
rect 0 27973 624 28021
rect 330 27849 438 27925
rect 0 27753 624 27801
rect 330 27595 438 27705
rect 0 27499 624 27547
rect 330 27375 438 27451
rect 0 27279 624 27327
rect 0 27183 624 27231
rect 330 27059 438 27135
rect 0 26963 624 27011
rect 330 26805 438 26915
rect 0 26709 624 26757
rect 330 26585 438 26661
rect 0 26489 624 26537
rect 0 26393 624 26441
rect 330 26269 438 26345
rect 0 26173 624 26221
rect 330 26015 438 26125
rect 0 25919 624 25967
rect 330 25795 438 25871
rect 0 25699 624 25747
rect 0 25603 624 25651
rect 330 25479 438 25555
rect 0 25383 624 25431
rect 330 25225 438 25335
rect 0 25129 624 25177
rect 330 25005 438 25081
rect 0 24909 624 24957
rect 0 24813 624 24861
rect 330 24689 438 24765
rect 0 24593 624 24641
rect 330 24435 438 24545
rect 0 24339 624 24387
rect 330 24215 438 24291
rect 0 24119 624 24167
rect 0 24023 624 24071
rect 330 23899 438 23975
rect 0 23803 624 23851
rect 330 23645 438 23755
rect 0 23549 624 23597
rect 330 23425 438 23501
rect 0 23329 624 23377
rect 0 23233 624 23281
rect 330 23109 438 23185
rect 0 23013 624 23061
rect 330 22855 438 22965
rect 0 22759 624 22807
rect 330 22635 438 22711
rect 0 22539 624 22587
rect 0 22443 624 22491
rect 330 22319 438 22395
rect 0 22223 624 22271
rect 330 22065 438 22175
rect 0 21969 624 22017
rect 330 21845 438 21921
rect 0 21749 624 21797
rect 0 21653 624 21701
rect 330 21529 438 21605
rect 0 21433 624 21481
rect 330 21275 438 21385
rect 0 21179 624 21227
rect 330 21055 438 21131
rect 0 20959 624 21007
rect 0 20863 624 20911
rect 330 20739 438 20815
rect 0 20643 624 20691
rect 330 20485 438 20595
rect 0 20389 624 20437
rect 330 20265 438 20341
rect 0 20169 624 20217
rect 0 20073 624 20121
rect 330 19949 438 20025
rect 0 19853 624 19901
rect 330 19695 438 19805
rect 0 19599 624 19647
rect 330 19475 438 19551
rect 0 19379 624 19427
rect 0 19283 624 19331
rect 330 19159 438 19235
rect 0 19063 624 19111
rect 330 18905 438 19015
rect 0 18809 624 18857
rect 330 18685 438 18761
rect 0 18589 624 18637
rect 0 18493 624 18541
rect 330 18369 438 18445
rect 0 18273 624 18321
rect 330 18115 438 18225
rect 0 18019 624 18067
rect 330 17895 438 17971
rect 0 17799 624 17847
rect 0 17703 624 17751
rect 330 17579 438 17655
rect 0 17483 624 17531
rect 330 17325 438 17435
rect 0 17229 624 17277
rect 330 17105 438 17181
rect 0 17009 624 17057
rect 0 16913 624 16961
rect 330 16789 438 16865
rect 0 16693 624 16741
rect 330 16535 438 16645
rect 0 16439 624 16487
rect 330 16315 438 16391
rect 0 16219 624 16267
rect 0 16123 624 16171
rect 330 15999 438 16075
rect 0 15903 624 15951
rect 330 15745 438 15855
rect 0 15649 624 15697
rect 330 15525 438 15601
rect 0 15429 624 15477
rect 0 15333 624 15381
rect 330 15209 438 15285
rect 0 15113 624 15161
rect 330 14955 438 15065
rect 0 14859 624 14907
rect 330 14735 438 14811
rect 0 14639 624 14687
rect 0 14543 624 14591
rect 330 14419 438 14495
rect 0 14323 624 14371
rect 330 14165 438 14275
rect 0 14069 624 14117
rect 330 13945 438 14021
rect 0 13849 624 13897
rect 0 13753 624 13801
rect 330 13629 438 13705
rect 0 13533 624 13581
rect 330 13375 438 13485
rect 0 13279 624 13327
rect 330 13155 438 13231
rect 0 13059 624 13107
rect 0 12963 624 13011
rect 330 12839 438 12915
rect 0 12743 624 12791
rect 330 12585 438 12695
rect 0 12489 624 12537
rect 330 12365 438 12441
rect 0 12269 624 12317
rect 0 12173 624 12221
rect 330 12049 438 12125
rect 0 11953 624 12001
rect 330 11795 438 11905
rect 0 11699 624 11747
rect 330 11575 438 11651
rect 0 11479 624 11527
rect 0 11383 624 11431
rect 330 11259 438 11335
rect 0 11163 624 11211
rect 330 11005 438 11115
rect 0 10909 624 10957
rect 330 10785 438 10861
rect 0 10689 624 10737
rect 0 10593 624 10641
rect 330 10469 438 10545
rect 0 10373 624 10421
rect 330 10215 438 10325
rect 0 10119 624 10167
rect 330 9995 438 10071
rect 0 9899 624 9947
rect 0 9803 624 9851
rect 330 9679 438 9755
rect 0 9583 624 9631
rect 330 9425 438 9535
rect 0 9329 624 9377
rect 330 9205 438 9281
rect 0 9109 624 9157
rect 0 9013 624 9061
rect 330 8889 438 8965
rect 0 8793 624 8841
rect 330 8635 438 8745
rect 0 8539 624 8587
rect 330 8415 438 8491
rect 0 8319 624 8367
rect 0 8223 624 8271
rect 330 8099 438 8175
rect 0 8003 624 8051
rect 330 7845 438 7955
rect 0 7749 624 7797
rect 330 7625 438 7701
rect 0 7529 624 7577
rect 0 7433 624 7481
rect 330 7309 438 7385
rect 0 7213 624 7261
rect 330 7055 438 7165
rect 0 6959 624 7007
rect 330 6835 438 6911
rect 0 6739 624 6787
rect 0 6643 624 6691
rect 330 6519 438 6595
rect 0 6423 624 6471
rect 330 6265 438 6375
rect 0 6169 624 6217
rect 330 6045 438 6121
rect 0 5949 624 5997
rect 0 5853 624 5901
rect 330 5729 438 5805
rect 0 5633 624 5681
rect 330 5475 438 5585
rect 0 5379 624 5427
rect 330 5255 438 5331
rect 0 5159 624 5207
rect 0 5063 624 5111
rect 330 4939 438 5015
rect 0 4843 624 4891
rect 330 4685 438 4795
rect 0 4589 624 4637
rect 330 4465 438 4541
rect 0 4369 624 4417
rect 0 4273 624 4321
rect 330 4149 438 4225
rect 0 4053 624 4101
rect 330 3895 438 4005
rect 0 3799 624 3847
rect 330 3675 438 3751
rect 0 3579 624 3627
rect 0 3483 624 3531
rect 330 3359 438 3435
rect 0 3263 624 3311
rect 330 3105 438 3215
rect 0 3009 624 3057
rect 330 2885 438 2961
rect 0 2789 624 2837
rect 0 2693 624 2741
rect 330 2569 438 2645
rect 0 2473 624 2521
rect 330 2315 438 2425
rect 0 2219 624 2267
rect 330 2095 438 2171
rect 0 1999 624 2047
rect 0 1903 624 1951
rect 330 1779 438 1855
rect 0 1683 624 1731
rect 330 1525 438 1635
rect 0 1429 624 1477
rect 330 1305 438 1381
rect 0 1209 624 1257
rect 0 1113 624 1161
rect 330 989 438 1065
rect 0 893 624 941
rect 330 735 438 845
rect 0 639 624 687
rect 330 515 438 591
rect 0 419 624 467
<< metal3 >>
rect 263 102422 361 102520
rect 263 180 361 278
use contact_9  contact_9_1
timestamp 1624494425
transform 1 0 279 0 1 192
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_1
timestamp 1624494425
transform -1 0 624 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_0
timestamp 1624494425
transform -1 0 624 0 -1 102700
box 0 0 624 474
use contact_9  contact_9_0
timestamp 1624494425
transform 1 0 279 0 1 102434
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_0
timestamp 1624494425
transform -1 0 624 0 1 101910
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_256
timestamp 1624494425
transform -1 0 624 0 -1 790
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_255
timestamp 1624494425
transform -1 0 624 0 1 790
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_254
timestamp 1624494425
transform -1 0 624 0 -1 1580
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_253
timestamp 1624494425
transform -1 0 624 0 1 1580
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_252
timestamp 1624494425
transform -1 0 624 0 -1 2370
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_251
timestamp 1624494425
transform -1 0 624 0 1 2370
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_250
timestamp 1624494425
transform -1 0 624 0 -1 3160
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_249
timestamp 1624494425
transform -1 0 624 0 1 3160
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_248
timestamp 1624494425
transform -1 0 624 0 -1 3950
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_247
timestamp 1624494425
transform -1 0 624 0 1 3950
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_246
timestamp 1624494425
transform -1 0 624 0 -1 4740
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_245
timestamp 1624494425
transform -1 0 624 0 1 4740
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_244
timestamp 1624494425
transform -1 0 624 0 -1 5530
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_243
timestamp 1624494425
transform -1 0 624 0 1 5530
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_242
timestamp 1624494425
transform -1 0 624 0 -1 6320
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_241
timestamp 1624494425
transform -1 0 624 0 1 6320
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_240
timestamp 1624494425
transform -1 0 624 0 -1 7110
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_239
timestamp 1624494425
transform -1 0 624 0 1 7110
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_238
timestamp 1624494425
transform -1 0 624 0 -1 7900
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_237
timestamp 1624494425
transform -1 0 624 0 1 7900
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_236
timestamp 1624494425
transform -1 0 624 0 -1 8690
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_235
timestamp 1624494425
transform -1 0 624 0 1 8690
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_234
timestamp 1624494425
transform -1 0 624 0 -1 9480
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_233
timestamp 1624494425
transform -1 0 624 0 1 9480
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_232
timestamp 1624494425
transform -1 0 624 0 -1 10270
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_231
timestamp 1624494425
transform -1 0 624 0 1 10270
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_230
timestamp 1624494425
transform -1 0 624 0 -1 11060
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_229
timestamp 1624494425
transform -1 0 624 0 1 11060
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_228
timestamp 1624494425
transform -1 0 624 0 -1 11850
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_227
timestamp 1624494425
transform -1 0 624 0 1 11850
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_226
timestamp 1624494425
transform -1 0 624 0 -1 12640
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_225
timestamp 1624494425
transform -1 0 624 0 1 12640
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_224
timestamp 1624494425
transform -1 0 624 0 -1 13430
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_223
timestamp 1624494425
transform -1 0 624 0 1 13430
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_222
timestamp 1624494425
transform -1 0 624 0 -1 14220
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_221
timestamp 1624494425
transform -1 0 624 0 1 14220
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_220
timestamp 1624494425
transform -1 0 624 0 -1 15010
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_219
timestamp 1624494425
transform -1 0 624 0 1 15010
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_218
timestamp 1624494425
transform -1 0 624 0 -1 15800
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_217
timestamp 1624494425
transform -1 0 624 0 1 15800
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_216
timestamp 1624494425
transform -1 0 624 0 -1 16590
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_215
timestamp 1624494425
transform -1 0 624 0 1 16590
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_214
timestamp 1624494425
transform -1 0 624 0 -1 17380
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_213
timestamp 1624494425
transform -1 0 624 0 1 17380
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_212
timestamp 1624494425
transform -1 0 624 0 -1 18170
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_211
timestamp 1624494425
transform -1 0 624 0 1 18170
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_210
timestamp 1624494425
transform -1 0 624 0 -1 18960
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_209
timestamp 1624494425
transform -1 0 624 0 1 18960
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_208
timestamp 1624494425
transform -1 0 624 0 -1 19750
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_207
timestamp 1624494425
transform -1 0 624 0 1 19750
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_206
timestamp 1624494425
transform -1 0 624 0 -1 20540
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_205
timestamp 1624494425
transform -1 0 624 0 1 20540
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_204
timestamp 1624494425
transform -1 0 624 0 -1 21330
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_203
timestamp 1624494425
transform -1 0 624 0 1 21330
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_202
timestamp 1624494425
transform -1 0 624 0 -1 22120
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_201
timestamp 1624494425
transform -1 0 624 0 1 22120
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_200
timestamp 1624494425
transform -1 0 624 0 -1 22910
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_199
timestamp 1624494425
transform -1 0 624 0 1 22910
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_198
timestamp 1624494425
transform -1 0 624 0 -1 23700
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_197
timestamp 1624494425
transform -1 0 624 0 1 23700
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_196
timestamp 1624494425
transform -1 0 624 0 -1 24490
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_195
timestamp 1624494425
transform -1 0 624 0 1 24490
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_194
timestamp 1624494425
transform -1 0 624 0 -1 25280
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_193
timestamp 1624494425
transform -1 0 624 0 1 25280
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_192
timestamp 1624494425
transform -1 0 624 0 -1 26070
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_191
timestamp 1624494425
transform -1 0 624 0 1 26070
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_190
timestamp 1624494425
transform -1 0 624 0 -1 26860
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_189
timestamp 1624494425
transform -1 0 624 0 1 26860
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_188
timestamp 1624494425
transform -1 0 624 0 -1 27650
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_187
timestamp 1624494425
transform -1 0 624 0 1 27650
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_186
timestamp 1624494425
transform -1 0 624 0 -1 28440
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_185
timestamp 1624494425
transform -1 0 624 0 1 28440
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_184
timestamp 1624494425
transform -1 0 624 0 -1 29230
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_183
timestamp 1624494425
transform -1 0 624 0 1 29230
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_182
timestamp 1624494425
transform -1 0 624 0 -1 30020
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_181
timestamp 1624494425
transform -1 0 624 0 1 30020
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_180
timestamp 1624494425
transform -1 0 624 0 -1 30810
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_179
timestamp 1624494425
transform -1 0 624 0 1 30810
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_178
timestamp 1624494425
transform -1 0 624 0 -1 31600
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_177
timestamp 1624494425
transform -1 0 624 0 1 31600
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_176
timestamp 1624494425
transform -1 0 624 0 -1 32390
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_175
timestamp 1624494425
transform -1 0 624 0 1 32390
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_174
timestamp 1624494425
transform -1 0 624 0 -1 33180
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_173
timestamp 1624494425
transform -1 0 624 0 1 33180
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_172
timestamp 1624494425
transform -1 0 624 0 -1 33970
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_171
timestamp 1624494425
transform -1 0 624 0 1 33970
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_170
timestamp 1624494425
transform -1 0 624 0 -1 34760
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_169
timestamp 1624494425
transform -1 0 624 0 1 34760
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_168
timestamp 1624494425
transform -1 0 624 0 -1 35550
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_167
timestamp 1624494425
transform -1 0 624 0 1 35550
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_166
timestamp 1624494425
transform -1 0 624 0 -1 36340
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_165
timestamp 1624494425
transform -1 0 624 0 1 36340
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_164
timestamp 1624494425
transform -1 0 624 0 -1 37130
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_163
timestamp 1624494425
transform -1 0 624 0 1 37130
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_162
timestamp 1624494425
transform -1 0 624 0 -1 37920
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_161
timestamp 1624494425
transform -1 0 624 0 1 37920
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_160
timestamp 1624494425
transform -1 0 624 0 -1 38710
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_159
timestamp 1624494425
transform -1 0 624 0 1 38710
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_158
timestamp 1624494425
transform -1 0 624 0 -1 39500
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_157
timestamp 1624494425
transform -1 0 624 0 1 39500
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_156
timestamp 1624494425
transform -1 0 624 0 -1 40290
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_155
timestamp 1624494425
transform -1 0 624 0 1 40290
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_154
timestamp 1624494425
transform -1 0 624 0 -1 41080
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_153
timestamp 1624494425
transform -1 0 624 0 1 41080
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_152
timestamp 1624494425
transform -1 0 624 0 -1 41870
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_151
timestamp 1624494425
transform -1 0 624 0 1 41870
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_150
timestamp 1624494425
transform -1 0 624 0 -1 42660
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_149
timestamp 1624494425
transform -1 0 624 0 1 42660
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_148
timestamp 1624494425
transform -1 0 624 0 -1 43450
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_147
timestamp 1624494425
transform -1 0 624 0 1 43450
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_146
timestamp 1624494425
transform -1 0 624 0 -1 44240
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_145
timestamp 1624494425
transform -1 0 624 0 1 44240
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_144
timestamp 1624494425
transform -1 0 624 0 -1 45030
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_143
timestamp 1624494425
transform -1 0 624 0 1 45030
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_142
timestamp 1624494425
transform -1 0 624 0 -1 45820
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_141
timestamp 1624494425
transform -1 0 624 0 1 45820
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_140
timestamp 1624494425
transform -1 0 624 0 -1 46610
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_139
timestamp 1624494425
transform -1 0 624 0 1 46610
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_138
timestamp 1624494425
transform -1 0 624 0 -1 47400
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_137
timestamp 1624494425
transform -1 0 624 0 1 47400
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_136
timestamp 1624494425
transform -1 0 624 0 -1 48190
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_135
timestamp 1624494425
transform -1 0 624 0 1 48190
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_134
timestamp 1624494425
transform -1 0 624 0 -1 48980
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_133
timestamp 1624494425
transform -1 0 624 0 1 48980
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_132
timestamp 1624494425
transform -1 0 624 0 -1 49770
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_131
timestamp 1624494425
transform -1 0 624 0 1 49770
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_130
timestamp 1624494425
transform -1 0 624 0 -1 50560
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_129
timestamp 1624494425
transform -1 0 624 0 1 50560
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_128
timestamp 1624494425
transform -1 0 624 0 -1 51350
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_127
timestamp 1624494425
transform -1 0 624 0 1 51350
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_126
timestamp 1624494425
transform -1 0 624 0 -1 52140
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_125
timestamp 1624494425
transform -1 0 624 0 1 52140
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_124
timestamp 1624494425
transform -1 0 624 0 -1 52930
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_123
timestamp 1624494425
transform -1 0 624 0 1 52930
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_122
timestamp 1624494425
transform -1 0 624 0 -1 53720
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_121
timestamp 1624494425
transform -1 0 624 0 1 53720
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_120
timestamp 1624494425
transform -1 0 624 0 -1 54510
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_119
timestamp 1624494425
transform -1 0 624 0 1 54510
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_118
timestamp 1624494425
transform -1 0 624 0 -1 55300
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_117
timestamp 1624494425
transform -1 0 624 0 1 55300
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_116
timestamp 1624494425
transform -1 0 624 0 -1 56090
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_115
timestamp 1624494425
transform -1 0 624 0 1 56090
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_114
timestamp 1624494425
transform -1 0 624 0 -1 56880
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_113
timestamp 1624494425
transform -1 0 624 0 1 56880
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_112
timestamp 1624494425
transform -1 0 624 0 -1 57670
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_111
timestamp 1624494425
transform -1 0 624 0 1 57670
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_110
timestamp 1624494425
transform -1 0 624 0 -1 58460
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_109
timestamp 1624494425
transform -1 0 624 0 1 58460
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_108
timestamp 1624494425
transform -1 0 624 0 -1 59250
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_107
timestamp 1624494425
transform -1 0 624 0 1 59250
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_106
timestamp 1624494425
transform -1 0 624 0 -1 60040
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_105
timestamp 1624494425
transform -1 0 624 0 1 60040
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_104
timestamp 1624494425
transform -1 0 624 0 -1 60830
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_103
timestamp 1624494425
transform -1 0 624 0 1 60830
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_102
timestamp 1624494425
transform -1 0 624 0 -1 61620
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_101
timestamp 1624494425
transform -1 0 624 0 1 61620
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_100
timestamp 1624494425
transform -1 0 624 0 -1 62410
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_99
timestamp 1624494425
transform -1 0 624 0 1 62410
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_98
timestamp 1624494425
transform -1 0 624 0 -1 63200
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_97
timestamp 1624494425
transform -1 0 624 0 1 63200
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_96
timestamp 1624494425
transform -1 0 624 0 -1 63990
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_95
timestamp 1624494425
transform -1 0 624 0 1 63990
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_94
timestamp 1624494425
transform -1 0 624 0 -1 64780
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_93
timestamp 1624494425
transform -1 0 624 0 1 64780
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_92
timestamp 1624494425
transform -1 0 624 0 -1 65570
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_91
timestamp 1624494425
transform -1 0 624 0 1 65570
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_90
timestamp 1624494425
transform -1 0 624 0 -1 66360
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_89
timestamp 1624494425
transform -1 0 624 0 1 66360
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_88
timestamp 1624494425
transform -1 0 624 0 -1 67150
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_87
timestamp 1624494425
transform -1 0 624 0 1 67150
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_86
timestamp 1624494425
transform -1 0 624 0 -1 67940
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_85
timestamp 1624494425
transform -1 0 624 0 1 67940
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_84
timestamp 1624494425
transform -1 0 624 0 -1 68730
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_83
timestamp 1624494425
transform -1 0 624 0 1 68730
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_82
timestamp 1624494425
transform -1 0 624 0 -1 69520
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_81
timestamp 1624494425
transform -1 0 624 0 1 69520
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_80
timestamp 1624494425
transform -1 0 624 0 -1 70310
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_79
timestamp 1624494425
transform -1 0 624 0 1 70310
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_78
timestamp 1624494425
transform -1 0 624 0 -1 71100
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_77
timestamp 1624494425
transform -1 0 624 0 1 71100
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_76
timestamp 1624494425
transform -1 0 624 0 -1 71890
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_75
timestamp 1624494425
transform -1 0 624 0 1 71890
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_74
timestamp 1624494425
transform -1 0 624 0 -1 72680
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_73
timestamp 1624494425
transform -1 0 624 0 1 72680
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_72
timestamp 1624494425
transform -1 0 624 0 -1 73470
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_71
timestamp 1624494425
transform -1 0 624 0 1 73470
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_70
timestamp 1624494425
transform -1 0 624 0 -1 74260
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_69
timestamp 1624494425
transform -1 0 624 0 1 74260
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_68
timestamp 1624494425
transform -1 0 624 0 -1 75050
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_67
timestamp 1624494425
transform -1 0 624 0 1 75050
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_66
timestamp 1624494425
transform -1 0 624 0 -1 75840
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_65
timestamp 1624494425
transform -1 0 624 0 1 75840
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_64
timestamp 1624494425
transform -1 0 624 0 -1 76630
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_63
timestamp 1624494425
transform -1 0 624 0 1 76630
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_62
timestamp 1624494425
transform -1 0 624 0 -1 77420
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_61
timestamp 1624494425
transform -1 0 624 0 1 77420
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_60
timestamp 1624494425
transform -1 0 624 0 -1 78210
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_59
timestamp 1624494425
transform -1 0 624 0 1 78210
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_58
timestamp 1624494425
transform -1 0 624 0 -1 79000
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_57
timestamp 1624494425
transform -1 0 624 0 1 79000
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_56
timestamp 1624494425
transform -1 0 624 0 -1 79790
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_55
timestamp 1624494425
transform -1 0 624 0 1 79790
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_54
timestamp 1624494425
transform -1 0 624 0 -1 80580
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_53
timestamp 1624494425
transform -1 0 624 0 1 80580
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_52
timestamp 1624494425
transform -1 0 624 0 -1 81370
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_51
timestamp 1624494425
transform -1 0 624 0 1 81370
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_50
timestamp 1624494425
transform -1 0 624 0 -1 82160
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_49
timestamp 1624494425
transform -1 0 624 0 1 82160
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_48
timestamp 1624494425
transform -1 0 624 0 -1 82950
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_47
timestamp 1624494425
transform -1 0 624 0 1 82950
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_46
timestamp 1624494425
transform -1 0 624 0 -1 83740
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_45
timestamp 1624494425
transform -1 0 624 0 1 83740
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_44
timestamp 1624494425
transform -1 0 624 0 -1 84530
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_43
timestamp 1624494425
transform -1 0 624 0 1 84530
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_42
timestamp 1624494425
transform -1 0 624 0 -1 85320
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_41
timestamp 1624494425
transform -1 0 624 0 1 85320
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_40
timestamp 1624494425
transform -1 0 624 0 -1 86110
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_39
timestamp 1624494425
transform -1 0 624 0 1 86110
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_38
timestamp 1624494425
transform -1 0 624 0 -1 86900
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_37
timestamp 1624494425
transform -1 0 624 0 1 86900
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_36
timestamp 1624494425
transform -1 0 624 0 -1 87690
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_35
timestamp 1624494425
transform -1 0 624 0 1 87690
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_34
timestamp 1624494425
transform -1 0 624 0 -1 88480
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_33
timestamp 1624494425
transform -1 0 624 0 1 88480
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_32
timestamp 1624494425
transform -1 0 624 0 -1 89270
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_31
timestamp 1624494425
transform -1 0 624 0 1 89270
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_30
timestamp 1624494425
transform -1 0 624 0 -1 90060
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_29
timestamp 1624494425
transform -1 0 624 0 1 90060
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_28
timestamp 1624494425
transform -1 0 624 0 -1 90850
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_27
timestamp 1624494425
transform -1 0 624 0 1 90850
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_26
timestamp 1624494425
transform -1 0 624 0 -1 91640
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_25
timestamp 1624494425
transform -1 0 624 0 1 91640
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_24
timestamp 1624494425
transform -1 0 624 0 -1 92430
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_23
timestamp 1624494425
transform -1 0 624 0 1 92430
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_22
timestamp 1624494425
transform -1 0 624 0 -1 93220
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_21
timestamp 1624494425
transform -1 0 624 0 1 93220
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_20
timestamp 1624494425
transform -1 0 624 0 -1 94010
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_19
timestamp 1624494425
transform -1 0 624 0 1 94010
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_18
timestamp 1624494425
transform -1 0 624 0 -1 94800
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_17
timestamp 1624494425
transform -1 0 624 0 1 94800
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_16
timestamp 1624494425
transform -1 0 624 0 -1 95590
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_15
timestamp 1624494425
transform -1 0 624 0 1 95590
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_14
timestamp 1624494425
transform -1 0 624 0 -1 96380
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_13
timestamp 1624494425
transform -1 0 624 0 1 96380
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_12
timestamp 1624494425
transform -1 0 624 0 -1 97170
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_11
timestamp 1624494425
transform -1 0 624 0 1 97170
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_10
timestamp 1624494425
transform -1 0 624 0 -1 97960
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_9
timestamp 1624494425
transform -1 0 624 0 1 97960
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_8
timestamp 1624494425
transform -1 0 624 0 -1 98750
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_7
timestamp 1624494425
transform -1 0 624 0 1 98750
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_6
timestamp 1624494425
transform -1 0 624 0 -1 99540
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_5
timestamp 1624494425
transform -1 0 624 0 1 99540
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_4
timestamp 1624494425
transform -1 0 624 0 -1 100330
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_3
timestamp 1624494425
transform -1 0 624 0 1 100330
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_2
timestamp 1624494425
transform -1 0 624 0 -1 101120
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_1
timestamp 1624494425
transform -1 0 624 0 1 101120
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_0
timestamp 1624494425
transform -1 0 624 0 -1 101910
box -42 -105 650 424
<< labels >>
rlabel metal1 s 510 0 546 102700 4 bl_0_0
rlabel metal1 s 438 0 474 102700 4 br_0_0
rlabel metal1 s 294 0 330 102700 4 bl_1_0
rlabel metal1 s 222 0 258 102700 4 br_1_0
rlabel metal2 s 0 419 624 467 4 wl_0_0
rlabel metal2 s 0 1113 624 1161 4 wl_0_1
rlabel metal2 s 0 1209 624 1257 4 wl_0_2
rlabel metal2 s 0 1903 624 1951 4 wl_0_3
rlabel metal2 s 0 1999 624 2047 4 wl_0_4
rlabel metal2 s 0 2693 624 2741 4 wl_0_5
rlabel metal2 s 0 2789 624 2837 4 wl_0_6
rlabel metal2 s 0 3483 624 3531 4 wl_0_7
rlabel metal2 s 0 3579 624 3627 4 wl_0_8
rlabel metal2 s 0 4273 624 4321 4 wl_0_9
rlabel metal2 s 0 4369 624 4417 4 wl_0_10
rlabel metal2 s 0 5063 624 5111 4 wl_0_11
rlabel metal2 s 0 5159 624 5207 4 wl_0_12
rlabel metal2 s 0 5853 624 5901 4 wl_0_13
rlabel metal2 s 0 5949 624 5997 4 wl_0_14
rlabel metal2 s 0 6643 624 6691 4 wl_0_15
rlabel metal2 s 0 6739 624 6787 4 wl_0_16
rlabel metal2 s 0 7433 624 7481 4 wl_0_17
rlabel metal2 s 0 7529 624 7577 4 wl_0_18
rlabel metal2 s 0 8223 624 8271 4 wl_0_19
rlabel metal2 s 0 8319 624 8367 4 wl_0_20
rlabel metal2 s 0 9013 624 9061 4 wl_0_21
rlabel metal2 s 0 9109 624 9157 4 wl_0_22
rlabel metal2 s 0 9803 624 9851 4 wl_0_23
rlabel metal2 s 0 9899 624 9947 4 wl_0_24
rlabel metal2 s 0 10593 624 10641 4 wl_0_25
rlabel metal2 s 0 10689 624 10737 4 wl_0_26
rlabel metal2 s 0 11383 624 11431 4 wl_0_27
rlabel metal2 s 0 11479 624 11527 4 wl_0_28
rlabel metal2 s 0 12173 624 12221 4 wl_0_29
rlabel metal2 s 0 12269 624 12317 4 wl_0_30
rlabel metal2 s 0 12963 624 13011 4 wl_0_31
rlabel metal2 s 0 13059 624 13107 4 wl_0_32
rlabel metal2 s 0 13753 624 13801 4 wl_0_33
rlabel metal2 s 0 13849 624 13897 4 wl_0_34
rlabel metal2 s 0 14543 624 14591 4 wl_0_35
rlabel metal2 s 0 14639 624 14687 4 wl_0_36
rlabel metal2 s 0 15333 624 15381 4 wl_0_37
rlabel metal2 s 0 15429 624 15477 4 wl_0_38
rlabel metal2 s 0 16123 624 16171 4 wl_0_39
rlabel metal2 s 0 16219 624 16267 4 wl_0_40
rlabel metal2 s 0 16913 624 16961 4 wl_0_41
rlabel metal2 s 0 17009 624 17057 4 wl_0_42
rlabel metal2 s 0 17703 624 17751 4 wl_0_43
rlabel metal2 s 0 17799 624 17847 4 wl_0_44
rlabel metal2 s 0 18493 624 18541 4 wl_0_45
rlabel metal2 s 0 18589 624 18637 4 wl_0_46
rlabel metal2 s 0 19283 624 19331 4 wl_0_47
rlabel metal2 s 0 19379 624 19427 4 wl_0_48
rlabel metal2 s 0 20073 624 20121 4 wl_0_49
rlabel metal2 s 0 20169 624 20217 4 wl_0_50
rlabel metal2 s 0 20863 624 20911 4 wl_0_51
rlabel metal2 s 0 20959 624 21007 4 wl_0_52
rlabel metal2 s 0 21653 624 21701 4 wl_0_53
rlabel metal2 s 0 21749 624 21797 4 wl_0_54
rlabel metal2 s 0 22443 624 22491 4 wl_0_55
rlabel metal2 s 0 22539 624 22587 4 wl_0_56
rlabel metal2 s 0 23233 624 23281 4 wl_0_57
rlabel metal2 s 0 23329 624 23377 4 wl_0_58
rlabel metal2 s 0 24023 624 24071 4 wl_0_59
rlabel metal2 s 0 24119 624 24167 4 wl_0_60
rlabel metal2 s 0 24813 624 24861 4 wl_0_61
rlabel metal2 s 0 24909 624 24957 4 wl_0_62
rlabel metal2 s 0 25603 624 25651 4 wl_0_63
rlabel metal2 s 0 25699 624 25747 4 wl_0_64
rlabel metal2 s 0 26393 624 26441 4 wl_0_65
rlabel metal2 s 0 26489 624 26537 4 wl_0_66
rlabel metal2 s 0 27183 624 27231 4 wl_0_67
rlabel metal2 s 0 27279 624 27327 4 wl_0_68
rlabel metal2 s 0 27973 624 28021 4 wl_0_69
rlabel metal2 s 0 28069 624 28117 4 wl_0_70
rlabel metal2 s 0 28763 624 28811 4 wl_0_71
rlabel metal2 s 0 28859 624 28907 4 wl_0_72
rlabel metal2 s 0 29553 624 29601 4 wl_0_73
rlabel metal2 s 0 29649 624 29697 4 wl_0_74
rlabel metal2 s 0 30343 624 30391 4 wl_0_75
rlabel metal2 s 0 30439 624 30487 4 wl_0_76
rlabel metal2 s 0 31133 624 31181 4 wl_0_77
rlabel metal2 s 0 31229 624 31277 4 wl_0_78
rlabel metal2 s 0 31923 624 31971 4 wl_0_79
rlabel metal2 s 0 32019 624 32067 4 wl_0_80
rlabel metal2 s 0 32713 624 32761 4 wl_0_81
rlabel metal2 s 0 32809 624 32857 4 wl_0_82
rlabel metal2 s 0 33503 624 33551 4 wl_0_83
rlabel metal2 s 0 33599 624 33647 4 wl_0_84
rlabel metal2 s 0 34293 624 34341 4 wl_0_85
rlabel metal2 s 0 34389 624 34437 4 wl_0_86
rlabel metal2 s 0 35083 624 35131 4 wl_0_87
rlabel metal2 s 0 35179 624 35227 4 wl_0_88
rlabel metal2 s 0 35873 624 35921 4 wl_0_89
rlabel metal2 s 0 35969 624 36017 4 wl_0_90
rlabel metal2 s 0 36663 624 36711 4 wl_0_91
rlabel metal2 s 0 36759 624 36807 4 wl_0_92
rlabel metal2 s 0 37453 624 37501 4 wl_0_93
rlabel metal2 s 0 37549 624 37597 4 wl_0_94
rlabel metal2 s 0 38243 624 38291 4 wl_0_95
rlabel metal2 s 0 38339 624 38387 4 wl_0_96
rlabel metal2 s 0 39033 624 39081 4 wl_0_97
rlabel metal2 s 0 39129 624 39177 4 wl_0_98
rlabel metal2 s 0 39823 624 39871 4 wl_0_99
rlabel metal2 s 0 39919 624 39967 4 wl_0_100
rlabel metal2 s 0 40613 624 40661 4 wl_0_101
rlabel metal2 s 0 40709 624 40757 4 wl_0_102
rlabel metal2 s 0 41403 624 41451 4 wl_0_103
rlabel metal2 s 0 41499 624 41547 4 wl_0_104
rlabel metal2 s 0 42193 624 42241 4 wl_0_105
rlabel metal2 s 0 42289 624 42337 4 wl_0_106
rlabel metal2 s 0 42983 624 43031 4 wl_0_107
rlabel metal2 s 0 43079 624 43127 4 wl_0_108
rlabel metal2 s 0 43773 624 43821 4 wl_0_109
rlabel metal2 s 0 43869 624 43917 4 wl_0_110
rlabel metal2 s 0 44563 624 44611 4 wl_0_111
rlabel metal2 s 0 44659 624 44707 4 wl_0_112
rlabel metal2 s 0 45353 624 45401 4 wl_0_113
rlabel metal2 s 0 45449 624 45497 4 wl_0_114
rlabel metal2 s 0 46143 624 46191 4 wl_0_115
rlabel metal2 s 0 46239 624 46287 4 wl_0_116
rlabel metal2 s 0 46933 624 46981 4 wl_0_117
rlabel metal2 s 0 47029 624 47077 4 wl_0_118
rlabel metal2 s 0 47723 624 47771 4 wl_0_119
rlabel metal2 s 0 47819 624 47867 4 wl_0_120
rlabel metal2 s 0 48513 624 48561 4 wl_0_121
rlabel metal2 s 0 48609 624 48657 4 wl_0_122
rlabel metal2 s 0 49303 624 49351 4 wl_0_123
rlabel metal2 s 0 49399 624 49447 4 wl_0_124
rlabel metal2 s 0 50093 624 50141 4 wl_0_125
rlabel metal2 s 0 50189 624 50237 4 wl_0_126
rlabel metal2 s 0 50883 624 50931 4 wl_0_127
rlabel metal2 s 0 50979 624 51027 4 wl_0_128
rlabel metal2 s 0 51673 624 51721 4 wl_0_129
rlabel metal2 s 0 51769 624 51817 4 wl_0_130
rlabel metal2 s 0 52463 624 52511 4 wl_0_131
rlabel metal2 s 0 52559 624 52607 4 wl_0_132
rlabel metal2 s 0 53253 624 53301 4 wl_0_133
rlabel metal2 s 0 53349 624 53397 4 wl_0_134
rlabel metal2 s 0 54043 624 54091 4 wl_0_135
rlabel metal2 s 0 54139 624 54187 4 wl_0_136
rlabel metal2 s 0 54833 624 54881 4 wl_0_137
rlabel metal2 s 0 54929 624 54977 4 wl_0_138
rlabel metal2 s 0 55623 624 55671 4 wl_0_139
rlabel metal2 s 0 55719 624 55767 4 wl_0_140
rlabel metal2 s 0 56413 624 56461 4 wl_0_141
rlabel metal2 s 0 56509 624 56557 4 wl_0_142
rlabel metal2 s 0 57203 624 57251 4 wl_0_143
rlabel metal2 s 0 57299 624 57347 4 wl_0_144
rlabel metal2 s 0 57993 624 58041 4 wl_0_145
rlabel metal2 s 0 58089 624 58137 4 wl_0_146
rlabel metal2 s 0 58783 624 58831 4 wl_0_147
rlabel metal2 s 0 58879 624 58927 4 wl_0_148
rlabel metal2 s 0 59573 624 59621 4 wl_0_149
rlabel metal2 s 0 59669 624 59717 4 wl_0_150
rlabel metal2 s 0 60363 624 60411 4 wl_0_151
rlabel metal2 s 0 60459 624 60507 4 wl_0_152
rlabel metal2 s 0 61153 624 61201 4 wl_0_153
rlabel metal2 s 0 61249 624 61297 4 wl_0_154
rlabel metal2 s 0 61943 624 61991 4 wl_0_155
rlabel metal2 s 0 62039 624 62087 4 wl_0_156
rlabel metal2 s 0 62733 624 62781 4 wl_0_157
rlabel metal2 s 0 62829 624 62877 4 wl_0_158
rlabel metal2 s 0 63523 624 63571 4 wl_0_159
rlabel metal2 s 0 63619 624 63667 4 wl_0_160
rlabel metal2 s 0 64313 624 64361 4 wl_0_161
rlabel metal2 s 0 64409 624 64457 4 wl_0_162
rlabel metal2 s 0 65103 624 65151 4 wl_0_163
rlabel metal2 s 0 65199 624 65247 4 wl_0_164
rlabel metal2 s 0 65893 624 65941 4 wl_0_165
rlabel metal2 s 0 65989 624 66037 4 wl_0_166
rlabel metal2 s 0 66683 624 66731 4 wl_0_167
rlabel metal2 s 0 66779 624 66827 4 wl_0_168
rlabel metal2 s 0 67473 624 67521 4 wl_0_169
rlabel metal2 s 0 67569 624 67617 4 wl_0_170
rlabel metal2 s 0 68263 624 68311 4 wl_0_171
rlabel metal2 s 0 68359 624 68407 4 wl_0_172
rlabel metal2 s 0 69053 624 69101 4 wl_0_173
rlabel metal2 s 0 69149 624 69197 4 wl_0_174
rlabel metal2 s 0 69843 624 69891 4 wl_0_175
rlabel metal2 s 0 69939 624 69987 4 wl_0_176
rlabel metal2 s 0 70633 624 70681 4 wl_0_177
rlabel metal2 s 0 70729 624 70777 4 wl_0_178
rlabel metal2 s 0 71423 624 71471 4 wl_0_179
rlabel metal2 s 0 71519 624 71567 4 wl_0_180
rlabel metal2 s 0 72213 624 72261 4 wl_0_181
rlabel metal2 s 0 72309 624 72357 4 wl_0_182
rlabel metal2 s 0 73003 624 73051 4 wl_0_183
rlabel metal2 s 0 73099 624 73147 4 wl_0_184
rlabel metal2 s 0 73793 624 73841 4 wl_0_185
rlabel metal2 s 0 73889 624 73937 4 wl_0_186
rlabel metal2 s 0 74583 624 74631 4 wl_0_187
rlabel metal2 s 0 74679 624 74727 4 wl_0_188
rlabel metal2 s 0 75373 624 75421 4 wl_0_189
rlabel metal2 s 0 75469 624 75517 4 wl_0_190
rlabel metal2 s 0 76163 624 76211 4 wl_0_191
rlabel metal2 s 0 76259 624 76307 4 wl_0_192
rlabel metal2 s 0 76953 624 77001 4 wl_0_193
rlabel metal2 s 0 77049 624 77097 4 wl_0_194
rlabel metal2 s 0 77743 624 77791 4 wl_0_195
rlabel metal2 s 0 77839 624 77887 4 wl_0_196
rlabel metal2 s 0 78533 624 78581 4 wl_0_197
rlabel metal2 s 0 78629 624 78677 4 wl_0_198
rlabel metal2 s 0 79323 624 79371 4 wl_0_199
rlabel metal2 s 0 79419 624 79467 4 wl_0_200
rlabel metal2 s 0 80113 624 80161 4 wl_0_201
rlabel metal2 s 0 80209 624 80257 4 wl_0_202
rlabel metal2 s 0 80903 624 80951 4 wl_0_203
rlabel metal2 s 0 80999 624 81047 4 wl_0_204
rlabel metal2 s 0 81693 624 81741 4 wl_0_205
rlabel metal2 s 0 81789 624 81837 4 wl_0_206
rlabel metal2 s 0 82483 624 82531 4 wl_0_207
rlabel metal2 s 0 82579 624 82627 4 wl_0_208
rlabel metal2 s 0 83273 624 83321 4 wl_0_209
rlabel metal2 s 0 83369 624 83417 4 wl_0_210
rlabel metal2 s 0 84063 624 84111 4 wl_0_211
rlabel metal2 s 0 84159 624 84207 4 wl_0_212
rlabel metal2 s 0 84853 624 84901 4 wl_0_213
rlabel metal2 s 0 84949 624 84997 4 wl_0_214
rlabel metal2 s 0 85643 624 85691 4 wl_0_215
rlabel metal2 s 0 85739 624 85787 4 wl_0_216
rlabel metal2 s 0 86433 624 86481 4 wl_0_217
rlabel metal2 s 0 86529 624 86577 4 wl_0_218
rlabel metal2 s 0 87223 624 87271 4 wl_0_219
rlabel metal2 s 0 87319 624 87367 4 wl_0_220
rlabel metal2 s 0 88013 624 88061 4 wl_0_221
rlabel metal2 s 0 88109 624 88157 4 wl_0_222
rlabel metal2 s 0 88803 624 88851 4 wl_0_223
rlabel metal2 s 0 88899 624 88947 4 wl_0_224
rlabel metal2 s 0 89593 624 89641 4 wl_0_225
rlabel metal2 s 0 89689 624 89737 4 wl_0_226
rlabel metal2 s 0 90383 624 90431 4 wl_0_227
rlabel metal2 s 0 90479 624 90527 4 wl_0_228
rlabel metal2 s 0 91173 624 91221 4 wl_0_229
rlabel metal2 s 0 91269 624 91317 4 wl_0_230
rlabel metal2 s 0 91963 624 92011 4 wl_0_231
rlabel metal2 s 0 92059 624 92107 4 wl_0_232
rlabel metal2 s 0 92753 624 92801 4 wl_0_233
rlabel metal2 s 0 92849 624 92897 4 wl_0_234
rlabel metal2 s 0 93543 624 93591 4 wl_0_235
rlabel metal2 s 0 93639 624 93687 4 wl_0_236
rlabel metal2 s 0 94333 624 94381 4 wl_0_237
rlabel metal2 s 0 94429 624 94477 4 wl_0_238
rlabel metal2 s 0 95123 624 95171 4 wl_0_239
rlabel metal2 s 0 95219 624 95267 4 wl_0_240
rlabel metal2 s 0 95913 624 95961 4 wl_0_241
rlabel metal2 s 0 96009 624 96057 4 wl_0_242
rlabel metal2 s 0 96703 624 96751 4 wl_0_243
rlabel metal2 s 0 96799 624 96847 4 wl_0_244
rlabel metal2 s 0 97493 624 97541 4 wl_0_245
rlabel metal2 s 0 97589 624 97637 4 wl_0_246
rlabel metal2 s 0 98283 624 98331 4 wl_0_247
rlabel metal2 s 0 98379 624 98427 4 wl_0_248
rlabel metal2 s 0 99073 624 99121 4 wl_0_249
rlabel metal2 s 0 99169 624 99217 4 wl_0_250
rlabel metal2 s 0 99863 624 99911 4 wl_0_251
rlabel metal2 s 0 99959 624 100007 4 wl_0_252
rlabel metal2 s 0 100653 624 100701 4 wl_0_253
rlabel metal2 s 0 100749 624 100797 4 wl_0_254
rlabel metal2 s 0 101443 624 101491 4 wl_0_255
rlabel metal2 s 0 101539 624 101587 4 wl_0_256
rlabel metal2 s 0 102233 624 102281 4 wl_0_257
rlabel metal2 s 0 639 624 687 4 wl_1_0
rlabel metal2 s 0 893 624 941 4 wl_1_1
rlabel metal2 s 0 1429 624 1477 4 wl_1_2
rlabel metal2 s 0 1683 624 1731 4 wl_1_3
rlabel metal2 s 0 2219 624 2267 4 wl_1_4
rlabel metal2 s 0 2473 624 2521 4 wl_1_5
rlabel metal2 s 0 3009 624 3057 4 wl_1_6
rlabel metal2 s 0 3263 624 3311 4 wl_1_7
rlabel metal2 s 0 3799 624 3847 4 wl_1_8
rlabel metal2 s 0 4053 624 4101 4 wl_1_9
rlabel metal2 s 0 4589 624 4637 4 wl_1_10
rlabel metal2 s 0 4843 624 4891 4 wl_1_11
rlabel metal2 s 0 5379 624 5427 4 wl_1_12
rlabel metal2 s 0 5633 624 5681 4 wl_1_13
rlabel metal2 s 0 6169 624 6217 4 wl_1_14
rlabel metal2 s 0 6423 624 6471 4 wl_1_15
rlabel metal2 s 0 6959 624 7007 4 wl_1_16
rlabel metal2 s 0 7213 624 7261 4 wl_1_17
rlabel metal2 s 0 7749 624 7797 4 wl_1_18
rlabel metal2 s 0 8003 624 8051 4 wl_1_19
rlabel metal2 s 0 8539 624 8587 4 wl_1_20
rlabel metal2 s 0 8793 624 8841 4 wl_1_21
rlabel metal2 s 0 9329 624 9377 4 wl_1_22
rlabel metal2 s 0 9583 624 9631 4 wl_1_23
rlabel metal2 s 0 10119 624 10167 4 wl_1_24
rlabel metal2 s 0 10373 624 10421 4 wl_1_25
rlabel metal2 s 0 10909 624 10957 4 wl_1_26
rlabel metal2 s 0 11163 624 11211 4 wl_1_27
rlabel metal2 s 0 11699 624 11747 4 wl_1_28
rlabel metal2 s 0 11953 624 12001 4 wl_1_29
rlabel metal2 s 0 12489 624 12537 4 wl_1_30
rlabel metal2 s 0 12743 624 12791 4 wl_1_31
rlabel metal2 s 0 13279 624 13327 4 wl_1_32
rlabel metal2 s 0 13533 624 13581 4 wl_1_33
rlabel metal2 s 0 14069 624 14117 4 wl_1_34
rlabel metal2 s 0 14323 624 14371 4 wl_1_35
rlabel metal2 s 0 14859 624 14907 4 wl_1_36
rlabel metal2 s 0 15113 624 15161 4 wl_1_37
rlabel metal2 s 0 15649 624 15697 4 wl_1_38
rlabel metal2 s 0 15903 624 15951 4 wl_1_39
rlabel metal2 s 0 16439 624 16487 4 wl_1_40
rlabel metal2 s 0 16693 624 16741 4 wl_1_41
rlabel metal2 s 0 17229 624 17277 4 wl_1_42
rlabel metal2 s 0 17483 624 17531 4 wl_1_43
rlabel metal2 s 0 18019 624 18067 4 wl_1_44
rlabel metal2 s 0 18273 624 18321 4 wl_1_45
rlabel metal2 s 0 18809 624 18857 4 wl_1_46
rlabel metal2 s 0 19063 624 19111 4 wl_1_47
rlabel metal2 s 0 19599 624 19647 4 wl_1_48
rlabel metal2 s 0 19853 624 19901 4 wl_1_49
rlabel metal2 s 0 20389 624 20437 4 wl_1_50
rlabel metal2 s 0 20643 624 20691 4 wl_1_51
rlabel metal2 s 0 21179 624 21227 4 wl_1_52
rlabel metal2 s 0 21433 624 21481 4 wl_1_53
rlabel metal2 s 0 21969 624 22017 4 wl_1_54
rlabel metal2 s 0 22223 624 22271 4 wl_1_55
rlabel metal2 s 0 22759 624 22807 4 wl_1_56
rlabel metal2 s 0 23013 624 23061 4 wl_1_57
rlabel metal2 s 0 23549 624 23597 4 wl_1_58
rlabel metal2 s 0 23803 624 23851 4 wl_1_59
rlabel metal2 s 0 24339 624 24387 4 wl_1_60
rlabel metal2 s 0 24593 624 24641 4 wl_1_61
rlabel metal2 s 0 25129 624 25177 4 wl_1_62
rlabel metal2 s 0 25383 624 25431 4 wl_1_63
rlabel metal2 s 0 25919 624 25967 4 wl_1_64
rlabel metal2 s 0 26173 624 26221 4 wl_1_65
rlabel metal2 s 0 26709 624 26757 4 wl_1_66
rlabel metal2 s 0 26963 624 27011 4 wl_1_67
rlabel metal2 s 0 27499 624 27547 4 wl_1_68
rlabel metal2 s 0 27753 624 27801 4 wl_1_69
rlabel metal2 s 0 28289 624 28337 4 wl_1_70
rlabel metal2 s 0 28543 624 28591 4 wl_1_71
rlabel metal2 s 0 29079 624 29127 4 wl_1_72
rlabel metal2 s 0 29333 624 29381 4 wl_1_73
rlabel metal2 s 0 29869 624 29917 4 wl_1_74
rlabel metal2 s 0 30123 624 30171 4 wl_1_75
rlabel metal2 s 0 30659 624 30707 4 wl_1_76
rlabel metal2 s 0 30913 624 30961 4 wl_1_77
rlabel metal2 s 0 31449 624 31497 4 wl_1_78
rlabel metal2 s 0 31703 624 31751 4 wl_1_79
rlabel metal2 s 0 32239 624 32287 4 wl_1_80
rlabel metal2 s 0 32493 624 32541 4 wl_1_81
rlabel metal2 s 0 33029 624 33077 4 wl_1_82
rlabel metal2 s 0 33283 624 33331 4 wl_1_83
rlabel metal2 s 0 33819 624 33867 4 wl_1_84
rlabel metal2 s 0 34073 624 34121 4 wl_1_85
rlabel metal2 s 0 34609 624 34657 4 wl_1_86
rlabel metal2 s 0 34863 624 34911 4 wl_1_87
rlabel metal2 s 0 35399 624 35447 4 wl_1_88
rlabel metal2 s 0 35653 624 35701 4 wl_1_89
rlabel metal2 s 0 36189 624 36237 4 wl_1_90
rlabel metal2 s 0 36443 624 36491 4 wl_1_91
rlabel metal2 s 0 36979 624 37027 4 wl_1_92
rlabel metal2 s 0 37233 624 37281 4 wl_1_93
rlabel metal2 s 0 37769 624 37817 4 wl_1_94
rlabel metal2 s 0 38023 624 38071 4 wl_1_95
rlabel metal2 s 0 38559 624 38607 4 wl_1_96
rlabel metal2 s 0 38813 624 38861 4 wl_1_97
rlabel metal2 s 0 39349 624 39397 4 wl_1_98
rlabel metal2 s 0 39603 624 39651 4 wl_1_99
rlabel metal2 s 0 40139 624 40187 4 wl_1_100
rlabel metal2 s 0 40393 624 40441 4 wl_1_101
rlabel metal2 s 0 40929 624 40977 4 wl_1_102
rlabel metal2 s 0 41183 624 41231 4 wl_1_103
rlabel metal2 s 0 41719 624 41767 4 wl_1_104
rlabel metal2 s 0 41973 624 42021 4 wl_1_105
rlabel metal2 s 0 42509 624 42557 4 wl_1_106
rlabel metal2 s 0 42763 624 42811 4 wl_1_107
rlabel metal2 s 0 43299 624 43347 4 wl_1_108
rlabel metal2 s 0 43553 624 43601 4 wl_1_109
rlabel metal2 s 0 44089 624 44137 4 wl_1_110
rlabel metal2 s 0 44343 624 44391 4 wl_1_111
rlabel metal2 s 0 44879 624 44927 4 wl_1_112
rlabel metal2 s 0 45133 624 45181 4 wl_1_113
rlabel metal2 s 0 45669 624 45717 4 wl_1_114
rlabel metal2 s 0 45923 624 45971 4 wl_1_115
rlabel metal2 s 0 46459 624 46507 4 wl_1_116
rlabel metal2 s 0 46713 624 46761 4 wl_1_117
rlabel metal2 s 0 47249 624 47297 4 wl_1_118
rlabel metal2 s 0 47503 624 47551 4 wl_1_119
rlabel metal2 s 0 48039 624 48087 4 wl_1_120
rlabel metal2 s 0 48293 624 48341 4 wl_1_121
rlabel metal2 s 0 48829 624 48877 4 wl_1_122
rlabel metal2 s 0 49083 624 49131 4 wl_1_123
rlabel metal2 s 0 49619 624 49667 4 wl_1_124
rlabel metal2 s 0 49873 624 49921 4 wl_1_125
rlabel metal2 s 0 50409 624 50457 4 wl_1_126
rlabel metal2 s 0 50663 624 50711 4 wl_1_127
rlabel metal2 s 0 51199 624 51247 4 wl_1_128
rlabel metal2 s 0 51453 624 51501 4 wl_1_129
rlabel metal2 s 0 51989 624 52037 4 wl_1_130
rlabel metal2 s 0 52243 624 52291 4 wl_1_131
rlabel metal2 s 0 52779 624 52827 4 wl_1_132
rlabel metal2 s 0 53033 624 53081 4 wl_1_133
rlabel metal2 s 0 53569 624 53617 4 wl_1_134
rlabel metal2 s 0 53823 624 53871 4 wl_1_135
rlabel metal2 s 0 54359 624 54407 4 wl_1_136
rlabel metal2 s 0 54613 624 54661 4 wl_1_137
rlabel metal2 s 0 55149 624 55197 4 wl_1_138
rlabel metal2 s 0 55403 624 55451 4 wl_1_139
rlabel metal2 s 0 55939 624 55987 4 wl_1_140
rlabel metal2 s 0 56193 624 56241 4 wl_1_141
rlabel metal2 s 0 56729 624 56777 4 wl_1_142
rlabel metal2 s 0 56983 624 57031 4 wl_1_143
rlabel metal2 s 0 57519 624 57567 4 wl_1_144
rlabel metal2 s 0 57773 624 57821 4 wl_1_145
rlabel metal2 s 0 58309 624 58357 4 wl_1_146
rlabel metal2 s 0 58563 624 58611 4 wl_1_147
rlabel metal2 s 0 59099 624 59147 4 wl_1_148
rlabel metal2 s 0 59353 624 59401 4 wl_1_149
rlabel metal2 s 0 59889 624 59937 4 wl_1_150
rlabel metal2 s 0 60143 624 60191 4 wl_1_151
rlabel metal2 s 0 60679 624 60727 4 wl_1_152
rlabel metal2 s 0 60933 624 60981 4 wl_1_153
rlabel metal2 s 0 61469 624 61517 4 wl_1_154
rlabel metal2 s 0 61723 624 61771 4 wl_1_155
rlabel metal2 s 0 62259 624 62307 4 wl_1_156
rlabel metal2 s 0 62513 624 62561 4 wl_1_157
rlabel metal2 s 0 63049 624 63097 4 wl_1_158
rlabel metal2 s 0 63303 624 63351 4 wl_1_159
rlabel metal2 s 0 63839 624 63887 4 wl_1_160
rlabel metal2 s 0 64093 624 64141 4 wl_1_161
rlabel metal2 s 0 64629 624 64677 4 wl_1_162
rlabel metal2 s 0 64883 624 64931 4 wl_1_163
rlabel metal2 s 0 65419 624 65467 4 wl_1_164
rlabel metal2 s 0 65673 624 65721 4 wl_1_165
rlabel metal2 s 0 66209 624 66257 4 wl_1_166
rlabel metal2 s 0 66463 624 66511 4 wl_1_167
rlabel metal2 s 0 66999 624 67047 4 wl_1_168
rlabel metal2 s 0 67253 624 67301 4 wl_1_169
rlabel metal2 s 0 67789 624 67837 4 wl_1_170
rlabel metal2 s 0 68043 624 68091 4 wl_1_171
rlabel metal2 s 0 68579 624 68627 4 wl_1_172
rlabel metal2 s 0 68833 624 68881 4 wl_1_173
rlabel metal2 s 0 69369 624 69417 4 wl_1_174
rlabel metal2 s 0 69623 624 69671 4 wl_1_175
rlabel metal2 s 0 70159 624 70207 4 wl_1_176
rlabel metal2 s 0 70413 624 70461 4 wl_1_177
rlabel metal2 s 0 70949 624 70997 4 wl_1_178
rlabel metal2 s 0 71203 624 71251 4 wl_1_179
rlabel metal2 s 0 71739 624 71787 4 wl_1_180
rlabel metal2 s 0 71993 624 72041 4 wl_1_181
rlabel metal2 s 0 72529 624 72577 4 wl_1_182
rlabel metal2 s 0 72783 624 72831 4 wl_1_183
rlabel metal2 s 0 73319 624 73367 4 wl_1_184
rlabel metal2 s 0 73573 624 73621 4 wl_1_185
rlabel metal2 s 0 74109 624 74157 4 wl_1_186
rlabel metal2 s 0 74363 624 74411 4 wl_1_187
rlabel metal2 s 0 74899 624 74947 4 wl_1_188
rlabel metal2 s 0 75153 624 75201 4 wl_1_189
rlabel metal2 s 0 75689 624 75737 4 wl_1_190
rlabel metal2 s 0 75943 624 75991 4 wl_1_191
rlabel metal2 s 0 76479 624 76527 4 wl_1_192
rlabel metal2 s 0 76733 624 76781 4 wl_1_193
rlabel metal2 s 0 77269 624 77317 4 wl_1_194
rlabel metal2 s 0 77523 624 77571 4 wl_1_195
rlabel metal2 s 0 78059 624 78107 4 wl_1_196
rlabel metal2 s 0 78313 624 78361 4 wl_1_197
rlabel metal2 s 0 78849 624 78897 4 wl_1_198
rlabel metal2 s 0 79103 624 79151 4 wl_1_199
rlabel metal2 s 0 79639 624 79687 4 wl_1_200
rlabel metal2 s 0 79893 624 79941 4 wl_1_201
rlabel metal2 s 0 80429 624 80477 4 wl_1_202
rlabel metal2 s 0 80683 624 80731 4 wl_1_203
rlabel metal2 s 0 81219 624 81267 4 wl_1_204
rlabel metal2 s 0 81473 624 81521 4 wl_1_205
rlabel metal2 s 0 82009 624 82057 4 wl_1_206
rlabel metal2 s 0 82263 624 82311 4 wl_1_207
rlabel metal2 s 0 82799 624 82847 4 wl_1_208
rlabel metal2 s 0 83053 624 83101 4 wl_1_209
rlabel metal2 s 0 83589 624 83637 4 wl_1_210
rlabel metal2 s 0 83843 624 83891 4 wl_1_211
rlabel metal2 s 0 84379 624 84427 4 wl_1_212
rlabel metal2 s 0 84633 624 84681 4 wl_1_213
rlabel metal2 s 0 85169 624 85217 4 wl_1_214
rlabel metal2 s 0 85423 624 85471 4 wl_1_215
rlabel metal2 s 0 85959 624 86007 4 wl_1_216
rlabel metal2 s 0 86213 624 86261 4 wl_1_217
rlabel metal2 s 0 86749 624 86797 4 wl_1_218
rlabel metal2 s 0 87003 624 87051 4 wl_1_219
rlabel metal2 s 0 87539 624 87587 4 wl_1_220
rlabel metal2 s 0 87793 624 87841 4 wl_1_221
rlabel metal2 s 0 88329 624 88377 4 wl_1_222
rlabel metal2 s 0 88583 624 88631 4 wl_1_223
rlabel metal2 s 0 89119 624 89167 4 wl_1_224
rlabel metal2 s 0 89373 624 89421 4 wl_1_225
rlabel metal2 s 0 89909 624 89957 4 wl_1_226
rlabel metal2 s 0 90163 624 90211 4 wl_1_227
rlabel metal2 s 0 90699 624 90747 4 wl_1_228
rlabel metal2 s 0 90953 624 91001 4 wl_1_229
rlabel metal2 s 0 91489 624 91537 4 wl_1_230
rlabel metal2 s 0 91743 624 91791 4 wl_1_231
rlabel metal2 s 0 92279 624 92327 4 wl_1_232
rlabel metal2 s 0 92533 624 92581 4 wl_1_233
rlabel metal2 s 0 93069 624 93117 4 wl_1_234
rlabel metal2 s 0 93323 624 93371 4 wl_1_235
rlabel metal2 s 0 93859 624 93907 4 wl_1_236
rlabel metal2 s 0 94113 624 94161 4 wl_1_237
rlabel metal2 s 0 94649 624 94697 4 wl_1_238
rlabel metal2 s 0 94903 624 94951 4 wl_1_239
rlabel metal2 s 0 95439 624 95487 4 wl_1_240
rlabel metal2 s 0 95693 624 95741 4 wl_1_241
rlabel metal2 s 0 96229 624 96277 4 wl_1_242
rlabel metal2 s 0 96483 624 96531 4 wl_1_243
rlabel metal2 s 0 97019 624 97067 4 wl_1_244
rlabel metal2 s 0 97273 624 97321 4 wl_1_245
rlabel metal2 s 0 97809 624 97857 4 wl_1_246
rlabel metal2 s 0 98063 624 98111 4 wl_1_247
rlabel metal2 s 0 98599 624 98647 4 wl_1_248
rlabel metal2 s 0 98853 624 98901 4 wl_1_249
rlabel metal2 s 0 99389 624 99437 4 wl_1_250
rlabel metal2 s 0 99643 624 99691 4 wl_1_251
rlabel metal2 s 0 100179 624 100227 4 wl_1_252
rlabel metal2 s 0 100433 624 100481 4 wl_1_253
rlabel metal2 s 0 100969 624 101017 4 wl_1_254
rlabel metal2 s 0 101223 624 101271 4 wl_1_255
rlabel metal2 s 0 101759 624 101807 4 wl_1_256
rlabel metal2 s 0 102013 624 102061 4 wl_1_257
rlabel metal1 s 366 869 402 1210 4 vdd
rlabel metal1 s 366 89640 402 89981 4 vdd
rlabel metal1 s 366 100409 402 100750 4 vdd
rlabel metal1 s 366 35920 402 36261 4 vdd
rlabel metal1 s 366 53799 402 54140 4 vdd
rlabel metal1 s 366 58830 402 59171 4 vdd
rlabel metal1 s 366 78289 402 78630 4 vdd
rlabel metal1 s 366 87769 402 88110 4 vdd
rlabel metal1 s 366 20619 402 20960 4 vdd
rlabel metal1 s 366 77499 402 77840 4 vdd
rlabel metal1 s 366 77000 402 77341 4 vdd
rlabel metal1 s 366 101989 402 102330 4 vdd
rlabel metal1 s 366 95170 402 95511 4 vdd
rlabel metal1 s 366 73050 402 73391 4 vdd
rlabel metal1 s 366 99910 402 100251 4 vdd
rlabel metal1 s 366 30099 402 30440 4 vdd
rlabel metal1 s 366 99619 402 99960 4 vdd
rlabel metal1 s 366 85690 402 86031 4 vdd
rlabel metal1 s 366 41949 402 42290 4 vdd
rlabel metal1 s 366 46689 402 47030 4 vdd
rlabel metal1 s 366 25650 402 25991 4 vdd
rlabel metal1 s 366 52510 402 52851 4 vdd
rlabel metal1 s 366 13509 402 13850 4 vdd
rlabel metal1 s 366 26440 402 26781 4 vdd
rlabel metal1 s 366 57749 402 58090 4 vdd
rlabel metal1 s 366 68310 402 68651 4 vdd
rlabel metal1 s 366 20120 402 20461 4 vdd
rlabel metal1 s 366 54589 402 54930 4 vdd
rlabel metal1 s 366 60410 402 60751 4 vdd
rlabel metal1 s 366 84110 402 84451 4 vdd
rlabel metal1 s 366 23280 402 23621 4 vdd
rlabel metal1 s 366 15380 402 15721 4 vdd
rlabel metal1 s 366 97540 402 97881 4 vdd
rlabel metal1 s 366 14590 402 14931 4 vdd
rlabel metal1 s 366 100700 402 101041 4 vdd
rlabel metal1 s 366 69890 402 70231 4 vdd
rlabel metal1 s 366 88850 402 89191 4 vdd
rlabel metal1 s 366 90430 402 90771 4 vdd
rlabel metal1 s 366 33550 402 33891 4 vdd
rlabel metal1 s 366 81740 402 82081 4 vdd
rlabel metal1 s 366 32760 402 33101 4 vdd
rlabel metal1 s 366 39579 402 39920 4 vdd
rlabel metal1 s 366 46190 402 46531 4 vdd
rlabel metal1 s 366 56169 402 56510 4 vdd
rlabel metal1 s 366 80950 402 81291 4 vdd
rlabel metal1 s 366 58040 402 58381 4 vdd
rlabel metal1 s 366 55379 402 55720 4 vdd
rlabel metal1 s 366 40369 402 40710 4 vdd
rlabel metal1 s 366 67520 402 67861 4 vdd
rlabel metal1 s 366 5110 402 5451 4 vdd
rlabel metal1 s 366 43030 402 43371 4 vdd
rlabel metal1 s 366 49849 402 50190 4 vdd
rlabel metal1 s 366 98330 402 98671 4 vdd
rlabel metal1 s 366 43820 402 44161 4 vdd
rlabel metal1 s 366 89349 402 89690 4 vdd
rlabel metal1 s 366 6690 402 7031 4 vdd
rlabel metal1 s 366 86979 402 87320 4 vdd
rlabel metal1 s 366 96750 402 97091 4 vdd
rlabel metal1 s 366 94380 402 94721 4 vdd
rlabel metal1 s 366 30390 402 30731 4 vdd
rlabel metal1 s 366 91719 402 92060 4 vdd
rlabel metal1 s 366 8270 402 8611 4 vdd
rlabel metal1 s 366 71969 402 72310 4 vdd
rlabel metal1 s 366 92800 402 93141 4 vdd
rlabel metal1 s 366 2449 402 2790 4 vdd
rlabel metal1 s 366 52219 402 52560 4 vdd
rlabel metal1 s 366 63570 402 63911 4 vdd
rlabel metal1 s 366 81449 402 81790 4 vdd
rlabel metal3 s 263 180 361 278 4 vdd
rlabel metal1 s 366 49350 402 49691 4 vdd
rlabel metal1 s 366 94879 402 95220 4 vdd
rlabel metal1 s 366 98829 402 99170 4 vdd
rlabel metal1 s 366 26939 402 27280 4 vdd
rlabel metal1 s 366 45109 402 45450 4 vdd
rlabel metal1 s 366 54880 402 55221 4 vdd
rlabel metal1 s 366 66730 402 67071 4 vdd
rlabel metal1 s 366 31679 402 32020 4 vdd
rlabel metal1 s 366 37500 402 37841 4 vdd
rlabel metal1 s 366 65150 402 65491 4 vdd
rlabel metal1 s 366 7189 402 7530 4 vdd
rlabel metal1 s 366 13800 402 14141 4 vdd
rlabel metal1 s 366 47479 402 47820 4 vdd
rlabel metal1 s 366 90139 402 90480 4 vdd
rlabel metal1 s 366 70680 402 71021 4 vdd
rlabel metal1 s 366 71179 402 71520 4 vdd
rlabel metal1 s 366 22490 402 22831 4 vdd
rlabel metal1 s 366 1659 402 2000 4 vdd
rlabel metal1 s 366 30889 402 31230 4 vdd
rlabel metal1 s 366 21700 402 22041 4 vdd
rlabel metal1 s 366 42240 402 42581 4 vdd
rlabel metal1 s 366 48560 402 48901 4 vdd
rlabel metal1 s 366 58539 402 58880 4 vdd
rlabel metal1 s 366 29600 402 29941 4 vdd
rlabel metal1 s 366 11929 402 12270 4 vdd
rlabel metal1 s 366 40660 402 41001 4 vdd
rlabel metal1 s 366 34340 402 34681 4 vdd
rlabel metal1 s 366 36710 402 37051 4 vdd
rlabel metal1 s 366 62780 402 63121 4 vdd
rlabel metal1 s 366 70389 402 70730 4 vdd
rlabel metal1 s 366 35130 402 35471 4 vdd
rlabel metal1 s 366 42739 402 43080 4 vdd
rlabel metal1 s 366 10349 402 10690 4 vdd
rlabel metal1 s 366 95669 402 96010 4 vdd
rlabel metal1 s 366 51429 402 51770 4 vdd
rlabel metal1 s 366 78580 402 78921 4 vdd
rlabel metal1 s 366 19829 402 20170 4 vdd
rlabel metal1 s 366 48269 402 48610 4 vdd
rlabel metal1 s 366 88559 402 88900 4 vdd
rlabel metal1 s 366 50639 402 50980 4 vdd
rlabel metal1 s 366 69599 402 69940 4 vdd
rlabel metal1 s 366 97249 402 97590 4 vdd
rlabel metal1 s 366 60909 402 61250 4 vdd
rlabel metal1 s 366 93299 402 93640 4 vdd
rlabel metal1 s 366 79869 402 80210 4 vdd
rlabel metal1 s 366 88060 402 88401 4 vdd
rlabel metal1 s 366 56460 402 56801 4 vdd
rlabel metal1 s 366 25359 402 25700 4 vdd
rlabel metal1 s 366 83029 402 83370 4 vdd
rlabel metal1 s 366 68809 402 69150 4 vdd
rlabel metal1 s 366 27230 402 27571 4 vdd
rlabel metal1 s 366 28020 402 28361 4 vdd
rlabel metal1 s 366 54090 402 54431 4 vdd
rlabel metal1 s 366 4029 402 4370 4 vdd
rlabel metal1 s 366 28810 402 29151 4 vdd
rlabel metal1 s 366 10640 402 10981 4 vdd
rlabel metal1 s 366 23779 402 24120 4 vdd
rlabel metal1 s 366 18249 402 18590 4 vdd
rlabel metal1 s 366 4819 402 5160 4 vdd
rlabel metal1 s 366 45899 402 46240 4 vdd
rlabel metal1 s 366 11139 402 11480 4 vdd
rlabel metal1 s 366 24070 402 24411 4 vdd
rlabel metal1 s 366 96459 402 96800 4 vdd
rlabel metal1 s 366 3239 402 3580 4 vdd
rlabel metal1 s 366 86189 402 86530 4 vdd
rlabel metal1 s 366 49059 402 49400 4 vdd
rlabel metal1 s 366 75129 402 75470 4 vdd
rlabel metal1 s 366 18540 402 18881 4 vdd
rlabel metal1 s 366 93590 402 93931 4 vdd
rlabel metal1 s 366 53300 402 53641 4 vdd
rlabel metal1 s 366 21409 402 21750 4 vdd
rlabel metal1 s 366 15879 402 16220 4 vdd
rlabel metal1 s 366 16960 402 17301 4 vdd
rlabel metal1 s 366 74339 402 74680 4 vdd
rlabel metal1 s 366 47770 402 48111 4 vdd
rlabel metal1 s 366 67229 402 67570 4 vdd
rlabel metal1 s 366 12719 402 13060 4 vdd
rlabel metal1 s 366 24860 402 25201 4 vdd
rlabel metal1 s 366 45400 402 45741 4 vdd
rlabel metal1 s 366 95960 402 96301 4 vdd
rlabel metal1 s 366 72759 402 73100 4 vdd
rlabel metal1 s 366 11430 402 11771 4 vdd
rlabel metal1 s 366 75420 402 75761 4 vdd
rlabel metal1 s 366 59620 402 59961 4 vdd
rlabel metal1 s 366 22199 402 22540 4 vdd
rlabel metal1 s 366 61699 402 62040 4 vdd
rlabel metal1 s 366 73840 402 74181 4 vdd
rlabel metal1 s 366 16669 402 17010 4 vdd
rlabel metal1 s 366 46980 402 47321 4 vdd
rlabel metal3 s 263 102422 361 102520 4 vdd
rlabel metal1 s 366 94089 402 94430 4 vdd
rlabel metal1 s 366 77790 402 78131 4 vdd
rlabel metal1 s 366 17459 402 17800 4 vdd
rlabel metal1 s 366 12220 402 12561 4 vdd
rlabel metal1 s 366 37209 402 37550 4 vdd
rlabel metal1 s 366 5609 402 5950 4 vdd
rlabel metal1 s 366 36419 402 36760 4 vdd
rlabel metal1 s 366 56959 402 57300 4 vdd
rlabel metal1 s 366 16170 402 16511 4 vdd
rlabel metal1 s 366 90929 402 91270 4 vdd
rlabel metal1 s 366 39080 402 39421 4 vdd
rlabel metal1 s 366 24569 402 24910 4 vdd
rlabel metal1 s 366 27729 402 28070 4 vdd
rlabel metal1 s 366 86480 402 86821 4 vdd
rlabel metal1 s 366 4320 402 4661 4 vdd
rlabel metal1 s 366 51720 402 52061 4 vdd
rlabel metal1 s 366 26149 402 26490 4 vdd
rlabel metal1 s 366 83320 402 83661 4 vdd
rlabel metal1 s 366 1160 402 1501 4 vdd
rlabel metal1 s 366 53009 402 53350 4 vdd
rlabel metal1 s 366 68019 402 68360 4 vdd
rlabel metal1 s 366 1950 402 2291 4 vdd
rlabel metal1 s 366 79370 402 79711 4 vdd
rlabel metal1 s 366 92010 402 92351 4 vdd
rlabel metal1 s 366 19330 402 19671 4 vdd
rlabel metal1 s 366 64069 402 64410 4 vdd
rlabel metal1 s 366 38789 402 39130 4 vdd
rlabel metal1 s 366 61200 402 61541 4 vdd
rlabel metal1 s 366 98039 402 98380 4 vdd
rlabel metal1 s 366 34049 402 34390 4 vdd
rlabel metal1 s 366 19039 402 19380 4 vdd
rlabel metal1 s 366 13010 402 13351 4 vdd
rlabel metal1 s 366 87270 402 87611 4 vdd
rlabel metal1 s 366 61990 402 62331 4 vdd
rlabel metal1 s 366 75919 402 76260 4 vdd
rlabel metal1 s 366 65649 402 65990 4 vdd
rlabel metal1 s 366 66439 402 66780 4 vdd
rlabel metal1 s 366 31180 402 31521 4 vdd
rlabel metal1 s 366 50930 402 51271 4 vdd
rlabel metal1 s 366 62489 402 62830 4 vdd
rlabel metal1 s 366 9060 402 9401 4 vdd
rlabel metal1 s 366 34839 402 35180 4 vdd
rlabel metal1 s 366 38290 402 38631 4 vdd
rlabel metal1 s 366 73549 402 73890 4 vdd
rlabel metal1 s 366 17750 402 18091 4 vdd
rlabel metal1 s 366 82239 402 82580 4 vdd
rlabel metal1 s 366 85399 402 85740 4 vdd
rlabel metal1 s 366 69100 402 69441 4 vdd
rlabel metal1 s 366 65940 402 66281 4 vdd
rlabel metal1 s 366 41450 402 41791 4 vdd
rlabel metal1 s 366 7979 402 8320 4 vdd
rlabel metal1 s 366 41159 402 41500 4 vdd
rlabel metal1 s 366 28519 402 28860 4 vdd
rlabel metal1 s 366 31970 402 32311 4 vdd
rlabel metal1 s 366 44610 402 44951 4 vdd
rlabel metal1 s 366 15089 402 15430 4 vdd
rlabel metal1 s 366 80160 402 80501 4 vdd
rlabel metal1 s 366 83819 402 84160 4 vdd
rlabel metal1 s 366 72260 402 72601 4 vdd
rlabel metal1 s 366 22989 402 23330 4 vdd
rlabel metal1 s 366 64360 402 64701 4 vdd
rlabel metal1 s 366 101199 402 101540 4 vdd
rlabel metal1 s 366 32469 402 32810 4 vdd
rlabel metal1 s 366 37999 402 38340 4 vdd
rlabel metal1 s 366 59329 402 59670 4 vdd
rlabel metal1 s 366 29309 402 29650 4 vdd
rlabel metal1 s 366 76210 402 76551 4 vdd
rlabel metal1 s 366 91220 402 91561 4 vdd
rlabel metal1 s 366 5900 402 6241 4 vdd
rlabel metal1 s 366 33259 402 33600 4 vdd
rlabel metal1 s 366 64859 402 65200 4 vdd
rlabel metal1 s 366 370 402 711 4 vdd
rlabel metal1 s 366 3530 402 3871 4 vdd
rlabel metal1 s 366 76709 402 77050 4 vdd
rlabel metal1 s 366 82530 402 82871 4 vdd
rlabel metal1 s 366 9850 402 10191 4 vdd
rlabel metal1 s 366 80659 402 81000 4 vdd
rlabel metal1 s 366 14299 402 14640 4 vdd
rlabel metal1 s 366 101490 402 101831 4 vdd
rlabel metal1 s 366 7480 402 7821 4 vdd
rlabel metal1 s 366 50140 402 50481 4 vdd
rlabel metal1 s 366 99120 402 99461 4 vdd
rlabel metal1 s 366 6399 402 6740 4 vdd
rlabel metal1 s 366 20910 402 21251 4 vdd
rlabel metal1 s 366 57250 402 57591 4 vdd
rlabel metal1 s 366 84900 402 85241 4 vdd
rlabel metal1 s 366 8769 402 9110 4 vdd
rlabel metal1 s 366 63279 402 63620 4 vdd
rlabel metal1 s 366 92509 402 92850 4 vdd
rlabel metal1 s 366 35629 402 35970 4 vdd
rlabel metal1 s 366 74630 402 74971 4 vdd
rlabel metal1 s 366 39870 402 40211 4 vdd
rlabel metal1 s 366 43529 402 43870 4 vdd
rlabel metal1 s 366 84609 402 84950 4 vdd
rlabel metal1 s 366 60119 402 60460 4 vdd
rlabel metal1 s 366 44319 402 44660 4 vdd
rlabel metal1 s 366 79079 402 79420 4 vdd
rlabel metal1 s 366 2740 402 3081 4 vdd
rlabel metal1 s 366 55670 402 56011 4 vdd
rlabel metal1 s 366 9559 402 9900 4 vdd
rlabel metal1 s 366 71470 402 71811 4 vdd
rlabel metal2 s 330 25225 438 25335 4 gnd
rlabel metal2 s 330 41595 438 41671 4 gnd
rlabel metal2 s 330 6045 438 6121 4 gnd
rlabel metal2 s 330 57869 438 57945 4 gnd
rlabel metal2 s 330 11259 438 11335 4 gnd
rlabel metal2 s 330 69245 438 69321 4 gnd
rlabel metal2 s 330 735 438 845 4 gnd
rlabel metal2 s 330 80525 438 80635 4 gnd
rlabel metal2 s 330 45765 438 45875 4 gnd
rlabel metal2 s 330 71615 438 71691 4 gnd
rlabel metal2 s 330 83939 438 84015 4 gnd
rlabel metal2 s 330 93955 438 94065 4 gnd
rlabel metal2 s 330 16535 438 16645 4 gnd
rlabel metal2 s 330 71045 438 71155 4 gnd
rlabel metal2 s 330 11575 438 11651 4 gnd
rlabel metal2 s 330 77619 438 77695 4 gnd
rlabel metal2 s 330 32115 438 32191 4 gnd
rlabel metal2 s 330 60775 438 60885 4 gnd
rlabel metal2 s 330 79199 438 79275 4 gnd
rlabel metal2 s 330 72625 438 72735 4 gnd
rlabel metal2 s 330 65295 438 65371 4 gnd
rlabel metal2 s 330 43649 438 43725 4 gnd
rlabel metal2 s 330 98695 438 98805 4 gnd
rlabel metal2 s 330 30219 438 30295 4 gnd
rlabel metal2 s 330 5729 438 5805 4 gnd
rlabel metal2 s 330 37645 438 37721 4 gnd
rlabel metal2 s 330 15745 438 15855 4 gnd
rlabel metal2 s 330 14955 438 15065 4 gnd
rlabel metal2 s 330 88995 438 89071 4 gnd
rlabel metal2 s 330 19949 438 20025 4 gnd
rlabel metal2 s 330 87099 438 87175 4 gnd
rlabel metal2 s 330 90005 438 90115 4 gnd
rlabel metal2 s 330 81885 438 81961 4 gnd
rlabel metal2 s 330 64505 438 64581 4 gnd
rlabel metal2 s 330 16315 438 16391 4 gnd
rlabel metal2 s 330 93419 438 93495 4 gnd
rlabel metal2 s 330 4149 438 4225 4 gnd
rlabel metal2 s 330 93735 438 93811 4 gnd
rlabel metal2 s 330 18369 438 18445 4 gnd
rlabel metal2 s 330 76575 438 76685 4 gnd
rlabel metal2 s 330 65769 438 65845 4 gnd
rlabel metal2 s 330 21845 438 21921 4 gnd
rlabel metal2 s 330 4685 438 4795 4 gnd
rlabel metal2 s 330 100055 438 100131 4 gnd
rlabel metal2 s 330 14165 438 14275 4 gnd
rlabel metal2 s 330 48925 438 49035 4 gnd
rlabel metal2 s 330 63715 438 63791 4 gnd
rlabel metal2 s 330 19159 438 19235 4 gnd
rlabel metal2 s 330 94525 438 94601 4 gnd
rlabel metal2 s 330 89469 438 89545 4 gnd
rlabel metal2 s 330 29965 438 30075 4 gnd
rlabel metal2 s 330 55815 438 55891 4 gnd
rlabel metal2 s 330 7845 438 7955 4 gnd
rlabel metal2 s 330 54455 438 54565 4 gnd
rlabel metal2 s 330 1779 438 1855 4 gnd
rlabel metal2 s 330 21275 438 21385 4 gnd
rlabel metal2 s 330 57615 438 57725 4 gnd
rlabel metal2 s 330 59985 438 60095 4 gnd
rlabel metal2 s 330 36539 438 36615 4 gnd
rlabel metal2 s 330 34959 438 35035 4 gnd
rlabel metal2 s 330 91839 438 91915 4 gnd
rlabel metal2 s 330 7055 438 7165 4 gnd
rlabel metal2 s 330 91049 438 91125 4 gnd
rlabel metal2 s 330 39225 438 39301 4 gnd
rlabel metal2 s 330 20265 438 20341 4 gnd
rlabel metal2 s 330 95315 438 95391 4 gnd
rlabel metal2 s 330 75785 438 75895 4 gnd
rlabel metal2 s 330 88425 438 88535 4 gnd
rlabel metal2 s 330 97369 438 97445 4 gnd
rlabel metal2 s 330 25795 438 25871 4 gnd
rlabel metal2 s 330 55245 438 55355 4 gnd
rlabel metal2 s 330 28385 438 28495 4 gnd
rlabel metal2 s 330 8415 438 8491 4 gnd
rlabel metal2 s 330 27595 438 27705 4 gnd
rlabel metal2 s 330 11005 438 11115 4 gnd
rlabel metal2 s 330 3359 438 3435 4 gnd
rlabel metal2 s 330 76829 438 76905 4 gnd
rlabel metal2 s 330 43965 438 44041 4 gnd
rlabel metal2 s 330 48389 438 48465 4 gnd
rlabel metal2 s 330 18905 438 19015 4 gnd
rlabel metal2 s 330 24215 438 24291 4 gnd
rlabel metal2 s 330 15525 438 15601 4 gnd
rlabel metal2 s 330 25479 438 25555 4 gnd
rlabel metal2 s 330 50759 438 50835 4 gnd
rlabel metal2 s 330 99265 438 99341 4 gnd
rlabel metal2 s 330 68139 438 68215 4 gnd
rlabel metal2 s 330 37865 438 37975 4 gnd
rlabel metal2 s 330 28165 438 28241 4 gnd
rlabel metal2 s 330 77365 438 77475 4 gnd
rlabel metal2 s 330 7625 438 7701 4 gnd
rlabel metal2 s 330 98475 438 98551 4 gnd
rlabel metal2 s 330 51865 438 51941 4 gnd
rlabel metal2 s 330 56289 438 56365 4 gnd
rlabel metal2 s 330 67095 438 67205 4 gnd
rlabel metal2 s 330 73415 438 73525 4 gnd
rlabel metal2 s 330 52085 438 52195 4 gnd
rlabel metal2 s 330 44185 438 44295 4 gnd
rlabel metal2 s 330 89215 438 89325 4 gnd
rlabel metal2 s 330 58659 438 58735 4 gnd
rlabel metal2 s 330 32589 438 32665 4 gnd
rlabel metal2 s 330 24689 438 24765 4 gnd
rlabel metal2 s 330 22635 438 22711 4 gnd
rlabel metal2 s 330 101065 438 101175 4 gnd
rlabel metal2 s 330 62355 438 62465 4 gnd
rlabel metal2 s 330 86309 438 86385 4 gnd
rlabel metal2 s 330 93165 438 93275 4 gnd
rlabel metal2 s 330 63145 438 63255 4 gnd
rlabel metal2 s 330 46335 438 46411 4 gnd
rlabel metal2 s 330 50285 438 50361 4 gnd
rlabel metal2 s 330 77935 438 78011 4 gnd
rlabel metal2 s 330 54235 438 54311 4 gnd
rlabel metal2 s 330 75565 438 75641 4 gnd
rlabel metal2 s 330 20739 438 20815 4 gnd
rlabel metal2 s 330 20485 438 20595 4 gnd
rlabel metal2 s 330 31009 438 31085 4 gnd
rlabel metal2 s 330 83685 438 83795 4 gnd
rlabel metal2 s 330 23425 438 23501 4 gnd
rlabel metal2 s 330 40235 438 40345 4 gnd
rlabel metal2 s 330 8635 438 8745 4 gnd
rlabel metal2 s 330 72089 438 72165 4 gnd
rlabel metal2 s 330 73669 438 73745 4 gnd
rlabel metal2 s 330 41815 438 41925 4 gnd
rlabel metal2 s 330 89785 438 89861 4 gnd
rlabel metal2 s 330 26015 438 26125 4 gnd
rlabel metal2 s 330 53665 438 53775 4 gnd
rlabel metal2 s 330 46555 438 46665 4 gnd
rlabel metal2 s 330 62925 438 63001 4 gnd
rlabel metal2 s 330 35749 438 35825 4 gnd
rlabel metal2 s 330 95535 438 95645 4 gnd
rlabel metal2 s 330 41279 438 41355 4 gnd
rlabel metal2 s 330 68929 438 69005 4 gnd
rlabel metal2 s 330 26805 438 26915 4 gnd
rlabel metal2 s 330 74205 438 74315 4 gnd
rlabel metal2 s 330 10469 438 10545 4 gnd
rlabel metal2 s 330 61345 438 61421 4 gnd
rlabel metal2 s 330 84255 438 84331 4 gnd
rlabel metal2 s 330 1525 438 1635 4 gnd
rlabel metal2 s 330 23899 438 23975 4 gnd
rlabel metal2 s 330 58185 438 58261 4 gnd
rlabel metal2 s 330 82675 438 82751 4 gnd
rlabel metal2 s 330 38909 438 38985 4 gnd
rlabel metal2 s 330 35275 438 35351 4 gnd
rlabel metal2 s 330 21529 438 21605 4 gnd
rlabel metal2 s 330 52655 438 52731 4 gnd
rlabel metal2 s 330 15999 438 16075 4 gnd
rlabel metal2 s 330 22855 438 22965 4 gnd
rlabel metal2 s 330 9425 438 9535 4 gnd
rlabel metal2 s 330 56035 438 56145 4 gnd
rlabel metal2 s 330 41025 438 41135 4 gnd
rlabel metal2 s 330 12049 438 12125 4 gnd
rlabel metal2 s 330 44975 438 45085 4 gnd
rlabel metal2 s 330 68455 438 68531 4 gnd
rlabel metal2 s 330 64979 438 65055 4 gnd
rlabel metal2 s 330 90575 438 90651 4 gnd
rlabel metal2 s 330 26269 438 26345 4 gnd
rlabel metal2 s 330 43395 438 43505 4 gnd
rlabel metal2 s 330 71835 438 71945 4 gnd
rlabel metal2 s 330 100845 438 100921 4 gnd
rlabel metal2 s 330 17895 438 17971 4 gnd
rlabel metal2 s 330 44755 438 44831 4 gnd
rlabel metal2 s 330 78725 438 78801 4 gnd
rlabel metal2 s 330 2095 438 2171 4 gnd
rlabel metal2 s 330 66305 438 66415 4 gnd
rlabel metal2 s 330 83465 438 83541 4 gnd
rlabel metal2 s 330 30535 438 30611 4 gnd
rlabel metal2 s 330 75249 438 75325 4 gnd
rlabel metal2 s 330 85045 438 85121 4 gnd
rlabel metal2 s 330 14419 438 14495 4 gnd
rlabel metal2 s 330 66085 438 66161 4 gnd
rlabel metal2 s 330 58975 438 59051 4 gnd
rlabel metal2 s 330 27849 438 27925 4 gnd
rlabel metal2 s 330 36855 438 36931 4 gnd
rlabel metal2 s 330 88679 438 88755 4 gnd
rlabel metal2 s 330 59765 438 59841 4 gnd
rlabel metal2 s 330 42605 438 42715 4 gnd
rlabel metal2 s 330 72405 438 72481 4 gnd
rlabel metal2 s 330 87635 438 87745 4 gnd
rlabel metal2 s 330 42385 438 42461 4 gnd
rlabel metal2 s 330 90795 438 90905 4 gnd
rlabel metal2 s 330 37075 438 37185 4 gnd
rlabel metal2 s 330 96325 438 96435 4 gnd
rlabel metal2 s 330 33125 438 33235 4 gnd
rlabel metal2 s 330 79989 438 80065 4 gnd
rlabel metal2 s 330 9995 438 10071 4 gnd
rlabel metal2 s 330 34169 438 34245 4 gnd
rlabel metal2 s 330 22319 438 22395 4 gnd
rlabel metal2 s 330 94999 438 95075 4 gnd
rlabel metal2 s 330 8099 438 8175 4 gnd
rlabel metal2 s 330 55025 438 55101 4 gnd
rlabel metal2 s 330 65515 438 65625 4 gnd
rlabel metal2 s 330 52339 438 52415 4 gnd
rlabel metal2 s 330 92155 438 92231 4 gnd
rlabel metal2 s 330 23109 438 23185 4 gnd
rlabel metal2 s 330 96105 438 96181 4 gnd
rlabel metal2 s 330 79735 438 79845 4 gnd
rlabel metal2 s 330 86055 438 86165 4 gnd
rlabel metal2 s 330 32335 438 32445 4 gnd
rlabel metal2 s 330 21055 438 21131 4 gnd
rlabel metal2 s 330 1305 438 1381 4 gnd
rlabel metal2 s 330 45545 438 45621 4 gnd
rlabel metal2 s 330 4939 438 5015 4 gnd
rlabel metal2 s 330 33379 438 33455 4 gnd
rlabel metal2 s 330 63935 438 64045 4 gnd
rlabel metal2 s 330 19695 438 19805 4 gnd
rlabel metal2 s 330 53445 438 53521 4 gnd
rlabel metal2 s 330 35495 438 35605 4 gnd
rlabel metal2 s 330 78409 438 78485 4 gnd
rlabel metal2 s 330 14735 438 14811 4 gnd
rlabel metal2 s 330 81095 438 81171 4 gnd
rlabel metal2 s 330 96579 438 96655 4 gnd
rlabel metal2 s 330 79515 438 79591 4 gnd
rlabel metal2 s 330 34705 438 34815 4 gnd
rlabel metal2 s 330 49179 438 49255 4 gnd
rlabel metal2 s 330 45229 438 45305 4 gnd
rlabel metal2 s 330 61819 438 61895 4 gnd
rlabel metal2 s 330 5475 438 5585 4 gnd
rlabel metal2 s 330 47915 438 47991 4 gnd
rlabel metal2 s 330 77145 438 77221 4 gnd
rlabel metal2 s 330 92945 438 93021 4 gnd
rlabel metal2 s 330 13375 438 13485 4 gnd
rlabel metal2 s 330 58405 438 58515 4 gnd
rlabel metal2 s 330 37329 438 37405 4 gnd
rlabel metal2 s 330 32905 438 32981 4 gnd
rlabel metal2 s 330 87889 438 87965 4 gnd
rlabel metal2 s 330 28639 438 28715 4 gnd
rlabel metal2 s 330 17105 438 17181 4 gnd
rlabel metal2 s 330 88205 438 88281 4 gnd
rlabel metal2 s 330 7309 438 7385 4 gnd
rlabel metal2 s 330 38655 438 38765 4 gnd
rlabel metal2 s 330 6519 438 6595 4 gnd
rlabel metal2 s 330 52875 438 52985 4 gnd
rlabel metal2 s 330 51295 438 51405 4 gnd
rlabel metal2 s 330 67885 438 67995 4 gnd
rlabel metal2 s 330 73195 438 73271 4 gnd
rlabel metal2 s 330 68675 438 68785 4 gnd
rlabel metal2 s 330 9205 438 9281 4 gnd
rlabel metal2 s 330 9679 438 9755 4 gnd
rlabel metal2 s 330 29175 438 29285 4 gnd
rlabel metal2 s 330 42859 438 42935 4 gnd
rlabel metal2 s 330 3105 438 3215 4 gnd
rlabel metal2 s 330 94745 438 94855 4 gnd
rlabel metal2 s 330 15209 438 15285 4 gnd
rlabel metal2 s 330 27375 438 27451 4 gnd
rlabel metal2 s 330 25005 438 25081 4 gnd
rlabel metal2 s 330 60555 438 60631 4 gnd
rlabel metal2 s 330 69465 438 69575 4 gnd
rlabel metal2 s 330 8889 438 8965 4 gnd
rlabel metal2 s 330 39699 438 39775 4 gnd
rlabel metal2 s 330 97115 438 97225 4 gnd
rlabel metal2 s 330 17579 438 17655 4 gnd
rlabel metal2 s 330 50505 438 50615 4 gnd
rlabel metal2 s 330 38435 438 38511 4 gnd
rlabel metal2 s 330 60239 438 60315 4 gnd
rlabel metal2 s 330 80305 438 80381 4 gnd
rlabel metal2 s 330 10215 438 10325 4 gnd
rlabel metal2 s 330 18685 438 18761 4 gnd
rlabel metal2 s 330 22065 438 22175 4 gnd
rlabel metal2 s 330 56605 438 56681 4 gnd
rlabel metal2 s 330 48135 438 48245 4 gnd
rlabel metal2 s 330 78945 438 79055 4 gnd
rlabel metal2 s 330 4465 438 4541 4 gnd
rlabel metal2 s 330 72879 438 72955 4 gnd
rlabel metal2 s 330 6835 438 6911 4 gnd
rlabel metal2 s 330 29745 438 29821 4 gnd
rlabel metal2 s 330 12839 438 12915 4 gnd
rlabel metal2 s 330 96895 438 96971 4 gnd
rlabel metal2 s 330 2885 438 2961 4 gnd
rlabel metal2 s 330 90259 438 90335 4 gnd
rlabel metal2 s 330 33915 438 34025 4 gnd
rlabel metal2 s 330 43175 438 43251 4 gnd
rlabel metal2 s 330 74775 438 74851 4 gnd
rlabel metal2 s 330 84475 438 84585 4 gnd
rlabel metal2 s 330 101855 438 101965 4 gnd
rlabel metal2 s 330 44439 438 44515 4 gnd
rlabel metal2 s 330 5255 438 5331 4 gnd
rlabel metal2 s 330 2315 438 2425 4 gnd
rlabel metal2 s 330 85265 438 85375 4 gnd
rlabel metal2 s 330 49495 438 49571 4 gnd
rlabel metal2 s 330 100275 438 100385 4 gnd
rlabel metal2 s 330 3675 438 3751 4 gnd
rlabel metal2 s 330 59195 438 59305 4 gnd
rlabel metal2 s 330 31545 438 31655 4 gnd
rlabel metal2 s 330 40015 438 40091 4 gnd
rlabel metal2 s 330 11795 438 11905 4 gnd
rlabel metal2 s 330 67665 438 67741 4 gnd
rlabel metal2 s 330 97905 438 98015 4 gnd
rlabel metal2 s 330 98949 438 99025 4 gnd
rlabel metal2 s 330 70825 438 70901 4 gnd
rlabel metal2 s 330 39445 438 39555 4 gnd
rlabel metal2 s 330 23645 438 23755 4 gnd
rlabel metal2 s 330 82359 438 82435 4 gnd
rlabel metal2 s 330 10785 438 10861 4 gnd
rlabel metal2 s 330 84729 438 84805 4 gnd
rlabel metal2 s 330 53129 438 53205 4 gnd
rlabel metal2 s 330 6265 438 6375 4 gnd
rlabel metal2 s 330 64725 438 64835 4 gnd
rlabel metal2 s 330 47599 438 47675 4 gnd
rlabel metal2 s 330 47125 438 47201 4 gnd
rlabel metal2 s 330 94209 438 94285 4 gnd
rlabel metal2 s 330 71299 438 71375 4 gnd
rlabel metal2 s 330 54709 438 54785 4 gnd
rlabel metal2 s 330 74995 438 75105 4 gnd
rlabel metal2 s 330 59449 438 59525 4 gnd
rlabel metal2 s 330 51549 438 51625 4 gnd
rlabel metal2 s 330 13155 438 13231 4 gnd
rlabel metal2 s 330 55499 438 55575 4 gnd
rlabel metal2 s 330 33695 438 33771 4 gnd
rlabel metal2 s 330 101319 438 101395 4 gnd
rlabel metal2 s 330 91585 438 91695 4 gnd
rlabel metal2 s 330 92375 438 92485 4 gnd
rlabel metal2 s 330 99485 438 99595 4 gnd
rlabel metal2 s 330 61565 438 61675 4 gnd
rlabel metal2 s 330 85519 438 85595 4 gnd
rlabel metal2 s 330 62135 438 62211 4 gnd
rlabel metal2 s 330 49715 438 49825 4 gnd
rlabel metal2 s 330 64189 438 64265 4 gnd
rlabel metal2 s 330 515 438 591 4 gnd
rlabel metal2 s 330 34485 438 34561 4 gnd
rlabel metal2 s 330 40805 438 40881 4 gnd
rlabel metal2 s 330 70255 438 70365 4 gnd
rlabel metal2 s 330 100529 438 100605 4 gnd
rlabel metal2 s 330 73985 438 74061 4 gnd
rlabel metal2 s 330 63399 438 63475 4 gnd
rlabel metal2 s 330 27059 438 27135 4 gnd
rlabel metal2 s 330 36065 438 36141 4 gnd
rlabel metal2 s 330 49969 438 50045 4 gnd
rlabel metal2 s 330 82895 438 83005 4 gnd
rlabel metal2 s 330 95789 438 95865 4 gnd
rlabel metal2 s 330 13629 438 13705 4 gnd
rlabel metal2 s 330 19475 438 19551 4 gnd
rlabel metal2 s 330 87415 438 87491 4 gnd
rlabel metal2 s 330 78155 438 78265 4 gnd
rlabel metal2 s 330 28955 438 29031 4 gnd
rlabel metal2 s 330 17325 438 17435 4 gnd
rlabel metal2 s 330 57395 438 57471 4 gnd
rlabel metal2 s 330 3895 438 4005 4 gnd
rlabel metal2 s 330 47345 438 47455 4 gnd
rlabel metal2 s 330 51075 438 51151 4 gnd
rlabel metal2 s 330 66875 438 66951 4 gnd
rlabel metal2 s 330 30755 438 30865 4 gnd
rlabel metal2 s 330 29429 438 29505 4 gnd
rlabel metal2 s 330 86625 438 86701 4 gnd
rlabel metal2 s 330 86845 438 86955 4 gnd
rlabel metal2 s 330 53919 438 53995 4 gnd
rlabel metal2 s 330 74459 438 74535 4 gnd
rlabel metal2 s 330 101635 438 101711 4 gnd
rlabel metal2 s 330 76355 438 76431 4 gnd
rlabel metal2 s 330 46809 438 46885 4 gnd
rlabel metal2 s 330 26585 438 26661 4 gnd
rlabel metal2 s 330 92629 438 92705 4 gnd
rlabel metal2 s 330 40489 438 40565 4 gnd
rlabel metal2 s 330 76039 438 76115 4 gnd
rlabel metal2 s 330 82105 438 82215 4 gnd
rlabel metal2 s 330 97685 438 97761 4 gnd
rlabel metal2 s 330 36285 438 36395 4 gnd
rlabel metal2 s 330 83149 438 83225 4 gnd
rlabel metal2 s 330 56825 438 56935 4 gnd
rlabel metal2 s 330 62609 438 62685 4 gnd
rlabel metal2 s 330 48705 438 48781 4 gnd
rlabel metal2 s 330 42069 438 42145 4 gnd
rlabel metal2 s 330 12585 438 12695 4 gnd
rlabel metal2 s 330 61029 438 61105 4 gnd
rlabel metal2 s 330 31799 438 31875 4 gnd
rlabel metal2 s 330 69719 438 69795 4 gnd
rlabel metal2 s 330 85835 438 85911 4 gnd
rlabel metal2 s 330 2569 438 2645 4 gnd
rlabel metal2 s 330 46019 438 46095 4 gnd
rlabel metal2 s 330 70035 438 70111 4 gnd
rlabel metal2 s 330 91365 438 91441 4 gnd
rlabel metal2 s 330 989 438 1065 4 gnd
rlabel metal2 s 330 81315 438 81425 4 gnd
rlabel metal2 s 330 98159 438 98235 4 gnd
rlabel metal2 s 330 31325 438 31401 4 gnd
rlabel metal2 s 330 66559 438 66635 4 gnd
rlabel metal2 s 330 102109 438 102185 4 gnd
rlabel metal2 s 330 18115 438 18225 4 gnd
rlabel metal2 s 330 70509 438 70585 4 gnd
rlabel metal2 s 330 67349 438 67425 4 gnd
rlabel metal2 s 330 38119 438 38195 4 gnd
rlabel metal2 s 330 13945 438 14021 4 gnd
rlabel metal2 s 330 12365 438 12441 4 gnd
rlabel metal2 s 330 57079 438 57155 4 gnd
rlabel metal2 s 330 99739 438 99815 4 gnd
rlabel metal2 s 330 16789 438 16865 4 gnd
rlabel metal2 s 330 80779 438 80855 4 gnd
rlabel metal2 s 330 81569 438 81645 4 gnd
rlabel metal2 s 330 24435 438 24545 4 gnd
<< properties >>
string FIXED_BBOX 0 0 624 102700
<< end >>
