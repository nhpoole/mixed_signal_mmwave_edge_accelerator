magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< error_p >>
rect -4187 -900 4187 900
<< nwell >>
rect -4187 -900 4187 900
<< pmoshvt >>
rect -4093 -800 -3693 800
rect -3635 -800 -3235 800
rect -3177 -800 -2777 800
rect -2719 -800 -2319 800
rect -2261 -800 -1861 800
rect -1803 -800 -1403 800
rect -1345 -800 -945 800
rect -887 -800 -487 800
rect -429 -800 -29 800
rect 29 -800 429 800
rect 487 -800 887 800
rect 945 -800 1345 800
rect 1403 -800 1803 800
rect 1861 -800 2261 800
rect 2319 -800 2719 800
rect 2777 -800 3177 800
rect 3235 -800 3635 800
rect 3693 -800 4093 800
<< pdiff >>
rect -4151 788 -4093 800
rect -4151 -788 -4139 788
rect -4105 -788 -4093 788
rect -4151 -800 -4093 -788
rect -3693 788 -3635 800
rect -3693 -788 -3681 788
rect -3647 -788 -3635 788
rect -3693 -800 -3635 -788
rect -3235 788 -3177 800
rect -3235 -788 -3223 788
rect -3189 -788 -3177 788
rect -3235 -800 -3177 -788
rect -2777 788 -2719 800
rect -2777 -788 -2765 788
rect -2731 -788 -2719 788
rect -2777 -800 -2719 -788
rect -2319 788 -2261 800
rect -2319 -788 -2307 788
rect -2273 -788 -2261 788
rect -2319 -800 -2261 -788
rect -1861 788 -1803 800
rect -1861 -788 -1849 788
rect -1815 -788 -1803 788
rect -1861 -800 -1803 -788
rect -1403 788 -1345 800
rect -1403 -788 -1391 788
rect -1357 -788 -1345 788
rect -1403 -800 -1345 -788
rect -945 788 -887 800
rect -945 -788 -933 788
rect -899 -788 -887 788
rect -945 -800 -887 -788
rect -487 788 -429 800
rect -487 -788 -475 788
rect -441 -788 -429 788
rect -487 -800 -429 -788
rect -29 788 29 800
rect -29 -788 -17 788
rect 17 -788 29 788
rect -29 -800 29 -788
rect 429 788 487 800
rect 429 -788 441 788
rect 475 -788 487 788
rect 429 -800 487 -788
rect 887 788 945 800
rect 887 -788 899 788
rect 933 -788 945 788
rect 887 -800 945 -788
rect 1345 788 1403 800
rect 1345 -788 1357 788
rect 1391 -788 1403 788
rect 1345 -800 1403 -788
rect 1803 788 1861 800
rect 1803 -788 1815 788
rect 1849 -788 1861 788
rect 1803 -800 1861 -788
rect 2261 788 2319 800
rect 2261 -788 2273 788
rect 2307 -788 2319 788
rect 2261 -800 2319 -788
rect 2719 788 2777 800
rect 2719 -788 2731 788
rect 2765 -788 2777 788
rect 2719 -800 2777 -788
rect 3177 788 3235 800
rect 3177 -788 3189 788
rect 3223 -788 3235 788
rect 3177 -800 3235 -788
rect 3635 788 3693 800
rect 3635 -788 3647 788
rect 3681 -788 3693 788
rect 3635 -800 3693 -788
rect 4093 788 4151 800
rect 4093 -788 4105 788
rect 4139 -788 4151 788
rect 4093 -800 4151 -788
<< pdiffc >>
rect -4139 -788 -4105 788
rect -3681 -788 -3647 788
rect -3223 -788 -3189 788
rect -2765 -788 -2731 788
rect -2307 -788 -2273 788
rect -1849 -788 -1815 788
rect -1391 -788 -1357 788
rect -933 -788 -899 788
rect -475 -788 -441 788
rect -17 -788 17 788
rect 441 -788 475 788
rect 899 -788 933 788
rect 1357 -788 1391 788
rect 1815 -788 1849 788
rect 2273 -788 2307 788
rect 2731 -788 2765 788
rect 3189 -788 3223 788
rect 3647 -788 3681 788
rect 4105 -788 4139 788
<< poly >>
rect -4019 881 -3767 897
rect -4019 864 -4003 881
rect -4093 847 -4003 864
rect -3783 864 -3767 881
rect -3561 881 -3309 897
rect -3561 864 -3545 881
rect -3783 847 -3693 864
rect -4093 800 -3693 847
rect -3635 847 -3545 864
rect -3325 864 -3309 881
rect -3103 881 -2851 897
rect -3103 864 -3087 881
rect -3325 847 -3235 864
rect -3635 800 -3235 847
rect -3177 847 -3087 864
rect -2867 864 -2851 881
rect -2645 881 -2393 897
rect -2645 864 -2629 881
rect -2867 847 -2777 864
rect -3177 800 -2777 847
rect -2719 847 -2629 864
rect -2409 864 -2393 881
rect -2187 881 -1935 897
rect -2187 864 -2171 881
rect -2409 847 -2319 864
rect -2719 800 -2319 847
rect -2261 847 -2171 864
rect -1951 864 -1935 881
rect -1729 881 -1477 897
rect -1729 864 -1713 881
rect -1951 847 -1861 864
rect -2261 800 -1861 847
rect -1803 847 -1713 864
rect -1493 864 -1477 881
rect -1271 881 -1019 897
rect -1271 864 -1255 881
rect -1493 847 -1403 864
rect -1803 800 -1403 847
rect -1345 847 -1255 864
rect -1035 864 -1019 881
rect -813 881 -561 897
rect -813 864 -797 881
rect -1035 847 -945 864
rect -1345 800 -945 847
rect -887 847 -797 864
rect -577 864 -561 881
rect -355 881 -103 897
rect -355 864 -339 881
rect -577 847 -487 864
rect -887 800 -487 847
rect -429 847 -339 864
rect -119 864 -103 881
rect 103 881 355 897
rect 103 864 119 881
rect -119 847 -29 864
rect -429 800 -29 847
rect 29 847 119 864
rect 339 864 355 881
rect 561 881 813 897
rect 561 864 577 881
rect 339 847 429 864
rect 29 800 429 847
rect 487 847 577 864
rect 797 864 813 881
rect 1019 881 1271 897
rect 1019 864 1035 881
rect 797 847 887 864
rect 487 800 887 847
rect 945 847 1035 864
rect 1255 864 1271 881
rect 1477 881 1729 897
rect 1477 864 1493 881
rect 1255 847 1345 864
rect 945 800 1345 847
rect 1403 847 1493 864
rect 1713 864 1729 881
rect 1935 881 2187 897
rect 1935 864 1951 881
rect 1713 847 1803 864
rect 1403 800 1803 847
rect 1861 847 1951 864
rect 2171 864 2187 881
rect 2393 881 2645 897
rect 2393 864 2409 881
rect 2171 847 2261 864
rect 1861 800 2261 847
rect 2319 847 2409 864
rect 2629 864 2645 881
rect 2851 881 3103 897
rect 2851 864 2867 881
rect 2629 847 2719 864
rect 2319 800 2719 847
rect 2777 847 2867 864
rect 3087 864 3103 881
rect 3309 881 3561 897
rect 3309 864 3325 881
rect 3087 847 3177 864
rect 2777 800 3177 847
rect 3235 847 3325 864
rect 3545 864 3561 881
rect 3767 881 4019 897
rect 3767 864 3783 881
rect 3545 847 3635 864
rect 3235 800 3635 847
rect 3693 847 3783 864
rect 4003 864 4019 881
rect 4003 847 4093 864
rect 3693 800 4093 847
rect -4093 -847 -3693 -800
rect -4093 -864 -4003 -847
rect -4019 -881 -4003 -864
rect -3783 -864 -3693 -847
rect -3635 -847 -3235 -800
rect -3635 -864 -3545 -847
rect -3783 -881 -3767 -864
rect -4019 -897 -3767 -881
rect -3561 -881 -3545 -864
rect -3325 -864 -3235 -847
rect -3177 -847 -2777 -800
rect -3177 -864 -3087 -847
rect -3325 -881 -3309 -864
rect -3561 -897 -3309 -881
rect -3103 -881 -3087 -864
rect -2867 -864 -2777 -847
rect -2719 -847 -2319 -800
rect -2719 -864 -2629 -847
rect -2867 -881 -2851 -864
rect -3103 -897 -2851 -881
rect -2645 -881 -2629 -864
rect -2409 -864 -2319 -847
rect -2261 -847 -1861 -800
rect -2261 -864 -2171 -847
rect -2409 -881 -2393 -864
rect -2645 -897 -2393 -881
rect -2187 -881 -2171 -864
rect -1951 -864 -1861 -847
rect -1803 -847 -1403 -800
rect -1803 -864 -1713 -847
rect -1951 -881 -1935 -864
rect -2187 -897 -1935 -881
rect -1729 -881 -1713 -864
rect -1493 -864 -1403 -847
rect -1345 -847 -945 -800
rect -1345 -864 -1255 -847
rect -1493 -881 -1477 -864
rect -1729 -897 -1477 -881
rect -1271 -881 -1255 -864
rect -1035 -864 -945 -847
rect -887 -847 -487 -800
rect -887 -864 -797 -847
rect -1035 -881 -1019 -864
rect -1271 -897 -1019 -881
rect -813 -881 -797 -864
rect -577 -864 -487 -847
rect -429 -847 -29 -800
rect -429 -864 -339 -847
rect -577 -881 -561 -864
rect -813 -897 -561 -881
rect -355 -881 -339 -864
rect -119 -864 -29 -847
rect 29 -847 429 -800
rect 29 -864 119 -847
rect -119 -881 -103 -864
rect -355 -897 -103 -881
rect 103 -881 119 -864
rect 339 -864 429 -847
rect 487 -847 887 -800
rect 487 -864 577 -847
rect 339 -881 355 -864
rect 103 -897 355 -881
rect 561 -881 577 -864
rect 797 -864 887 -847
rect 945 -847 1345 -800
rect 945 -864 1035 -847
rect 797 -881 813 -864
rect 561 -897 813 -881
rect 1019 -881 1035 -864
rect 1255 -864 1345 -847
rect 1403 -847 1803 -800
rect 1403 -864 1493 -847
rect 1255 -881 1271 -864
rect 1019 -897 1271 -881
rect 1477 -881 1493 -864
rect 1713 -864 1803 -847
rect 1861 -847 2261 -800
rect 1861 -864 1951 -847
rect 1713 -881 1729 -864
rect 1477 -897 1729 -881
rect 1935 -881 1951 -864
rect 2171 -864 2261 -847
rect 2319 -847 2719 -800
rect 2319 -864 2409 -847
rect 2171 -881 2187 -864
rect 1935 -897 2187 -881
rect 2393 -881 2409 -864
rect 2629 -864 2719 -847
rect 2777 -847 3177 -800
rect 2777 -864 2867 -847
rect 2629 -881 2645 -864
rect 2393 -897 2645 -881
rect 2851 -881 2867 -864
rect 3087 -864 3177 -847
rect 3235 -847 3635 -800
rect 3235 -864 3325 -847
rect 3087 -881 3103 -864
rect 2851 -897 3103 -881
rect 3309 -881 3325 -864
rect 3545 -864 3635 -847
rect 3693 -847 4093 -800
rect 3693 -864 3783 -847
rect 3545 -881 3561 -864
rect 3309 -897 3561 -881
rect 3767 -881 3783 -864
rect 4003 -864 4093 -847
rect 4003 -881 4019 -864
rect 3767 -897 4019 -881
<< polycont >>
rect -4003 847 -3783 881
rect -3545 847 -3325 881
rect -3087 847 -2867 881
rect -2629 847 -2409 881
rect -2171 847 -1951 881
rect -1713 847 -1493 881
rect -1255 847 -1035 881
rect -797 847 -577 881
rect -339 847 -119 881
rect 119 847 339 881
rect 577 847 797 881
rect 1035 847 1255 881
rect 1493 847 1713 881
rect 1951 847 2171 881
rect 2409 847 2629 881
rect 2867 847 3087 881
rect 3325 847 3545 881
rect 3783 847 4003 881
rect -4003 -881 -3783 -847
rect -3545 -881 -3325 -847
rect -3087 -881 -2867 -847
rect -2629 -881 -2409 -847
rect -2171 -881 -1951 -847
rect -1713 -881 -1493 -847
rect -1255 -881 -1035 -847
rect -797 -881 -577 -847
rect -339 -881 -119 -847
rect 119 -881 339 -847
rect 577 -881 797 -847
rect 1035 -881 1255 -847
rect 1493 -881 1713 -847
rect 1951 -881 2171 -847
rect 2409 -881 2629 -847
rect 2867 -881 3087 -847
rect 3325 -881 3545 -847
rect 3783 -881 4003 -847
<< locali >>
rect -4019 847 -4003 881
rect -3783 847 -3767 881
rect -3561 847 -3545 881
rect -3325 847 -3309 881
rect -3103 847 -3087 881
rect -2867 847 -2851 881
rect -2645 847 -2629 881
rect -2409 847 -2393 881
rect -2187 847 -2171 881
rect -1951 847 -1935 881
rect -1729 847 -1713 881
rect -1493 847 -1477 881
rect -1271 847 -1255 881
rect -1035 847 -1019 881
rect -813 847 -797 881
rect -577 847 -561 881
rect -355 847 -339 881
rect -119 847 -103 881
rect 103 847 119 881
rect 339 847 355 881
rect 561 847 577 881
rect 797 847 813 881
rect 1019 847 1035 881
rect 1255 847 1271 881
rect 1477 847 1493 881
rect 1713 847 1729 881
rect 1935 847 1951 881
rect 2171 847 2187 881
rect 2393 847 2409 881
rect 2629 847 2645 881
rect 2851 847 2867 881
rect 3087 847 3103 881
rect 3309 847 3325 881
rect 3545 847 3561 881
rect 3767 847 3783 881
rect 4003 847 4019 881
rect -4139 788 -4105 804
rect -4139 -804 -4105 -788
rect -3681 788 -3647 804
rect -3681 -804 -3647 -788
rect -3223 788 -3189 804
rect -3223 -804 -3189 -788
rect -2765 788 -2731 804
rect -2765 -804 -2731 -788
rect -2307 788 -2273 804
rect -2307 -804 -2273 -788
rect -1849 788 -1815 804
rect -1849 -804 -1815 -788
rect -1391 788 -1357 804
rect -1391 -804 -1357 -788
rect -933 788 -899 804
rect -933 -804 -899 -788
rect -475 788 -441 804
rect -475 -804 -441 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 441 788 475 804
rect 441 -804 475 -788
rect 899 788 933 804
rect 899 -804 933 -788
rect 1357 788 1391 804
rect 1357 -804 1391 -788
rect 1815 788 1849 804
rect 1815 -804 1849 -788
rect 2273 788 2307 804
rect 2273 -804 2307 -788
rect 2731 788 2765 804
rect 2731 -804 2765 -788
rect 3189 788 3223 804
rect 3189 -804 3223 -788
rect 3647 788 3681 804
rect 3647 -804 3681 -788
rect 4105 788 4139 804
rect 4105 -804 4139 -788
rect -4019 -881 -4003 -847
rect -3783 -881 -3767 -847
rect -3561 -881 -3545 -847
rect -3325 -881 -3309 -847
rect -3103 -881 -3087 -847
rect -2867 -881 -2851 -847
rect -2645 -881 -2629 -847
rect -2409 -881 -2393 -847
rect -2187 -881 -2171 -847
rect -1951 -881 -1935 -847
rect -1729 -881 -1713 -847
rect -1493 -881 -1477 -847
rect -1271 -881 -1255 -847
rect -1035 -881 -1019 -847
rect -813 -881 -797 -847
rect -577 -881 -561 -847
rect -355 -881 -339 -847
rect -119 -881 -103 -847
rect 103 -881 119 -847
rect 339 -881 355 -847
rect 561 -881 577 -847
rect 797 -881 813 -847
rect 1019 -881 1035 -847
rect 1255 -881 1271 -847
rect 1477 -881 1493 -847
rect 1713 -881 1729 -847
rect 1935 -881 1951 -847
rect 2171 -881 2187 -847
rect 2393 -881 2409 -847
rect 2629 -881 2645 -847
rect 2851 -881 2867 -847
rect 3087 -881 3103 -847
rect 3309 -881 3325 -847
rect 3545 -881 3561 -847
rect 3767 -881 3783 -847
rect 4003 -881 4019 -847
<< viali >>
rect -3985 847 -3801 881
rect -3527 847 -3343 881
rect -3069 847 -2885 881
rect -2611 847 -2427 881
rect -2153 847 -1969 881
rect -1695 847 -1511 881
rect -1237 847 -1053 881
rect -779 847 -595 881
rect -321 847 -137 881
rect 137 847 321 881
rect 595 847 779 881
rect 1053 847 1237 881
rect 1511 847 1695 881
rect 1969 847 2153 881
rect 2427 847 2611 881
rect 2885 847 3069 881
rect 3343 847 3527 881
rect 3801 847 3985 881
rect -4139 -788 -4105 788
rect -3681 -788 -3647 788
rect -3223 -788 -3189 788
rect -2765 -788 -2731 788
rect -2307 -788 -2273 788
rect -1849 -788 -1815 788
rect -1391 -788 -1357 788
rect -933 -788 -899 788
rect -475 -788 -441 788
rect -17 -788 17 788
rect 441 -788 475 788
rect 899 -788 933 788
rect 1357 -788 1391 788
rect 1815 -788 1849 788
rect 2273 -788 2307 788
rect 2731 -788 2765 788
rect 3189 -788 3223 788
rect 3647 -788 3681 788
rect 4105 -788 4139 788
rect -3985 -881 -3801 -847
rect -3527 -881 -3343 -847
rect -3069 -881 -2885 -847
rect -2611 -881 -2427 -847
rect -2153 -881 -1969 -847
rect -1695 -881 -1511 -847
rect -1237 -881 -1053 -847
rect -779 -881 -595 -847
rect -321 -881 -137 -847
rect 137 -881 321 -847
rect 595 -881 779 -847
rect 1053 -881 1237 -847
rect 1511 -881 1695 -847
rect 1969 -881 2153 -847
rect 2427 -881 2611 -847
rect 2885 -881 3069 -847
rect 3343 -881 3527 -847
rect 3801 -881 3985 -847
<< metal1 >>
rect -3997 881 -3789 887
rect -3997 847 -3985 881
rect -3801 847 -3789 881
rect -3997 841 -3789 847
rect -3539 881 -3331 887
rect -3539 847 -3527 881
rect -3343 847 -3331 881
rect -3539 841 -3331 847
rect -3081 881 -2873 887
rect -3081 847 -3069 881
rect -2885 847 -2873 881
rect -3081 841 -2873 847
rect -2623 881 -2415 887
rect -2623 847 -2611 881
rect -2427 847 -2415 881
rect -2623 841 -2415 847
rect -2165 881 -1957 887
rect -2165 847 -2153 881
rect -1969 847 -1957 881
rect -2165 841 -1957 847
rect -1707 881 -1499 887
rect -1707 847 -1695 881
rect -1511 847 -1499 881
rect -1707 841 -1499 847
rect -1249 881 -1041 887
rect -1249 847 -1237 881
rect -1053 847 -1041 881
rect -1249 841 -1041 847
rect -791 881 -583 887
rect -791 847 -779 881
rect -595 847 -583 881
rect -791 841 -583 847
rect -333 881 -125 887
rect -333 847 -321 881
rect -137 847 -125 881
rect -333 841 -125 847
rect 125 881 333 887
rect 125 847 137 881
rect 321 847 333 881
rect 125 841 333 847
rect 583 881 791 887
rect 583 847 595 881
rect 779 847 791 881
rect 583 841 791 847
rect 1041 881 1249 887
rect 1041 847 1053 881
rect 1237 847 1249 881
rect 1041 841 1249 847
rect 1499 881 1707 887
rect 1499 847 1511 881
rect 1695 847 1707 881
rect 1499 841 1707 847
rect 1957 881 2165 887
rect 1957 847 1969 881
rect 2153 847 2165 881
rect 1957 841 2165 847
rect 2415 881 2623 887
rect 2415 847 2427 881
rect 2611 847 2623 881
rect 2415 841 2623 847
rect 2873 881 3081 887
rect 2873 847 2885 881
rect 3069 847 3081 881
rect 2873 841 3081 847
rect 3331 881 3539 887
rect 3331 847 3343 881
rect 3527 847 3539 881
rect 3331 841 3539 847
rect 3789 881 3997 887
rect 3789 847 3801 881
rect 3985 847 3997 881
rect 3789 841 3997 847
rect -4145 788 -4099 800
rect -4145 -788 -4139 788
rect -4105 -788 -4099 788
rect -4145 -800 -4099 -788
rect -3687 788 -3641 800
rect -3687 -788 -3681 788
rect -3647 -788 -3641 788
rect -3687 -800 -3641 -788
rect -3229 788 -3183 800
rect -3229 -788 -3223 788
rect -3189 -788 -3183 788
rect -3229 -800 -3183 -788
rect -2771 788 -2725 800
rect -2771 -788 -2765 788
rect -2731 -788 -2725 788
rect -2771 -800 -2725 -788
rect -2313 788 -2267 800
rect -2313 -788 -2307 788
rect -2273 -788 -2267 788
rect -2313 -800 -2267 -788
rect -1855 788 -1809 800
rect -1855 -788 -1849 788
rect -1815 -788 -1809 788
rect -1855 -800 -1809 -788
rect -1397 788 -1351 800
rect -1397 -788 -1391 788
rect -1357 -788 -1351 788
rect -1397 -800 -1351 -788
rect -939 788 -893 800
rect -939 -788 -933 788
rect -899 -788 -893 788
rect -939 -800 -893 -788
rect -481 788 -435 800
rect -481 -788 -475 788
rect -441 -788 -435 788
rect -481 -800 -435 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 435 788 481 800
rect 435 -788 441 788
rect 475 -788 481 788
rect 435 -800 481 -788
rect 893 788 939 800
rect 893 -788 899 788
rect 933 -788 939 788
rect 893 -800 939 -788
rect 1351 788 1397 800
rect 1351 -788 1357 788
rect 1391 -788 1397 788
rect 1351 -800 1397 -788
rect 1809 788 1855 800
rect 1809 -788 1815 788
rect 1849 -788 1855 788
rect 1809 -800 1855 -788
rect 2267 788 2313 800
rect 2267 -788 2273 788
rect 2307 -788 2313 788
rect 2267 -800 2313 -788
rect 2725 788 2771 800
rect 2725 -788 2731 788
rect 2765 -788 2771 788
rect 2725 -800 2771 -788
rect 3183 788 3229 800
rect 3183 -788 3189 788
rect 3223 -788 3229 788
rect 3183 -800 3229 -788
rect 3641 788 3687 800
rect 3641 -788 3647 788
rect 3681 -788 3687 788
rect 3641 -800 3687 -788
rect 4099 788 4145 800
rect 4099 -788 4105 788
rect 4139 -788 4145 788
rect 4099 -800 4145 -788
rect -3997 -847 -3789 -841
rect -3997 -881 -3985 -847
rect -3801 -881 -3789 -847
rect -3997 -887 -3789 -881
rect -3539 -847 -3331 -841
rect -3539 -881 -3527 -847
rect -3343 -881 -3331 -847
rect -3539 -887 -3331 -881
rect -3081 -847 -2873 -841
rect -3081 -881 -3069 -847
rect -2885 -881 -2873 -847
rect -3081 -887 -2873 -881
rect -2623 -847 -2415 -841
rect -2623 -881 -2611 -847
rect -2427 -881 -2415 -847
rect -2623 -887 -2415 -881
rect -2165 -847 -1957 -841
rect -2165 -881 -2153 -847
rect -1969 -881 -1957 -847
rect -2165 -887 -1957 -881
rect -1707 -847 -1499 -841
rect -1707 -881 -1695 -847
rect -1511 -881 -1499 -847
rect -1707 -887 -1499 -881
rect -1249 -847 -1041 -841
rect -1249 -881 -1237 -847
rect -1053 -881 -1041 -847
rect -1249 -887 -1041 -881
rect -791 -847 -583 -841
rect -791 -881 -779 -847
rect -595 -881 -583 -847
rect -791 -887 -583 -881
rect -333 -847 -125 -841
rect -333 -881 -321 -847
rect -137 -881 -125 -847
rect -333 -887 -125 -881
rect 125 -847 333 -841
rect 125 -881 137 -847
rect 321 -881 333 -847
rect 125 -887 333 -881
rect 583 -847 791 -841
rect 583 -881 595 -847
rect 779 -881 791 -847
rect 583 -887 791 -881
rect 1041 -847 1249 -841
rect 1041 -881 1053 -847
rect 1237 -881 1249 -847
rect 1041 -887 1249 -881
rect 1499 -847 1707 -841
rect 1499 -881 1511 -847
rect 1695 -881 1707 -847
rect 1499 -887 1707 -881
rect 1957 -847 2165 -841
rect 1957 -881 1969 -847
rect 2153 -881 2165 -847
rect 1957 -887 2165 -881
rect 2415 -847 2623 -841
rect 2415 -881 2427 -847
rect 2611 -881 2623 -847
rect 2415 -887 2623 -881
rect 2873 -847 3081 -841
rect 2873 -881 2885 -847
rect 3069 -881 3081 -847
rect 2873 -887 3081 -881
rect 3331 -847 3539 -841
rect 3331 -881 3343 -847
rect 3527 -881 3539 -847
rect 3331 -887 3539 -881
rect 3789 -847 3997 -841
rect 3789 -881 3801 -847
rect 3985 -881 3997 -847
rect 3789 -887 3997 -881
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_hvt
string parameters w 8 l 2 m 1 nf 18 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
