magic
tech sky130A
timestamp 1626486988
<< checkpaint >>
rect -885 -720 885 720
<< metal4 >>
rect -255 59 255 90
rect -255 -59 -219 59
rect -101 -59 -59 59
rect 59 -59 101 59
rect 219 -59 255 59
rect -255 -90 255 -59
<< via4 >>
rect -219 -59 -101 59
rect -59 -59 59 59
rect 101 -59 219 59
<< metal5 >>
rect -255 59 255 90
rect -255 -59 -219 59
rect -101 -59 -59 59
rect 59 -59 101 59
rect 219 -59 255 59
rect -255 -90 255 -59
<< end >>
