magic
tech sky130A
timestamp 1626486988
<< checkpaint >>
rect -720 -817 720 817
<< metal4 >>
rect -90 139 90 187
rect -90 21 -59 139
rect 59 21 90 139
rect -90 -21 90 21
rect -90 -139 -59 -21
rect 59 -139 90 -21
rect -90 -187 90 -139
<< via4 >>
rect -59 21 59 139
rect -59 -139 59 -21
<< metal5 >>
rect -90 139 90 187
rect -90 21 -59 139
rect 59 21 90 139
rect -90 -21 90 21
rect -90 -139 -59 -21
rect 59 -139 90 -21
rect -90 -187 90 -139
<< end >>
