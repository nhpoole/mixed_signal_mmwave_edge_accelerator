magic
tech sky130A
magscale 1 2
timestamp 1622079483
<< nwell >>
rect 10 157 1834 478
<< pwell >>
rect 752 53 934 97
rect 1242 53 1795 99
rect 49 -83 1795 53
rect 77 -121 111 -83
<< scnmos >>
rect 127 -57 157 27
rect 211 -57 241 27
rect 399 -57 429 27
rect 511 -57 541 15
rect 610 -57 640 15
rect 709 -57 739 27
rect 828 -57 858 71
rect 929 -57 959 15
rect 1035 -57 1065 15
rect 1130 -57 1160 27
rect 1320 -57 1350 73
rect 1404 -57 1434 73
rect 1592 -57 1622 27
rect 1687 -57 1717 73
<< scpmoshvt >>
rect 127 259 157 387
rect 211 259 241 387
rect 399 309 429 393
rect 484 309 514 393
rect 579 309 609 393
rect 682 309 712 393
rect 814 243 844 393
rect 909 309 939 393
rect 993 309 1023 393
rect 1107 309 1137 393
rect 1318 193 1348 393
rect 1402 193 1432 393
rect 1590 265 1620 393
rect 1687 193 1717 393
<< ndiff >>
rect 75 15 127 27
rect 75 -19 83 15
rect 117 -19 127 15
rect 75 -57 127 -19
rect 157 -11 211 27
rect 157 -45 167 -11
rect 201 -45 211 -11
rect 157 -57 211 -45
rect 241 15 293 27
rect 241 -19 251 15
rect 285 -19 293 15
rect 241 -57 293 -19
rect 347 -11 399 27
rect 347 -45 355 -11
rect 389 -45 399 -11
rect 347 -57 399 -45
rect 429 15 479 27
rect 778 27 828 71
rect 659 15 709 27
rect 429 3 511 15
rect 429 -31 440 3
rect 474 -31 511 3
rect 429 -57 511 -31
rect 541 3 610 15
rect 541 -31 551 3
rect 585 -31 610 3
rect 541 -57 610 -31
rect 640 -57 709 15
rect 739 -3 828 27
rect 739 -37 750 -3
rect 784 -37 828 -3
rect 739 -57 828 -37
rect 858 15 908 71
rect 1268 58 1320 73
rect 1080 15 1130 27
rect 858 3 929 15
rect 858 -31 869 3
rect 903 -31 929 3
rect 858 -57 929 -31
rect 959 3 1035 15
rect 959 -31 972 3
rect 1006 -31 1035 3
rect 959 -57 1035 -31
rect 1065 -57 1130 15
rect 1160 3 1212 27
rect 1160 -31 1170 3
rect 1204 -31 1212 3
rect 1160 -57 1212 -31
rect 1268 24 1276 58
rect 1310 24 1320 58
rect 1268 -10 1320 24
rect 1268 -44 1276 -10
rect 1310 -44 1320 -10
rect 1268 -57 1320 -44
rect 1350 19 1404 73
rect 1350 -15 1360 19
rect 1394 -15 1404 19
rect 1350 -57 1404 -15
rect 1434 60 1486 73
rect 1434 26 1444 60
rect 1478 26 1486 60
rect 1637 27 1687 73
rect 1434 -8 1486 26
rect 1434 -42 1444 -8
rect 1478 -42 1486 -8
rect 1434 -57 1486 -42
rect 1540 15 1592 27
rect 1540 -19 1548 15
rect 1582 -19 1592 15
rect 1540 -57 1592 -19
rect 1622 -11 1687 27
rect 1622 -45 1643 -11
rect 1677 -45 1687 -11
rect 1622 -57 1687 -45
rect 1717 27 1769 73
rect 1717 -7 1727 27
rect 1761 -7 1769 27
rect 1717 -57 1769 -7
<< pdiff >>
rect 75 373 127 387
rect 75 339 83 373
rect 117 339 127 373
rect 75 305 127 339
rect 75 271 83 305
rect 117 271 127 305
rect 75 259 127 271
rect 157 357 211 387
rect 157 323 167 357
rect 201 323 211 357
rect 157 259 211 323
rect 241 373 293 387
rect 241 339 251 373
rect 285 339 293 373
rect 241 305 293 339
rect 347 381 399 393
rect 347 347 355 381
rect 389 347 399 381
rect 347 309 399 347
rect 429 373 484 393
rect 429 339 439 373
rect 473 339 484 373
rect 429 309 484 339
rect 514 368 579 393
rect 514 334 531 368
rect 565 334 579 368
rect 514 309 579 334
rect 609 309 682 393
rect 712 381 814 393
rect 712 347 770 381
rect 804 347 814 381
rect 712 313 814 347
rect 712 309 770 313
rect 241 271 251 305
rect 285 271 293 305
rect 241 259 293 271
rect 727 279 770 309
rect 804 279 814 313
rect 727 243 814 279
rect 844 373 909 393
rect 844 339 854 373
rect 888 339 909 373
rect 844 309 909 339
rect 939 363 993 393
rect 939 329 949 363
rect 983 329 993 363
rect 939 309 993 329
rect 1023 309 1107 393
rect 1137 373 1190 393
rect 1137 339 1148 373
rect 1182 339 1190 373
rect 1137 309 1190 339
rect 1264 381 1318 393
rect 1264 347 1272 381
rect 1306 347 1318 381
rect 1264 310 1318 347
rect 844 243 894 309
rect 1264 276 1272 310
rect 1306 276 1318 310
rect 1264 239 1318 276
rect 1264 205 1272 239
rect 1306 205 1318 239
rect 1264 193 1318 205
rect 1348 351 1402 393
rect 1348 317 1358 351
rect 1392 317 1402 351
rect 1348 271 1402 317
rect 1348 237 1358 271
rect 1392 237 1402 271
rect 1348 193 1402 237
rect 1432 375 1484 393
rect 1432 341 1442 375
rect 1476 341 1484 375
rect 1432 307 1484 341
rect 1432 273 1442 307
rect 1476 273 1484 307
rect 1432 239 1484 273
rect 1538 381 1590 393
rect 1538 347 1546 381
rect 1580 347 1590 381
rect 1538 313 1590 347
rect 1538 279 1546 313
rect 1580 279 1590 313
rect 1538 265 1590 279
rect 1620 381 1687 393
rect 1620 347 1643 381
rect 1677 347 1687 381
rect 1620 313 1687 347
rect 1620 279 1643 313
rect 1677 279 1687 313
rect 1620 265 1687 279
rect 1432 205 1442 239
rect 1476 205 1484 239
rect 1432 193 1484 205
rect 1635 245 1687 265
rect 1635 211 1643 245
rect 1677 211 1687 245
rect 1635 193 1687 211
rect 1717 381 1769 393
rect 1717 347 1727 381
rect 1761 347 1769 381
rect 1717 310 1769 347
rect 1717 276 1727 310
rect 1761 276 1769 310
rect 1717 239 1769 276
rect 1717 205 1727 239
rect 1761 205 1769 239
rect 1717 193 1769 205
<< ndiffc >>
rect 83 -19 117 15
rect 167 -45 201 -11
rect 251 -19 285 15
rect 355 -45 389 -11
rect 440 -31 474 3
rect 551 -31 585 3
rect 750 -37 784 -3
rect 869 -31 903 3
rect 972 -31 1006 3
rect 1170 -31 1204 3
rect 1276 24 1310 58
rect 1276 -44 1310 -10
rect 1360 -15 1394 19
rect 1444 26 1478 60
rect 1444 -42 1478 -8
rect 1548 -19 1582 15
rect 1643 -45 1677 -11
rect 1727 -7 1761 27
<< pdiffc >>
rect 83 339 117 373
rect 83 271 117 305
rect 167 323 201 357
rect 251 339 285 373
rect 355 347 389 381
rect 439 339 473 373
rect 531 334 565 368
rect 770 347 804 381
rect 251 271 285 305
rect 770 279 804 313
rect 854 339 888 373
rect 949 329 983 363
rect 1148 339 1182 373
rect 1272 347 1306 381
rect 1272 276 1306 310
rect 1272 205 1306 239
rect 1358 317 1392 351
rect 1358 237 1392 271
rect 1442 341 1476 375
rect 1442 273 1476 307
rect 1546 347 1580 381
rect 1546 279 1580 313
rect 1643 347 1677 381
rect 1643 279 1677 313
rect 1442 205 1476 239
rect 1643 211 1677 245
rect 1727 347 1761 381
rect 1727 276 1761 310
rect 1727 205 1761 239
<< poly >>
rect 127 387 157 413
rect 211 387 241 413
rect 399 393 429 419
rect 484 393 514 419
rect 579 393 609 419
rect 682 393 712 419
rect 814 393 844 419
rect 909 393 939 419
rect 993 393 1023 419
rect 1107 393 1137 419
rect 1318 393 1348 419
rect 1402 393 1432 419
rect 1590 393 1620 419
rect 1687 393 1717 419
rect 127 244 157 259
rect 94 214 157 244
rect 94 161 124 214
rect 211 170 241 259
rect 399 229 429 309
rect 70 145 124 161
rect 70 111 80 145
rect 114 111 124 145
rect 166 160 241 170
rect 334 213 429 229
rect 334 179 344 213
rect 378 179 429 213
rect 484 193 514 309
rect 579 277 609 309
rect 579 261 640 277
rect 579 227 596 261
rect 630 227 640 261
rect 579 211 640 227
rect 334 163 429 179
rect 166 126 182 160
rect 216 126 241 160
rect 166 116 241 126
rect 70 95 124 111
rect 94 72 124 95
rect 94 42 157 72
rect 127 27 157 42
rect 211 27 241 116
rect 399 27 429 163
rect 471 183 537 193
rect 471 149 487 183
rect 521 169 537 183
rect 521 149 640 169
rect 471 139 640 149
rect 491 87 557 97
rect 491 53 507 87
rect 541 53 557 87
rect 491 43 557 53
rect 511 15 541 43
rect 610 15 640 139
rect 682 109 712 309
rect 814 205 844 243
rect 909 211 939 309
rect 993 271 1023 309
rect 1107 277 1137 309
rect 992 261 1058 271
rect 992 227 1008 261
rect 1042 227 1058 261
rect 992 217 1058 227
rect 1107 261 1188 277
rect 1107 227 1144 261
rect 1178 227 1188 261
rect 1107 211 1188 227
rect 754 195 844 205
rect 754 161 770 195
rect 804 161 844 195
rect 754 151 844 161
rect 814 116 844 151
rect 896 195 950 211
rect 896 161 906 195
rect 940 175 950 195
rect 940 161 1065 175
rect 896 145 1065 161
rect 682 99 756 109
rect 682 65 706 99
rect 740 65 756 99
rect 814 86 858 116
rect 828 71 858 86
rect 929 87 993 103
rect 682 55 756 65
rect 709 27 739 55
rect 929 53 949 87
rect 983 53 993 87
rect 929 37 993 53
rect 929 15 959 37
rect 1035 15 1065 145
rect 1130 27 1160 211
rect 1590 229 1620 265
rect 1581 199 1620 229
rect 1318 161 1348 193
rect 1402 161 1432 193
rect 1581 161 1611 199
rect 1687 161 1717 193
rect 1208 145 1350 161
rect 1208 111 1218 145
rect 1252 111 1350 145
rect 1208 95 1350 111
rect 1392 145 1611 161
rect 1392 111 1402 145
rect 1436 111 1611 145
rect 1392 95 1611 111
rect 1653 145 1717 161
rect 1653 111 1663 145
rect 1697 111 1717 145
rect 1653 95 1717 111
rect 1320 73 1350 95
rect 1404 73 1434 95
rect 1581 66 1611 95
rect 1687 73 1717 95
rect 1581 42 1622 66
rect 1592 27 1622 42
rect 127 -83 157 -57
rect 211 -83 241 -57
rect 399 -83 429 -57
rect 511 -83 541 -57
rect 610 -83 640 -57
rect 709 -83 739 -57
rect 828 -83 858 -57
rect 929 -83 959 -57
rect 1035 -83 1065 -57
rect 1130 -83 1160 -57
rect 1320 -83 1350 -57
rect 1404 -83 1434 -57
rect 1592 -83 1622 -57
rect 1687 -83 1717 -57
<< polycont >>
rect 80 111 114 145
rect 344 179 378 213
rect 596 227 630 261
rect 182 126 216 160
rect 487 149 521 183
rect 507 53 541 87
rect 1008 227 1042 261
rect 1144 227 1178 261
rect 770 161 804 195
rect 906 161 940 195
rect 706 65 740 99
rect 949 53 983 87
rect 1218 111 1252 145
rect 1402 111 1436 145
rect 1663 111 1697 145
<< locali >>
rect 48 423 77 457
rect 111 423 169 457
rect 203 423 261 457
rect 295 423 353 457
rect 387 423 445 457
rect 479 423 537 457
rect 571 423 629 457
rect 663 423 721 457
rect 755 423 813 457
rect 847 423 905 457
rect 939 423 997 457
rect 1031 423 1089 457
rect 1123 423 1181 457
rect 1215 423 1273 457
rect 1307 423 1365 457
rect 1399 423 1457 457
rect 1491 423 1549 457
rect 1583 423 1641 457
rect 1675 423 1733 457
rect 1767 423 1796 457
rect 83 373 117 389
rect 83 305 117 339
rect 151 357 217 423
rect 151 323 167 357
rect 201 323 217 357
rect 251 373 288 389
rect 285 339 288 373
rect 251 305 288 339
rect 336 381 389 423
rect 336 347 355 381
rect 336 331 389 347
rect 423 373 473 389
rect 423 339 439 373
rect 770 381 804 423
rect 117 287 216 289
rect 117 271 174 287
rect 83 255 174 271
rect 170 253 174 255
rect 208 253 216 287
rect 66 164 136 221
rect 66 111 80 164
rect 128 116 136 164
rect 114 111 136 116
rect 66 91 136 111
rect 170 160 216 253
rect 170 126 182 160
rect 170 57 216 126
rect 83 23 216 57
rect 285 271 288 305
rect 423 304 473 339
rect 515 334 531 368
rect 565 334 736 368
rect 251 219 288 271
rect 412 278 473 304
rect 562 287 668 300
rect 251 185 253 219
rect 287 185 288 219
rect 83 15 117 23
rect 251 15 288 185
rect 322 213 378 229
rect 322 179 344 213
rect 322 134 378 179
rect 322 86 326 134
rect 374 86 378 134
rect 322 39 378 86
rect 412 57 446 278
rect 562 253 594 287
rect 628 261 668 287
rect 480 219 528 240
rect 480 185 491 219
rect 525 185 528 219
rect 480 183 528 185
rect 480 149 487 183
rect 521 149 528 183
rect 480 121 528 149
rect 562 87 596 253
rect 630 227 668 261
rect 702 211 736 334
rect 770 313 804 347
rect 770 263 804 279
rect 838 373 888 389
rect 838 339 854 373
rect 1146 373 1209 423
rect 838 323 888 339
rect 933 329 949 363
rect 983 329 1110 363
rect 702 195 804 211
rect 702 193 770 195
rect 412 31 457 57
rect 491 53 507 87
rect 541 53 596 87
rect 491 43 596 53
rect 630 161 770 193
rect 630 159 804 161
rect 83 -35 117 -19
rect 151 -45 167 -11
rect 201 -45 217 -11
rect 285 -19 288 15
rect 251 -35 288 -19
rect 339 -11 389 5
rect 151 -87 217 -45
rect 339 -45 355 -11
rect 423 3 457 31
rect 630 3 664 159
rect 770 145 804 159
rect 706 109 746 115
rect 838 109 872 323
rect 906 287 944 289
rect 906 253 908 287
rect 942 253 944 287
rect 906 195 944 253
rect 940 161 944 195
rect 906 145 944 161
rect 978 261 1042 295
rect 978 227 1008 261
rect 978 219 1042 227
rect 978 185 995 219
rect 1029 185 1042 219
rect 706 99 872 109
rect 978 103 1042 185
rect 740 65 872 99
rect 706 49 872 65
rect 423 -31 440 3
rect 474 -31 490 3
rect 529 -31 551 3
rect 585 -31 664 3
rect 728 -3 802 13
rect 339 -87 389 -45
rect 728 -37 750 -3
rect 784 -37 802 -3
rect 838 3 872 49
rect 949 87 1042 103
rect 983 53 1042 87
rect 949 37 1042 53
rect 1076 161 1110 329
rect 1146 339 1148 373
rect 1182 339 1209 373
rect 1146 323 1209 339
rect 1256 381 1324 389
rect 1256 347 1272 381
rect 1306 347 1324 381
rect 1256 310 1324 347
rect 1256 277 1272 310
rect 1144 276 1272 277
rect 1306 276 1324 310
rect 1144 261 1324 276
rect 1178 239 1324 261
rect 1178 227 1272 239
rect 1144 205 1272 227
rect 1306 205 1324 239
rect 1358 351 1392 423
rect 1530 381 1596 385
rect 1358 271 1392 317
rect 1358 221 1392 237
rect 1426 375 1492 380
rect 1426 341 1442 375
rect 1476 341 1492 375
rect 1426 307 1492 341
rect 1426 273 1442 307
rect 1476 273 1492 307
rect 1426 239 1492 273
rect 1530 347 1546 381
rect 1580 347 1596 381
rect 1530 313 1596 347
rect 1530 279 1546 313
rect 1580 279 1596 313
rect 1530 239 1596 279
rect 1144 202 1324 205
rect 1286 161 1324 202
rect 1426 205 1442 239
rect 1476 211 1492 239
rect 1476 205 1508 211
rect 1426 195 1508 205
rect 1461 185 1508 195
rect 1076 145 1252 161
rect 1076 111 1218 145
rect 1076 95 1252 111
rect 1286 145 1436 161
rect 1286 111 1402 145
rect 1286 95 1436 111
rect 1076 3 1110 95
rect 1286 61 1326 95
rect 1470 69 1508 185
rect 1459 61 1508 69
rect 1260 58 1326 61
rect 1260 24 1276 58
rect 1310 24 1326 58
rect 1428 60 1508 61
rect 1428 44 1444 60
rect 1478 44 1508 60
rect 1542 161 1596 239
rect 1634 381 1677 423
rect 1634 347 1643 381
rect 1634 313 1677 347
rect 1634 279 1643 313
rect 1634 245 1677 279
rect 1634 211 1643 245
rect 1634 195 1677 211
rect 1711 381 1778 389
rect 1711 347 1727 381
rect 1761 347 1778 381
rect 1711 310 1778 347
rect 1711 276 1727 310
rect 1761 276 1778 310
rect 1711 256 1778 276
rect 1711 208 1718 256
rect 1766 208 1778 256
rect 1711 205 1727 208
rect 1761 205 1778 208
rect 1711 192 1778 205
rect 1542 145 1697 161
rect 1542 111 1663 145
rect 1542 95 1697 111
rect 838 -31 869 3
rect 903 -31 919 3
rect 953 -31 972 3
rect 1006 -31 1110 3
rect 1165 3 1207 19
rect 1165 -31 1170 3
rect 1204 -31 1207 3
rect 728 -87 802 -37
rect 1165 -87 1207 -31
rect 1260 -10 1326 24
rect 1260 -44 1276 -10
rect 1310 -44 1326 -10
rect 1360 19 1394 35
rect 1360 -87 1394 -15
rect 1428 -4 1434 44
rect 1482 -4 1494 44
rect 1542 19 1582 95
rect 1731 78 1778 192
rect 1428 -8 1494 -4
rect 1428 -42 1444 -8
rect 1478 -42 1494 -8
rect 1532 15 1582 19
rect 1532 -19 1548 15
rect 1727 27 1778 78
rect 1532 -35 1582 -19
rect 1629 -11 1693 5
rect 1428 -43 1494 -42
rect 1629 -45 1643 -11
rect 1677 -45 1693 -11
rect 1629 -87 1693 -45
rect 1761 -7 1778 27
rect 1727 -53 1778 -7
rect 48 -121 77 -87
rect 111 -121 169 -87
rect 203 -121 261 -87
rect 295 -121 353 -87
rect 387 -121 445 -87
rect 479 -121 537 -87
rect 571 -121 629 -87
rect 663 -121 721 -87
rect 755 -121 813 -87
rect 847 -121 905 -87
rect 939 -121 997 -87
rect 1031 -121 1089 -87
rect 1123 -121 1181 -87
rect 1215 -121 1273 -87
rect 1307 -121 1365 -87
rect 1399 -121 1457 -87
rect 1491 -121 1549 -87
rect 1583 -121 1641 -87
rect 1675 -121 1733 -87
rect 1767 -121 1796 -87
<< viali >>
rect 77 423 111 457
rect 169 423 203 457
rect 261 423 295 457
rect 353 423 387 457
rect 445 423 479 457
rect 537 423 571 457
rect 629 423 663 457
rect 721 423 755 457
rect 813 423 847 457
rect 905 423 939 457
rect 997 423 1031 457
rect 1089 423 1123 457
rect 1181 423 1215 457
rect 1273 423 1307 457
rect 1365 423 1399 457
rect 1457 423 1491 457
rect 1549 423 1583 457
rect 1641 423 1675 457
rect 1733 423 1767 457
rect 174 253 208 287
rect 80 145 128 164
rect 80 116 114 145
rect 114 116 128 145
rect 253 185 287 219
rect 326 86 374 134
rect 594 261 628 287
rect 594 253 596 261
rect 596 253 628 261
rect 491 185 525 219
rect 908 253 942 287
rect 995 185 1029 219
rect 1718 239 1766 256
rect 1718 208 1727 239
rect 1727 208 1761 239
rect 1761 208 1766 239
rect 1434 26 1444 44
rect 1444 26 1478 44
rect 1478 26 1482 44
rect 1434 -4 1482 26
rect 77 -121 111 -87
rect 169 -121 203 -87
rect 261 -121 295 -87
rect 353 -121 387 -87
rect 445 -121 479 -87
rect 537 -121 571 -87
rect 629 -121 663 -87
rect 721 -121 755 -87
rect 813 -121 847 -87
rect 905 -121 939 -87
rect 997 -121 1031 -87
rect 1089 -121 1123 -87
rect 1181 -121 1215 -87
rect 1273 -121 1307 -87
rect 1365 -121 1399 -87
rect 1457 -121 1491 -87
rect 1549 -121 1583 -87
rect 1641 -121 1675 -87
rect 1733 -121 1767 -87
<< metal1 >>
rect -154 457 1796 488
rect -154 423 77 457
rect 111 423 169 457
rect 203 423 261 457
rect 295 423 353 457
rect 387 423 445 457
rect 479 423 537 457
rect 571 423 629 457
rect 663 423 721 457
rect 755 423 813 457
rect 847 423 905 457
rect 939 423 997 457
rect 1031 423 1089 457
rect 1123 423 1181 457
rect 1215 423 1273 457
rect 1307 423 1365 457
rect 1399 423 1457 457
rect 1491 423 1549 457
rect 1583 423 1641 457
rect 1675 423 1733 457
rect 1767 423 1796 457
rect -154 392 1796 423
rect 162 287 220 293
rect 162 253 174 287
rect 208 284 220 287
rect 582 287 640 293
rect 582 284 594 287
rect 208 256 594 284
rect 208 253 220 256
rect 162 247 220 253
rect 582 253 594 256
rect 628 284 640 287
rect 896 287 954 293
rect 896 284 908 287
rect 628 256 908 284
rect 628 253 640 256
rect 582 247 640 253
rect 896 253 908 256
rect 942 253 954 287
rect 896 247 954 253
rect 1706 256 1992 262
rect 241 219 299 225
rect 241 185 253 219
rect 287 216 299 219
rect 479 219 537 225
rect 479 216 491 219
rect 287 188 491 216
rect 287 185 299 188
rect 241 179 299 185
rect 479 185 491 188
rect 525 216 537 219
rect 983 219 1041 225
rect 983 216 995 219
rect 525 188 995 216
rect 525 185 537 188
rect 479 179 537 185
rect 983 185 995 188
rect 1029 185 1041 219
rect 1706 208 1718 256
rect 1766 208 1992 256
rect 1706 202 1992 208
rect 983 179 1041 185
rect -66 164 140 170
rect -66 116 80 164
rect 128 116 140 164
rect -66 110 140 116
rect 314 134 386 140
rect 314 86 326 134
rect 374 86 386 134
rect 314 80 386 86
rect 314 60 380 80
rect -164 0 380 60
rect 1422 44 1878 50
rect 1422 -4 1434 44
rect 1482 -4 1878 44
rect 1422 -10 1878 -4
rect -134 -87 1796 -56
rect -134 -121 77 -87
rect 111 -121 169 -87
rect 203 -121 261 -87
rect 295 -121 353 -87
rect 387 -121 445 -87
rect 479 -121 537 -87
rect 571 -121 629 -87
rect 663 -121 721 -87
rect 755 -121 813 -87
rect 847 -121 905 -87
rect 939 -121 997 -87
rect 1031 -121 1089 -87
rect 1123 -121 1181 -87
rect 1215 -121 1273 -87
rect 1307 -121 1365 -87
rect 1399 -121 1457 -87
rect 1491 -121 1549 -87
rect 1583 -121 1641 -87
rect 1675 -121 1733 -87
rect 1767 -121 1796 -87
rect -134 -152 1796 -121
<< labels >>
flabel metal1 -26 128 -20 136 1 FreeSans 480 0 0 0 CLK
port 2 n
flabel metal1 -126 20 -120 28 1 FreeSans 480 0 0 0 D
port 1 n
flabel metal1 -60 -106 -56 -100 1 FreeSans 480 0 0 0 VSS
port 6 n ground bidirectional
flabel metal1 -90 436 -88 440 1 FreeSans 480 0 0 0 VDD
port 5 n power bidirectional
flabel metal1 1932 226 1936 230 1 FreeSans 480 0 0 0 QB
port 4 n
flabel metal1 1840 22 1842 24 1 FreeSans 480 0 0 0 Q
port 3 n
flabel metal1 77 -121 111 -87 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VGND
flabel metal1 77 423 111 457 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VPWR
flabel locali 1733 200 1767 234 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/Q_N
flabel locali 337 117 371 151 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/D
flabel locali 77 117 111 151 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/CLK
flabel locali 1438 -19 1472 15 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/Q
flabel pwell 77 -121 111 -87 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VNB
flabel pwell 94 -104 94 -104 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VNB
flabel nwell 77 423 111 457 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VPB
flabel nwell 94 440 94 440 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VPB
rlabel comment 48 -104 48 -104 4 sky130_fd_sc_hd__dfxbp_1_0/dfxbp_1
<< end >>
