magic
tech sky130A
timestamp 1626486988
<< checkpaint >>
rect -1038 -798 1038 798
<< metal4 >>
rect -408 139 408 168
rect -408 -139 -379 139
rect 379 -139 408 139
rect -408 -168 408 -139
<< via4 >>
rect -379 -139 379 139
<< metal5 >>
rect -408 139 408 168
rect -408 -139 -379 139
rect 379 -139 408 139
rect -408 -168 408 -139
<< end >>
