magic
tech sky130A
magscale 1 2
timestamp 1623920776
<< metal1 >>
rect -30 100 30 157
rect -30 -157 30 -100
<< rmetal1 >>
rect -30 -100 30 100
<< properties >>
string gencell sky130_fd_pr__res_generic_m1
string parameters w 0.30 l 1 m 1 nx 1 wmin 0.14 lmin 0.14 rho 0.125 val 416.666m dummy 0 dw 0.0 term 0.0 roverlap 0
string library sky130
<< end >>
