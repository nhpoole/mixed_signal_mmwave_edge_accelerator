magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -2099 -1560 2099 1560
<< nwell >>
rect -839 -300 839 300
<< pmoshvt >>
rect -745 -200 -545 200
rect -487 -200 -287 200
rect -229 -200 -29 200
rect 29 -200 229 200
rect 287 -200 487 200
rect 545 -200 745 200
<< pdiff >>
rect -803 187 -745 200
rect -803 153 -791 187
rect -757 153 -745 187
rect -803 119 -745 153
rect -803 85 -791 119
rect -757 85 -745 119
rect -803 51 -745 85
rect -803 17 -791 51
rect -757 17 -745 51
rect -803 -17 -745 17
rect -803 -51 -791 -17
rect -757 -51 -745 -17
rect -803 -85 -745 -51
rect -803 -119 -791 -85
rect -757 -119 -745 -85
rect -803 -153 -745 -119
rect -803 -187 -791 -153
rect -757 -187 -745 -153
rect -803 -200 -745 -187
rect -545 187 -487 200
rect -545 153 -533 187
rect -499 153 -487 187
rect -545 119 -487 153
rect -545 85 -533 119
rect -499 85 -487 119
rect -545 51 -487 85
rect -545 17 -533 51
rect -499 17 -487 51
rect -545 -17 -487 17
rect -545 -51 -533 -17
rect -499 -51 -487 -17
rect -545 -85 -487 -51
rect -545 -119 -533 -85
rect -499 -119 -487 -85
rect -545 -153 -487 -119
rect -545 -187 -533 -153
rect -499 -187 -487 -153
rect -545 -200 -487 -187
rect -287 187 -229 200
rect -287 153 -275 187
rect -241 153 -229 187
rect -287 119 -229 153
rect -287 85 -275 119
rect -241 85 -229 119
rect -287 51 -229 85
rect -287 17 -275 51
rect -241 17 -229 51
rect -287 -17 -229 17
rect -287 -51 -275 -17
rect -241 -51 -229 -17
rect -287 -85 -229 -51
rect -287 -119 -275 -85
rect -241 -119 -229 -85
rect -287 -153 -229 -119
rect -287 -187 -275 -153
rect -241 -187 -229 -153
rect -287 -200 -229 -187
rect -29 187 29 200
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -200 29 -187
rect 229 187 287 200
rect 229 153 241 187
rect 275 153 287 187
rect 229 119 287 153
rect 229 85 241 119
rect 275 85 287 119
rect 229 51 287 85
rect 229 17 241 51
rect 275 17 287 51
rect 229 -17 287 17
rect 229 -51 241 -17
rect 275 -51 287 -17
rect 229 -85 287 -51
rect 229 -119 241 -85
rect 275 -119 287 -85
rect 229 -153 287 -119
rect 229 -187 241 -153
rect 275 -187 287 -153
rect 229 -200 287 -187
rect 487 187 545 200
rect 487 153 499 187
rect 533 153 545 187
rect 487 119 545 153
rect 487 85 499 119
rect 533 85 545 119
rect 487 51 545 85
rect 487 17 499 51
rect 533 17 545 51
rect 487 -17 545 17
rect 487 -51 499 -17
rect 533 -51 545 -17
rect 487 -85 545 -51
rect 487 -119 499 -85
rect 533 -119 545 -85
rect 487 -153 545 -119
rect 487 -187 499 -153
rect 533 -187 545 -153
rect 487 -200 545 -187
rect 745 187 803 200
rect 745 153 757 187
rect 791 153 803 187
rect 745 119 803 153
rect 745 85 757 119
rect 791 85 803 119
rect 745 51 803 85
rect 745 17 757 51
rect 791 17 803 51
rect 745 -17 803 17
rect 745 -51 757 -17
rect 791 -51 803 -17
rect 745 -85 803 -51
rect 745 -119 757 -85
rect 791 -119 803 -85
rect 745 -153 803 -119
rect 745 -187 757 -153
rect 791 -187 803 -153
rect 745 -200 803 -187
<< pdiffc >>
rect -791 153 -757 187
rect -791 85 -757 119
rect -791 17 -757 51
rect -791 -51 -757 -17
rect -791 -119 -757 -85
rect -791 -187 -757 -153
rect -533 153 -499 187
rect -533 85 -499 119
rect -533 17 -499 51
rect -533 -51 -499 -17
rect -533 -119 -499 -85
rect -533 -187 -499 -153
rect -275 153 -241 187
rect -275 85 -241 119
rect -275 17 -241 51
rect -275 -51 -241 -17
rect -275 -119 -241 -85
rect -275 -187 -241 -153
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect 241 153 275 187
rect 241 85 275 119
rect 241 17 275 51
rect 241 -51 275 -17
rect 241 -119 275 -85
rect 241 -187 275 -153
rect 499 153 533 187
rect 499 85 533 119
rect 499 17 533 51
rect 499 -51 533 -17
rect 499 -119 533 -85
rect 499 -187 533 -153
rect 757 153 791 187
rect 757 85 791 119
rect 757 17 791 51
rect 757 -51 791 -17
rect 757 -119 791 -85
rect 757 -187 791 -153
<< poly >>
rect -711 281 -579 297
rect -711 264 -662 281
rect -745 247 -662 264
rect -628 264 -579 281
rect -453 281 -321 297
rect -453 264 -404 281
rect -628 247 -545 264
rect -745 200 -545 247
rect -487 247 -404 264
rect -370 264 -321 281
rect -195 281 -63 297
rect -195 264 -146 281
rect -370 247 -287 264
rect -487 200 -287 247
rect -229 247 -146 264
rect -112 264 -63 281
rect 63 281 195 297
rect 63 264 112 281
rect -112 247 -29 264
rect -229 200 -29 247
rect 29 247 112 264
rect 146 264 195 281
rect 321 281 453 297
rect 321 264 370 281
rect 146 247 229 264
rect 29 200 229 247
rect 287 247 370 264
rect 404 264 453 281
rect 579 281 711 297
rect 579 264 628 281
rect 404 247 487 264
rect 287 200 487 247
rect 545 247 628 264
rect 662 264 711 281
rect 662 247 745 264
rect 545 200 745 247
rect -745 -247 -545 -200
rect -745 -264 -662 -247
rect -711 -281 -662 -264
rect -628 -264 -545 -247
rect -487 -247 -287 -200
rect -487 -264 -404 -247
rect -628 -281 -579 -264
rect -711 -297 -579 -281
rect -453 -281 -404 -264
rect -370 -264 -287 -247
rect -229 -247 -29 -200
rect -229 -264 -146 -247
rect -370 -281 -321 -264
rect -453 -297 -321 -281
rect -195 -281 -146 -264
rect -112 -264 -29 -247
rect 29 -247 229 -200
rect 29 -264 112 -247
rect -112 -281 -63 -264
rect -195 -297 -63 -281
rect 63 -281 112 -264
rect 146 -264 229 -247
rect 287 -247 487 -200
rect 287 -264 370 -247
rect 146 -281 195 -264
rect 63 -297 195 -281
rect 321 -281 370 -264
rect 404 -264 487 -247
rect 545 -247 745 -200
rect 545 -264 628 -247
rect 404 -281 453 -264
rect 321 -297 453 -281
rect 579 -281 628 -264
rect 662 -264 745 -247
rect 662 -281 711 -264
rect 579 -297 711 -281
<< polycont >>
rect -662 247 -628 281
rect -404 247 -370 281
rect -146 247 -112 281
rect 112 247 146 281
rect 370 247 404 281
rect 628 247 662 281
rect -662 -281 -628 -247
rect -404 -281 -370 -247
rect -146 -281 -112 -247
rect 112 -281 146 -247
rect 370 -281 404 -247
rect 628 -281 662 -247
<< locali >>
rect -711 247 -662 281
rect -628 247 -579 281
rect -453 247 -404 281
rect -370 247 -321 281
rect -195 247 -146 281
rect -112 247 -63 281
rect 63 247 112 281
rect 146 247 195 281
rect 321 247 370 281
rect 404 247 453 281
rect 579 247 628 281
rect 662 247 711 281
rect -791 187 -757 204
rect -791 119 -757 127
rect -791 51 -757 55
rect -791 -55 -757 -51
rect -791 -127 -757 -119
rect -791 -204 -757 -187
rect -533 187 -499 204
rect -533 119 -499 127
rect -533 51 -499 55
rect -533 -55 -499 -51
rect -533 -127 -499 -119
rect -533 -204 -499 -187
rect -275 187 -241 204
rect -275 119 -241 127
rect -275 51 -241 55
rect -275 -55 -241 -51
rect -275 -127 -241 -119
rect -275 -204 -241 -187
rect -17 187 17 204
rect -17 119 17 127
rect -17 51 17 55
rect -17 -55 17 -51
rect -17 -127 17 -119
rect -17 -204 17 -187
rect 241 187 275 204
rect 241 119 275 127
rect 241 51 275 55
rect 241 -55 275 -51
rect 241 -127 275 -119
rect 241 -204 275 -187
rect 499 187 533 204
rect 499 119 533 127
rect 499 51 533 55
rect 499 -55 533 -51
rect 499 -127 533 -119
rect 499 -204 533 -187
rect 757 187 791 204
rect 757 119 791 127
rect 757 51 791 55
rect 757 -55 791 -51
rect 757 -127 791 -119
rect 757 -204 791 -187
rect -711 -281 -662 -247
rect -628 -281 -579 -247
rect -453 -281 -404 -247
rect -370 -281 -321 -247
rect -195 -281 -146 -247
rect -112 -281 -63 -247
rect 63 -281 112 -247
rect 146 -281 195 -247
rect 321 -281 370 -247
rect 404 -281 453 -247
rect 579 -281 628 -247
rect 662 -281 711 -247
<< viali >>
rect -662 247 -628 281
rect -404 247 -370 281
rect -146 247 -112 281
rect 112 247 146 281
rect 370 247 404 281
rect 628 247 662 281
rect -791 153 -757 161
rect -791 127 -757 153
rect -791 85 -757 89
rect -791 55 -757 85
rect -791 -17 -757 17
rect -791 -85 -757 -55
rect -791 -89 -757 -85
rect -791 -153 -757 -127
rect -791 -161 -757 -153
rect -533 153 -499 161
rect -533 127 -499 153
rect -533 85 -499 89
rect -533 55 -499 85
rect -533 -17 -499 17
rect -533 -85 -499 -55
rect -533 -89 -499 -85
rect -533 -153 -499 -127
rect -533 -161 -499 -153
rect -275 153 -241 161
rect -275 127 -241 153
rect -275 85 -241 89
rect -275 55 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -55
rect -275 -89 -241 -85
rect -275 -153 -241 -127
rect -275 -161 -241 -153
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect 241 153 275 161
rect 241 127 275 153
rect 241 85 275 89
rect 241 55 275 85
rect 241 -17 275 17
rect 241 -85 275 -55
rect 241 -89 275 -85
rect 241 -153 275 -127
rect 241 -161 275 -153
rect 499 153 533 161
rect 499 127 533 153
rect 499 85 533 89
rect 499 55 533 85
rect 499 -17 533 17
rect 499 -85 533 -55
rect 499 -89 533 -85
rect 499 -153 533 -127
rect 499 -161 533 -153
rect 757 153 791 161
rect 757 127 791 153
rect 757 85 791 89
rect 757 55 791 85
rect 757 -17 791 17
rect 757 -85 791 -55
rect 757 -89 791 -85
rect 757 -153 791 -127
rect 757 -161 791 -153
rect -662 -281 -628 -247
rect -404 -281 -370 -247
rect -146 -281 -112 -247
rect 112 -281 146 -247
rect 370 -281 404 -247
rect 628 -281 662 -247
<< metal1 >>
rect -699 281 -591 287
rect -699 247 -662 281
rect -628 247 -591 281
rect -699 241 -591 247
rect -441 281 -333 287
rect -441 247 -404 281
rect -370 247 -333 281
rect -441 241 -333 247
rect -183 281 -75 287
rect -183 247 -146 281
rect -112 247 -75 281
rect -183 241 -75 247
rect 75 281 183 287
rect 75 247 112 281
rect 146 247 183 281
rect 75 241 183 247
rect 333 281 441 287
rect 333 247 370 281
rect 404 247 441 281
rect 333 241 441 247
rect 591 281 699 287
rect 591 247 628 281
rect 662 247 699 281
rect 591 241 699 247
rect -797 161 -751 200
rect -797 127 -791 161
rect -757 127 -751 161
rect -797 89 -751 127
rect -797 55 -791 89
rect -757 55 -751 89
rect -797 17 -751 55
rect -797 -17 -791 17
rect -757 -17 -751 17
rect -797 -55 -751 -17
rect -797 -89 -791 -55
rect -757 -89 -751 -55
rect -797 -127 -751 -89
rect -797 -161 -791 -127
rect -757 -161 -751 -127
rect -797 -200 -751 -161
rect -539 161 -493 200
rect -539 127 -533 161
rect -499 127 -493 161
rect -539 89 -493 127
rect -539 55 -533 89
rect -499 55 -493 89
rect -539 17 -493 55
rect -539 -17 -533 17
rect -499 -17 -493 17
rect -539 -55 -493 -17
rect -539 -89 -533 -55
rect -499 -89 -493 -55
rect -539 -127 -493 -89
rect -539 -161 -533 -127
rect -499 -161 -493 -127
rect -539 -200 -493 -161
rect -281 161 -235 200
rect -281 127 -275 161
rect -241 127 -235 161
rect -281 89 -235 127
rect -281 55 -275 89
rect -241 55 -235 89
rect -281 17 -235 55
rect -281 -17 -275 17
rect -241 -17 -235 17
rect -281 -55 -235 -17
rect -281 -89 -275 -55
rect -241 -89 -235 -55
rect -281 -127 -235 -89
rect -281 -161 -275 -127
rect -241 -161 -235 -127
rect -281 -200 -235 -161
rect -23 161 23 200
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -200 23 -161
rect 235 161 281 200
rect 235 127 241 161
rect 275 127 281 161
rect 235 89 281 127
rect 235 55 241 89
rect 275 55 281 89
rect 235 17 281 55
rect 235 -17 241 17
rect 275 -17 281 17
rect 235 -55 281 -17
rect 235 -89 241 -55
rect 275 -89 281 -55
rect 235 -127 281 -89
rect 235 -161 241 -127
rect 275 -161 281 -127
rect 235 -200 281 -161
rect 493 161 539 200
rect 493 127 499 161
rect 533 127 539 161
rect 493 89 539 127
rect 493 55 499 89
rect 533 55 539 89
rect 493 17 539 55
rect 493 -17 499 17
rect 533 -17 539 17
rect 493 -55 539 -17
rect 493 -89 499 -55
rect 533 -89 539 -55
rect 493 -127 539 -89
rect 493 -161 499 -127
rect 533 -161 539 -127
rect 493 -200 539 -161
rect 751 161 797 200
rect 751 127 757 161
rect 791 127 797 161
rect 751 89 797 127
rect 751 55 757 89
rect 791 55 797 89
rect 751 17 797 55
rect 751 -17 757 17
rect 791 -17 797 17
rect 751 -55 797 -17
rect 751 -89 757 -55
rect 791 -89 797 -55
rect 751 -127 797 -89
rect 751 -161 757 -127
rect 791 -161 797 -127
rect 751 -200 797 -161
rect -699 -247 -591 -241
rect -699 -281 -662 -247
rect -628 -281 -591 -247
rect -699 -287 -591 -281
rect -441 -247 -333 -241
rect -441 -281 -404 -247
rect -370 -281 -333 -247
rect -441 -287 -333 -281
rect -183 -247 -75 -241
rect -183 -281 -146 -247
rect -112 -281 -75 -247
rect -183 -287 -75 -281
rect 75 -247 183 -241
rect 75 -281 112 -247
rect 146 -281 183 -247
rect 75 -287 183 -281
rect 333 -247 441 -241
rect 333 -281 370 -247
rect 404 -281 441 -247
rect 333 -287 441 -281
rect 591 -247 699 -241
rect 591 -281 628 -247
rect 662 -281 699 -247
rect 591 -287 699 -281
<< end >>
