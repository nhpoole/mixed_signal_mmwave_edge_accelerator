magic
tech sky130A
magscale 1 2
timestamp 1622100421
<< nmoslvt >>
rect -358 -100 -158 100
rect -100 -100 100 100
rect 158 -100 358 100
<< ndiff >>
rect -416 88 -358 100
rect -416 -88 -404 88
rect -370 -88 -358 88
rect -416 -100 -358 -88
rect -158 88 -100 100
rect -158 -88 -146 88
rect -112 -88 -100 88
rect -158 -100 -100 -88
rect 100 88 158 100
rect 100 -88 112 88
rect 146 -88 158 88
rect 100 -100 158 -88
rect 358 88 416 100
rect 358 -88 370 88
rect 404 -88 416 88
rect 358 -100 416 -88
<< ndiffc >>
rect -404 -88 -370 88
rect -146 -88 -112 88
rect 112 -88 146 88
rect 370 -88 404 88
<< poly >>
rect -324 172 -192 188
rect -324 155 -308 172
rect -358 138 -308 155
rect -208 155 -192 172
rect -66 172 66 188
rect -66 155 -50 172
rect -208 138 -158 155
rect -358 100 -158 138
rect -100 138 -50 155
rect 50 155 66 172
rect 192 172 324 188
rect 192 155 208 172
rect 50 138 100 155
rect -100 100 100 138
rect 158 138 208 155
rect 308 155 324 172
rect 308 138 358 155
rect 158 100 358 138
rect -358 -138 -158 -100
rect -358 -155 -308 -138
rect -324 -172 -308 -155
rect -208 -155 -158 -138
rect -100 -138 100 -100
rect -100 -155 -50 -138
rect -208 -172 -192 -155
rect -324 -188 -192 -172
rect -66 -172 -50 -155
rect 50 -155 100 -138
rect 158 -138 358 -100
rect 158 -155 208 -138
rect 50 -172 66 -155
rect -66 -188 66 -172
rect 192 -172 208 -155
rect 308 -155 358 -138
rect 308 -172 324 -155
rect 192 -188 324 -172
<< polycont >>
rect -308 138 -208 172
rect -50 138 50 172
rect 208 138 308 172
rect -308 -172 -208 -138
rect -50 -172 50 -138
rect 208 -172 308 -138
<< locali >>
rect -324 138 -308 172
rect -208 138 -192 172
rect -66 138 -50 172
rect 50 138 66 172
rect 192 138 208 172
rect 308 138 324 172
rect -404 88 -370 104
rect -404 -104 -370 -88
rect -146 88 -112 104
rect -146 -104 -112 -88
rect 112 88 146 104
rect 112 -104 146 -88
rect 370 88 404 104
rect 370 -104 404 -88
rect -324 -172 -308 -138
rect -208 -172 -192 -138
rect -66 -172 -50 -138
rect 50 -172 66 -138
rect 192 -172 208 -138
rect 308 -172 324 -138
<< viali >>
rect -300 138 -216 172
rect -42 138 42 172
rect 216 138 300 172
rect -404 -88 -370 88
rect -146 -88 -112 88
rect 112 -88 146 88
rect 370 -88 404 88
rect -300 -172 -216 -138
rect -42 -172 42 -138
rect 216 -172 300 -138
<< metal1 >>
rect -312 172 -204 178
rect -312 138 -300 172
rect -216 138 -204 172
rect -312 132 -204 138
rect -54 172 54 178
rect -54 138 -42 172
rect 42 138 54 172
rect -54 132 54 138
rect 204 172 312 178
rect 204 138 216 172
rect 300 138 312 172
rect 204 132 312 138
rect -410 88 -364 100
rect -410 -88 -404 88
rect -370 -88 -364 88
rect -410 -100 -364 -88
rect -152 88 -106 100
rect -152 -88 -146 88
rect -112 -88 -106 88
rect -152 -100 -106 -88
rect 106 88 152 100
rect 106 -88 112 88
rect 146 -88 152 88
rect 106 -100 152 -88
rect 364 88 410 100
rect 364 -88 370 88
rect 404 -88 410 88
rect 364 -100 410 -88
rect -312 -138 -204 -132
rect -312 -172 -300 -138
rect -216 -172 -204 -138
rect -312 -178 -204 -172
rect -54 -138 54 -132
rect -54 -172 -42 -138
rect 42 -172 54 -138
rect -54 -178 54 -172
rect 204 -138 312 -132
rect 204 -172 216 -138
rect 300 -172 312 -138
rect 204 -178 312 -172
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string parameters w 1 l 1 m 1 nf 3 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
