magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -1309 -1309 3850 2731
<< locali >>
rect 0 1396 2554 1432
rect 0 -18 2554 18
<< metal1 >>
rect -32 1388 32 1440
rect -32 -26 32 26
<< metal2 >>
rect -28 1390 28 1438
rect 137 538 203 590
rect -28 -24 28 24
rect 369 0 397 1414
rect 1858 871 1886 899
rect 2364 489 2392 517
<< metal3 >>
rect -49 1365 49 1463
rect -49 -49 49 49
use sky130_sram_2kbyte_1rw1r_32x512_8_dff_buf_0  sky130_sram_2kbyte_1rw1r_32x512_8_dff_buf_0_0
timestamp 1626486988
transform 1 0 0 0 1 0
box -36 -43 2590 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_0
timestamp 1626486988
transform 1 0 -33 0 1 -37
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_0
timestamp 1626486988
transform 1 0 -32 0 1 -32
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_0
timestamp 1626486988
transform 1 0 -29 0 1 -33
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_1
timestamp 1626486988
transform 1 0 -33 0 1 1377
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_1
timestamp 1626486988
transform 1 0 -32 0 1 1382
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1
timestamp 1626486988
transform 1 0 -29 0 1 1381
box 0 0 58 66
<< labels >>
rlabel metal3 s -49 1365 49 1463 4 vdd
rlabel metal3 s -49 -49 49 49 4 gnd
rlabel metal2 s 137 538 203 590 4 din_0
rlabel metal2 s 2364 489 2392 517 4 dout_0
rlabel metal2 s 1858 871 1886 899 4 dout_bar_0
rlabel metal2 s 369 0 397 1414 4 clk
<< properties >>
string FIXED_BBOX 0 0 2554 1414
<< end >>
