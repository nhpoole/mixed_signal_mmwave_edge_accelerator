magic
tech sky130A
magscale 1 2
timestamp 1620700822
<< error_p >>
rect -2589 2550 -2529 4950
rect -2509 2550 -2449 4950
rect -70 2550 -10 4950
rect 10 2550 70 4950
rect 2449 2550 2509 4950
rect 2529 2550 2589 4950
rect -2589 50 -2529 2450
rect -2509 50 -2449 2450
rect -70 50 -10 2450
rect 10 50 70 2450
rect 2449 50 2509 2450
rect 2529 50 2589 2450
rect -2589 -2450 -2529 -50
rect -2509 -2450 -2449 -50
rect -70 -2450 -10 -50
rect 10 -2450 70 -50
rect 2449 -2450 2509 -50
rect 2529 -2450 2589 -50
rect -2589 -4950 -2529 -2550
rect -2509 -4950 -2449 -2550
rect -70 -4950 -10 -2550
rect 10 -4950 70 -2550
rect 2449 -4950 2509 -2550
rect 2529 -4950 2589 -2550
<< metal3 >>
rect -5028 4922 -2529 4950
rect -5028 2578 -2613 4922
rect -2549 2578 -2529 4922
rect -5028 2550 -2529 2578
rect -2509 4922 -10 4950
rect -2509 2578 -94 4922
rect -30 2578 -10 4922
rect -2509 2550 -10 2578
rect 10 4922 2509 4950
rect 10 2578 2425 4922
rect 2489 2578 2509 4922
rect 10 2550 2509 2578
rect 2529 4922 5028 4950
rect 2529 2578 4944 4922
rect 5008 2578 5028 4922
rect 2529 2550 5028 2578
rect -5028 2422 -2529 2450
rect -5028 78 -2613 2422
rect -2549 78 -2529 2422
rect -5028 50 -2529 78
rect -2509 2422 -10 2450
rect -2509 78 -94 2422
rect -30 78 -10 2422
rect -2509 50 -10 78
rect 10 2422 2509 2450
rect 10 78 2425 2422
rect 2489 78 2509 2422
rect 10 50 2509 78
rect 2529 2422 5028 2450
rect 2529 78 4944 2422
rect 5008 78 5028 2422
rect 2529 50 5028 78
rect -5028 -78 -2529 -50
rect -5028 -2422 -2613 -78
rect -2549 -2422 -2529 -78
rect -5028 -2450 -2529 -2422
rect -2509 -78 -10 -50
rect -2509 -2422 -94 -78
rect -30 -2422 -10 -78
rect -2509 -2450 -10 -2422
rect 10 -78 2509 -50
rect 10 -2422 2425 -78
rect 2489 -2422 2509 -78
rect 10 -2450 2509 -2422
rect 2529 -78 5028 -50
rect 2529 -2422 4944 -78
rect 5008 -2422 5028 -78
rect 2529 -2450 5028 -2422
rect -5028 -2578 -2529 -2550
rect -5028 -4922 -2613 -2578
rect -2549 -4922 -2529 -2578
rect -5028 -4950 -2529 -4922
rect -2509 -2578 -10 -2550
rect -2509 -4922 -94 -2578
rect -30 -4922 -10 -2578
rect -2509 -4950 -10 -4922
rect 10 -2578 2509 -2550
rect 10 -4922 2425 -2578
rect 2489 -4922 2509 -2578
rect 10 -4950 2509 -4922
rect 2529 -2578 5028 -2550
rect 2529 -4922 4944 -2578
rect 5008 -4922 5028 -2578
rect 2529 -4950 5028 -4922
<< via3 >>
rect -2613 2578 -2549 4922
rect -94 2578 -30 4922
rect 2425 2578 2489 4922
rect 4944 2578 5008 4922
rect -2613 78 -2549 2422
rect -94 78 -30 2422
rect 2425 78 2489 2422
rect 4944 78 5008 2422
rect -2613 -2422 -2549 -78
rect -94 -2422 -30 -78
rect 2425 -2422 2489 -78
rect 4944 -2422 5008 -78
rect -2613 -4922 -2549 -2578
rect -94 -4922 -30 -2578
rect 2425 -4922 2489 -2578
rect 4944 -4922 5008 -2578
<< mimcap >>
rect -4928 4810 -2728 4850
rect -4928 2690 -4888 4810
rect -2768 2690 -2728 4810
rect -4928 2650 -2728 2690
rect -2409 4810 -209 4850
rect -2409 2690 -2369 4810
rect -249 2690 -209 4810
rect -2409 2650 -209 2690
rect 110 4810 2310 4850
rect 110 2690 150 4810
rect 2270 2690 2310 4810
rect 110 2650 2310 2690
rect 2629 4810 4829 4850
rect 2629 2690 2669 4810
rect 4789 2690 4829 4810
rect 2629 2650 4829 2690
rect -4928 2310 -2728 2350
rect -4928 190 -4888 2310
rect -2768 190 -2728 2310
rect -4928 150 -2728 190
rect -2409 2310 -209 2350
rect -2409 190 -2369 2310
rect -249 190 -209 2310
rect -2409 150 -209 190
rect 110 2310 2310 2350
rect 110 190 150 2310
rect 2270 190 2310 2310
rect 110 150 2310 190
rect 2629 2310 4829 2350
rect 2629 190 2669 2310
rect 4789 190 4829 2310
rect 2629 150 4829 190
rect -4928 -190 -2728 -150
rect -4928 -2310 -4888 -190
rect -2768 -2310 -2728 -190
rect -4928 -2350 -2728 -2310
rect -2409 -190 -209 -150
rect -2409 -2310 -2369 -190
rect -249 -2310 -209 -190
rect -2409 -2350 -209 -2310
rect 110 -190 2310 -150
rect 110 -2310 150 -190
rect 2270 -2310 2310 -190
rect 110 -2350 2310 -2310
rect 2629 -190 4829 -150
rect 2629 -2310 2669 -190
rect 4789 -2310 4829 -190
rect 2629 -2350 4829 -2310
rect -4928 -2690 -2728 -2650
rect -4928 -4810 -4888 -2690
rect -2768 -4810 -2728 -2690
rect -4928 -4850 -2728 -4810
rect -2409 -2690 -209 -2650
rect -2409 -4810 -2369 -2690
rect -249 -4810 -209 -2690
rect -2409 -4850 -209 -4810
rect 110 -2690 2310 -2650
rect 110 -4810 150 -2690
rect 2270 -4810 2310 -2690
rect 110 -4850 2310 -4810
rect 2629 -2690 4829 -2650
rect 2629 -4810 2669 -2690
rect 4789 -4810 4829 -2690
rect 2629 -4850 4829 -4810
<< mimcapcontact >>
rect -4888 2690 -2768 4810
rect -2369 2690 -249 4810
rect 150 2690 2270 4810
rect 2669 2690 4789 4810
rect -4888 190 -2768 2310
rect -2369 190 -249 2310
rect 150 190 2270 2310
rect 2669 190 4789 2310
rect -4888 -2310 -2768 -190
rect -2369 -2310 -249 -190
rect 150 -2310 2270 -190
rect 2669 -2310 4789 -190
rect -4888 -4810 -2768 -2690
rect -2369 -4810 -249 -2690
rect 150 -4810 2270 -2690
rect 2669 -4810 4789 -2690
<< metal4 >>
rect -3880 4811 -3776 5000
rect -2660 4938 -2556 5000
rect -2660 4922 -2533 4938
rect -4889 4810 -2767 4811
rect -4889 2690 -4888 4810
rect -2768 2690 -2767 4810
rect -4889 2689 -2767 2690
rect -3880 2311 -3776 2689
rect -2660 2578 -2613 4922
rect -2549 2578 -2533 4922
rect -1361 4811 -1257 5000
rect -141 4938 -37 5000
rect -141 4922 -14 4938
rect -2370 4810 -248 4811
rect -2370 2690 -2369 4810
rect -249 2690 -248 4810
rect -2370 2689 -248 2690
rect -2660 2562 -2533 2578
rect -2660 2438 -2556 2562
rect -2660 2422 -2533 2438
rect -4889 2310 -2767 2311
rect -4889 190 -4888 2310
rect -2768 190 -2767 2310
rect -4889 189 -2767 190
rect -3880 -189 -3776 189
rect -2660 78 -2613 2422
rect -2549 78 -2533 2422
rect -1361 2311 -1257 2689
rect -141 2578 -94 4922
rect -30 2578 -14 4922
rect 1158 4811 1262 5000
rect 2378 4938 2482 5000
rect 2378 4922 2505 4938
rect 149 4810 2271 4811
rect 149 2690 150 4810
rect 2270 2690 2271 4810
rect 149 2689 2271 2690
rect -141 2562 -14 2578
rect -141 2438 -37 2562
rect -141 2422 -14 2438
rect -2370 2310 -248 2311
rect -2370 190 -2369 2310
rect -249 190 -248 2310
rect -2370 189 -248 190
rect -2660 62 -2533 78
rect -2660 -62 -2556 62
rect -2660 -78 -2533 -62
rect -4889 -190 -2767 -189
rect -4889 -2310 -4888 -190
rect -2768 -2310 -2767 -190
rect -4889 -2311 -2767 -2310
rect -3880 -2689 -3776 -2311
rect -2660 -2422 -2613 -78
rect -2549 -2422 -2533 -78
rect -1361 -189 -1257 189
rect -141 78 -94 2422
rect -30 78 -14 2422
rect 1158 2311 1262 2689
rect 2378 2578 2425 4922
rect 2489 2578 2505 4922
rect 3677 4811 3781 5000
rect 4897 4938 5001 5000
rect 4897 4922 5024 4938
rect 2668 4810 4790 4811
rect 2668 2690 2669 4810
rect 4789 2690 4790 4810
rect 2668 2689 4790 2690
rect 2378 2562 2505 2578
rect 2378 2438 2482 2562
rect 2378 2422 2505 2438
rect 149 2310 2271 2311
rect 149 190 150 2310
rect 2270 190 2271 2310
rect 149 189 2271 190
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -2370 -190 -248 -189
rect -2370 -2310 -2369 -190
rect -249 -2310 -248 -190
rect -2370 -2311 -248 -2310
rect -2660 -2438 -2533 -2422
rect -2660 -2562 -2556 -2438
rect -2660 -2578 -2533 -2562
rect -4889 -2690 -2767 -2689
rect -4889 -4810 -4888 -2690
rect -2768 -4810 -2767 -2690
rect -4889 -4811 -2767 -4810
rect -3880 -5000 -3776 -4811
rect -2660 -4922 -2613 -2578
rect -2549 -4922 -2533 -2578
rect -1361 -2689 -1257 -2311
rect -141 -2422 -94 -78
rect -30 -2422 -14 -78
rect 1158 -189 1262 189
rect 2378 78 2425 2422
rect 2489 78 2505 2422
rect 3677 2311 3781 2689
rect 4897 2578 4944 4922
rect 5008 2578 5024 4922
rect 4897 2562 5024 2578
rect 4897 2438 5001 2562
rect 4897 2422 5024 2438
rect 2668 2310 4790 2311
rect 2668 190 2669 2310
rect 4789 190 4790 2310
rect 2668 189 4790 190
rect 2378 62 2505 78
rect 2378 -62 2482 62
rect 2378 -78 2505 -62
rect 149 -190 2271 -189
rect 149 -2310 150 -190
rect 2270 -2310 2271 -190
rect 149 -2311 2271 -2310
rect -141 -2438 -14 -2422
rect -141 -2562 -37 -2438
rect -141 -2578 -14 -2562
rect -2370 -2690 -248 -2689
rect -2370 -4810 -2369 -2690
rect -249 -4810 -248 -2690
rect -2370 -4811 -248 -4810
rect -2660 -4938 -2533 -4922
rect -2660 -5000 -2556 -4938
rect -1361 -5000 -1257 -4811
rect -141 -4922 -94 -2578
rect -30 -4922 -14 -2578
rect 1158 -2689 1262 -2311
rect 2378 -2422 2425 -78
rect 2489 -2422 2505 -78
rect 3677 -189 3781 189
rect 4897 78 4944 2422
rect 5008 78 5024 2422
rect 4897 62 5024 78
rect 4897 -62 5001 62
rect 4897 -78 5024 -62
rect 2668 -190 4790 -189
rect 2668 -2310 2669 -190
rect 4789 -2310 4790 -190
rect 2668 -2311 4790 -2310
rect 2378 -2438 2505 -2422
rect 2378 -2562 2482 -2438
rect 2378 -2578 2505 -2562
rect 149 -2690 2271 -2689
rect 149 -4810 150 -2690
rect 2270 -4810 2271 -2690
rect 149 -4811 2271 -4810
rect -141 -4938 -14 -4922
rect -141 -5000 -37 -4938
rect 1158 -5000 1262 -4811
rect 2378 -4922 2425 -2578
rect 2489 -4922 2505 -2578
rect 3677 -2689 3781 -2311
rect 4897 -2422 4944 -78
rect 5008 -2422 5024 -78
rect 4897 -2438 5024 -2422
rect 4897 -2562 5001 -2438
rect 4897 -2578 5024 -2562
rect 2668 -2690 4790 -2689
rect 2668 -4810 2669 -2690
rect 4789 -4810 4790 -2690
rect 2668 -4811 4790 -4810
rect 2378 -4938 2505 -4922
rect 2378 -5000 2482 -4938
rect 3677 -5000 3781 -4811
rect 4897 -4922 4944 -2578
rect 5008 -4922 5024 -2578
rect 4897 -4938 5024 -4922
rect 4897 -5000 5001 -4938
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 2529 2550 4929 4950
string parameters w 11.0 l 11.0 val 128.479 carea 1.00 cperi 0.17 nx 4 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
