magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -9469 -1660 9469 1660
<< nwell >>
rect -8209 -400 8209 400
<< pmoslvt >>
rect -8115 -300 -7155 300
rect -7097 -300 -6137 300
rect -6079 -300 -5119 300
rect -5061 -300 -4101 300
rect -4043 -300 -3083 300
rect -3025 -300 -2065 300
rect -2007 -300 -1047 300
rect -989 -300 -29 300
rect 29 -300 989 300
rect 1047 -300 2007 300
rect 2065 -300 3025 300
rect 3083 -300 4043 300
rect 4101 -300 5061 300
rect 5119 -300 6079 300
rect 6137 -300 7097 300
rect 7155 -300 8115 300
<< pdiff >>
rect -8173 255 -8115 300
rect -8173 221 -8161 255
rect -8127 221 -8115 255
rect -8173 187 -8115 221
rect -8173 153 -8161 187
rect -8127 153 -8115 187
rect -8173 119 -8115 153
rect -8173 85 -8161 119
rect -8127 85 -8115 119
rect -8173 51 -8115 85
rect -8173 17 -8161 51
rect -8127 17 -8115 51
rect -8173 -17 -8115 17
rect -8173 -51 -8161 -17
rect -8127 -51 -8115 -17
rect -8173 -85 -8115 -51
rect -8173 -119 -8161 -85
rect -8127 -119 -8115 -85
rect -8173 -153 -8115 -119
rect -8173 -187 -8161 -153
rect -8127 -187 -8115 -153
rect -8173 -221 -8115 -187
rect -8173 -255 -8161 -221
rect -8127 -255 -8115 -221
rect -8173 -300 -8115 -255
rect -7155 255 -7097 300
rect -7155 221 -7143 255
rect -7109 221 -7097 255
rect -7155 187 -7097 221
rect -7155 153 -7143 187
rect -7109 153 -7097 187
rect -7155 119 -7097 153
rect -7155 85 -7143 119
rect -7109 85 -7097 119
rect -7155 51 -7097 85
rect -7155 17 -7143 51
rect -7109 17 -7097 51
rect -7155 -17 -7097 17
rect -7155 -51 -7143 -17
rect -7109 -51 -7097 -17
rect -7155 -85 -7097 -51
rect -7155 -119 -7143 -85
rect -7109 -119 -7097 -85
rect -7155 -153 -7097 -119
rect -7155 -187 -7143 -153
rect -7109 -187 -7097 -153
rect -7155 -221 -7097 -187
rect -7155 -255 -7143 -221
rect -7109 -255 -7097 -221
rect -7155 -300 -7097 -255
rect -6137 255 -6079 300
rect -6137 221 -6125 255
rect -6091 221 -6079 255
rect -6137 187 -6079 221
rect -6137 153 -6125 187
rect -6091 153 -6079 187
rect -6137 119 -6079 153
rect -6137 85 -6125 119
rect -6091 85 -6079 119
rect -6137 51 -6079 85
rect -6137 17 -6125 51
rect -6091 17 -6079 51
rect -6137 -17 -6079 17
rect -6137 -51 -6125 -17
rect -6091 -51 -6079 -17
rect -6137 -85 -6079 -51
rect -6137 -119 -6125 -85
rect -6091 -119 -6079 -85
rect -6137 -153 -6079 -119
rect -6137 -187 -6125 -153
rect -6091 -187 -6079 -153
rect -6137 -221 -6079 -187
rect -6137 -255 -6125 -221
rect -6091 -255 -6079 -221
rect -6137 -300 -6079 -255
rect -5119 255 -5061 300
rect -5119 221 -5107 255
rect -5073 221 -5061 255
rect -5119 187 -5061 221
rect -5119 153 -5107 187
rect -5073 153 -5061 187
rect -5119 119 -5061 153
rect -5119 85 -5107 119
rect -5073 85 -5061 119
rect -5119 51 -5061 85
rect -5119 17 -5107 51
rect -5073 17 -5061 51
rect -5119 -17 -5061 17
rect -5119 -51 -5107 -17
rect -5073 -51 -5061 -17
rect -5119 -85 -5061 -51
rect -5119 -119 -5107 -85
rect -5073 -119 -5061 -85
rect -5119 -153 -5061 -119
rect -5119 -187 -5107 -153
rect -5073 -187 -5061 -153
rect -5119 -221 -5061 -187
rect -5119 -255 -5107 -221
rect -5073 -255 -5061 -221
rect -5119 -300 -5061 -255
rect -4101 255 -4043 300
rect -4101 221 -4089 255
rect -4055 221 -4043 255
rect -4101 187 -4043 221
rect -4101 153 -4089 187
rect -4055 153 -4043 187
rect -4101 119 -4043 153
rect -4101 85 -4089 119
rect -4055 85 -4043 119
rect -4101 51 -4043 85
rect -4101 17 -4089 51
rect -4055 17 -4043 51
rect -4101 -17 -4043 17
rect -4101 -51 -4089 -17
rect -4055 -51 -4043 -17
rect -4101 -85 -4043 -51
rect -4101 -119 -4089 -85
rect -4055 -119 -4043 -85
rect -4101 -153 -4043 -119
rect -4101 -187 -4089 -153
rect -4055 -187 -4043 -153
rect -4101 -221 -4043 -187
rect -4101 -255 -4089 -221
rect -4055 -255 -4043 -221
rect -4101 -300 -4043 -255
rect -3083 255 -3025 300
rect -3083 221 -3071 255
rect -3037 221 -3025 255
rect -3083 187 -3025 221
rect -3083 153 -3071 187
rect -3037 153 -3025 187
rect -3083 119 -3025 153
rect -3083 85 -3071 119
rect -3037 85 -3025 119
rect -3083 51 -3025 85
rect -3083 17 -3071 51
rect -3037 17 -3025 51
rect -3083 -17 -3025 17
rect -3083 -51 -3071 -17
rect -3037 -51 -3025 -17
rect -3083 -85 -3025 -51
rect -3083 -119 -3071 -85
rect -3037 -119 -3025 -85
rect -3083 -153 -3025 -119
rect -3083 -187 -3071 -153
rect -3037 -187 -3025 -153
rect -3083 -221 -3025 -187
rect -3083 -255 -3071 -221
rect -3037 -255 -3025 -221
rect -3083 -300 -3025 -255
rect -2065 255 -2007 300
rect -2065 221 -2053 255
rect -2019 221 -2007 255
rect -2065 187 -2007 221
rect -2065 153 -2053 187
rect -2019 153 -2007 187
rect -2065 119 -2007 153
rect -2065 85 -2053 119
rect -2019 85 -2007 119
rect -2065 51 -2007 85
rect -2065 17 -2053 51
rect -2019 17 -2007 51
rect -2065 -17 -2007 17
rect -2065 -51 -2053 -17
rect -2019 -51 -2007 -17
rect -2065 -85 -2007 -51
rect -2065 -119 -2053 -85
rect -2019 -119 -2007 -85
rect -2065 -153 -2007 -119
rect -2065 -187 -2053 -153
rect -2019 -187 -2007 -153
rect -2065 -221 -2007 -187
rect -2065 -255 -2053 -221
rect -2019 -255 -2007 -221
rect -2065 -300 -2007 -255
rect -1047 255 -989 300
rect -1047 221 -1035 255
rect -1001 221 -989 255
rect -1047 187 -989 221
rect -1047 153 -1035 187
rect -1001 153 -989 187
rect -1047 119 -989 153
rect -1047 85 -1035 119
rect -1001 85 -989 119
rect -1047 51 -989 85
rect -1047 17 -1035 51
rect -1001 17 -989 51
rect -1047 -17 -989 17
rect -1047 -51 -1035 -17
rect -1001 -51 -989 -17
rect -1047 -85 -989 -51
rect -1047 -119 -1035 -85
rect -1001 -119 -989 -85
rect -1047 -153 -989 -119
rect -1047 -187 -1035 -153
rect -1001 -187 -989 -153
rect -1047 -221 -989 -187
rect -1047 -255 -1035 -221
rect -1001 -255 -989 -221
rect -1047 -300 -989 -255
rect -29 255 29 300
rect -29 221 -17 255
rect 17 221 29 255
rect -29 187 29 221
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -221 29 -187
rect -29 -255 -17 -221
rect 17 -255 29 -221
rect -29 -300 29 -255
rect 989 255 1047 300
rect 989 221 1001 255
rect 1035 221 1047 255
rect 989 187 1047 221
rect 989 153 1001 187
rect 1035 153 1047 187
rect 989 119 1047 153
rect 989 85 1001 119
rect 1035 85 1047 119
rect 989 51 1047 85
rect 989 17 1001 51
rect 1035 17 1047 51
rect 989 -17 1047 17
rect 989 -51 1001 -17
rect 1035 -51 1047 -17
rect 989 -85 1047 -51
rect 989 -119 1001 -85
rect 1035 -119 1047 -85
rect 989 -153 1047 -119
rect 989 -187 1001 -153
rect 1035 -187 1047 -153
rect 989 -221 1047 -187
rect 989 -255 1001 -221
rect 1035 -255 1047 -221
rect 989 -300 1047 -255
rect 2007 255 2065 300
rect 2007 221 2019 255
rect 2053 221 2065 255
rect 2007 187 2065 221
rect 2007 153 2019 187
rect 2053 153 2065 187
rect 2007 119 2065 153
rect 2007 85 2019 119
rect 2053 85 2065 119
rect 2007 51 2065 85
rect 2007 17 2019 51
rect 2053 17 2065 51
rect 2007 -17 2065 17
rect 2007 -51 2019 -17
rect 2053 -51 2065 -17
rect 2007 -85 2065 -51
rect 2007 -119 2019 -85
rect 2053 -119 2065 -85
rect 2007 -153 2065 -119
rect 2007 -187 2019 -153
rect 2053 -187 2065 -153
rect 2007 -221 2065 -187
rect 2007 -255 2019 -221
rect 2053 -255 2065 -221
rect 2007 -300 2065 -255
rect 3025 255 3083 300
rect 3025 221 3037 255
rect 3071 221 3083 255
rect 3025 187 3083 221
rect 3025 153 3037 187
rect 3071 153 3083 187
rect 3025 119 3083 153
rect 3025 85 3037 119
rect 3071 85 3083 119
rect 3025 51 3083 85
rect 3025 17 3037 51
rect 3071 17 3083 51
rect 3025 -17 3083 17
rect 3025 -51 3037 -17
rect 3071 -51 3083 -17
rect 3025 -85 3083 -51
rect 3025 -119 3037 -85
rect 3071 -119 3083 -85
rect 3025 -153 3083 -119
rect 3025 -187 3037 -153
rect 3071 -187 3083 -153
rect 3025 -221 3083 -187
rect 3025 -255 3037 -221
rect 3071 -255 3083 -221
rect 3025 -300 3083 -255
rect 4043 255 4101 300
rect 4043 221 4055 255
rect 4089 221 4101 255
rect 4043 187 4101 221
rect 4043 153 4055 187
rect 4089 153 4101 187
rect 4043 119 4101 153
rect 4043 85 4055 119
rect 4089 85 4101 119
rect 4043 51 4101 85
rect 4043 17 4055 51
rect 4089 17 4101 51
rect 4043 -17 4101 17
rect 4043 -51 4055 -17
rect 4089 -51 4101 -17
rect 4043 -85 4101 -51
rect 4043 -119 4055 -85
rect 4089 -119 4101 -85
rect 4043 -153 4101 -119
rect 4043 -187 4055 -153
rect 4089 -187 4101 -153
rect 4043 -221 4101 -187
rect 4043 -255 4055 -221
rect 4089 -255 4101 -221
rect 4043 -300 4101 -255
rect 5061 255 5119 300
rect 5061 221 5073 255
rect 5107 221 5119 255
rect 5061 187 5119 221
rect 5061 153 5073 187
rect 5107 153 5119 187
rect 5061 119 5119 153
rect 5061 85 5073 119
rect 5107 85 5119 119
rect 5061 51 5119 85
rect 5061 17 5073 51
rect 5107 17 5119 51
rect 5061 -17 5119 17
rect 5061 -51 5073 -17
rect 5107 -51 5119 -17
rect 5061 -85 5119 -51
rect 5061 -119 5073 -85
rect 5107 -119 5119 -85
rect 5061 -153 5119 -119
rect 5061 -187 5073 -153
rect 5107 -187 5119 -153
rect 5061 -221 5119 -187
rect 5061 -255 5073 -221
rect 5107 -255 5119 -221
rect 5061 -300 5119 -255
rect 6079 255 6137 300
rect 6079 221 6091 255
rect 6125 221 6137 255
rect 6079 187 6137 221
rect 6079 153 6091 187
rect 6125 153 6137 187
rect 6079 119 6137 153
rect 6079 85 6091 119
rect 6125 85 6137 119
rect 6079 51 6137 85
rect 6079 17 6091 51
rect 6125 17 6137 51
rect 6079 -17 6137 17
rect 6079 -51 6091 -17
rect 6125 -51 6137 -17
rect 6079 -85 6137 -51
rect 6079 -119 6091 -85
rect 6125 -119 6137 -85
rect 6079 -153 6137 -119
rect 6079 -187 6091 -153
rect 6125 -187 6137 -153
rect 6079 -221 6137 -187
rect 6079 -255 6091 -221
rect 6125 -255 6137 -221
rect 6079 -300 6137 -255
rect 7097 255 7155 300
rect 7097 221 7109 255
rect 7143 221 7155 255
rect 7097 187 7155 221
rect 7097 153 7109 187
rect 7143 153 7155 187
rect 7097 119 7155 153
rect 7097 85 7109 119
rect 7143 85 7155 119
rect 7097 51 7155 85
rect 7097 17 7109 51
rect 7143 17 7155 51
rect 7097 -17 7155 17
rect 7097 -51 7109 -17
rect 7143 -51 7155 -17
rect 7097 -85 7155 -51
rect 7097 -119 7109 -85
rect 7143 -119 7155 -85
rect 7097 -153 7155 -119
rect 7097 -187 7109 -153
rect 7143 -187 7155 -153
rect 7097 -221 7155 -187
rect 7097 -255 7109 -221
rect 7143 -255 7155 -221
rect 7097 -300 7155 -255
rect 8115 255 8173 300
rect 8115 221 8127 255
rect 8161 221 8173 255
rect 8115 187 8173 221
rect 8115 153 8127 187
rect 8161 153 8173 187
rect 8115 119 8173 153
rect 8115 85 8127 119
rect 8161 85 8173 119
rect 8115 51 8173 85
rect 8115 17 8127 51
rect 8161 17 8173 51
rect 8115 -17 8173 17
rect 8115 -51 8127 -17
rect 8161 -51 8173 -17
rect 8115 -85 8173 -51
rect 8115 -119 8127 -85
rect 8161 -119 8173 -85
rect 8115 -153 8173 -119
rect 8115 -187 8127 -153
rect 8161 -187 8173 -153
rect 8115 -221 8173 -187
rect 8115 -255 8127 -221
rect 8161 -255 8173 -221
rect 8115 -300 8173 -255
<< pdiffc >>
rect -8161 221 -8127 255
rect -8161 153 -8127 187
rect -8161 85 -8127 119
rect -8161 17 -8127 51
rect -8161 -51 -8127 -17
rect -8161 -119 -8127 -85
rect -8161 -187 -8127 -153
rect -8161 -255 -8127 -221
rect -7143 221 -7109 255
rect -7143 153 -7109 187
rect -7143 85 -7109 119
rect -7143 17 -7109 51
rect -7143 -51 -7109 -17
rect -7143 -119 -7109 -85
rect -7143 -187 -7109 -153
rect -7143 -255 -7109 -221
rect -6125 221 -6091 255
rect -6125 153 -6091 187
rect -6125 85 -6091 119
rect -6125 17 -6091 51
rect -6125 -51 -6091 -17
rect -6125 -119 -6091 -85
rect -6125 -187 -6091 -153
rect -6125 -255 -6091 -221
rect -5107 221 -5073 255
rect -5107 153 -5073 187
rect -5107 85 -5073 119
rect -5107 17 -5073 51
rect -5107 -51 -5073 -17
rect -5107 -119 -5073 -85
rect -5107 -187 -5073 -153
rect -5107 -255 -5073 -221
rect -4089 221 -4055 255
rect -4089 153 -4055 187
rect -4089 85 -4055 119
rect -4089 17 -4055 51
rect -4089 -51 -4055 -17
rect -4089 -119 -4055 -85
rect -4089 -187 -4055 -153
rect -4089 -255 -4055 -221
rect -3071 221 -3037 255
rect -3071 153 -3037 187
rect -3071 85 -3037 119
rect -3071 17 -3037 51
rect -3071 -51 -3037 -17
rect -3071 -119 -3037 -85
rect -3071 -187 -3037 -153
rect -3071 -255 -3037 -221
rect -2053 221 -2019 255
rect -2053 153 -2019 187
rect -2053 85 -2019 119
rect -2053 17 -2019 51
rect -2053 -51 -2019 -17
rect -2053 -119 -2019 -85
rect -2053 -187 -2019 -153
rect -2053 -255 -2019 -221
rect -1035 221 -1001 255
rect -1035 153 -1001 187
rect -1035 85 -1001 119
rect -1035 17 -1001 51
rect -1035 -51 -1001 -17
rect -1035 -119 -1001 -85
rect -1035 -187 -1001 -153
rect -1035 -255 -1001 -221
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect 1001 221 1035 255
rect 1001 153 1035 187
rect 1001 85 1035 119
rect 1001 17 1035 51
rect 1001 -51 1035 -17
rect 1001 -119 1035 -85
rect 1001 -187 1035 -153
rect 1001 -255 1035 -221
rect 2019 221 2053 255
rect 2019 153 2053 187
rect 2019 85 2053 119
rect 2019 17 2053 51
rect 2019 -51 2053 -17
rect 2019 -119 2053 -85
rect 2019 -187 2053 -153
rect 2019 -255 2053 -221
rect 3037 221 3071 255
rect 3037 153 3071 187
rect 3037 85 3071 119
rect 3037 17 3071 51
rect 3037 -51 3071 -17
rect 3037 -119 3071 -85
rect 3037 -187 3071 -153
rect 3037 -255 3071 -221
rect 4055 221 4089 255
rect 4055 153 4089 187
rect 4055 85 4089 119
rect 4055 17 4089 51
rect 4055 -51 4089 -17
rect 4055 -119 4089 -85
rect 4055 -187 4089 -153
rect 4055 -255 4089 -221
rect 5073 221 5107 255
rect 5073 153 5107 187
rect 5073 85 5107 119
rect 5073 17 5107 51
rect 5073 -51 5107 -17
rect 5073 -119 5107 -85
rect 5073 -187 5107 -153
rect 5073 -255 5107 -221
rect 6091 221 6125 255
rect 6091 153 6125 187
rect 6091 85 6125 119
rect 6091 17 6125 51
rect 6091 -51 6125 -17
rect 6091 -119 6125 -85
rect 6091 -187 6125 -153
rect 6091 -255 6125 -221
rect 7109 221 7143 255
rect 7109 153 7143 187
rect 7109 85 7143 119
rect 7109 17 7143 51
rect 7109 -51 7143 -17
rect 7109 -119 7143 -85
rect 7109 -187 7143 -153
rect 7109 -255 7143 -221
rect 8127 221 8161 255
rect 8127 153 8161 187
rect 8127 85 8161 119
rect 8127 17 8161 51
rect 8127 -51 8161 -17
rect 8127 -119 8161 -85
rect 8127 -187 8161 -153
rect 8127 -255 8161 -221
<< poly >>
rect -7929 381 -7341 397
rect -7929 364 -7890 381
rect -8115 347 -7890 364
rect -7856 347 -7822 381
rect -7788 347 -7754 381
rect -7720 347 -7686 381
rect -7652 347 -7618 381
rect -7584 347 -7550 381
rect -7516 347 -7482 381
rect -7448 347 -7414 381
rect -7380 364 -7341 381
rect -6911 381 -6323 397
rect -6911 364 -6872 381
rect -7380 347 -7155 364
rect -8115 300 -7155 347
rect -7097 347 -6872 364
rect -6838 347 -6804 381
rect -6770 347 -6736 381
rect -6702 347 -6668 381
rect -6634 347 -6600 381
rect -6566 347 -6532 381
rect -6498 347 -6464 381
rect -6430 347 -6396 381
rect -6362 364 -6323 381
rect -5893 381 -5305 397
rect -5893 364 -5854 381
rect -6362 347 -6137 364
rect -7097 300 -6137 347
rect -6079 347 -5854 364
rect -5820 347 -5786 381
rect -5752 347 -5718 381
rect -5684 347 -5650 381
rect -5616 347 -5582 381
rect -5548 347 -5514 381
rect -5480 347 -5446 381
rect -5412 347 -5378 381
rect -5344 364 -5305 381
rect -4875 381 -4287 397
rect -4875 364 -4836 381
rect -5344 347 -5119 364
rect -6079 300 -5119 347
rect -5061 347 -4836 364
rect -4802 347 -4768 381
rect -4734 347 -4700 381
rect -4666 347 -4632 381
rect -4598 347 -4564 381
rect -4530 347 -4496 381
rect -4462 347 -4428 381
rect -4394 347 -4360 381
rect -4326 364 -4287 381
rect -3857 381 -3269 397
rect -3857 364 -3818 381
rect -4326 347 -4101 364
rect -5061 300 -4101 347
rect -4043 347 -3818 364
rect -3784 347 -3750 381
rect -3716 347 -3682 381
rect -3648 347 -3614 381
rect -3580 347 -3546 381
rect -3512 347 -3478 381
rect -3444 347 -3410 381
rect -3376 347 -3342 381
rect -3308 364 -3269 381
rect -2839 381 -2251 397
rect -2839 364 -2800 381
rect -3308 347 -3083 364
rect -4043 300 -3083 347
rect -3025 347 -2800 364
rect -2766 347 -2732 381
rect -2698 347 -2664 381
rect -2630 347 -2596 381
rect -2562 347 -2528 381
rect -2494 347 -2460 381
rect -2426 347 -2392 381
rect -2358 347 -2324 381
rect -2290 364 -2251 381
rect -1821 381 -1233 397
rect -1821 364 -1782 381
rect -2290 347 -2065 364
rect -3025 300 -2065 347
rect -2007 347 -1782 364
rect -1748 347 -1714 381
rect -1680 347 -1646 381
rect -1612 347 -1578 381
rect -1544 347 -1510 381
rect -1476 347 -1442 381
rect -1408 347 -1374 381
rect -1340 347 -1306 381
rect -1272 364 -1233 381
rect -803 381 -215 397
rect -803 364 -764 381
rect -1272 347 -1047 364
rect -2007 300 -1047 347
rect -989 347 -764 364
rect -730 347 -696 381
rect -662 347 -628 381
rect -594 347 -560 381
rect -526 347 -492 381
rect -458 347 -424 381
rect -390 347 -356 381
rect -322 347 -288 381
rect -254 364 -215 381
rect 215 381 803 397
rect 215 364 254 381
rect -254 347 -29 364
rect -989 300 -29 347
rect 29 347 254 364
rect 288 347 322 381
rect 356 347 390 381
rect 424 347 458 381
rect 492 347 526 381
rect 560 347 594 381
rect 628 347 662 381
rect 696 347 730 381
rect 764 364 803 381
rect 1233 381 1821 397
rect 1233 364 1272 381
rect 764 347 989 364
rect 29 300 989 347
rect 1047 347 1272 364
rect 1306 347 1340 381
rect 1374 347 1408 381
rect 1442 347 1476 381
rect 1510 347 1544 381
rect 1578 347 1612 381
rect 1646 347 1680 381
rect 1714 347 1748 381
rect 1782 364 1821 381
rect 2251 381 2839 397
rect 2251 364 2290 381
rect 1782 347 2007 364
rect 1047 300 2007 347
rect 2065 347 2290 364
rect 2324 347 2358 381
rect 2392 347 2426 381
rect 2460 347 2494 381
rect 2528 347 2562 381
rect 2596 347 2630 381
rect 2664 347 2698 381
rect 2732 347 2766 381
rect 2800 364 2839 381
rect 3269 381 3857 397
rect 3269 364 3308 381
rect 2800 347 3025 364
rect 2065 300 3025 347
rect 3083 347 3308 364
rect 3342 347 3376 381
rect 3410 347 3444 381
rect 3478 347 3512 381
rect 3546 347 3580 381
rect 3614 347 3648 381
rect 3682 347 3716 381
rect 3750 347 3784 381
rect 3818 364 3857 381
rect 4287 381 4875 397
rect 4287 364 4326 381
rect 3818 347 4043 364
rect 3083 300 4043 347
rect 4101 347 4326 364
rect 4360 347 4394 381
rect 4428 347 4462 381
rect 4496 347 4530 381
rect 4564 347 4598 381
rect 4632 347 4666 381
rect 4700 347 4734 381
rect 4768 347 4802 381
rect 4836 364 4875 381
rect 5305 381 5893 397
rect 5305 364 5344 381
rect 4836 347 5061 364
rect 4101 300 5061 347
rect 5119 347 5344 364
rect 5378 347 5412 381
rect 5446 347 5480 381
rect 5514 347 5548 381
rect 5582 347 5616 381
rect 5650 347 5684 381
rect 5718 347 5752 381
rect 5786 347 5820 381
rect 5854 364 5893 381
rect 6323 381 6911 397
rect 6323 364 6362 381
rect 5854 347 6079 364
rect 5119 300 6079 347
rect 6137 347 6362 364
rect 6396 347 6430 381
rect 6464 347 6498 381
rect 6532 347 6566 381
rect 6600 347 6634 381
rect 6668 347 6702 381
rect 6736 347 6770 381
rect 6804 347 6838 381
rect 6872 364 6911 381
rect 7341 381 7929 397
rect 7341 364 7380 381
rect 6872 347 7097 364
rect 6137 300 7097 347
rect 7155 347 7380 364
rect 7414 347 7448 381
rect 7482 347 7516 381
rect 7550 347 7584 381
rect 7618 347 7652 381
rect 7686 347 7720 381
rect 7754 347 7788 381
rect 7822 347 7856 381
rect 7890 364 7929 381
rect 7890 347 8115 364
rect 7155 300 8115 347
rect -8115 -347 -7155 -300
rect -8115 -364 -7890 -347
rect -7929 -381 -7890 -364
rect -7856 -381 -7822 -347
rect -7788 -381 -7754 -347
rect -7720 -381 -7686 -347
rect -7652 -381 -7618 -347
rect -7584 -381 -7550 -347
rect -7516 -381 -7482 -347
rect -7448 -381 -7414 -347
rect -7380 -364 -7155 -347
rect -7097 -347 -6137 -300
rect -7097 -364 -6872 -347
rect -7380 -381 -7341 -364
rect -7929 -397 -7341 -381
rect -6911 -381 -6872 -364
rect -6838 -381 -6804 -347
rect -6770 -381 -6736 -347
rect -6702 -381 -6668 -347
rect -6634 -381 -6600 -347
rect -6566 -381 -6532 -347
rect -6498 -381 -6464 -347
rect -6430 -381 -6396 -347
rect -6362 -364 -6137 -347
rect -6079 -347 -5119 -300
rect -6079 -364 -5854 -347
rect -6362 -381 -6323 -364
rect -6911 -397 -6323 -381
rect -5893 -381 -5854 -364
rect -5820 -381 -5786 -347
rect -5752 -381 -5718 -347
rect -5684 -381 -5650 -347
rect -5616 -381 -5582 -347
rect -5548 -381 -5514 -347
rect -5480 -381 -5446 -347
rect -5412 -381 -5378 -347
rect -5344 -364 -5119 -347
rect -5061 -347 -4101 -300
rect -5061 -364 -4836 -347
rect -5344 -381 -5305 -364
rect -5893 -397 -5305 -381
rect -4875 -381 -4836 -364
rect -4802 -381 -4768 -347
rect -4734 -381 -4700 -347
rect -4666 -381 -4632 -347
rect -4598 -381 -4564 -347
rect -4530 -381 -4496 -347
rect -4462 -381 -4428 -347
rect -4394 -381 -4360 -347
rect -4326 -364 -4101 -347
rect -4043 -347 -3083 -300
rect -4043 -364 -3818 -347
rect -4326 -381 -4287 -364
rect -4875 -397 -4287 -381
rect -3857 -381 -3818 -364
rect -3784 -381 -3750 -347
rect -3716 -381 -3682 -347
rect -3648 -381 -3614 -347
rect -3580 -381 -3546 -347
rect -3512 -381 -3478 -347
rect -3444 -381 -3410 -347
rect -3376 -381 -3342 -347
rect -3308 -364 -3083 -347
rect -3025 -347 -2065 -300
rect -3025 -364 -2800 -347
rect -3308 -381 -3269 -364
rect -3857 -397 -3269 -381
rect -2839 -381 -2800 -364
rect -2766 -381 -2732 -347
rect -2698 -381 -2664 -347
rect -2630 -381 -2596 -347
rect -2562 -381 -2528 -347
rect -2494 -381 -2460 -347
rect -2426 -381 -2392 -347
rect -2358 -381 -2324 -347
rect -2290 -364 -2065 -347
rect -2007 -347 -1047 -300
rect -2007 -364 -1782 -347
rect -2290 -381 -2251 -364
rect -2839 -397 -2251 -381
rect -1821 -381 -1782 -364
rect -1748 -381 -1714 -347
rect -1680 -381 -1646 -347
rect -1612 -381 -1578 -347
rect -1544 -381 -1510 -347
rect -1476 -381 -1442 -347
rect -1408 -381 -1374 -347
rect -1340 -381 -1306 -347
rect -1272 -364 -1047 -347
rect -989 -347 -29 -300
rect -989 -364 -764 -347
rect -1272 -381 -1233 -364
rect -1821 -397 -1233 -381
rect -803 -381 -764 -364
rect -730 -381 -696 -347
rect -662 -381 -628 -347
rect -594 -381 -560 -347
rect -526 -381 -492 -347
rect -458 -381 -424 -347
rect -390 -381 -356 -347
rect -322 -381 -288 -347
rect -254 -364 -29 -347
rect 29 -347 989 -300
rect 29 -364 254 -347
rect -254 -381 -215 -364
rect -803 -397 -215 -381
rect 215 -381 254 -364
rect 288 -381 322 -347
rect 356 -381 390 -347
rect 424 -381 458 -347
rect 492 -381 526 -347
rect 560 -381 594 -347
rect 628 -381 662 -347
rect 696 -381 730 -347
rect 764 -364 989 -347
rect 1047 -347 2007 -300
rect 1047 -364 1272 -347
rect 764 -381 803 -364
rect 215 -397 803 -381
rect 1233 -381 1272 -364
rect 1306 -381 1340 -347
rect 1374 -381 1408 -347
rect 1442 -381 1476 -347
rect 1510 -381 1544 -347
rect 1578 -381 1612 -347
rect 1646 -381 1680 -347
rect 1714 -381 1748 -347
rect 1782 -364 2007 -347
rect 2065 -347 3025 -300
rect 2065 -364 2290 -347
rect 1782 -381 1821 -364
rect 1233 -397 1821 -381
rect 2251 -381 2290 -364
rect 2324 -381 2358 -347
rect 2392 -381 2426 -347
rect 2460 -381 2494 -347
rect 2528 -381 2562 -347
rect 2596 -381 2630 -347
rect 2664 -381 2698 -347
rect 2732 -381 2766 -347
rect 2800 -364 3025 -347
rect 3083 -347 4043 -300
rect 3083 -364 3308 -347
rect 2800 -381 2839 -364
rect 2251 -397 2839 -381
rect 3269 -381 3308 -364
rect 3342 -381 3376 -347
rect 3410 -381 3444 -347
rect 3478 -381 3512 -347
rect 3546 -381 3580 -347
rect 3614 -381 3648 -347
rect 3682 -381 3716 -347
rect 3750 -381 3784 -347
rect 3818 -364 4043 -347
rect 4101 -347 5061 -300
rect 4101 -364 4326 -347
rect 3818 -381 3857 -364
rect 3269 -397 3857 -381
rect 4287 -381 4326 -364
rect 4360 -381 4394 -347
rect 4428 -381 4462 -347
rect 4496 -381 4530 -347
rect 4564 -381 4598 -347
rect 4632 -381 4666 -347
rect 4700 -381 4734 -347
rect 4768 -381 4802 -347
rect 4836 -364 5061 -347
rect 5119 -347 6079 -300
rect 5119 -364 5344 -347
rect 4836 -381 4875 -364
rect 4287 -397 4875 -381
rect 5305 -381 5344 -364
rect 5378 -381 5412 -347
rect 5446 -381 5480 -347
rect 5514 -381 5548 -347
rect 5582 -381 5616 -347
rect 5650 -381 5684 -347
rect 5718 -381 5752 -347
rect 5786 -381 5820 -347
rect 5854 -364 6079 -347
rect 6137 -347 7097 -300
rect 6137 -364 6362 -347
rect 5854 -381 5893 -364
rect 5305 -397 5893 -381
rect 6323 -381 6362 -364
rect 6396 -381 6430 -347
rect 6464 -381 6498 -347
rect 6532 -381 6566 -347
rect 6600 -381 6634 -347
rect 6668 -381 6702 -347
rect 6736 -381 6770 -347
rect 6804 -381 6838 -347
rect 6872 -364 7097 -347
rect 7155 -347 8115 -300
rect 7155 -364 7380 -347
rect 6872 -381 6911 -364
rect 6323 -397 6911 -381
rect 7341 -381 7380 -364
rect 7414 -381 7448 -347
rect 7482 -381 7516 -347
rect 7550 -381 7584 -347
rect 7618 -381 7652 -347
rect 7686 -381 7720 -347
rect 7754 -381 7788 -347
rect 7822 -381 7856 -347
rect 7890 -364 8115 -347
rect 7890 -381 7929 -364
rect 7341 -397 7929 -381
<< polycont >>
rect -7890 347 -7856 381
rect -7822 347 -7788 381
rect -7754 347 -7720 381
rect -7686 347 -7652 381
rect -7618 347 -7584 381
rect -7550 347 -7516 381
rect -7482 347 -7448 381
rect -7414 347 -7380 381
rect -6872 347 -6838 381
rect -6804 347 -6770 381
rect -6736 347 -6702 381
rect -6668 347 -6634 381
rect -6600 347 -6566 381
rect -6532 347 -6498 381
rect -6464 347 -6430 381
rect -6396 347 -6362 381
rect -5854 347 -5820 381
rect -5786 347 -5752 381
rect -5718 347 -5684 381
rect -5650 347 -5616 381
rect -5582 347 -5548 381
rect -5514 347 -5480 381
rect -5446 347 -5412 381
rect -5378 347 -5344 381
rect -4836 347 -4802 381
rect -4768 347 -4734 381
rect -4700 347 -4666 381
rect -4632 347 -4598 381
rect -4564 347 -4530 381
rect -4496 347 -4462 381
rect -4428 347 -4394 381
rect -4360 347 -4326 381
rect -3818 347 -3784 381
rect -3750 347 -3716 381
rect -3682 347 -3648 381
rect -3614 347 -3580 381
rect -3546 347 -3512 381
rect -3478 347 -3444 381
rect -3410 347 -3376 381
rect -3342 347 -3308 381
rect -2800 347 -2766 381
rect -2732 347 -2698 381
rect -2664 347 -2630 381
rect -2596 347 -2562 381
rect -2528 347 -2494 381
rect -2460 347 -2426 381
rect -2392 347 -2358 381
rect -2324 347 -2290 381
rect -1782 347 -1748 381
rect -1714 347 -1680 381
rect -1646 347 -1612 381
rect -1578 347 -1544 381
rect -1510 347 -1476 381
rect -1442 347 -1408 381
rect -1374 347 -1340 381
rect -1306 347 -1272 381
rect -764 347 -730 381
rect -696 347 -662 381
rect -628 347 -594 381
rect -560 347 -526 381
rect -492 347 -458 381
rect -424 347 -390 381
rect -356 347 -322 381
rect -288 347 -254 381
rect 254 347 288 381
rect 322 347 356 381
rect 390 347 424 381
rect 458 347 492 381
rect 526 347 560 381
rect 594 347 628 381
rect 662 347 696 381
rect 730 347 764 381
rect 1272 347 1306 381
rect 1340 347 1374 381
rect 1408 347 1442 381
rect 1476 347 1510 381
rect 1544 347 1578 381
rect 1612 347 1646 381
rect 1680 347 1714 381
rect 1748 347 1782 381
rect 2290 347 2324 381
rect 2358 347 2392 381
rect 2426 347 2460 381
rect 2494 347 2528 381
rect 2562 347 2596 381
rect 2630 347 2664 381
rect 2698 347 2732 381
rect 2766 347 2800 381
rect 3308 347 3342 381
rect 3376 347 3410 381
rect 3444 347 3478 381
rect 3512 347 3546 381
rect 3580 347 3614 381
rect 3648 347 3682 381
rect 3716 347 3750 381
rect 3784 347 3818 381
rect 4326 347 4360 381
rect 4394 347 4428 381
rect 4462 347 4496 381
rect 4530 347 4564 381
rect 4598 347 4632 381
rect 4666 347 4700 381
rect 4734 347 4768 381
rect 4802 347 4836 381
rect 5344 347 5378 381
rect 5412 347 5446 381
rect 5480 347 5514 381
rect 5548 347 5582 381
rect 5616 347 5650 381
rect 5684 347 5718 381
rect 5752 347 5786 381
rect 5820 347 5854 381
rect 6362 347 6396 381
rect 6430 347 6464 381
rect 6498 347 6532 381
rect 6566 347 6600 381
rect 6634 347 6668 381
rect 6702 347 6736 381
rect 6770 347 6804 381
rect 6838 347 6872 381
rect 7380 347 7414 381
rect 7448 347 7482 381
rect 7516 347 7550 381
rect 7584 347 7618 381
rect 7652 347 7686 381
rect 7720 347 7754 381
rect 7788 347 7822 381
rect 7856 347 7890 381
rect -7890 -381 -7856 -347
rect -7822 -381 -7788 -347
rect -7754 -381 -7720 -347
rect -7686 -381 -7652 -347
rect -7618 -381 -7584 -347
rect -7550 -381 -7516 -347
rect -7482 -381 -7448 -347
rect -7414 -381 -7380 -347
rect -6872 -381 -6838 -347
rect -6804 -381 -6770 -347
rect -6736 -381 -6702 -347
rect -6668 -381 -6634 -347
rect -6600 -381 -6566 -347
rect -6532 -381 -6498 -347
rect -6464 -381 -6430 -347
rect -6396 -381 -6362 -347
rect -5854 -381 -5820 -347
rect -5786 -381 -5752 -347
rect -5718 -381 -5684 -347
rect -5650 -381 -5616 -347
rect -5582 -381 -5548 -347
rect -5514 -381 -5480 -347
rect -5446 -381 -5412 -347
rect -5378 -381 -5344 -347
rect -4836 -381 -4802 -347
rect -4768 -381 -4734 -347
rect -4700 -381 -4666 -347
rect -4632 -381 -4598 -347
rect -4564 -381 -4530 -347
rect -4496 -381 -4462 -347
rect -4428 -381 -4394 -347
rect -4360 -381 -4326 -347
rect -3818 -381 -3784 -347
rect -3750 -381 -3716 -347
rect -3682 -381 -3648 -347
rect -3614 -381 -3580 -347
rect -3546 -381 -3512 -347
rect -3478 -381 -3444 -347
rect -3410 -381 -3376 -347
rect -3342 -381 -3308 -347
rect -2800 -381 -2766 -347
rect -2732 -381 -2698 -347
rect -2664 -381 -2630 -347
rect -2596 -381 -2562 -347
rect -2528 -381 -2494 -347
rect -2460 -381 -2426 -347
rect -2392 -381 -2358 -347
rect -2324 -381 -2290 -347
rect -1782 -381 -1748 -347
rect -1714 -381 -1680 -347
rect -1646 -381 -1612 -347
rect -1578 -381 -1544 -347
rect -1510 -381 -1476 -347
rect -1442 -381 -1408 -347
rect -1374 -381 -1340 -347
rect -1306 -381 -1272 -347
rect -764 -381 -730 -347
rect -696 -381 -662 -347
rect -628 -381 -594 -347
rect -560 -381 -526 -347
rect -492 -381 -458 -347
rect -424 -381 -390 -347
rect -356 -381 -322 -347
rect -288 -381 -254 -347
rect 254 -381 288 -347
rect 322 -381 356 -347
rect 390 -381 424 -347
rect 458 -381 492 -347
rect 526 -381 560 -347
rect 594 -381 628 -347
rect 662 -381 696 -347
rect 730 -381 764 -347
rect 1272 -381 1306 -347
rect 1340 -381 1374 -347
rect 1408 -381 1442 -347
rect 1476 -381 1510 -347
rect 1544 -381 1578 -347
rect 1612 -381 1646 -347
rect 1680 -381 1714 -347
rect 1748 -381 1782 -347
rect 2290 -381 2324 -347
rect 2358 -381 2392 -347
rect 2426 -381 2460 -347
rect 2494 -381 2528 -347
rect 2562 -381 2596 -347
rect 2630 -381 2664 -347
rect 2698 -381 2732 -347
rect 2766 -381 2800 -347
rect 3308 -381 3342 -347
rect 3376 -381 3410 -347
rect 3444 -381 3478 -347
rect 3512 -381 3546 -347
rect 3580 -381 3614 -347
rect 3648 -381 3682 -347
rect 3716 -381 3750 -347
rect 3784 -381 3818 -347
rect 4326 -381 4360 -347
rect 4394 -381 4428 -347
rect 4462 -381 4496 -347
rect 4530 -381 4564 -347
rect 4598 -381 4632 -347
rect 4666 -381 4700 -347
rect 4734 -381 4768 -347
rect 4802 -381 4836 -347
rect 5344 -381 5378 -347
rect 5412 -381 5446 -347
rect 5480 -381 5514 -347
rect 5548 -381 5582 -347
rect 5616 -381 5650 -347
rect 5684 -381 5718 -347
rect 5752 -381 5786 -347
rect 5820 -381 5854 -347
rect 6362 -381 6396 -347
rect 6430 -381 6464 -347
rect 6498 -381 6532 -347
rect 6566 -381 6600 -347
rect 6634 -381 6668 -347
rect 6702 -381 6736 -347
rect 6770 -381 6804 -347
rect 6838 -381 6872 -347
rect 7380 -381 7414 -347
rect 7448 -381 7482 -347
rect 7516 -381 7550 -347
rect 7584 -381 7618 -347
rect 7652 -381 7686 -347
rect 7720 -381 7754 -347
rect 7788 -381 7822 -347
rect 7856 -381 7890 -347
<< locali >>
rect -7929 347 -7890 381
rect -7856 347 -7832 381
rect -7788 347 -7760 381
rect -7720 347 -7688 381
rect -7652 347 -7618 381
rect -7582 347 -7550 381
rect -7510 347 -7482 381
rect -7438 347 -7414 381
rect -7380 347 -7341 381
rect -6911 347 -6872 381
rect -6838 347 -6814 381
rect -6770 347 -6742 381
rect -6702 347 -6670 381
rect -6634 347 -6600 381
rect -6564 347 -6532 381
rect -6492 347 -6464 381
rect -6420 347 -6396 381
rect -6362 347 -6323 381
rect -5893 347 -5854 381
rect -5820 347 -5796 381
rect -5752 347 -5724 381
rect -5684 347 -5652 381
rect -5616 347 -5582 381
rect -5546 347 -5514 381
rect -5474 347 -5446 381
rect -5402 347 -5378 381
rect -5344 347 -5305 381
rect -4875 347 -4836 381
rect -4802 347 -4778 381
rect -4734 347 -4706 381
rect -4666 347 -4634 381
rect -4598 347 -4564 381
rect -4528 347 -4496 381
rect -4456 347 -4428 381
rect -4384 347 -4360 381
rect -4326 347 -4287 381
rect -3857 347 -3818 381
rect -3784 347 -3760 381
rect -3716 347 -3688 381
rect -3648 347 -3616 381
rect -3580 347 -3546 381
rect -3510 347 -3478 381
rect -3438 347 -3410 381
rect -3366 347 -3342 381
rect -3308 347 -3269 381
rect -2839 347 -2800 381
rect -2766 347 -2742 381
rect -2698 347 -2670 381
rect -2630 347 -2598 381
rect -2562 347 -2528 381
rect -2492 347 -2460 381
rect -2420 347 -2392 381
rect -2348 347 -2324 381
rect -2290 347 -2251 381
rect -1821 347 -1782 381
rect -1748 347 -1724 381
rect -1680 347 -1652 381
rect -1612 347 -1580 381
rect -1544 347 -1510 381
rect -1474 347 -1442 381
rect -1402 347 -1374 381
rect -1330 347 -1306 381
rect -1272 347 -1233 381
rect -803 347 -764 381
rect -730 347 -706 381
rect -662 347 -634 381
rect -594 347 -562 381
rect -526 347 -492 381
rect -456 347 -424 381
rect -384 347 -356 381
rect -312 347 -288 381
rect -254 347 -215 381
rect 215 347 254 381
rect 288 347 312 381
rect 356 347 384 381
rect 424 347 456 381
rect 492 347 526 381
rect 562 347 594 381
rect 634 347 662 381
rect 706 347 730 381
rect 764 347 803 381
rect 1233 347 1272 381
rect 1306 347 1330 381
rect 1374 347 1402 381
rect 1442 347 1474 381
rect 1510 347 1544 381
rect 1580 347 1612 381
rect 1652 347 1680 381
rect 1724 347 1748 381
rect 1782 347 1821 381
rect 2251 347 2290 381
rect 2324 347 2348 381
rect 2392 347 2420 381
rect 2460 347 2492 381
rect 2528 347 2562 381
rect 2598 347 2630 381
rect 2670 347 2698 381
rect 2742 347 2766 381
rect 2800 347 2839 381
rect 3269 347 3308 381
rect 3342 347 3366 381
rect 3410 347 3438 381
rect 3478 347 3510 381
rect 3546 347 3580 381
rect 3616 347 3648 381
rect 3688 347 3716 381
rect 3760 347 3784 381
rect 3818 347 3857 381
rect 4287 347 4326 381
rect 4360 347 4384 381
rect 4428 347 4456 381
rect 4496 347 4528 381
rect 4564 347 4598 381
rect 4634 347 4666 381
rect 4706 347 4734 381
rect 4778 347 4802 381
rect 4836 347 4875 381
rect 5305 347 5344 381
rect 5378 347 5402 381
rect 5446 347 5474 381
rect 5514 347 5546 381
rect 5582 347 5616 381
rect 5652 347 5684 381
rect 5724 347 5752 381
rect 5796 347 5820 381
rect 5854 347 5893 381
rect 6323 347 6362 381
rect 6396 347 6420 381
rect 6464 347 6492 381
rect 6532 347 6564 381
rect 6600 347 6634 381
rect 6670 347 6702 381
rect 6742 347 6770 381
rect 6814 347 6838 381
rect 6872 347 6911 381
rect 7341 347 7380 381
rect 7414 347 7438 381
rect 7482 347 7510 381
rect 7550 347 7582 381
rect 7618 347 7652 381
rect 7688 347 7720 381
rect 7760 347 7788 381
rect 7832 347 7856 381
rect 7890 347 7929 381
rect -8161 269 -8127 304
rect -8161 197 -8127 221
rect -8161 125 -8127 153
rect -8161 53 -8127 85
rect -8161 -17 -8127 17
rect -8161 -85 -8127 -53
rect -8161 -153 -8127 -125
rect -8161 -221 -8127 -197
rect -8161 -304 -8127 -269
rect -7143 269 -7109 304
rect -7143 197 -7109 221
rect -7143 125 -7109 153
rect -7143 53 -7109 85
rect -7143 -17 -7109 17
rect -7143 -85 -7109 -53
rect -7143 -153 -7109 -125
rect -7143 -221 -7109 -197
rect -7143 -304 -7109 -269
rect -6125 269 -6091 304
rect -6125 197 -6091 221
rect -6125 125 -6091 153
rect -6125 53 -6091 85
rect -6125 -17 -6091 17
rect -6125 -85 -6091 -53
rect -6125 -153 -6091 -125
rect -6125 -221 -6091 -197
rect -6125 -304 -6091 -269
rect -5107 269 -5073 304
rect -5107 197 -5073 221
rect -5107 125 -5073 153
rect -5107 53 -5073 85
rect -5107 -17 -5073 17
rect -5107 -85 -5073 -53
rect -5107 -153 -5073 -125
rect -5107 -221 -5073 -197
rect -5107 -304 -5073 -269
rect -4089 269 -4055 304
rect -4089 197 -4055 221
rect -4089 125 -4055 153
rect -4089 53 -4055 85
rect -4089 -17 -4055 17
rect -4089 -85 -4055 -53
rect -4089 -153 -4055 -125
rect -4089 -221 -4055 -197
rect -4089 -304 -4055 -269
rect -3071 269 -3037 304
rect -3071 197 -3037 221
rect -3071 125 -3037 153
rect -3071 53 -3037 85
rect -3071 -17 -3037 17
rect -3071 -85 -3037 -53
rect -3071 -153 -3037 -125
rect -3071 -221 -3037 -197
rect -3071 -304 -3037 -269
rect -2053 269 -2019 304
rect -2053 197 -2019 221
rect -2053 125 -2019 153
rect -2053 53 -2019 85
rect -2053 -17 -2019 17
rect -2053 -85 -2019 -53
rect -2053 -153 -2019 -125
rect -2053 -221 -2019 -197
rect -2053 -304 -2019 -269
rect -1035 269 -1001 304
rect -1035 197 -1001 221
rect -1035 125 -1001 153
rect -1035 53 -1001 85
rect -1035 -17 -1001 17
rect -1035 -85 -1001 -53
rect -1035 -153 -1001 -125
rect -1035 -221 -1001 -197
rect -1035 -304 -1001 -269
rect -17 269 17 304
rect -17 197 17 221
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -221 17 -197
rect -17 -304 17 -269
rect 1001 269 1035 304
rect 1001 197 1035 221
rect 1001 125 1035 153
rect 1001 53 1035 85
rect 1001 -17 1035 17
rect 1001 -85 1035 -53
rect 1001 -153 1035 -125
rect 1001 -221 1035 -197
rect 1001 -304 1035 -269
rect 2019 269 2053 304
rect 2019 197 2053 221
rect 2019 125 2053 153
rect 2019 53 2053 85
rect 2019 -17 2053 17
rect 2019 -85 2053 -53
rect 2019 -153 2053 -125
rect 2019 -221 2053 -197
rect 2019 -304 2053 -269
rect 3037 269 3071 304
rect 3037 197 3071 221
rect 3037 125 3071 153
rect 3037 53 3071 85
rect 3037 -17 3071 17
rect 3037 -85 3071 -53
rect 3037 -153 3071 -125
rect 3037 -221 3071 -197
rect 3037 -304 3071 -269
rect 4055 269 4089 304
rect 4055 197 4089 221
rect 4055 125 4089 153
rect 4055 53 4089 85
rect 4055 -17 4089 17
rect 4055 -85 4089 -53
rect 4055 -153 4089 -125
rect 4055 -221 4089 -197
rect 4055 -304 4089 -269
rect 5073 269 5107 304
rect 5073 197 5107 221
rect 5073 125 5107 153
rect 5073 53 5107 85
rect 5073 -17 5107 17
rect 5073 -85 5107 -53
rect 5073 -153 5107 -125
rect 5073 -221 5107 -197
rect 5073 -304 5107 -269
rect 6091 269 6125 304
rect 6091 197 6125 221
rect 6091 125 6125 153
rect 6091 53 6125 85
rect 6091 -17 6125 17
rect 6091 -85 6125 -53
rect 6091 -153 6125 -125
rect 6091 -221 6125 -197
rect 6091 -304 6125 -269
rect 7109 269 7143 304
rect 7109 197 7143 221
rect 7109 125 7143 153
rect 7109 53 7143 85
rect 7109 -17 7143 17
rect 7109 -85 7143 -53
rect 7109 -153 7143 -125
rect 7109 -221 7143 -197
rect 7109 -304 7143 -269
rect 8127 269 8161 304
rect 8127 197 8161 221
rect 8127 125 8161 153
rect 8127 53 8161 85
rect 8127 -17 8161 17
rect 8127 -85 8161 -53
rect 8127 -153 8161 -125
rect 8127 -221 8161 -197
rect 8127 -304 8161 -269
rect -7929 -381 -7890 -347
rect -7856 -381 -7832 -347
rect -7788 -381 -7760 -347
rect -7720 -381 -7688 -347
rect -7652 -381 -7618 -347
rect -7582 -381 -7550 -347
rect -7510 -381 -7482 -347
rect -7438 -381 -7414 -347
rect -7380 -381 -7341 -347
rect -6911 -381 -6872 -347
rect -6838 -381 -6814 -347
rect -6770 -381 -6742 -347
rect -6702 -381 -6670 -347
rect -6634 -381 -6600 -347
rect -6564 -381 -6532 -347
rect -6492 -381 -6464 -347
rect -6420 -381 -6396 -347
rect -6362 -381 -6323 -347
rect -5893 -381 -5854 -347
rect -5820 -381 -5796 -347
rect -5752 -381 -5724 -347
rect -5684 -381 -5652 -347
rect -5616 -381 -5582 -347
rect -5546 -381 -5514 -347
rect -5474 -381 -5446 -347
rect -5402 -381 -5378 -347
rect -5344 -381 -5305 -347
rect -4875 -381 -4836 -347
rect -4802 -381 -4778 -347
rect -4734 -381 -4706 -347
rect -4666 -381 -4634 -347
rect -4598 -381 -4564 -347
rect -4528 -381 -4496 -347
rect -4456 -381 -4428 -347
rect -4384 -381 -4360 -347
rect -4326 -381 -4287 -347
rect -3857 -381 -3818 -347
rect -3784 -381 -3760 -347
rect -3716 -381 -3688 -347
rect -3648 -381 -3616 -347
rect -3580 -381 -3546 -347
rect -3510 -381 -3478 -347
rect -3438 -381 -3410 -347
rect -3366 -381 -3342 -347
rect -3308 -381 -3269 -347
rect -2839 -381 -2800 -347
rect -2766 -381 -2742 -347
rect -2698 -381 -2670 -347
rect -2630 -381 -2598 -347
rect -2562 -381 -2528 -347
rect -2492 -381 -2460 -347
rect -2420 -381 -2392 -347
rect -2348 -381 -2324 -347
rect -2290 -381 -2251 -347
rect -1821 -381 -1782 -347
rect -1748 -381 -1724 -347
rect -1680 -381 -1652 -347
rect -1612 -381 -1580 -347
rect -1544 -381 -1510 -347
rect -1474 -381 -1442 -347
rect -1402 -381 -1374 -347
rect -1330 -381 -1306 -347
rect -1272 -381 -1233 -347
rect -803 -381 -764 -347
rect -730 -381 -706 -347
rect -662 -381 -634 -347
rect -594 -381 -562 -347
rect -526 -381 -492 -347
rect -456 -381 -424 -347
rect -384 -381 -356 -347
rect -312 -381 -288 -347
rect -254 -381 -215 -347
rect 215 -381 254 -347
rect 288 -381 312 -347
rect 356 -381 384 -347
rect 424 -381 456 -347
rect 492 -381 526 -347
rect 562 -381 594 -347
rect 634 -381 662 -347
rect 706 -381 730 -347
rect 764 -381 803 -347
rect 1233 -381 1272 -347
rect 1306 -381 1330 -347
rect 1374 -381 1402 -347
rect 1442 -381 1474 -347
rect 1510 -381 1544 -347
rect 1580 -381 1612 -347
rect 1652 -381 1680 -347
rect 1724 -381 1748 -347
rect 1782 -381 1821 -347
rect 2251 -381 2290 -347
rect 2324 -381 2348 -347
rect 2392 -381 2420 -347
rect 2460 -381 2492 -347
rect 2528 -381 2562 -347
rect 2598 -381 2630 -347
rect 2670 -381 2698 -347
rect 2742 -381 2766 -347
rect 2800 -381 2839 -347
rect 3269 -381 3308 -347
rect 3342 -381 3366 -347
rect 3410 -381 3438 -347
rect 3478 -381 3510 -347
rect 3546 -381 3580 -347
rect 3616 -381 3648 -347
rect 3688 -381 3716 -347
rect 3760 -381 3784 -347
rect 3818 -381 3857 -347
rect 4287 -381 4326 -347
rect 4360 -381 4384 -347
rect 4428 -381 4456 -347
rect 4496 -381 4528 -347
rect 4564 -381 4598 -347
rect 4634 -381 4666 -347
rect 4706 -381 4734 -347
rect 4778 -381 4802 -347
rect 4836 -381 4875 -347
rect 5305 -381 5344 -347
rect 5378 -381 5402 -347
rect 5446 -381 5474 -347
rect 5514 -381 5546 -347
rect 5582 -381 5616 -347
rect 5652 -381 5684 -347
rect 5724 -381 5752 -347
rect 5796 -381 5820 -347
rect 5854 -381 5893 -347
rect 6323 -381 6362 -347
rect 6396 -381 6420 -347
rect 6464 -381 6492 -347
rect 6532 -381 6564 -347
rect 6600 -381 6634 -347
rect 6670 -381 6702 -347
rect 6742 -381 6770 -347
rect 6814 -381 6838 -347
rect 6872 -381 6911 -347
rect 7341 -381 7380 -347
rect 7414 -381 7438 -347
rect 7482 -381 7510 -347
rect 7550 -381 7582 -347
rect 7618 -381 7652 -347
rect 7688 -381 7720 -347
rect 7760 -381 7788 -347
rect 7832 -381 7856 -347
rect 7890 -381 7929 -347
<< viali >>
rect -7832 347 -7822 381
rect -7822 347 -7798 381
rect -7760 347 -7754 381
rect -7754 347 -7726 381
rect -7688 347 -7686 381
rect -7686 347 -7654 381
rect -7616 347 -7584 381
rect -7584 347 -7582 381
rect -7544 347 -7516 381
rect -7516 347 -7510 381
rect -7472 347 -7448 381
rect -7448 347 -7438 381
rect -6814 347 -6804 381
rect -6804 347 -6780 381
rect -6742 347 -6736 381
rect -6736 347 -6708 381
rect -6670 347 -6668 381
rect -6668 347 -6636 381
rect -6598 347 -6566 381
rect -6566 347 -6564 381
rect -6526 347 -6498 381
rect -6498 347 -6492 381
rect -6454 347 -6430 381
rect -6430 347 -6420 381
rect -5796 347 -5786 381
rect -5786 347 -5762 381
rect -5724 347 -5718 381
rect -5718 347 -5690 381
rect -5652 347 -5650 381
rect -5650 347 -5618 381
rect -5580 347 -5548 381
rect -5548 347 -5546 381
rect -5508 347 -5480 381
rect -5480 347 -5474 381
rect -5436 347 -5412 381
rect -5412 347 -5402 381
rect -4778 347 -4768 381
rect -4768 347 -4744 381
rect -4706 347 -4700 381
rect -4700 347 -4672 381
rect -4634 347 -4632 381
rect -4632 347 -4600 381
rect -4562 347 -4530 381
rect -4530 347 -4528 381
rect -4490 347 -4462 381
rect -4462 347 -4456 381
rect -4418 347 -4394 381
rect -4394 347 -4384 381
rect -3760 347 -3750 381
rect -3750 347 -3726 381
rect -3688 347 -3682 381
rect -3682 347 -3654 381
rect -3616 347 -3614 381
rect -3614 347 -3582 381
rect -3544 347 -3512 381
rect -3512 347 -3510 381
rect -3472 347 -3444 381
rect -3444 347 -3438 381
rect -3400 347 -3376 381
rect -3376 347 -3366 381
rect -2742 347 -2732 381
rect -2732 347 -2708 381
rect -2670 347 -2664 381
rect -2664 347 -2636 381
rect -2598 347 -2596 381
rect -2596 347 -2564 381
rect -2526 347 -2494 381
rect -2494 347 -2492 381
rect -2454 347 -2426 381
rect -2426 347 -2420 381
rect -2382 347 -2358 381
rect -2358 347 -2348 381
rect -1724 347 -1714 381
rect -1714 347 -1690 381
rect -1652 347 -1646 381
rect -1646 347 -1618 381
rect -1580 347 -1578 381
rect -1578 347 -1546 381
rect -1508 347 -1476 381
rect -1476 347 -1474 381
rect -1436 347 -1408 381
rect -1408 347 -1402 381
rect -1364 347 -1340 381
rect -1340 347 -1330 381
rect -706 347 -696 381
rect -696 347 -672 381
rect -634 347 -628 381
rect -628 347 -600 381
rect -562 347 -560 381
rect -560 347 -528 381
rect -490 347 -458 381
rect -458 347 -456 381
rect -418 347 -390 381
rect -390 347 -384 381
rect -346 347 -322 381
rect -322 347 -312 381
rect 312 347 322 381
rect 322 347 346 381
rect 384 347 390 381
rect 390 347 418 381
rect 456 347 458 381
rect 458 347 490 381
rect 528 347 560 381
rect 560 347 562 381
rect 600 347 628 381
rect 628 347 634 381
rect 672 347 696 381
rect 696 347 706 381
rect 1330 347 1340 381
rect 1340 347 1364 381
rect 1402 347 1408 381
rect 1408 347 1436 381
rect 1474 347 1476 381
rect 1476 347 1508 381
rect 1546 347 1578 381
rect 1578 347 1580 381
rect 1618 347 1646 381
rect 1646 347 1652 381
rect 1690 347 1714 381
rect 1714 347 1724 381
rect 2348 347 2358 381
rect 2358 347 2382 381
rect 2420 347 2426 381
rect 2426 347 2454 381
rect 2492 347 2494 381
rect 2494 347 2526 381
rect 2564 347 2596 381
rect 2596 347 2598 381
rect 2636 347 2664 381
rect 2664 347 2670 381
rect 2708 347 2732 381
rect 2732 347 2742 381
rect 3366 347 3376 381
rect 3376 347 3400 381
rect 3438 347 3444 381
rect 3444 347 3472 381
rect 3510 347 3512 381
rect 3512 347 3544 381
rect 3582 347 3614 381
rect 3614 347 3616 381
rect 3654 347 3682 381
rect 3682 347 3688 381
rect 3726 347 3750 381
rect 3750 347 3760 381
rect 4384 347 4394 381
rect 4394 347 4418 381
rect 4456 347 4462 381
rect 4462 347 4490 381
rect 4528 347 4530 381
rect 4530 347 4562 381
rect 4600 347 4632 381
rect 4632 347 4634 381
rect 4672 347 4700 381
rect 4700 347 4706 381
rect 4744 347 4768 381
rect 4768 347 4778 381
rect 5402 347 5412 381
rect 5412 347 5436 381
rect 5474 347 5480 381
rect 5480 347 5508 381
rect 5546 347 5548 381
rect 5548 347 5580 381
rect 5618 347 5650 381
rect 5650 347 5652 381
rect 5690 347 5718 381
rect 5718 347 5724 381
rect 5762 347 5786 381
rect 5786 347 5796 381
rect 6420 347 6430 381
rect 6430 347 6454 381
rect 6492 347 6498 381
rect 6498 347 6526 381
rect 6564 347 6566 381
rect 6566 347 6598 381
rect 6636 347 6668 381
rect 6668 347 6670 381
rect 6708 347 6736 381
rect 6736 347 6742 381
rect 6780 347 6804 381
rect 6804 347 6814 381
rect 7438 347 7448 381
rect 7448 347 7472 381
rect 7510 347 7516 381
rect 7516 347 7544 381
rect 7582 347 7584 381
rect 7584 347 7616 381
rect 7654 347 7686 381
rect 7686 347 7688 381
rect 7726 347 7754 381
rect 7754 347 7760 381
rect 7798 347 7822 381
rect 7822 347 7832 381
rect -8161 255 -8127 269
rect -8161 235 -8127 255
rect -8161 187 -8127 197
rect -8161 163 -8127 187
rect -8161 119 -8127 125
rect -8161 91 -8127 119
rect -8161 51 -8127 53
rect -8161 19 -8127 51
rect -8161 -51 -8127 -19
rect -8161 -53 -8127 -51
rect -8161 -119 -8127 -91
rect -8161 -125 -8127 -119
rect -8161 -187 -8127 -163
rect -8161 -197 -8127 -187
rect -8161 -255 -8127 -235
rect -8161 -269 -8127 -255
rect -7143 255 -7109 269
rect -7143 235 -7109 255
rect -7143 187 -7109 197
rect -7143 163 -7109 187
rect -7143 119 -7109 125
rect -7143 91 -7109 119
rect -7143 51 -7109 53
rect -7143 19 -7109 51
rect -7143 -51 -7109 -19
rect -7143 -53 -7109 -51
rect -7143 -119 -7109 -91
rect -7143 -125 -7109 -119
rect -7143 -187 -7109 -163
rect -7143 -197 -7109 -187
rect -7143 -255 -7109 -235
rect -7143 -269 -7109 -255
rect -6125 255 -6091 269
rect -6125 235 -6091 255
rect -6125 187 -6091 197
rect -6125 163 -6091 187
rect -6125 119 -6091 125
rect -6125 91 -6091 119
rect -6125 51 -6091 53
rect -6125 19 -6091 51
rect -6125 -51 -6091 -19
rect -6125 -53 -6091 -51
rect -6125 -119 -6091 -91
rect -6125 -125 -6091 -119
rect -6125 -187 -6091 -163
rect -6125 -197 -6091 -187
rect -6125 -255 -6091 -235
rect -6125 -269 -6091 -255
rect -5107 255 -5073 269
rect -5107 235 -5073 255
rect -5107 187 -5073 197
rect -5107 163 -5073 187
rect -5107 119 -5073 125
rect -5107 91 -5073 119
rect -5107 51 -5073 53
rect -5107 19 -5073 51
rect -5107 -51 -5073 -19
rect -5107 -53 -5073 -51
rect -5107 -119 -5073 -91
rect -5107 -125 -5073 -119
rect -5107 -187 -5073 -163
rect -5107 -197 -5073 -187
rect -5107 -255 -5073 -235
rect -5107 -269 -5073 -255
rect -4089 255 -4055 269
rect -4089 235 -4055 255
rect -4089 187 -4055 197
rect -4089 163 -4055 187
rect -4089 119 -4055 125
rect -4089 91 -4055 119
rect -4089 51 -4055 53
rect -4089 19 -4055 51
rect -4089 -51 -4055 -19
rect -4089 -53 -4055 -51
rect -4089 -119 -4055 -91
rect -4089 -125 -4055 -119
rect -4089 -187 -4055 -163
rect -4089 -197 -4055 -187
rect -4089 -255 -4055 -235
rect -4089 -269 -4055 -255
rect -3071 255 -3037 269
rect -3071 235 -3037 255
rect -3071 187 -3037 197
rect -3071 163 -3037 187
rect -3071 119 -3037 125
rect -3071 91 -3037 119
rect -3071 51 -3037 53
rect -3071 19 -3037 51
rect -3071 -51 -3037 -19
rect -3071 -53 -3037 -51
rect -3071 -119 -3037 -91
rect -3071 -125 -3037 -119
rect -3071 -187 -3037 -163
rect -3071 -197 -3037 -187
rect -3071 -255 -3037 -235
rect -3071 -269 -3037 -255
rect -2053 255 -2019 269
rect -2053 235 -2019 255
rect -2053 187 -2019 197
rect -2053 163 -2019 187
rect -2053 119 -2019 125
rect -2053 91 -2019 119
rect -2053 51 -2019 53
rect -2053 19 -2019 51
rect -2053 -51 -2019 -19
rect -2053 -53 -2019 -51
rect -2053 -119 -2019 -91
rect -2053 -125 -2019 -119
rect -2053 -187 -2019 -163
rect -2053 -197 -2019 -187
rect -2053 -255 -2019 -235
rect -2053 -269 -2019 -255
rect -1035 255 -1001 269
rect -1035 235 -1001 255
rect -1035 187 -1001 197
rect -1035 163 -1001 187
rect -1035 119 -1001 125
rect -1035 91 -1001 119
rect -1035 51 -1001 53
rect -1035 19 -1001 51
rect -1035 -51 -1001 -19
rect -1035 -53 -1001 -51
rect -1035 -119 -1001 -91
rect -1035 -125 -1001 -119
rect -1035 -187 -1001 -163
rect -1035 -197 -1001 -187
rect -1035 -255 -1001 -235
rect -1035 -269 -1001 -255
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect 1001 255 1035 269
rect 1001 235 1035 255
rect 1001 187 1035 197
rect 1001 163 1035 187
rect 1001 119 1035 125
rect 1001 91 1035 119
rect 1001 51 1035 53
rect 1001 19 1035 51
rect 1001 -51 1035 -19
rect 1001 -53 1035 -51
rect 1001 -119 1035 -91
rect 1001 -125 1035 -119
rect 1001 -187 1035 -163
rect 1001 -197 1035 -187
rect 1001 -255 1035 -235
rect 1001 -269 1035 -255
rect 2019 255 2053 269
rect 2019 235 2053 255
rect 2019 187 2053 197
rect 2019 163 2053 187
rect 2019 119 2053 125
rect 2019 91 2053 119
rect 2019 51 2053 53
rect 2019 19 2053 51
rect 2019 -51 2053 -19
rect 2019 -53 2053 -51
rect 2019 -119 2053 -91
rect 2019 -125 2053 -119
rect 2019 -187 2053 -163
rect 2019 -197 2053 -187
rect 2019 -255 2053 -235
rect 2019 -269 2053 -255
rect 3037 255 3071 269
rect 3037 235 3071 255
rect 3037 187 3071 197
rect 3037 163 3071 187
rect 3037 119 3071 125
rect 3037 91 3071 119
rect 3037 51 3071 53
rect 3037 19 3071 51
rect 3037 -51 3071 -19
rect 3037 -53 3071 -51
rect 3037 -119 3071 -91
rect 3037 -125 3071 -119
rect 3037 -187 3071 -163
rect 3037 -197 3071 -187
rect 3037 -255 3071 -235
rect 3037 -269 3071 -255
rect 4055 255 4089 269
rect 4055 235 4089 255
rect 4055 187 4089 197
rect 4055 163 4089 187
rect 4055 119 4089 125
rect 4055 91 4089 119
rect 4055 51 4089 53
rect 4055 19 4089 51
rect 4055 -51 4089 -19
rect 4055 -53 4089 -51
rect 4055 -119 4089 -91
rect 4055 -125 4089 -119
rect 4055 -187 4089 -163
rect 4055 -197 4089 -187
rect 4055 -255 4089 -235
rect 4055 -269 4089 -255
rect 5073 255 5107 269
rect 5073 235 5107 255
rect 5073 187 5107 197
rect 5073 163 5107 187
rect 5073 119 5107 125
rect 5073 91 5107 119
rect 5073 51 5107 53
rect 5073 19 5107 51
rect 5073 -51 5107 -19
rect 5073 -53 5107 -51
rect 5073 -119 5107 -91
rect 5073 -125 5107 -119
rect 5073 -187 5107 -163
rect 5073 -197 5107 -187
rect 5073 -255 5107 -235
rect 5073 -269 5107 -255
rect 6091 255 6125 269
rect 6091 235 6125 255
rect 6091 187 6125 197
rect 6091 163 6125 187
rect 6091 119 6125 125
rect 6091 91 6125 119
rect 6091 51 6125 53
rect 6091 19 6125 51
rect 6091 -51 6125 -19
rect 6091 -53 6125 -51
rect 6091 -119 6125 -91
rect 6091 -125 6125 -119
rect 6091 -187 6125 -163
rect 6091 -197 6125 -187
rect 6091 -255 6125 -235
rect 6091 -269 6125 -255
rect 7109 255 7143 269
rect 7109 235 7143 255
rect 7109 187 7143 197
rect 7109 163 7143 187
rect 7109 119 7143 125
rect 7109 91 7143 119
rect 7109 51 7143 53
rect 7109 19 7143 51
rect 7109 -51 7143 -19
rect 7109 -53 7143 -51
rect 7109 -119 7143 -91
rect 7109 -125 7143 -119
rect 7109 -187 7143 -163
rect 7109 -197 7143 -187
rect 7109 -255 7143 -235
rect 7109 -269 7143 -255
rect 8127 255 8161 269
rect 8127 235 8161 255
rect 8127 187 8161 197
rect 8127 163 8161 187
rect 8127 119 8161 125
rect 8127 91 8161 119
rect 8127 51 8161 53
rect 8127 19 8161 51
rect 8127 -51 8161 -19
rect 8127 -53 8161 -51
rect 8127 -119 8161 -91
rect 8127 -125 8161 -119
rect 8127 -187 8161 -163
rect 8127 -197 8161 -187
rect 8127 -255 8161 -235
rect 8127 -269 8161 -255
rect -7832 -381 -7822 -347
rect -7822 -381 -7798 -347
rect -7760 -381 -7754 -347
rect -7754 -381 -7726 -347
rect -7688 -381 -7686 -347
rect -7686 -381 -7654 -347
rect -7616 -381 -7584 -347
rect -7584 -381 -7582 -347
rect -7544 -381 -7516 -347
rect -7516 -381 -7510 -347
rect -7472 -381 -7448 -347
rect -7448 -381 -7438 -347
rect -6814 -381 -6804 -347
rect -6804 -381 -6780 -347
rect -6742 -381 -6736 -347
rect -6736 -381 -6708 -347
rect -6670 -381 -6668 -347
rect -6668 -381 -6636 -347
rect -6598 -381 -6566 -347
rect -6566 -381 -6564 -347
rect -6526 -381 -6498 -347
rect -6498 -381 -6492 -347
rect -6454 -381 -6430 -347
rect -6430 -381 -6420 -347
rect -5796 -381 -5786 -347
rect -5786 -381 -5762 -347
rect -5724 -381 -5718 -347
rect -5718 -381 -5690 -347
rect -5652 -381 -5650 -347
rect -5650 -381 -5618 -347
rect -5580 -381 -5548 -347
rect -5548 -381 -5546 -347
rect -5508 -381 -5480 -347
rect -5480 -381 -5474 -347
rect -5436 -381 -5412 -347
rect -5412 -381 -5402 -347
rect -4778 -381 -4768 -347
rect -4768 -381 -4744 -347
rect -4706 -381 -4700 -347
rect -4700 -381 -4672 -347
rect -4634 -381 -4632 -347
rect -4632 -381 -4600 -347
rect -4562 -381 -4530 -347
rect -4530 -381 -4528 -347
rect -4490 -381 -4462 -347
rect -4462 -381 -4456 -347
rect -4418 -381 -4394 -347
rect -4394 -381 -4384 -347
rect -3760 -381 -3750 -347
rect -3750 -381 -3726 -347
rect -3688 -381 -3682 -347
rect -3682 -381 -3654 -347
rect -3616 -381 -3614 -347
rect -3614 -381 -3582 -347
rect -3544 -381 -3512 -347
rect -3512 -381 -3510 -347
rect -3472 -381 -3444 -347
rect -3444 -381 -3438 -347
rect -3400 -381 -3376 -347
rect -3376 -381 -3366 -347
rect -2742 -381 -2732 -347
rect -2732 -381 -2708 -347
rect -2670 -381 -2664 -347
rect -2664 -381 -2636 -347
rect -2598 -381 -2596 -347
rect -2596 -381 -2564 -347
rect -2526 -381 -2494 -347
rect -2494 -381 -2492 -347
rect -2454 -381 -2426 -347
rect -2426 -381 -2420 -347
rect -2382 -381 -2358 -347
rect -2358 -381 -2348 -347
rect -1724 -381 -1714 -347
rect -1714 -381 -1690 -347
rect -1652 -381 -1646 -347
rect -1646 -381 -1618 -347
rect -1580 -381 -1578 -347
rect -1578 -381 -1546 -347
rect -1508 -381 -1476 -347
rect -1476 -381 -1474 -347
rect -1436 -381 -1408 -347
rect -1408 -381 -1402 -347
rect -1364 -381 -1340 -347
rect -1340 -381 -1330 -347
rect -706 -381 -696 -347
rect -696 -381 -672 -347
rect -634 -381 -628 -347
rect -628 -381 -600 -347
rect -562 -381 -560 -347
rect -560 -381 -528 -347
rect -490 -381 -458 -347
rect -458 -381 -456 -347
rect -418 -381 -390 -347
rect -390 -381 -384 -347
rect -346 -381 -322 -347
rect -322 -381 -312 -347
rect 312 -381 322 -347
rect 322 -381 346 -347
rect 384 -381 390 -347
rect 390 -381 418 -347
rect 456 -381 458 -347
rect 458 -381 490 -347
rect 528 -381 560 -347
rect 560 -381 562 -347
rect 600 -381 628 -347
rect 628 -381 634 -347
rect 672 -381 696 -347
rect 696 -381 706 -347
rect 1330 -381 1340 -347
rect 1340 -381 1364 -347
rect 1402 -381 1408 -347
rect 1408 -381 1436 -347
rect 1474 -381 1476 -347
rect 1476 -381 1508 -347
rect 1546 -381 1578 -347
rect 1578 -381 1580 -347
rect 1618 -381 1646 -347
rect 1646 -381 1652 -347
rect 1690 -381 1714 -347
rect 1714 -381 1724 -347
rect 2348 -381 2358 -347
rect 2358 -381 2382 -347
rect 2420 -381 2426 -347
rect 2426 -381 2454 -347
rect 2492 -381 2494 -347
rect 2494 -381 2526 -347
rect 2564 -381 2596 -347
rect 2596 -381 2598 -347
rect 2636 -381 2664 -347
rect 2664 -381 2670 -347
rect 2708 -381 2732 -347
rect 2732 -381 2742 -347
rect 3366 -381 3376 -347
rect 3376 -381 3400 -347
rect 3438 -381 3444 -347
rect 3444 -381 3472 -347
rect 3510 -381 3512 -347
rect 3512 -381 3544 -347
rect 3582 -381 3614 -347
rect 3614 -381 3616 -347
rect 3654 -381 3682 -347
rect 3682 -381 3688 -347
rect 3726 -381 3750 -347
rect 3750 -381 3760 -347
rect 4384 -381 4394 -347
rect 4394 -381 4418 -347
rect 4456 -381 4462 -347
rect 4462 -381 4490 -347
rect 4528 -381 4530 -347
rect 4530 -381 4562 -347
rect 4600 -381 4632 -347
rect 4632 -381 4634 -347
rect 4672 -381 4700 -347
rect 4700 -381 4706 -347
rect 4744 -381 4768 -347
rect 4768 -381 4778 -347
rect 5402 -381 5412 -347
rect 5412 -381 5436 -347
rect 5474 -381 5480 -347
rect 5480 -381 5508 -347
rect 5546 -381 5548 -347
rect 5548 -381 5580 -347
rect 5618 -381 5650 -347
rect 5650 -381 5652 -347
rect 5690 -381 5718 -347
rect 5718 -381 5724 -347
rect 5762 -381 5786 -347
rect 5786 -381 5796 -347
rect 6420 -381 6430 -347
rect 6430 -381 6454 -347
rect 6492 -381 6498 -347
rect 6498 -381 6526 -347
rect 6564 -381 6566 -347
rect 6566 -381 6598 -347
rect 6636 -381 6668 -347
rect 6668 -381 6670 -347
rect 6708 -381 6736 -347
rect 6736 -381 6742 -347
rect 6780 -381 6804 -347
rect 6804 -381 6814 -347
rect 7438 -381 7448 -347
rect 7448 -381 7472 -347
rect 7510 -381 7516 -347
rect 7516 -381 7544 -347
rect 7582 -381 7584 -347
rect 7584 -381 7616 -347
rect 7654 -381 7686 -347
rect 7686 -381 7688 -347
rect 7726 -381 7754 -347
rect 7754 -381 7760 -347
rect 7798 -381 7822 -347
rect 7822 -381 7832 -347
<< metal1 >>
rect -7879 381 -7391 387
rect -7879 347 -7832 381
rect -7798 347 -7760 381
rect -7726 347 -7688 381
rect -7654 347 -7616 381
rect -7582 347 -7544 381
rect -7510 347 -7472 381
rect -7438 347 -7391 381
rect -7879 341 -7391 347
rect -6861 381 -6373 387
rect -6861 347 -6814 381
rect -6780 347 -6742 381
rect -6708 347 -6670 381
rect -6636 347 -6598 381
rect -6564 347 -6526 381
rect -6492 347 -6454 381
rect -6420 347 -6373 381
rect -6861 341 -6373 347
rect -5843 381 -5355 387
rect -5843 347 -5796 381
rect -5762 347 -5724 381
rect -5690 347 -5652 381
rect -5618 347 -5580 381
rect -5546 347 -5508 381
rect -5474 347 -5436 381
rect -5402 347 -5355 381
rect -5843 341 -5355 347
rect -4825 381 -4337 387
rect -4825 347 -4778 381
rect -4744 347 -4706 381
rect -4672 347 -4634 381
rect -4600 347 -4562 381
rect -4528 347 -4490 381
rect -4456 347 -4418 381
rect -4384 347 -4337 381
rect -4825 341 -4337 347
rect -3807 381 -3319 387
rect -3807 347 -3760 381
rect -3726 347 -3688 381
rect -3654 347 -3616 381
rect -3582 347 -3544 381
rect -3510 347 -3472 381
rect -3438 347 -3400 381
rect -3366 347 -3319 381
rect -3807 341 -3319 347
rect -2789 381 -2301 387
rect -2789 347 -2742 381
rect -2708 347 -2670 381
rect -2636 347 -2598 381
rect -2564 347 -2526 381
rect -2492 347 -2454 381
rect -2420 347 -2382 381
rect -2348 347 -2301 381
rect -2789 341 -2301 347
rect -1771 381 -1283 387
rect -1771 347 -1724 381
rect -1690 347 -1652 381
rect -1618 347 -1580 381
rect -1546 347 -1508 381
rect -1474 347 -1436 381
rect -1402 347 -1364 381
rect -1330 347 -1283 381
rect -1771 341 -1283 347
rect -753 381 -265 387
rect -753 347 -706 381
rect -672 347 -634 381
rect -600 347 -562 381
rect -528 347 -490 381
rect -456 347 -418 381
rect -384 347 -346 381
rect -312 347 -265 381
rect -753 341 -265 347
rect 265 381 753 387
rect 265 347 312 381
rect 346 347 384 381
rect 418 347 456 381
rect 490 347 528 381
rect 562 347 600 381
rect 634 347 672 381
rect 706 347 753 381
rect 265 341 753 347
rect 1283 381 1771 387
rect 1283 347 1330 381
rect 1364 347 1402 381
rect 1436 347 1474 381
rect 1508 347 1546 381
rect 1580 347 1618 381
rect 1652 347 1690 381
rect 1724 347 1771 381
rect 1283 341 1771 347
rect 2301 381 2789 387
rect 2301 347 2348 381
rect 2382 347 2420 381
rect 2454 347 2492 381
rect 2526 347 2564 381
rect 2598 347 2636 381
rect 2670 347 2708 381
rect 2742 347 2789 381
rect 2301 341 2789 347
rect 3319 381 3807 387
rect 3319 347 3366 381
rect 3400 347 3438 381
rect 3472 347 3510 381
rect 3544 347 3582 381
rect 3616 347 3654 381
rect 3688 347 3726 381
rect 3760 347 3807 381
rect 3319 341 3807 347
rect 4337 381 4825 387
rect 4337 347 4384 381
rect 4418 347 4456 381
rect 4490 347 4528 381
rect 4562 347 4600 381
rect 4634 347 4672 381
rect 4706 347 4744 381
rect 4778 347 4825 381
rect 4337 341 4825 347
rect 5355 381 5843 387
rect 5355 347 5402 381
rect 5436 347 5474 381
rect 5508 347 5546 381
rect 5580 347 5618 381
rect 5652 347 5690 381
rect 5724 347 5762 381
rect 5796 347 5843 381
rect 5355 341 5843 347
rect 6373 381 6861 387
rect 6373 347 6420 381
rect 6454 347 6492 381
rect 6526 347 6564 381
rect 6598 347 6636 381
rect 6670 347 6708 381
rect 6742 347 6780 381
rect 6814 347 6861 381
rect 6373 341 6861 347
rect 7391 381 7879 387
rect 7391 347 7438 381
rect 7472 347 7510 381
rect 7544 347 7582 381
rect 7616 347 7654 381
rect 7688 347 7726 381
rect 7760 347 7798 381
rect 7832 347 7879 381
rect 7391 341 7879 347
rect -8167 269 -8121 300
rect -8167 235 -8161 269
rect -8127 235 -8121 269
rect -8167 197 -8121 235
rect -8167 163 -8161 197
rect -8127 163 -8121 197
rect -8167 125 -8121 163
rect -8167 91 -8161 125
rect -8127 91 -8121 125
rect -8167 53 -8121 91
rect -8167 19 -8161 53
rect -8127 19 -8121 53
rect -8167 -19 -8121 19
rect -8167 -53 -8161 -19
rect -8127 -53 -8121 -19
rect -8167 -91 -8121 -53
rect -8167 -125 -8161 -91
rect -8127 -125 -8121 -91
rect -8167 -163 -8121 -125
rect -8167 -197 -8161 -163
rect -8127 -197 -8121 -163
rect -8167 -235 -8121 -197
rect -8167 -269 -8161 -235
rect -8127 -269 -8121 -235
rect -8167 -300 -8121 -269
rect -7149 269 -7103 300
rect -7149 235 -7143 269
rect -7109 235 -7103 269
rect -7149 197 -7103 235
rect -7149 163 -7143 197
rect -7109 163 -7103 197
rect -7149 125 -7103 163
rect -7149 91 -7143 125
rect -7109 91 -7103 125
rect -7149 53 -7103 91
rect -7149 19 -7143 53
rect -7109 19 -7103 53
rect -7149 -19 -7103 19
rect -7149 -53 -7143 -19
rect -7109 -53 -7103 -19
rect -7149 -91 -7103 -53
rect -7149 -125 -7143 -91
rect -7109 -125 -7103 -91
rect -7149 -163 -7103 -125
rect -7149 -197 -7143 -163
rect -7109 -197 -7103 -163
rect -7149 -235 -7103 -197
rect -7149 -269 -7143 -235
rect -7109 -269 -7103 -235
rect -7149 -300 -7103 -269
rect -6131 269 -6085 300
rect -6131 235 -6125 269
rect -6091 235 -6085 269
rect -6131 197 -6085 235
rect -6131 163 -6125 197
rect -6091 163 -6085 197
rect -6131 125 -6085 163
rect -6131 91 -6125 125
rect -6091 91 -6085 125
rect -6131 53 -6085 91
rect -6131 19 -6125 53
rect -6091 19 -6085 53
rect -6131 -19 -6085 19
rect -6131 -53 -6125 -19
rect -6091 -53 -6085 -19
rect -6131 -91 -6085 -53
rect -6131 -125 -6125 -91
rect -6091 -125 -6085 -91
rect -6131 -163 -6085 -125
rect -6131 -197 -6125 -163
rect -6091 -197 -6085 -163
rect -6131 -235 -6085 -197
rect -6131 -269 -6125 -235
rect -6091 -269 -6085 -235
rect -6131 -300 -6085 -269
rect -5113 269 -5067 300
rect -5113 235 -5107 269
rect -5073 235 -5067 269
rect -5113 197 -5067 235
rect -5113 163 -5107 197
rect -5073 163 -5067 197
rect -5113 125 -5067 163
rect -5113 91 -5107 125
rect -5073 91 -5067 125
rect -5113 53 -5067 91
rect -5113 19 -5107 53
rect -5073 19 -5067 53
rect -5113 -19 -5067 19
rect -5113 -53 -5107 -19
rect -5073 -53 -5067 -19
rect -5113 -91 -5067 -53
rect -5113 -125 -5107 -91
rect -5073 -125 -5067 -91
rect -5113 -163 -5067 -125
rect -5113 -197 -5107 -163
rect -5073 -197 -5067 -163
rect -5113 -235 -5067 -197
rect -5113 -269 -5107 -235
rect -5073 -269 -5067 -235
rect -5113 -300 -5067 -269
rect -4095 269 -4049 300
rect -4095 235 -4089 269
rect -4055 235 -4049 269
rect -4095 197 -4049 235
rect -4095 163 -4089 197
rect -4055 163 -4049 197
rect -4095 125 -4049 163
rect -4095 91 -4089 125
rect -4055 91 -4049 125
rect -4095 53 -4049 91
rect -4095 19 -4089 53
rect -4055 19 -4049 53
rect -4095 -19 -4049 19
rect -4095 -53 -4089 -19
rect -4055 -53 -4049 -19
rect -4095 -91 -4049 -53
rect -4095 -125 -4089 -91
rect -4055 -125 -4049 -91
rect -4095 -163 -4049 -125
rect -4095 -197 -4089 -163
rect -4055 -197 -4049 -163
rect -4095 -235 -4049 -197
rect -4095 -269 -4089 -235
rect -4055 -269 -4049 -235
rect -4095 -300 -4049 -269
rect -3077 269 -3031 300
rect -3077 235 -3071 269
rect -3037 235 -3031 269
rect -3077 197 -3031 235
rect -3077 163 -3071 197
rect -3037 163 -3031 197
rect -3077 125 -3031 163
rect -3077 91 -3071 125
rect -3037 91 -3031 125
rect -3077 53 -3031 91
rect -3077 19 -3071 53
rect -3037 19 -3031 53
rect -3077 -19 -3031 19
rect -3077 -53 -3071 -19
rect -3037 -53 -3031 -19
rect -3077 -91 -3031 -53
rect -3077 -125 -3071 -91
rect -3037 -125 -3031 -91
rect -3077 -163 -3031 -125
rect -3077 -197 -3071 -163
rect -3037 -197 -3031 -163
rect -3077 -235 -3031 -197
rect -3077 -269 -3071 -235
rect -3037 -269 -3031 -235
rect -3077 -300 -3031 -269
rect -2059 269 -2013 300
rect -2059 235 -2053 269
rect -2019 235 -2013 269
rect -2059 197 -2013 235
rect -2059 163 -2053 197
rect -2019 163 -2013 197
rect -2059 125 -2013 163
rect -2059 91 -2053 125
rect -2019 91 -2013 125
rect -2059 53 -2013 91
rect -2059 19 -2053 53
rect -2019 19 -2013 53
rect -2059 -19 -2013 19
rect -2059 -53 -2053 -19
rect -2019 -53 -2013 -19
rect -2059 -91 -2013 -53
rect -2059 -125 -2053 -91
rect -2019 -125 -2013 -91
rect -2059 -163 -2013 -125
rect -2059 -197 -2053 -163
rect -2019 -197 -2013 -163
rect -2059 -235 -2013 -197
rect -2059 -269 -2053 -235
rect -2019 -269 -2013 -235
rect -2059 -300 -2013 -269
rect -1041 269 -995 300
rect -1041 235 -1035 269
rect -1001 235 -995 269
rect -1041 197 -995 235
rect -1041 163 -1035 197
rect -1001 163 -995 197
rect -1041 125 -995 163
rect -1041 91 -1035 125
rect -1001 91 -995 125
rect -1041 53 -995 91
rect -1041 19 -1035 53
rect -1001 19 -995 53
rect -1041 -19 -995 19
rect -1041 -53 -1035 -19
rect -1001 -53 -995 -19
rect -1041 -91 -995 -53
rect -1041 -125 -1035 -91
rect -1001 -125 -995 -91
rect -1041 -163 -995 -125
rect -1041 -197 -1035 -163
rect -1001 -197 -995 -163
rect -1041 -235 -995 -197
rect -1041 -269 -1035 -235
rect -1001 -269 -995 -235
rect -1041 -300 -995 -269
rect -23 269 23 300
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -300 23 -269
rect 995 269 1041 300
rect 995 235 1001 269
rect 1035 235 1041 269
rect 995 197 1041 235
rect 995 163 1001 197
rect 1035 163 1041 197
rect 995 125 1041 163
rect 995 91 1001 125
rect 1035 91 1041 125
rect 995 53 1041 91
rect 995 19 1001 53
rect 1035 19 1041 53
rect 995 -19 1041 19
rect 995 -53 1001 -19
rect 1035 -53 1041 -19
rect 995 -91 1041 -53
rect 995 -125 1001 -91
rect 1035 -125 1041 -91
rect 995 -163 1041 -125
rect 995 -197 1001 -163
rect 1035 -197 1041 -163
rect 995 -235 1041 -197
rect 995 -269 1001 -235
rect 1035 -269 1041 -235
rect 995 -300 1041 -269
rect 2013 269 2059 300
rect 2013 235 2019 269
rect 2053 235 2059 269
rect 2013 197 2059 235
rect 2013 163 2019 197
rect 2053 163 2059 197
rect 2013 125 2059 163
rect 2013 91 2019 125
rect 2053 91 2059 125
rect 2013 53 2059 91
rect 2013 19 2019 53
rect 2053 19 2059 53
rect 2013 -19 2059 19
rect 2013 -53 2019 -19
rect 2053 -53 2059 -19
rect 2013 -91 2059 -53
rect 2013 -125 2019 -91
rect 2053 -125 2059 -91
rect 2013 -163 2059 -125
rect 2013 -197 2019 -163
rect 2053 -197 2059 -163
rect 2013 -235 2059 -197
rect 2013 -269 2019 -235
rect 2053 -269 2059 -235
rect 2013 -300 2059 -269
rect 3031 269 3077 300
rect 3031 235 3037 269
rect 3071 235 3077 269
rect 3031 197 3077 235
rect 3031 163 3037 197
rect 3071 163 3077 197
rect 3031 125 3077 163
rect 3031 91 3037 125
rect 3071 91 3077 125
rect 3031 53 3077 91
rect 3031 19 3037 53
rect 3071 19 3077 53
rect 3031 -19 3077 19
rect 3031 -53 3037 -19
rect 3071 -53 3077 -19
rect 3031 -91 3077 -53
rect 3031 -125 3037 -91
rect 3071 -125 3077 -91
rect 3031 -163 3077 -125
rect 3031 -197 3037 -163
rect 3071 -197 3077 -163
rect 3031 -235 3077 -197
rect 3031 -269 3037 -235
rect 3071 -269 3077 -235
rect 3031 -300 3077 -269
rect 4049 269 4095 300
rect 4049 235 4055 269
rect 4089 235 4095 269
rect 4049 197 4095 235
rect 4049 163 4055 197
rect 4089 163 4095 197
rect 4049 125 4095 163
rect 4049 91 4055 125
rect 4089 91 4095 125
rect 4049 53 4095 91
rect 4049 19 4055 53
rect 4089 19 4095 53
rect 4049 -19 4095 19
rect 4049 -53 4055 -19
rect 4089 -53 4095 -19
rect 4049 -91 4095 -53
rect 4049 -125 4055 -91
rect 4089 -125 4095 -91
rect 4049 -163 4095 -125
rect 4049 -197 4055 -163
rect 4089 -197 4095 -163
rect 4049 -235 4095 -197
rect 4049 -269 4055 -235
rect 4089 -269 4095 -235
rect 4049 -300 4095 -269
rect 5067 269 5113 300
rect 5067 235 5073 269
rect 5107 235 5113 269
rect 5067 197 5113 235
rect 5067 163 5073 197
rect 5107 163 5113 197
rect 5067 125 5113 163
rect 5067 91 5073 125
rect 5107 91 5113 125
rect 5067 53 5113 91
rect 5067 19 5073 53
rect 5107 19 5113 53
rect 5067 -19 5113 19
rect 5067 -53 5073 -19
rect 5107 -53 5113 -19
rect 5067 -91 5113 -53
rect 5067 -125 5073 -91
rect 5107 -125 5113 -91
rect 5067 -163 5113 -125
rect 5067 -197 5073 -163
rect 5107 -197 5113 -163
rect 5067 -235 5113 -197
rect 5067 -269 5073 -235
rect 5107 -269 5113 -235
rect 5067 -300 5113 -269
rect 6085 269 6131 300
rect 6085 235 6091 269
rect 6125 235 6131 269
rect 6085 197 6131 235
rect 6085 163 6091 197
rect 6125 163 6131 197
rect 6085 125 6131 163
rect 6085 91 6091 125
rect 6125 91 6131 125
rect 6085 53 6131 91
rect 6085 19 6091 53
rect 6125 19 6131 53
rect 6085 -19 6131 19
rect 6085 -53 6091 -19
rect 6125 -53 6131 -19
rect 6085 -91 6131 -53
rect 6085 -125 6091 -91
rect 6125 -125 6131 -91
rect 6085 -163 6131 -125
rect 6085 -197 6091 -163
rect 6125 -197 6131 -163
rect 6085 -235 6131 -197
rect 6085 -269 6091 -235
rect 6125 -269 6131 -235
rect 6085 -300 6131 -269
rect 7103 269 7149 300
rect 7103 235 7109 269
rect 7143 235 7149 269
rect 7103 197 7149 235
rect 7103 163 7109 197
rect 7143 163 7149 197
rect 7103 125 7149 163
rect 7103 91 7109 125
rect 7143 91 7149 125
rect 7103 53 7149 91
rect 7103 19 7109 53
rect 7143 19 7149 53
rect 7103 -19 7149 19
rect 7103 -53 7109 -19
rect 7143 -53 7149 -19
rect 7103 -91 7149 -53
rect 7103 -125 7109 -91
rect 7143 -125 7149 -91
rect 7103 -163 7149 -125
rect 7103 -197 7109 -163
rect 7143 -197 7149 -163
rect 7103 -235 7149 -197
rect 7103 -269 7109 -235
rect 7143 -269 7149 -235
rect 7103 -300 7149 -269
rect 8121 269 8167 300
rect 8121 235 8127 269
rect 8161 235 8167 269
rect 8121 197 8167 235
rect 8121 163 8127 197
rect 8161 163 8167 197
rect 8121 125 8167 163
rect 8121 91 8127 125
rect 8161 91 8167 125
rect 8121 53 8167 91
rect 8121 19 8127 53
rect 8161 19 8167 53
rect 8121 -19 8167 19
rect 8121 -53 8127 -19
rect 8161 -53 8167 -19
rect 8121 -91 8167 -53
rect 8121 -125 8127 -91
rect 8161 -125 8167 -91
rect 8121 -163 8167 -125
rect 8121 -197 8127 -163
rect 8161 -197 8167 -163
rect 8121 -235 8167 -197
rect 8121 -269 8127 -235
rect 8161 -269 8167 -235
rect 8121 -300 8167 -269
rect -7879 -347 -7391 -341
rect -7879 -381 -7832 -347
rect -7798 -381 -7760 -347
rect -7726 -381 -7688 -347
rect -7654 -381 -7616 -347
rect -7582 -381 -7544 -347
rect -7510 -381 -7472 -347
rect -7438 -381 -7391 -347
rect -7879 -387 -7391 -381
rect -6861 -347 -6373 -341
rect -6861 -381 -6814 -347
rect -6780 -381 -6742 -347
rect -6708 -381 -6670 -347
rect -6636 -381 -6598 -347
rect -6564 -381 -6526 -347
rect -6492 -381 -6454 -347
rect -6420 -381 -6373 -347
rect -6861 -387 -6373 -381
rect -5843 -347 -5355 -341
rect -5843 -381 -5796 -347
rect -5762 -381 -5724 -347
rect -5690 -381 -5652 -347
rect -5618 -381 -5580 -347
rect -5546 -381 -5508 -347
rect -5474 -381 -5436 -347
rect -5402 -381 -5355 -347
rect -5843 -387 -5355 -381
rect -4825 -347 -4337 -341
rect -4825 -381 -4778 -347
rect -4744 -381 -4706 -347
rect -4672 -381 -4634 -347
rect -4600 -381 -4562 -347
rect -4528 -381 -4490 -347
rect -4456 -381 -4418 -347
rect -4384 -381 -4337 -347
rect -4825 -387 -4337 -381
rect -3807 -347 -3319 -341
rect -3807 -381 -3760 -347
rect -3726 -381 -3688 -347
rect -3654 -381 -3616 -347
rect -3582 -381 -3544 -347
rect -3510 -381 -3472 -347
rect -3438 -381 -3400 -347
rect -3366 -381 -3319 -347
rect -3807 -387 -3319 -381
rect -2789 -347 -2301 -341
rect -2789 -381 -2742 -347
rect -2708 -381 -2670 -347
rect -2636 -381 -2598 -347
rect -2564 -381 -2526 -347
rect -2492 -381 -2454 -347
rect -2420 -381 -2382 -347
rect -2348 -381 -2301 -347
rect -2789 -387 -2301 -381
rect -1771 -347 -1283 -341
rect -1771 -381 -1724 -347
rect -1690 -381 -1652 -347
rect -1618 -381 -1580 -347
rect -1546 -381 -1508 -347
rect -1474 -381 -1436 -347
rect -1402 -381 -1364 -347
rect -1330 -381 -1283 -347
rect -1771 -387 -1283 -381
rect -753 -347 -265 -341
rect -753 -381 -706 -347
rect -672 -381 -634 -347
rect -600 -381 -562 -347
rect -528 -381 -490 -347
rect -456 -381 -418 -347
rect -384 -381 -346 -347
rect -312 -381 -265 -347
rect -753 -387 -265 -381
rect 265 -347 753 -341
rect 265 -381 312 -347
rect 346 -381 384 -347
rect 418 -381 456 -347
rect 490 -381 528 -347
rect 562 -381 600 -347
rect 634 -381 672 -347
rect 706 -381 753 -347
rect 265 -387 753 -381
rect 1283 -347 1771 -341
rect 1283 -381 1330 -347
rect 1364 -381 1402 -347
rect 1436 -381 1474 -347
rect 1508 -381 1546 -347
rect 1580 -381 1618 -347
rect 1652 -381 1690 -347
rect 1724 -381 1771 -347
rect 1283 -387 1771 -381
rect 2301 -347 2789 -341
rect 2301 -381 2348 -347
rect 2382 -381 2420 -347
rect 2454 -381 2492 -347
rect 2526 -381 2564 -347
rect 2598 -381 2636 -347
rect 2670 -381 2708 -347
rect 2742 -381 2789 -347
rect 2301 -387 2789 -381
rect 3319 -347 3807 -341
rect 3319 -381 3366 -347
rect 3400 -381 3438 -347
rect 3472 -381 3510 -347
rect 3544 -381 3582 -347
rect 3616 -381 3654 -347
rect 3688 -381 3726 -347
rect 3760 -381 3807 -347
rect 3319 -387 3807 -381
rect 4337 -347 4825 -341
rect 4337 -381 4384 -347
rect 4418 -381 4456 -347
rect 4490 -381 4528 -347
rect 4562 -381 4600 -347
rect 4634 -381 4672 -347
rect 4706 -381 4744 -347
rect 4778 -381 4825 -347
rect 4337 -387 4825 -381
rect 5355 -347 5843 -341
rect 5355 -381 5402 -347
rect 5436 -381 5474 -347
rect 5508 -381 5546 -347
rect 5580 -381 5618 -347
rect 5652 -381 5690 -347
rect 5724 -381 5762 -347
rect 5796 -381 5843 -347
rect 5355 -387 5843 -381
rect 6373 -347 6861 -341
rect 6373 -381 6420 -347
rect 6454 -381 6492 -347
rect 6526 -381 6564 -347
rect 6598 -381 6636 -347
rect 6670 -381 6708 -347
rect 6742 -381 6780 -347
rect 6814 -381 6861 -347
rect 6373 -387 6861 -381
rect 7391 -347 7879 -341
rect 7391 -381 7438 -347
rect 7472 -381 7510 -347
rect 7544 -381 7582 -347
rect 7616 -381 7654 -347
rect 7688 -381 7726 -347
rect 7760 -381 7798 -347
rect 7832 -381 7879 -347
rect 7391 -387 7879 -381
<< end >>
