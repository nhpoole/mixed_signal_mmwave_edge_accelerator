magic
tech sky130A
timestamp 1626065694
<< checkpaint >>
rect -630 -630 662 656
<< metal1 >>
rect 0 0 3 26
rect 29 0 32 26
<< via1 >>
rect 3 0 29 26
<< metal2 >>
rect 0 0 3 26
rect 29 0 32 26
<< properties >>
string FIXED_BBOX 0 0 32 26
<< end >>
