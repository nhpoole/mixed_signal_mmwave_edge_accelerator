magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< error_p >>
rect -2319 -100 -2261 100
rect -1861 -100 -1803 100
rect -1403 -100 -1345 100
rect -945 -100 -887 100
rect -487 -100 -429 100
rect -29 -100 29 100
rect 429 -100 487 100
rect 887 -100 945 100
rect 1345 -100 1403 100
rect 1803 -100 1861 100
rect 2261 -100 2319 100
<< nmos >>
rect -2261 -100 -1861 100
rect -1803 -100 -1403 100
rect -1345 -100 -945 100
rect -887 -100 -487 100
rect -429 -100 -29 100
rect 29 -100 429 100
rect 487 -100 887 100
rect 945 -100 1345 100
rect 1403 -100 1803 100
rect 1861 -100 2261 100
<< ndiff >>
rect -2319 88 -2261 100
rect -2319 -88 -2307 88
rect -2273 -88 -2261 88
rect -2319 -100 -2261 -88
rect -1861 88 -1803 100
rect -1861 -88 -1849 88
rect -1815 -88 -1803 88
rect -1861 -100 -1803 -88
rect -1403 88 -1345 100
rect -1403 -88 -1391 88
rect -1357 -88 -1345 88
rect -1403 -100 -1345 -88
rect -945 88 -887 100
rect -945 -88 -933 88
rect -899 -88 -887 88
rect -945 -100 -887 -88
rect -487 88 -429 100
rect -487 -88 -475 88
rect -441 -88 -429 88
rect -487 -100 -429 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 429 88 487 100
rect 429 -88 441 88
rect 475 -88 487 88
rect 429 -100 487 -88
rect 887 88 945 100
rect 887 -88 899 88
rect 933 -88 945 88
rect 887 -100 945 -88
rect 1345 88 1403 100
rect 1345 -88 1357 88
rect 1391 -88 1403 88
rect 1345 -100 1403 -88
rect 1803 88 1861 100
rect 1803 -88 1815 88
rect 1849 -88 1861 88
rect 1803 -100 1861 -88
rect 2261 88 2319 100
rect 2261 -88 2273 88
rect 2307 -88 2319 88
rect 2261 -100 2319 -88
<< ndiffc >>
rect -2307 -88 -2273 88
rect -1849 -88 -1815 88
rect -1391 -88 -1357 88
rect -933 -88 -899 88
rect -475 -88 -441 88
rect -17 -88 17 88
rect 441 -88 475 88
rect 899 -88 933 88
rect 1357 -88 1391 88
rect 1815 -88 1849 88
rect 2273 -88 2307 88
<< poly >>
rect -2187 172 -1935 188
rect -2187 155 -2171 172
rect -2261 138 -2171 155
rect -1951 155 -1935 172
rect -1729 172 -1477 188
rect -1729 155 -1713 172
rect -1951 138 -1861 155
rect -2261 100 -1861 138
rect -1803 138 -1713 155
rect -1493 155 -1477 172
rect -1271 172 -1019 188
rect -1271 155 -1255 172
rect -1493 138 -1403 155
rect -1803 100 -1403 138
rect -1345 138 -1255 155
rect -1035 155 -1019 172
rect -813 172 -561 188
rect -813 155 -797 172
rect -1035 138 -945 155
rect -1345 100 -945 138
rect -887 138 -797 155
rect -577 155 -561 172
rect -355 172 -103 188
rect -355 155 -339 172
rect -577 138 -487 155
rect -887 100 -487 138
rect -429 138 -339 155
rect -119 155 -103 172
rect 103 172 355 188
rect 103 155 119 172
rect -119 138 -29 155
rect -429 100 -29 138
rect 29 138 119 155
rect 339 155 355 172
rect 561 172 813 188
rect 561 155 577 172
rect 339 138 429 155
rect 29 100 429 138
rect 487 138 577 155
rect 797 155 813 172
rect 1019 172 1271 188
rect 1019 155 1035 172
rect 797 138 887 155
rect 487 100 887 138
rect 945 138 1035 155
rect 1255 155 1271 172
rect 1477 172 1729 188
rect 1477 155 1493 172
rect 1255 138 1345 155
rect 945 100 1345 138
rect 1403 138 1493 155
rect 1713 155 1729 172
rect 1935 172 2187 188
rect 1935 155 1951 172
rect 1713 138 1803 155
rect 1403 100 1803 138
rect 1861 138 1951 155
rect 2171 155 2187 172
rect 2171 138 2261 155
rect 1861 100 2261 138
rect -2261 -138 -1861 -100
rect -2261 -155 -2171 -138
rect -2187 -172 -2171 -155
rect -1951 -155 -1861 -138
rect -1803 -138 -1403 -100
rect -1803 -155 -1713 -138
rect -1951 -172 -1935 -155
rect -2187 -188 -1935 -172
rect -1729 -172 -1713 -155
rect -1493 -155 -1403 -138
rect -1345 -138 -945 -100
rect -1345 -155 -1255 -138
rect -1493 -172 -1477 -155
rect -1729 -188 -1477 -172
rect -1271 -172 -1255 -155
rect -1035 -155 -945 -138
rect -887 -138 -487 -100
rect -887 -155 -797 -138
rect -1035 -172 -1019 -155
rect -1271 -188 -1019 -172
rect -813 -172 -797 -155
rect -577 -155 -487 -138
rect -429 -138 -29 -100
rect -429 -155 -339 -138
rect -577 -172 -561 -155
rect -813 -188 -561 -172
rect -355 -172 -339 -155
rect -119 -155 -29 -138
rect 29 -138 429 -100
rect 29 -155 119 -138
rect -119 -172 -103 -155
rect -355 -188 -103 -172
rect 103 -172 119 -155
rect 339 -155 429 -138
rect 487 -138 887 -100
rect 487 -155 577 -138
rect 339 -172 355 -155
rect 103 -188 355 -172
rect 561 -172 577 -155
rect 797 -155 887 -138
rect 945 -138 1345 -100
rect 945 -155 1035 -138
rect 797 -172 813 -155
rect 561 -188 813 -172
rect 1019 -172 1035 -155
rect 1255 -155 1345 -138
rect 1403 -138 1803 -100
rect 1403 -155 1493 -138
rect 1255 -172 1271 -155
rect 1019 -188 1271 -172
rect 1477 -172 1493 -155
rect 1713 -155 1803 -138
rect 1861 -138 2261 -100
rect 1861 -155 1951 -138
rect 1713 -172 1729 -155
rect 1477 -188 1729 -172
rect 1935 -172 1951 -155
rect 2171 -155 2261 -138
rect 2171 -172 2187 -155
rect 1935 -188 2187 -172
<< polycont >>
rect -2171 138 -1951 172
rect -1713 138 -1493 172
rect -1255 138 -1035 172
rect -797 138 -577 172
rect -339 138 -119 172
rect 119 138 339 172
rect 577 138 797 172
rect 1035 138 1255 172
rect 1493 138 1713 172
rect 1951 138 2171 172
rect -2171 -172 -1951 -138
rect -1713 -172 -1493 -138
rect -1255 -172 -1035 -138
rect -797 -172 -577 -138
rect -339 -172 -119 -138
rect 119 -172 339 -138
rect 577 -172 797 -138
rect 1035 -172 1255 -138
rect 1493 -172 1713 -138
rect 1951 -172 2171 -138
<< locali >>
rect -2187 138 -2171 172
rect -1951 138 -1935 172
rect -1729 138 -1713 172
rect -1493 138 -1477 172
rect -1271 138 -1255 172
rect -1035 138 -1019 172
rect -813 138 -797 172
rect -577 138 -561 172
rect -355 138 -339 172
rect -119 138 -103 172
rect 103 138 119 172
rect 339 138 355 172
rect 561 138 577 172
rect 797 138 813 172
rect 1019 138 1035 172
rect 1255 138 1271 172
rect 1477 138 1493 172
rect 1713 138 1729 172
rect 1935 138 1951 172
rect 2171 138 2187 172
rect -2307 88 -2273 104
rect -2307 -104 -2273 -88
rect -1849 88 -1815 104
rect -1849 -104 -1815 -88
rect -1391 88 -1357 104
rect -1391 -104 -1357 -88
rect -933 88 -899 104
rect -933 -104 -899 -88
rect -475 88 -441 104
rect -475 -104 -441 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 441 88 475 104
rect 441 -104 475 -88
rect 899 88 933 104
rect 899 -104 933 -88
rect 1357 88 1391 104
rect 1357 -104 1391 -88
rect 1815 88 1849 104
rect 1815 -104 1849 -88
rect 2273 88 2307 104
rect 2273 -104 2307 -88
rect -2187 -172 -2171 -138
rect -1951 -172 -1935 -138
rect -1729 -172 -1713 -138
rect -1493 -172 -1477 -138
rect -1271 -172 -1255 -138
rect -1035 -172 -1019 -138
rect -813 -172 -797 -138
rect -577 -172 -561 -138
rect -355 -172 -339 -138
rect -119 -172 -103 -138
rect 103 -172 119 -138
rect 339 -172 355 -138
rect 561 -172 577 -138
rect 797 -172 813 -138
rect 1019 -172 1035 -138
rect 1255 -172 1271 -138
rect 1477 -172 1493 -138
rect 1713 -172 1729 -138
rect 1935 -172 1951 -138
rect 2171 -172 2187 -138
<< viali >>
rect -2153 138 -1969 172
rect -1695 138 -1511 172
rect -1237 138 -1053 172
rect -779 138 -595 172
rect -321 138 -137 172
rect 137 138 321 172
rect 595 138 779 172
rect 1053 138 1237 172
rect 1511 138 1695 172
rect 1969 138 2153 172
rect -2307 -88 -2273 88
rect -1849 -88 -1815 88
rect -1391 -88 -1357 88
rect -933 -88 -899 88
rect -475 -88 -441 88
rect -17 -88 17 88
rect 441 -88 475 88
rect 899 -88 933 88
rect 1357 -88 1391 88
rect 1815 -88 1849 88
rect 2273 -88 2307 88
rect -2153 -172 -1969 -138
rect -1695 -172 -1511 -138
rect -1237 -172 -1053 -138
rect -779 -172 -595 -138
rect -321 -172 -137 -138
rect 137 -172 321 -138
rect 595 -172 779 -138
rect 1053 -172 1237 -138
rect 1511 -172 1695 -138
rect 1969 -172 2153 -138
<< metal1 >>
rect -2165 172 -1957 178
rect -2165 138 -2153 172
rect -1969 138 -1957 172
rect -2165 132 -1957 138
rect -1707 172 -1499 178
rect -1707 138 -1695 172
rect -1511 138 -1499 172
rect -1707 132 -1499 138
rect -1249 172 -1041 178
rect -1249 138 -1237 172
rect -1053 138 -1041 172
rect -1249 132 -1041 138
rect -791 172 -583 178
rect -791 138 -779 172
rect -595 138 -583 172
rect -791 132 -583 138
rect -333 172 -125 178
rect -333 138 -321 172
rect -137 138 -125 172
rect -333 132 -125 138
rect 125 172 333 178
rect 125 138 137 172
rect 321 138 333 172
rect 125 132 333 138
rect 583 172 791 178
rect 583 138 595 172
rect 779 138 791 172
rect 583 132 791 138
rect 1041 172 1249 178
rect 1041 138 1053 172
rect 1237 138 1249 172
rect 1041 132 1249 138
rect 1499 172 1707 178
rect 1499 138 1511 172
rect 1695 138 1707 172
rect 1499 132 1707 138
rect 1957 172 2165 178
rect 1957 138 1969 172
rect 2153 138 2165 172
rect 1957 132 2165 138
rect -2313 88 -2267 100
rect -2313 -88 -2307 88
rect -2273 -88 -2267 88
rect -2313 -100 -2267 -88
rect -1855 88 -1809 100
rect -1855 -88 -1849 88
rect -1815 -88 -1809 88
rect -1855 -100 -1809 -88
rect -1397 88 -1351 100
rect -1397 -88 -1391 88
rect -1357 -88 -1351 88
rect -1397 -100 -1351 -88
rect -939 88 -893 100
rect -939 -88 -933 88
rect -899 -88 -893 88
rect -939 -100 -893 -88
rect -481 88 -435 100
rect -481 -88 -475 88
rect -441 -88 -435 88
rect -481 -100 -435 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 435 88 481 100
rect 435 -88 441 88
rect 475 -88 481 88
rect 435 -100 481 -88
rect 893 88 939 100
rect 893 -88 899 88
rect 933 -88 939 88
rect 893 -100 939 -88
rect 1351 88 1397 100
rect 1351 -88 1357 88
rect 1391 -88 1397 88
rect 1351 -100 1397 -88
rect 1809 88 1855 100
rect 1809 -88 1815 88
rect 1849 -88 1855 88
rect 1809 -100 1855 -88
rect 2267 88 2313 100
rect 2267 -88 2273 88
rect 2307 -88 2313 88
rect 2267 -100 2313 -88
rect -2165 -138 -1957 -132
rect -2165 -172 -2153 -138
rect -1969 -172 -1957 -138
rect -2165 -178 -1957 -172
rect -1707 -138 -1499 -132
rect -1707 -172 -1695 -138
rect -1511 -172 -1499 -138
rect -1707 -178 -1499 -172
rect -1249 -138 -1041 -132
rect -1249 -172 -1237 -138
rect -1053 -172 -1041 -138
rect -1249 -178 -1041 -172
rect -791 -138 -583 -132
rect -791 -172 -779 -138
rect -595 -172 -583 -138
rect -791 -178 -583 -172
rect -333 -138 -125 -132
rect -333 -172 -321 -138
rect -137 -172 -125 -138
rect -333 -178 -125 -172
rect 125 -138 333 -132
rect 125 -172 137 -138
rect 321 -172 333 -138
rect 125 -178 333 -172
rect 583 -138 791 -132
rect 583 -172 595 -138
rect 779 -172 791 -138
rect 583 -178 791 -172
rect 1041 -138 1249 -132
rect 1041 -172 1053 -138
rect 1237 -172 1249 -138
rect 1041 -178 1249 -172
rect 1499 -138 1707 -132
rect 1499 -172 1511 -138
rect 1695 -172 1707 -138
rect 1499 -178 1707 -172
rect 1957 -138 2165 -132
rect 1957 -172 1969 -138
rect 2153 -172 2165 -138
rect 1957 -178 2165 -172
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 1 l 2 m 1 nf 10 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
