../results/deconv_kernel_estimator_top_level.lef