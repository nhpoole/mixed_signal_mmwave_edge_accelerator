magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -1814 -1679 1814 1679
<< nwell >>
rect -554 -419 554 419
<< pmoslvt >>
rect -358 -200 -158 200
rect -100 -200 100 200
rect 158 -200 358 200
<< pdiff >>
rect -416 187 -358 200
rect -416 153 -404 187
rect -370 153 -358 187
rect -416 119 -358 153
rect -416 85 -404 119
rect -370 85 -358 119
rect -416 51 -358 85
rect -416 17 -404 51
rect -370 17 -358 51
rect -416 -17 -358 17
rect -416 -51 -404 -17
rect -370 -51 -358 -17
rect -416 -85 -358 -51
rect -416 -119 -404 -85
rect -370 -119 -358 -85
rect -416 -153 -358 -119
rect -416 -187 -404 -153
rect -370 -187 -358 -153
rect -416 -200 -358 -187
rect -158 187 -100 200
rect -158 153 -146 187
rect -112 153 -100 187
rect -158 119 -100 153
rect -158 85 -146 119
rect -112 85 -100 119
rect -158 51 -100 85
rect -158 17 -146 51
rect -112 17 -100 51
rect -158 -17 -100 17
rect -158 -51 -146 -17
rect -112 -51 -100 -17
rect -158 -85 -100 -51
rect -158 -119 -146 -85
rect -112 -119 -100 -85
rect -158 -153 -100 -119
rect -158 -187 -146 -153
rect -112 -187 -100 -153
rect -158 -200 -100 -187
rect 100 187 158 200
rect 100 153 112 187
rect 146 153 158 187
rect 100 119 158 153
rect 100 85 112 119
rect 146 85 158 119
rect 100 51 158 85
rect 100 17 112 51
rect 146 17 158 51
rect 100 -17 158 17
rect 100 -51 112 -17
rect 146 -51 158 -17
rect 100 -85 158 -51
rect 100 -119 112 -85
rect 146 -119 158 -85
rect 100 -153 158 -119
rect 100 -187 112 -153
rect 146 -187 158 -153
rect 100 -200 158 -187
rect 358 187 416 200
rect 358 153 370 187
rect 404 153 416 187
rect 358 119 416 153
rect 358 85 370 119
rect 404 85 416 119
rect 358 51 416 85
rect 358 17 370 51
rect 404 17 416 51
rect 358 -17 416 17
rect 358 -51 370 -17
rect 404 -51 416 -17
rect 358 -85 416 -51
rect 358 -119 370 -85
rect 404 -119 416 -85
rect 358 -153 416 -119
rect 358 -187 370 -153
rect 404 -187 416 -153
rect 358 -200 416 -187
<< pdiffc >>
rect -404 153 -370 187
rect -404 85 -370 119
rect -404 17 -370 51
rect -404 -51 -370 -17
rect -404 -119 -370 -85
rect -404 -187 -370 -153
rect -146 153 -112 187
rect -146 85 -112 119
rect -146 17 -112 51
rect -146 -51 -112 -17
rect -146 -119 -112 -85
rect -146 -187 -112 -153
rect 112 153 146 187
rect 112 85 146 119
rect 112 17 146 51
rect 112 -51 146 -17
rect 112 -119 146 -85
rect 112 -187 146 -153
rect 370 153 404 187
rect 370 85 404 119
rect 370 17 404 51
rect 370 -51 404 -17
rect 370 -119 404 -85
rect 370 -187 404 -153
<< nsubdiff >>
rect -518 349 -391 383
rect -357 349 -323 383
rect -289 349 -255 383
rect -221 349 -187 383
rect -153 349 -119 383
rect -85 349 -51 383
rect -17 349 17 383
rect 51 349 85 383
rect 119 349 153 383
rect 187 349 221 383
rect 255 349 289 383
rect 323 349 357 383
rect 391 349 518 383
rect -518 255 -484 349
rect -518 187 -484 221
rect 484 255 518 349
rect -518 119 -484 153
rect -518 51 -484 85
rect -518 -17 -484 17
rect -518 -85 -484 -51
rect -518 -153 -484 -119
rect -518 -221 -484 -187
rect 484 187 518 221
rect 484 119 518 153
rect 484 51 518 85
rect 484 -17 518 17
rect 484 -85 518 -51
rect 484 -153 518 -119
rect -518 -349 -484 -255
rect 484 -221 518 -187
rect 484 -349 518 -255
rect -518 -383 -391 -349
rect -357 -383 -323 -349
rect -289 -383 -255 -349
rect -221 -383 -187 -349
rect -153 -383 -119 -349
rect -85 -383 -51 -349
rect -17 -383 17 -349
rect 51 -383 85 -349
rect 119 -383 153 -349
rect 187 -383 221 -349
rect 255 -383 289 -349
rect 323 -383 357 -349
rect 391 -383 518 -349
<< nsubdiffcont >>
rect -391 349 -357 383
rect -323 349 -289 383
rect -255 349 -221 383
rect -187 349 -153 383
rect -119 349 -85 383
rect -51 349 -17 383
rect 17 349 51 383
rect 85 349 119 383
rect 153 349 187 383
rect 221 349 255 383
rect 289 349 323 383
rect 357 349 391 383
rect -518 221 -484 255
rect 484 221 518 255
rect -518 153 -484 187
rect -518 85 -484 119
rect -518 17 -484 51
rect -518 -51 -484 -17
rect -518 -119 -484 -85
rect -518 -187 -484 -153
rect 484 153 518 187
rect 484 85 518 119
rect 484 17 518 51
rect 484 -51 518 -17
rect 484 -119 518 -85
rect 484 -187 518 -153
rect -518 -255 -484 -221
rect 484 -255 518 -221
rect -391 -383 -357 -349
rect -323 -383 -289 -349
rect -255 -383 -221 -349
rect -187 -383 -153 -349
rect -119 -383 -85 -349
rect -51 -383 -17 -349
rect 17 -383 51 -349
rect 85 -383 119 -349
rect 153 -383 187 -349
rect 221 -383 255 -349
rect 289 -383 323 -349
rect 357 -383 391 -349
<< poly >>
rect -324 281 -192 297
rect -324 264 -275 281
rect -358 247 -275 264
rect -241 264 -192 281
rect -66 281 66 297
rect -66 264 -17 281
rect -241 247 -158 264
rect -358 200 -158 247
rect -100 247 -17 264
rect 17 264 66 281
rect 192 281 324 297
rect 192 264 241 281
rect 17 247 100 264
rect -100 200 100 247
rect 158 247 241 264
rect 275 264 324 281
rect 275 247 358 264
rect 158 200 358 247
rect -358 -247 -158 -200
rect -358 -264 -275 -247
rect -324 -281 -275 -264
rect -241 -264 -158 -247
rect -100 -247 100 -200
rect -100 -264 -17 -247
rect -241 -281 -192 -264
rect -324 -297 -192 -281
rect -66 -281 -17 -264
rect 17 -264 100 -247
rect 158 -247 358 -200
rect 158 -264 241 -247
rect 17 -281 66 -264
rect -66 -297 66 -281
rect 192 -281 241 -264
rect 275 -264 358 -247
rect 275 -281 324 -264
rect 192 -297 324 -281
<< polycont >>
rect -275 247 -241 281
rect -17 247 17 281
rect 241 247 275 281
rect -275 -281 -241 -247
rect -17 -281 17 -247
rect 241 -281 275 -247
<< locali >>
rect -518 349 -391 383
rect -357 349 -323 383
rect -289 349 -255 383
rect -221 349 -187 383
rect -153 349 -119 383
rect -85 349 -51 383
rect -17 349 17 383
rect 51 349 85 383
rect 119 349 153 383
rect 187 349 221 383
rect 255 349 289 383
rect 323 349 357 383
rect 391 349 518 383
rect -518 255 -484 349
rect -324 247 -275 281
rect -241 247 -192 281
rect -66 247 -17 281
rect 17 247 66 281
rect 192 247 241 281
rect 275 247 324 281
rect 484 255 518 349
rect -518 187 -484 221
rect -518 119 -484 153
rect -518 51 -484 85
rect -518 -17 -484 17
rect -518 -85 -484 -51
rect -518 -153 -484 -119
rect -518 -221 -484 -187
rect -404 187 -370 204
rect -404 119 -370 127
rect -404 51 -370 55
rect -404 -55 -370 -51
rect -404 -127 -370 -119
rect -404 -204 -370 -187
rect -146 187 -112 204
rect -146 119 -112 127
rect -146 51 -112 55
rect -146 -55 -112 -51
rect -146 -127 -112 -119
rect -146 -204 -112 -187
rect 112 187 146 204
rect 112 119 146 127
rect 112 51 146 55
rect 112 -55 146 -51
rect 112 -127 146 -119
rect 112 -204 146 -187
rect 370 187 404 204
rect 370 119 404 127
rect 370 51 404 55
rect 370 -55 404 -51
rect 370 -127 404 -119
rect 370 -204 404 -187
rect 484 187 518 221
rect 484 119 518 153
rect 484 51 518 85
rect 484 -17 518 17
rect 484 -85 518 -51
rect 484 -153 518 -119
rect 484 -221 518 -187
rect -518 -349 -484 -255
rect -324 -281 -275 -247
rect -241 -281 -192 -247
rect -66 -281 -17 -247
rect 17 -281 66 -247
rect 192 -281 241 -247
rect 275 -281 324 -247
rect 484 -349 518 -255
rect -518 -383 -391 -349
rect -357 -383 -323 -349
rect -289 -383 -255 -349
rect -221 -383 -187 -349
rect -153 -383 -119 -349
rect -85 -383 -51 -349
rect -17 -383 17 -349
rect 51 -383 85 -349
rect 119 -383 153 -349
rect 187 -383 221 -349
rect 255 -383 289 -349
rect 323 -383 357 -349
rect 391 -383 518 -349
<< viali >>
rect -275 247 -241 281
rect -17 247 17 281
rect 241 247 275 281
rect -404 153 -370 161
rect -404 127 -370 153
rect -404 85 -370 89
rect -404 55 -370 85
rect -404 -17 -370 17
rect -404 -85 -370 -55
rect -404 -89 -370 -85
rect -404 -153 -370 -127
rect -404 -161 -370 -153
rect -146 153 -112 161
rect -146 127 -112 153
rect -146 85 -112 89
rect -146 55 -112 85
rect -146 -17 -112 17
rect -146 -85 -112 -55
rect -146 -89 -112 -85
rect -146 -153 -112 -127
rect -146 -161 -112 -153
rect 112 153 146 161
rect 112 127 146 153
rect 112 85 146 89
rect 112 55 146 85
rect 112 -17 146 17
rect 112 -85 146 -55
rect 112 -89 146 -85
rect 112 -153 146 -127
rect 112 -161 146 -153
rect 370 153 404 161
rect 370 127 404 153
rect 370 85 404 89
rect 370 55 404 85
rect 370 -17 404 17
rect 370 -85 404 -55
rect 370 -89 404 -85
rect 370 -153 404 -127
rect 370 -161 404 -153
rect -275 -281 -241 -247
rect -17 -281 17 -247
rect 241 -281 275 -247
<< metal1 >>
rect -312 281 -204 287
rect -312 247 -275 281
rect -241 247 -204 281
rect -312 241 -204 247
rect -54 281 54 287
rect -54 247 -17 281
rect 17 247 54 281
rect -54 241 54 247
rect 204 281 312 287
rect 204 247 241 281
rect 275 247 312 281
rect 204 241 312 247
rect -410 161 -364 200
rect -410 127 -404 161
rect -370 127 -364 161
rect -410 89 -364 127
rect -410 55 -404 89
rect -370 55 -364 89
rect -410 17 -364 55
rect -410 -17 -404 17
rect -370 -17 -364 17
rect -410 -55 -364 -17
rect -410 -89 -404 -55
rect -370 -89 -364 -55
rect -410 -127 -364 -89
rect -410 -161 -404 -127
rect -370 -161 -364 -127
rect -410 -200 -364 -161
rect -152 161 -106 200
rect -152 127 -146 161
rect -112 127 -106 161
rect -152 89 -106 127
rect -152 55 -146 89
rect -112 55 -106 89
rect -152 17 -106 55
rect -152 -17 -146 17
rect -112 -17 -106 17
rect -152 -55 -106 -17
rect -152 -89 -146 -55
rect -112 -89 -106 -55
rect -152 -127 -106 -89
rect -152 -161 -146 -127
rect -112 -161 -106 -127
rect -152 -200 -106 -161
rect 106 161 152 200
rect 106 127 112 161
rect 146 127 152 161
rect 106 89 152 127
rect 106 55 112 89
rect 146 55 152 89
rect 106 17 152 55
rect 106 -17 112 17
rect 146 -17 152 17
rect 106 -55 152 -17
rect 106 -89 112 -55
rect 146 -89 152 -55
rect 106 -127 152 -89
rect 106 -161 112 -127
rect 146 -161 152 -127
rect 106 -200 152 -161
rect 364 161 410 200
rect 364 127 370 161
rect 404 127 410 161
rect 364 89 410 127
rect 364 55 370 89
rect 404 55 410 89
rect 364 17 410 55
rect 364 -17 370 17
rect 404 -17 410 17
rect 364 -55 410 -17
rect 364 -89 370 -55
rect 404 -89 410 -55
rect 364 -127 410 -89
rect 364 -161 370 -127
rect 404 -161 410 -127
rect 364 -200 410 -161
rect -312 -247 -204 -241
rect -312 -281 -275 -247
rect -241 -281 -204 -247
rect -312 -287 -204 -281
rect -54 -247 54 -241
rect -54 -281 -17 -247
rect 17 -281 54 -247
rect -54 -287 54 -281
rect 204 -247 312 -241
rect 204 -281 241 -247
rect 275 -281 312 -247
rect 204 -287 312 -281
<< properties >>
string FIXED_BBOX -501 -366 501 366
<< end >>
