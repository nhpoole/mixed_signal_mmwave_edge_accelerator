../../6-testbench/outputs/testbench.sv