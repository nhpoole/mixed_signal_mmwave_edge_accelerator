magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -16428 -28508 26260 5660
<< nwell >>
rect 342 -10384 24858 4358
<< pwell >>
rect -12348 -11304 24948 -11152
rect -12348 -27096 -12196 -11304
rect -9222 -18864 50 -12486
rect 2544 -14858 23014 -14206
rect 2544 -16090 23014 -15438
rect 2542 -17324 23012 -16672
rect 2542 -18558 23012 -17906
rect 2542 -19790 23012 -19138
rect 2542 -21024 23012 -20372
rect 2542 -22258 23012 -21606
rect 2542 -23490 23012 -22838
rect 2542 -24724 23012 -24072
rect 24796 -27096 24948 -11304
rect -12348 -27248 24948 -27096
<< nmos >>
rect 2628 -14832 3588 -14232
rect 3646 -14832 4606 -14232
rect 4664 -14832 5624 -14232
rect 5682 -14832 6642 -14232
rect 6700 -14832 7660 -14232
rect 7718 -14832 8678 -14232
rect 8736 -14832 9696 -14232
rect 9754 -14832 10714 -14232
rect 10772 -14832 11732 -14232
rect 11790 -14832 12750 -14232
rect 12808 -14832 13768 -14232
rect 13826 -14832 14786 -14232
rect 14844 -14832 15804 -14232
rect 15862 -14832 16822 -14232
rect 16880 -14832 17840 -14232
rect 17898 -14832 18858 -14232
rect 18916 -14832 19876 -14232
rect 19934 -14832 20894 -14232
rect 20952 -14832 21912 -14232
rect 21970 -14832 22930 -14232
rect 2628 -16064 3588 -15464
rect 3646 -16064 4606 -15464
rect 4664 -16064 5624 -15464
rect 5682 -16064 6642 -15464
rect 6700 -16064 7660 -15464
rect 7718 -16064 8678 -15464
rect 8736 -16064 9696 -15464
rect 9754 -16064 10714 -15464
rect 10772 -16064 11732 -15464
rect 11790 -16064 12750 -15464
rect 12808 -16064 13768 -15464
rect 13826 -16064 14786 -15464
rect 14844 -16064 15804 -15464
rect 15862 -16064 16822 -15464
rect 16880 -16064 17840 -15464
rect 17898 -16064 18858 -15464
rect 18916 -16064 19876 -15464
rect 19934 -16064 20894 -15464
rect 20952 -16064 21912 -15464
rect 21970 -16064 22930 -15464
rect 2626 -17298 3586 -16698
rect 3644 -17298 4604 -16698
rect 4662 -17298 5622 -16698
rect 5680 -17298 6640 -16698
rect 6698 -17298 7658 -16698
rect 7716 -17298 8676 -16698
rect 8734 -17298 9694 -16698
rect 9752 -17298 10712 -16698
rect 10770 -17298 11730 -16698
rect 11788 -17298 12748 -16698
rect 12806 -17298 13766 -16698
rect 13824 -17298 14784 -16698
rect 14842 -17298 15802 -16698
rect 15860 -17298 16820 -16698
rect 16878 -17298 17838 -16698
rect 17896 -17298 18856 -16698
rect 18914 -17298 19874 -16698
rect 19932 -17298 20892 -16698
rect 20950 -17298 21910 -16698
rect 21968 -17298 22928 -16698
rect 2626 -18532 3586 -17932
rect 3644 -18532 4604 -17932
rect 4662 -18532 5622 -17932
rect 5680 -18532 6640 -17932
rect 6698 -18532 7658 -17932
rect 7716 -18532 8676 -17932
rect 8734 -18532 9694 -17932
rect 9752 -18532 10712 -17932
rect 10770 -18532 11730 -17932
rect 11788 -18532 12748 -17932
rect 12806 -18532 13766 -17932
rect 13824 -18532 14784 -17932
rect 14842 -18532 15802 -17932
rect 15860 -18532 16820 -17932
rect 16878 -18532 17838 -17932
rect 17896 -18532 18856 -17932
rect 18914 -18532 19874 -17932
rect 19932 -18532 20892 -17932
rect 20950 -18532 21910 -17932
rect 21968 -18532 22928 -17932
rect 2626 -19764 3586 -19164
rect 3644 -19764 4604 -19164
rect 4662 -19764 5622 -19164
rect 5680 -19764 6640 -19164
rect 6698 -19764 7658 -19164
rect 7716 -19764 8676 -19164
rect 8734 -19764 9694 -19164
rect 9752 -19764 10712 -19164
rect 10770 -19764 11730 -19164
rect 11788 -19764 12748 -19164
rect 12806 -19764 13766 -19164
rect 13824 -19764 14784 -19164
rect 14842 -19764 15802 -19164
rect 15860 -19764 16820 -19164
rect 16878 -19764 17838 -19164
rect 17896 -19764 18856 -19164
rect 18914 -19764 19874 -19164
rect 19932 -19764 20892 -19164
rect 20950 -19764 21910 -19164
rect 21968 -19764 22928 -19164
rect 2626 -20998 3586 -20398
rect 3644 -20998 4604 -20398
rect 4662 -20998 5622 -20398
rect 5680 -20998 6640 -20398
rect 6698 -20998 7658 -20398
rect 7716 -20998 8676 -20398
rect 8734 -20998 9694 -20398
rect 9752 -20998 10712 -20398
rect 10770 -20998 11730 -20398
rect 11788 -20998 12748 -20398
rect 12806 -20998 13766 -20398
rect 13824 -20998 14784 -20398
rect 14842 -20998 15802 -20398
rect 15860 -20998 16820 -20398
rect 16878 -20998 17838 -20398
rect 17896 -20998 18856 -20398
rect 18914 -20998 19874 -20398
rect 19932 -20998 20892 -20398
rect 20950 -20998 21910 -20398
rect 21968 -20998 22928 -20398
rect 2626 -22232 3586 -21632
rect 3644 -22232 4604 -21632
rect 4662 -22232 5622 -21632
rect 5680 -22232 6640 -21632
rect 6698 -22232 7658 -21632
rect 7716 -22232 8676 -21632
rect 8734 -22232 9694 -21632
rect 9752 -22232 10712 -21632
rect 10770 -22232 11730 -21632
rect 11788 -22232 12748 -21632
rect 12806 -22232 13766 -21632
rect 13824 -22232 14784 -21632
rect 14842 -22232 15802 -21632
rect 15860 -22232 16820 -21632
rect 16878 -22232 17838 -21632
rect 17896 -22232 18856 -21632
rect 18914 -22232 19874 -21632
rect 19932 -22232 20892 -21632
rect 20950 -22232 21910 -21632
rect 21968 -22232 22928 -21632
rect 2626 -23464 3586 -22864
rect 3644 -23464 4604 -22864
rect 4662 -23464 5622 -22864
rect 5680 -23464 6640 -22864
rect 6698 -23464 7658 -22864
rect 7716 -23464 8676 -22864
rect 8734 -23464 9694 -22864
rect 9752 -23464 10712 -22864
rect 10770 -23464 11730 -22864
rect 11788 -23464 12748 -22864
rect 12806 -23464 13766 -22864
rect 13824 -23464 14784 -22864
rect 14842 -23464 15802 -22864
rect 15860 -23464 16820 -22864
rect 16878 -23464 17838 -22864
rect 17896 -23464 18856 -22864
rect 18914 -23464 19874 -22864
rect 19932 -23464 20892 -22864
rect 20950 -23464 21910 -22864
rect 21968 -23464 22928 -22864
rect 2626 -24698 3586 -24098
rect 3644 -24698 4604 -24098
rect 4662 -24698 5622 -24098
rect 5680 -24698 6640 -24098
rect 6698 -24698 7658 -24098
rect 7716 -24698 8676 -24098
rect 8734 -24698 9694 -24098
rect 9752 -24698 10712 -24098
rect 10770 -24698 11730 -24098
rect 11788 -24698 12748 -24098
rect 12806 -24698 13766 -24098
rect 13824 -24698 14784 -24098
rect 14842 -24698 15802 -24098
rect 15860 -24698 16820 -24098
rect 16878 -24698 17838 -24098
rect 17896 -24698 18856 -24098
rect 18914 -24698 19874 -24098
rect 19932 -24698 20892 -24098
rect 20950 -24698 21910 -24098
rect 21968 -24698 22928 -24098
<< nmoslvt >>
rect -9138 -13112 -8178 -12512
rect -8120 -13112 -7160 -12512
rect -7102 -13112 -6142 -12512
rect -6084 -13112 -5124 -12512
rect -5066 -13112 -4106 -12512
rect -4048 -13112 -3088 -12512
rect -3030 -13112 -2070 -12512
rect -2012 -13112 -1052 -12512
rect -994 -13112 -34 -12512
rect -9138 -13930 -8178 -13330
rect -8120 -13930 -7160 -13330
rect -7102 -13930 -6142 -13330
rect -6084 -13930 -5124 -13330
rect -5066 -13930 -4106 -13330
rect -4048 -13930 -3088 -13330
rect -3030 -13930 -2070 -13330
rect -2012 -13930 -1052 -13330
rect -994 -13930 -34 -13330
rect -9138 -14748 -8178 -14148
rect -8120 -14748 -7160 -14148
rect -7102 -14748 -6142 -14148
rect -6084 -14748 -5124 -14148
rect -5066 -14748 -4106 -14148
rect -4048 -14748 -3088 -14148
rect -3030 -14748 -2070 -14148
rect -2012 -14748 -1052 -14148
rect -994 -14748 -34 -14148
rect -9138 -15566 -8178 -14966
rect -8120 -15566 -7160 -14966
rect -7102 -15566 -6142 -14966
rect -6084 -15566 -5124 -14966
rect -5066 -15566 -4106 -14966
rect -4048 -15566 -3088 -14966
rect -3030 -15566 -2070 -14966
rect -2012 -15566 -1052 -14966
rect -994 -15566 -34 -14966
rect -9138 -16384 -8178 -15784
rect -8120 -16384 -7160 -15784
rect -7102 -16384 -6142 -15784
rect -6084 -16384 -5124 -15784
rect -5066 -16384 -4106 -15784
rect -4048 -16384 -3088 -15784
rect -3030 -16384 -2070 -15784
rect -2012 -16384 -1052 -15784
rect -994 -16384 -34 -15784
rect -9138 -17202 -8178 -16602
rect -8120 -17202 -7160 -16602
rect -7102 -17202 -6142 -16602
rect -6084 -17202 -5124 -16602
rect -5066 -17202 -4106 -16602
rect -4048 -17202 -3088 -16602
rect -3030 -17202 -2070 -16602
rect -2012 -17202 -1052 -16602
rect -994 -17202 -34 -16602
rect -9138 -18020 -8178 -17420
rect -8120 -18020 -7160 -17420
rect -7102 -18020 -6142 -17420
rect -6084 -18020 -5124 -17420
rect -5066 -18020 -4106 -17420
rect -4048 -18020 -3088 -17420
rect -3030 -18020 -2070 -17420
rect -2012 -18020 -1052 -17420
rect -994 -18020 -34 -17420
rect -9138 -18838 -8178 -18238
rect -8120 -18838 -7160 -18238
rect -7102 -18838 -6142 -18238
rect -6084 -18838 -5124 -18238
rect -5066 -18838 -4106 -18238
rect -4048 -18838 -3088 -18238
rect -3030 -18838 -2070 -18238
rect -2012 -18838 -1052 -18238
rect -994 -18838 -34 -18238
<< ndiff >>
rect -9196 -12557 -9138 -12512
rect -9196 -12591 -9184 -12557
rect -9150 -12591 -9138 -12557
rect -9196 -12625 -9138 -12591
rect -9196 -12659 -9184 -12625
rect -9150 -12659 -9138 -12625
rect -9196 -12693 -9138 -12659
rect -9196 -12727 -9184 -12693
rect -9150 -12727 -9138 -12693
rect -9196 -12761 -9138 -12727
rect -9196 -12795 -9184 -12761
rect -9150 -12795 -9138 -12761
rect -9196 -12829 -9138 -12795
rect -9196 -12863 -9184 -12829
rect -9150 -12863 -9138 -12829
rect -9196 -12897 -9138 -12863
rect -9196 -12931 -9184 -12897
rect -9150 -12931 -9138 -12897
rect -9196 -12965 -9138 -12931
rect -9196 -12999 -9184 -12965
rect -9150 -12999 -9138 -12965
rect -9196 -13033 -9138 -12999
rect -9196 -13067 -9184 -13033
rect -9150 -13067 -9138 -13033
rect -9196 -13112 -9138 -13067
rect -8178 -12557 -8120 -12512
rect -8178 -12591 -8166 -12557
rect -8132 -12591 -8120 -12557
rect -8178 -12625 -8120 -12591
rect -8178 -12659 -8166 -12625
rect -8132 -12659 -8120 -12625
rect -8178 -12693 -8120 -12659
rect -8178 -12727 -8166 -12693
rect -8132 -12727 -8120 -12693
rect -8178 -12761 -8120 -12727
rect -8178 -12795 -8166 -12761
rect -8132 -12795 -8120 -12761
rect -8178 -12829 -8120 -12795
rect -8178 -12863 -8166 -12829
rect -8132 -12863 -8120 -12829
rect -8178 -12897 -8120 -12863
rect -8178 -12931 -8166 -12897
rect -8132 -12931 -8120 -12897
rect -8178 -12965 -8120 -12931
rect -8178 -12999 -8166 -12965
rect -8132 -12999 -8120 -12965
rect -8178 -13033 -8120 -12999
rect -8178 -13067 -8166 -13033
rect -8132 -13067 -8120 -13033
rect -8178 -13112 -8120 -13067
rect -7160 -12557 -7102 -12512
rect -7160 -12591 -7148 -12557
rect -7114 -12591 -7102 -12557
rect -7160 -12625 -7102 -12591
rect -7160 -12659 -7148 -12625
rect -7114 -12659 -7102 -12625
rect -7160 -12693 -7102 -12659
rect -7160 -12727 -7148 -12693
rect -7114 -12727 -7102 -12693
rect -7160 -12761 -7102 -12727
rect -7160 -12795 -7148 -12761
rect -7114 -12795 -7102 -12761
rect -7160 -12829 -7102 -12795
rect -7160 -12863 -7148 -12829
rect -7114 -12863 -7102 -12829
rect -7160 -12897 -7102 -12863
rect -7160 -12931 -7148 -12897
rect -7114 -12931 -7102 -12897
rect -7160 -12965 -7102 -12931
rect -7160 -12999 -7148 -12965
rect -7114 -12999 -7102 -12965
rect -7160 -13033 -7102 -12999
rect -7160 -13067 -7148 -13033
rect -7114 -13067 -7102 -13033
rect -7160 -13112 -7102 -13067
rect -6142 -12557 -6084 -12512
rect -6142 -12591 -6130 -12557
rect -6096 -12591 -6084 -12557
rect -6142 -12625 -6084 -12591
rect -6142 -12659 -6130 -12625
rect -6096 -12659 -6084 -12625
rect -6142 -12693 -6084 -12659
rect -6142 -12727 -6130 -12693
rect -6096 -12727 -6084 -12693
rect -6142 -12761 -6084 -12727
rect -6142 -12795 -6130 -12761
rect -6096 -12795 -6084 -12761
rect -6142 -12829 -6084 -12795
rect -6142 -12863 -6130 -12829
rect -6096 -12863 -6084 -12829
rect -6142 -12897 -6084 -12863
rect -6142 -12931 -6130 -12897
rect -6096 -12931 -6084 -12897
rect -6142 -12965 -6084 -12931
rect -6142 -12999 -6130 -12965
rect -6096 -12999 -6084 -12965
rect -6142 -13033 -6084 -12999
rect -6142 -13067 -6130 -13033
rect -6096 -13067 -6084 -13033
rect -6142 -13112 -6084 -13067
rect -5124 -12557 -5066 -12512
rect -5124 -12591 -5112 -12557
rect -5078 -12591 -5066 -12557
rect -5124 -12625 -5066 -12591
rect -5124 -12659 -5112 -12625
rect -5078 -12659 -5066 -12625
rect -5124 -12693 -5066 -12659
rect -5124 -12727 -5112 -12693
rect -5078 -12727 -5066 -12693
rect -5124 -12761 -5066 -12727
rect -5124 -12795 -5112 -12761
rect -5078 -12795 -5066 -12761
rect -5124 -12829 -5066 -12795
rect -5124 -12863 -5112 -12829
rect -5078 -12863 -5066 -12829
rect -5124 -12897 -5066 -12863
rect -5124 -12931 -5112 -12897
rect -5078 -12931 -5066 -12897
rect -5124 -12965 -5066 -12931
rect -5124 -12999 -5112 -12965
rect -5078 -12999 -5066 -12965
rect -5124 -13033 -5066 -12999
rect -5124 -13067 -5112 -13033
rect -5078 -13067 -5066 -13033
rect -5124 -13112 -5066 -13067
rect -4106 -12557 -4048 -12512
rect -4106 -12591 -4094 -12557
rect -4060 -12591 -4048 -12557
rect -4106 -12625 -4048 -12591
rect -4106 -12659 -4094 -12625
rect -4060 -12659 -4048 -12625
rect -4106 -12693 -4048 -12659
rect -4106 -12727 -4094 -12693
rect -4060 -12727 -4048 -12693
rect -4106 -12761 -4048 -12727
rect -4106 -12795 -4094 -12761
rect -4060 -12795 -4048 -12761
rect -4106 -12829 -4048 -12795
rect -4106 -12863 -4094 -12829
rect -4060 -12863 -4048 -12829
rect -4106 -12897 -4048 -12863
rect -4106 -12931 -4094 -12897
rect -4060 -12931 -4048 -12897
rect -4106 -12965 -4048 -12931
rect -4106 -12999 -4094 -12965
rect -4060 -12999 -4048 -12965
rect -4106 -13033 -4048 -12999
rect -4106 -13067 -4094 -13033
rect -4060 -13067 -4048 -13033
rect -4106 -13112 -4048 -13067
rect -3088 -12557 -3030 -12512
rect -3088 -12591 -3076 -12557
rect -3042 -12591 -3030 -12557
rect -3088 -12625 -3030 -12591
rect -3088 -12659 -3076 -12625
rect -3042 -12659 -3030 -12625
rect -3088 -12693 -3030 -12659
rect -3088 -12727 -3076 -12693
rect -3042 -12727 -3030 -12693
rect -3088 -12761 -3030 -12727
rect -3088 -12795 -3076 -12761
rect -3042 -12795 -3030 -12761
rect -3088 -12829 -3030 -12795
rect -3088 -12863 -3076 -12829
rect -3042 -12863 -3030 -12829
rect -3088 -12897 -3030 -12863
rect -3088 -12931 -3076 -12897
rect -3042 -12931 -3030 -12897
rect -3088 -12965 -3030 -12931
rect -3088 -12999 -3076 -12965
rect -3042 -12999 -3030 -12965
rect -3088 -13033 -3030 -12999
rect -3088 -13067 -3076 -13033
rect -3042 -13067 -3030 -13033
rect -3088 -13112 -3030 -13067
rect -2070 -12557 -2012 -12512
rect -2070 -12591 -2058 -12557
rect -2024 -12591 -2012 -12557
rect -2070 -12625 -2012 -12591
rect -2070 -12659 -2058 -12625
rect -2024 -12659 -2012 -12625
rect -2070 -12693 -2012 -12659
rect -2070 -12727 -2058 -12693
rect -2024 -12727 -2012 -12693
rect -2070 -12761 -2012 -12727
rect -2070 -12795 -2058 -12761
rect -2024 -12795 -2012 -12761
rect -2070 -12829 -2012 -12795
rect -2070 -12863 -2058 -12829
rect -2024 -12863 -2012 -12829
rect -2070 -12897 -2012 -12863
rect -2070 -12931 -2058 -12897
rect -2024 -12931 -2012 -12897
rect -2070 -12965 -2012 -12931
rect -2070 -12999 -2058 -12965
rect -2024 -12999 -2012 -12965
rect -2070 -13033 -2012 -12999
rect -2070 -13067 -2058 -13033
rect -2024 -13067 -2012 -13033
rect -2070 -13112 -2012 -13067
rect -1052 -12557 -994 -12512
rect -1052 -12591 -1040 -12557
rect -1006 -12591 -994 -12557
rect -1052 -12625 -994 -12591
rect -1052 -12659 -1040 -12625
rect -1006 -12659 -994 -12625
rect -1052 -12693 -994 -12659
rect -1052 -12727 -1040 -12693
rect -1006 -12727 -994 -12693
rect -1052 -12761 -994 -12727
rect -1052 -12795 -1040 -12761
rect -1006 -12795 -994 -12761
rect -1052 -12829 -994 -12795
rect -1052 -12863 -1040 -12829
rect -1006 -12863 -994 -12829
rect -1052 -12897 -994 -12863
rect -1052 -12931 -1040 -12897
rect -1006 -12931 -994 -12897
rect -1052 -12965 -994 -12931
rect -1052 -12999 -1040 -12965
rect -1006 -12999 -994 -12965
rect -1052 -13033 -994 -12999
rect -1052 -13067 -1040 -13033
rect -1006 -13067 -994 -13033
rect -1052 -13112 -994 -13067
rect -34 -12557 24 -12512
rect -34 -12591 -22 -12557
rect 12 -12591 24 -12557
rect -34 -12625 24 -12591
rect -34 -12659 -22 -12625
rect 12 -12659 24 -12625
rect -34 -12693 24 -12659
rect -34 -12727 -22 -12693
rect 12 -12727 24 -12693
rect -34 -12761 24 -12727
rect -34 -12795 -22 -12761
rect 12 -12795 24 -12761
rect -34 -12829 24 -12795
rect -34 -12863 -22 -12829
rect 12 -12863 24 -12829
rect -34 -12897 24 -12863
rect -34 -12931 -22 -12897
rect 12 -12931 24 -12897
rect -34 -12965 24 -12931
rect -34 -12999 -22 -12965
rect 12 -12999 24 -12965
rect -34 -13033 24 -12999
rect -34 -13067 -22 -13033
rect 12 -13067 24 -13033
rect -34 -13112 24 -13067
rect -9196 -13375 -9138 -13330
rect -9196 -13409 -9184 -13375
rect -9150 -13409 -9138 -13375
rect -9196 -13443 -9138 -13409
rect -9196 -13477 -9184 -13443
rect -9150 -13477 -9138 -13443
rect -9196 -13511 -9138 -13477
rect -9196 -13545 -9184 -13511
rect -9150 -13545 -9138 -13511
rect -9196 -13579 -9138 -13545
rect -9196 -13613 -9184 -13579
rect -9150 -13613 -9138 -13579
rect -9196 -13647 -9138 -13613
rect -9196 -13681 -9184 -13647
rect -9150 -13681 -9138 -13647
rect -9196 -13715 -9138 -13681
rect -9196 -13749 -9184 -13715
rect -9150 -13749 -9138 -13715
rect -9196 -13783 -9138 -13749
rect -9196 -13817 -9184 -13783
rect -9150 -13817 -9138 -13783
rect -9196 -13851 -9138 -13817
rect -9196 -13885 -9184 -13851
rect -9150 -13885 -9138 -13851
rect -9196 -13930 -9138 -13885
rect -8178 -13375 -8120 -13330
rect -8178 -13409 -8166 -13375
rect -8132 -13409 -8120 -13375
rect -8178 -13443 -8120 -13409
rect -8178 -13477 -8166 -13443
rect -8132 -13477 -8120 -13443
rect -8178 -13511 -8120 -13477
rect -8178 -13545 -8166 -13511
rect -8132 -13545 -8120 -13511
rect -8178 -13579 -8120 -13545
rect -8178 -13613 -8166 -13579
rect -8132 -13613 -8120 -13579
rect -8178 -13647 -8120 -13613
rect -8178 -13681 -8166 -13647
rect -8132 -13681 -8120 -13647
rect -8178 -13715 -8120 -13681
rect -8178 -13749 -8166 -13715
rect -8132 -13749 -8120 -13715
rect -8178 -13783 -8120 -13749
rect -8178 -13817 -8166 -13783
rect -8132 -13817 -8120 -13783
rect -8178 -13851 -8120 -13817
rect -8178 -13885 -8166 -13851
rect -8132 -13885 -8120 -13851
rect -8178 -13930 -8120 -13885
rect -7160 -13375 -7102 -13330
rect -7160 -13409 -7148 -13375
rect -7114 -13409 -7102 -13375
rect -7160 -13443 -7102 -13409
rect -7160 -13477 -7148 -13443
rect -7114 -13477 -7102 -13443
rect -7160 -13511 -7102 -13477
rect -7160 -13545 -7148 -13511
rect -7114 -13545 -7102 -13511
rect -7160 -13579 -7102 -13545
rect -7160 -13613 -7148 -13579
rect -7114 -13613 -7102 -13579
rect -7160 -13647 -7102 -13613
rect -7160 -13681 -7148 -13647
rect -7114 -13681 -7102 -13647
rect -7160 -13715 -7102 -13681
rect -7160 -13749 -7148 -13715
rect -7114 -13749 -7102 -13715
rect -7160 -13783 -7102 -13749
rect -7160 -13817 -7148 -13783
rect -7114 -13817 -7102 -13783
rect -7160 -13851 -7102 -13817
rect -7160 -13885 -7148 -13851
rect -7114 -13885 -7102 -13851
rect -7160 -13930 -7102 -13885
rect -6142 -13375 -6084 -13330
rect -6142 -13409 -6130 -13375
rect -6096 -13409 -6084 -13375
rect -6142 -13443 -6084 -13409
rect -6142 -13477 -6130 -13443
rect -6096 -13477 -6084 -13443
rect -6142 -13511 -6084 -13477
rect -6142 -13545 -6130 -13511
rect -6096 -13545 -6084 -13511
rect -6142 -13579 -6084 -13545
rect -6142 -13613 -6130 -13579
rect -6096 -13613 -6084 -13579
rect -6142 -13647 -6084 -13613
rect -6142 -13681 -6130 -13647
rect -6096 -13681 -6084 -13647
rect -6142 -13715 -6084 -13681
rect -6142 -13749 -6130 -13715
rect -6096 -13749 -6084 -13715
rect -6142 -13783 -6084 -13749
rect -6142 -13817 -6130 -13783
rect -6096 -13817 -6084 -13783
rect -6142 -13851 -6084 -13817
rect -6142 -13885 -6130 -13851
rect -6096 -13885 -6084 -13851
rect -6142 -13930 -6084 -13885
rect -5124 -13375 -5066 -13330
rect -5124 -13409 -5112 -13375
rect -5078 -13409 -5066 -13375
rect -5124 -13443 -5066 -13409
rect -5124 -13477 -5112 -13443
rect -5078 -13477 -5066 -13443
rect -5124 -13511 -5066 -13477
rect -5124 -13545 -5112 -13511
rect -5078 -13545 -5066 -13511
rect -5124 -13579 -5066 -13545
rect -5124 -13613 -5112 -13579
rect -5078 -13613 -5066 -13579
rect -5124 -13647 -5066 -13613
rect -5124 -13681 -5112 -13647
rect -5078 -13681 -5066 -13647
rect -5124 -13715 -5066 -13681
rect -5124 -13749 -5112 -13715
rect -5078 -13749 -5066 -13715
rect -5124 -13783 -5066 -13749
rect -5124 -13817 -5112 -13783
rect -5078 -13817 -5066 -13783
rect -5124 -13851 -5066 -13817
rect -5124 -13885 -5112 -13851
rect -5078 -13885 -5066 -13851
rect -5124 -13930 -5066 -13885
rect -4106 -13375 -4048 -13330
rect -4106 -13409 -4094 -13375
rect -4060 -13409 -4048 -13375
rect -4106 -13443 -4048 -13409
rect -4106 -13477 -4094 -13443
rect -4060 -13477 -4048 -13443
rect -4106 -13511 -4048 -13477
rect -4106 -13545 -4094 -13511
rect -4060 -13545 -4048 -13511
rect -4106 -13579 -4048 -13545
rect -4106 -13613 -4094 -13579
rect -4060 -13613 -4048 -13579
rect -4106 -13647 -4048 -13613
rect -4106 -13681 -4094 -13647
rect -4060 -13681 -4048 -13647
rect -4106 -13715 -4048 -13681
rect -4106 -13749 -4094 -13715
rect -4060 -13749 -4048 -13715
rect -4106 -13783 -4048 -13749
rect -4106 -13817 -4094 -13783
rect -4060 -13817 -4048 -13783
rect -4106 -13851 -4048 -13817
rect -4106 -13885 -4094 -13851
rect -4060 -13885 -4048 -13851
rect -4106 -13930 -4048 -13885
rect -3088 -13375 -3030 -13330
rect -3088 -13409 -3076 -13375
rect -3042 -13409 -3030 -13375
rect -3088 -13443 -3030 -13409
rect -3088 -13477 -3076 -13443
rect -3042 -13477 -3030 -13443
rect -3088 -13511 -3030 -13477
rect -3088 -13545 -3076 -13511
rect -3042 -13545 -3030 -13511
rect -3088 -13579 -3030 -13545
rect -3088 -13613 -3076 -13579
rect -3042 -13613 -3030 -13579
rect -3088 -13647 -3030 -13613
rect -3088 -13681 -3076 -13647
rect -3042 -13681 -3030 -13647
rect -3088 -13715 -3030 -13681
rect -3088 -13749 -3076 -13715
rect -3042 -13749 -3030 -13715
rect -3088 -13783 -3030 -13749
rect -3088 -13817 -3076 -13783
rect -3042 -13817 -3030 -13783
rect -3088 -13851 -3030 -13817
rect -3088 -13885 -3076 -13851
rect -3042 -13885 -3030 -13851
rect -3088 -13930 -3030 -13885
rect -2070 -13375 -2012 -13330
rect -2070 -13409 -2058 -13375
rect -2024 -13409 -2012 -13375
rect -2070 -13443 -2012 -13409
rect -2070 -13477 -2058 -13443
rect -2024 -13477 -2012 -13443
rect -2070 -13511 -2012 -13477
rect -2070 -13545 -2058 -13511
rect -2024 -13545 -2012 -13511
rect -2070 -13579 -2012 -13545
rect -2070 -13613 -2058 -13579
rect -2024 -13613 -2012 -13579
rect -2070 -13647 -2012 -13613
rect -2070 -13681 -2058 -13647
rect -2024 -13681 -2012 -13647
rect -2070 -13715 -2012 -13681
rect -2070 -13749 -2058 -13715
rect -2024 -13749 -2012 -13715
rect -2070 -13783 -2012 -13749
rect -2070 -13817 -2058 -13783
rect -2024 -13817 -2012 -13783
rect -2070 -13851 -2012 -13817
rect -2070 -13885 -2058 -13851
rect -2024 -13885 -2012 -13851
rect -2070 -13930 -2012 -13885
rect -1052 -13375 -994 -13330
rect -1052 -13409 -1040 -13375
rect -1006 -13409 -994 -13375
rect -1052 -13443 -994 -13409
rect -1052 -13477 -1040 -13443
rect -1006 -13477 -994 -13443
rect -1052 -13511 -994 -13477
rect -1052 -13545 -1040 -13511
rect -1006 -13545 -994 -13511
rect -1052 -13579 -994 -13545
rect -1052 -13613 -1040 -13579
rect -1006 -13613 -994 -13579
rect -1052 -13647 -994 -13613
rect -1052 -13681 -1040 -13647
rect -1006 -13681 -994 -13647
rect -1052 -13715 -994 -13681
rect -1052 -13749 -1040 -13715
rect -1006 -13749 -994 -13715
rect -1052 -13783 -994 -13749
rect -1052 -13817 -1040 -13783
rect -1006 -13817 -994 -13783
rect -1052 -13851 -994 -13817
rect -1052 -13885 -1040 -13851
rect -1006 -13885 -994 -13851
rect -1052 -13930 -994 -13885
rect -34 -13375 24 -13330
rect -34 -13409 -22 -13375
rect 12 -13409 24 -13375
rect -34 -13443 24 -13409
rect -34 -13477 -22 -13443
rect 12 -13477 24 -13443
rect -34 -13511 24 -13477
rect -34 -13545 -22 -13511
rect 12 -13545 24 -13511
rect -34 -13579 24 -13545
rect -34 -13613 -22 -13579
rect 12 -13613 24 -13579
rect -34 -13647 24 -13613
rect -34 -13681 -22 -13647
rect 12 -13681 24 -13647
rect -34 -13715 24 -13681
rect -34 -13749 -22 -13715
rect 12 -13749 24 -13715
rect -34 -13783 24 -13749
rect -34 -13817 -22 -13783
rect 12 -13817 24 -13783
rect -34 -13851 24 -13817
rect -34 -13885 -22 -13851
rect 12 -13885 24 -13851
rect -34 -13930 24 -13885
rect -9196 -14193 -9138 -14148
rect -9196 -14227 -9184 -14193
rect -9150 -14227 -9138 -14193
rect -9196 -14261 -9138 -14227
rect -9196 -14295 -9184 -14261
rect -9150 -14295 -9138 -14261
rect -9196 -14329 -9138 -14295
rect -9196 -14363 -9184 -14329
rect -9150 -14363 -9138 -14329
rect -9196 -14397 -9138 -14363
rect -9196 -14431 -9184 -14397
rect -9150 -14431 -9138 -14397
rect -9196 -14465 -9138 -14431
rect -9196 -14499 -9184 -14465
rect -9150 -14499 -9138 -14465
rect -9196 -14533 -9138 -14499
rect -9196 -14567 -9184 -14533
rect -9150 -14567 -9138 -14533
rect -9196 -14601 -9138 -14567
rect -9196 -14635 -9184 -14601
rect -9150 -14635 -9138 -14601
rect -9196 -14669 -9138 -14635
rect -9196 -14703 -9184 -14669
rect -9150 -14703 -9138 -14669
rect -9196 -14748 -9138 -14703
rect -8178 -14193 -8120 -14148
rect -8178 -14227 -8166 -14193
rect -8132 -14227 -8120 -14193
rect -8178 -14261 -8120 -14227
rect -8178 -14295 -8166 -14261
rect -8132 -14295 -8120 -14261
rect -8178 -14329 -8120 -14295
rect -8178 -14363 -8166 -14329
rect -8132 -14363 -8120 -14329
rect -8178 -14397 -8120 -14363
rect -8178 -14431 -8166 -14397
rect -8132 -14431 -8120 -14397
rect -8178 -14465 -8120 -14431
rect -8178 -14499 -8166 -14465
rect -8132 -14499 -8120 -14465
rect -8178 -14533 -8120 -14499
rect -8178 -14567 -8166 -14533
rect -8132 -14567 -8120 -14533
rect -8178 -14601 -8120 -14567
rect -8178 -14635 -8166 -14601
rect -8132 -14635 -8120 -14601
rect -8178 -14669 -8120 -14635
rect -8178 -14703 -8166 -14669
rect -8132 -14703 -8120 -14669
rect -8178 -14748 -8120 -14703
rect -7160 -14193 -7102 -14148
rect -7160 -14227 -7148 -14193
rect -7114 -14227 -7102 -14193
rect -7160 -14261 -7102 -14227
rect -7160 -14295 -7148 -14261
rect -7114 -14295 -7102 -14261
rect -7160 -14329 -7102 -14295
rect -7160 -14363 -7148 -14329
rect -7114 -14363 -7102 -14329
rect -7160 -14397 -7102 -14363
rect -7160 -14431 -7148 -14397
rect -7114 -14431 -7102 -14397
rect -7160 -14465 -7102 -14431
rect -7160 -14499 -7148 -14465
rect -7114 -14499 -7102 -14465
rect -7160 -14533 -7102 -14499
rect -7160 -14567 -7148 -14533
rect -7114 -14567 -7102 -14533
rect -7160 -14601 -7102 -14567
rect -7160 -14635 -7148 -14601
rect -7114 -14635 -7102 -14601
rect -7160 -14669 -7102 -14635
rect -7160 -14703 -7148 -14669
rect -7114 -14703 -7102 -14669
rect -7160 -14748 -7102 -14703
rect -6142 -14193 -6084 -14148
rect -6142 -14227 -6130 -14193
rect -6096 -14227 -6084 -14193
rect -6142 -14261 -6084 -14227
rect -6142 -14295 -6130 -14261
rect -6096 -14295 -6084 -14261
rect -6142 -14329 -6084 -14295
rect -6142 -14363 -6130 -14329
rect -6096 -14363 -6084 -14329
rect -6142 -14397 -6084 -14363
rect -6142 -14431 -6130 -14397
rect -6096 -14431 -6084 -14397
rect -6142 -14465 -6084 -14431
rect -6142 -14499 -6130 -14465
rect -6096 -14499 -6084 -14465
rect -6142 -14533 -6084 -14499
rect -6142 -14567 -6130 -14533
rect -6096 -14567 -6084 -14533
rect -6142 -14601 -6084 -14567
rect -6142 -14635 -6130 -14601
rect -6096 -14635 -6084 -14601
rect -6142 -14669 -6084 -14635
rect -6142 -14703 -6130 -14669
rect -6096 -14703 -6084 -14669
rect -6142 -14748 -6084 -14703
rect -5124 -14193 -5066 -14148
rect -5124 -14227 -5112 -14193
rect -5078 -14227 -5066 -14193
rect -5124 -14261 -5066 -14227
rect -5124 -14295 -5112 -14261
rect -5078 -14295 -5066 -14261
rect -5124 -14329 -5066 -14295
rect -5124 -14363 -5112 -14329
rect -5078 -14363 -5066 -14329
rect -5124 -14397 -5066 -14363
rect -5124 -14431 -5112 -14397
rect -5078 -14431 -5066 -14397
rect -5124 -14465 -5066 -14431
rect -5124 -14499 -5112 -14465
rect -5078 -14499 -5066 -14465
rect -5124 -14533 -5066 -14499
rect -5124 -14567 -5112 -14533
rect -5078 -14567 -5066 -14533
rect -5124 -14601 -5066 -14567
rect -5124 -14635 -5112 -14601
rect -5078 -14635 -5066 -14601
rect -5124 -14669 -5066 -14635
rect -5124 -14703 -5112 -14669
rect -5078 -14703 -5066 -14669
rect -5124 -14748 -5066 -14703
rect -4106 -14193 -4048 -14148
rect -4106 -14227 -4094 -14193
rect -4060 -14227 -4048 -14193
rect -4106 -14261 -4048 -14227
rect -4106 -14295 -4094 -14261
rect -4060 -14295 -4048 -14261
rect -4106 -14329 -4048 -14295
rect -4106 -14363 -4094 -14329
rect -4060 -14363 -4048 -14329
rect -4106 -14397 -4048 -14363
rect -4106 -14431 -4094 -14397
rect -4060 -14431 -4048 -14397
rect -4106 -14465 -4048 -14431
rect -4106 -14499 -4094 -14465
rect -4060 -14499 -4048 -14465
rect -4106 -14533 -4048 -14499
rect -4106 -14567 -4094 -14533
rect -4060 -14567 -4048 -14533
rect -4106 -14601 -4048 -14567
rect -4106 -14635 -4094 -14601
rect -4060 -14635 -4048 -14601
rect -4106 -14669 -4048 -14635
rect -4106 -14703 -4094 -14669
rect -4060 -14703 -4048 -14669
rect -4106 -14748 -4048 -14703
rect -3088 -14193 -3030 -14148
rect -3088 -14227 -3076 -14193
rect -3042 -14227 -3030 -14193
rect -3088 -14261 -3030 -14227
rect -3088 -14295 -3076 -14261
rect -3042 -14295 -3030 -14261
rect -3088 -14329 -3030 -14295
rect -3088 -14363 -3076 -14329
rect -3042 -14363 -3030 -14329
rect -3088 -14397 -3030 -14363
rect -3088 -14431 -3076 -14397
rect -3042 -14431 -3030 -14397
rect -3088 -14465 -3030 -14431
rect -3088 -14499 -3076 -14465
rect -3042 -14499 -3030 -14465
rect -3088 -14533 -3030 -14499
rect -3088 -14567 -3076 -14533
rect -3042 -14567 -3030 -14533
rect -3088 -14601 -3030 -14567
rect -3088 -14635 -3076 -14601
rect -3042 -14635 -3030 -14601
rect -3088 -14669 -3030 -14635
rect -3088 -14703 -3076 -14669
rect -3042 -14703 -3030 -14669
rect -3088 -14748 -3030 -14703
rect -2070 -14193 -2012 -14148
rect -2070 -14227 -2058 -14193
rect -2024 -14227 -2012 -14193
rect -2070 -14261 -2012 -14227
rect -2070 -14295 -2058 -14261
rect -2024 -14295 -2012 -14261
rect -2070 -14329 -2012 -14295
rect -2070 -14363 -2058 -14329
rect -2024 -14363 -2012 -14329
rect -2070 -14397 -2012 -14363
rect -2070 -14431 -2058 -14397
rect -2024 -14431 -2012 -14397
rect -2070 -14465 -2012 -14431
rect -2070 -14499 -2058 -14465
rect -2024 -14499 -2012 -14465
rect -2070 -14533 -2012 -14499
rect -2070 -14567 -2058 -14533
rect -2024 -14567 -2012 -14533
rect -2070 -14601 -2012 -14567
rect -2070 -14635 -2058 -14601
rect -2024 -14635 -2012 -14601
rect -2070 -14669 -2012 -14635
rect -2070 -14703 -2058 -14669
rect -2024 -14703 -2012 -14669
rect -2070 -14748 -2012 -14703
rect -1052 -14193 -994 -14148
rect -1052 -14227 -1040 -14193
rect -1006 -14227 -994 -14193
rect -1052 -14261 -994 -14227
rect -1052 -14295 -1040 -14261
rect -1006 -14295 -994 -14261
rect -1052 -14329 -994 -14295
rect -1052 -14363 -1040 -14329
rect -1006 -14363 -994 -14329
rect -1052 -14397 -994 -14363
rect -1052 -14431 -1040 -14397
rect -1006 -14431 -994 -14397
rect -1052 -14465 -994 -14431
rect -1052 -14499 -1040 -14465
rect -1006 -14499 -994 -14465
rect -1052 -14533 -994 -14499
rect -1052 -14567 -1040 -14533
rect -1006 -14567 -994 -14533
rect -1052 -14601 -994 -14567
rect -1052 -14635 -1040 -14601
rect -1006 -14635 -994 -14601
rect -1052 -14669 -994 -14635
rect -1052 -14703 -1040 -14669
rect -1006 -14703 -994 -14669
rect -1052 -14748 -994 -14703
rect -34 -14193 24 -14148
rect -34 -14227 -22 -14193
rect 12 -14227 24 -14193
rect -34 -14261 24 -14227
rect -34 -14295 -22 -14261
rect 12 -14295 24 -14261
rect -34 -14329 24 -14295
rect -34 -14363 -22 -14329
rect 12 -14363 24 -14329
rect -34 -14397 24 -14363
rect -34 -14431 -22 -14397
rect 12 -14431 24 -14397
rect -34 -14465 24 -14431
rect -34 -14499 -22 -14465
rect 12 -14499 24 -14465
rect -34 -14533 24 -14499
rect -34 -14567 -22 -14533
rect 12 -14567 24 -14533
rect -34 -14601 24 -14567
rect -34 -14635 -22 -14601
rect 12 -14635 24 -14601
rect -34 -14669 24 -14635
rect -34 -14703 -22 -14669
rect 12 -14703 24 -14669
rect -34 -14748 24 -14703
rect 2570 -14277 2628 -14232
rect 2570 -14311 2582 -14277
rect 2616 -14311 2628 -14277
rect 2570 -14345 2628 -14311
rect 2570 -14379 2582 -14345
rect 2616 -14379 2628 -14345
rect 2570 -14413 2628 -14379
rect 2570 -14447 2582 -14413
rect 2616 -14447 2628 -14413
rect 2570 -14481 2628 -14447
rect 2570 -14515 2582 -14481
rect 2616 -14515 2628 -14481
rect 2570 -14549 2628 -14515
rect 2570 -14583 2582 -14549
rect 2616 -14583 2628 -14549
rect 2570 -14617 2628 -14583
rect 2570 -14651 2582 -14617
rect 2616 -14651 2628 -14617
rect 2570 -14685 2628 -14651
rect 2570 -14719 2582 -14685
rect 2616 -14719 2628 -14685
rect 2570 -14753 2628 -14719
rect 2570 -14787 2582 -14753
rect 2616 -14787 2628 -14753
rect 2570 -14832 2628 -14787
rect 3588 -14277 3646 -14232
rect 3588 -14311 3600 -14277
rect 3634 -14311 3646 -14277
rect 3588 -14345 3646 -14311
rect 3588 -14379 3600 -14345
rect 3634 -14379 3646 -14345
rect 3588 -14413 3646 -14379
rect 3588 -14447 3600 -14413
rect 3634 -14447 3646 -14413
rect 3588 -14481 3646 -14447
rect 3588 -14515 3600 -14481
rect 3634 -14515 3646 -14481
rect 3588 -14549 3646 -14515
rect 3588 -14583 3600 -14549
rect 3634 -14583 3646 -14549
rect 3588 -14617 3646 -14583
rect 3588 -14651 3600 -14617
rect 3634 -14651 3646 -14617
rect 3588 -14685 3646 -14651
rect 3588 -14719 3600 -14685
rect 3634 -14719 3646 -14685
rect 3588 -14753 3646 -14719
rect 3588 -14787 3600 -14753
rect 3634 -14787 3646 -14753
rect 3588 -14832 3646 -14787
rect 4606 -14277 4664 -14232
rect 4606 -14311 4618 -14277
rect 4652 -14311 4664 -14277
rect 4606 -14345 4664 -14311
rect 4606 -14379 4618 -14345
rect 4652 -14379 4664 -14345
rect 4606 -14413 4664 -14379
rect 4606 -14447 4618 -14413
rect 4652 -14447 4664 -14413
rect 4606 -14481 4664 -14447
rect 4606 -14515 4618 -14481
rect 4652 -14515 4664 -14481
rect 4606 -14549 4664 -14515
rect 4606 -14583 4618 -14549
rect 4652 -14583 4664 -14549
rect 4606 -14617 4664 -14583
rect 4606 -14651 4618 -14617
rect 4652 -14651 4664 -14617
rect 4606 -14685 4664 -14651
rect 4606 -14719 4618 -14685
rect 4652 -14719 4664 -14685
rect 4606 -14753 4664 -14719
rect 4606 -14787 4618 -14753
rect 4652 -14787 4664 -14753
rect 4606 -14832 4664 -14787
rect 5624 -14277 5682 -14232
rect 5624 -14311 5636 -14277
rect 5670 -14311 5682 -14277
rect 5624 -14345 5682 -14311
rect 5624 -14379 5636 -14345
rect 5670 -14379 5682 -14345
rect 5624 -14413 5682 -14379
rect 5624 -14447 5636 -14413
rect 5670 -14447 5682 -14413
rect 5624 -14481 5682 -14447
rect 5624 -14515 5636 -14481
rect 5670 -14515 5682 -14481
rect 5624 -14549 5682 -14515
rect 5624 -14583 5636 -14549
rect 5670 -14583 5682 -14549
rect 5624 -14617 5682 -14583
rect 5624 -14651 5636 -14617
rect 5670 -14651 5682 -14617
rect 5624 -14685 5682 -14651
rect 5624 -14719 5636 -14685
rect 5670 -14719 5682 -14685
rect 5624 -14753 5682 -14719
rect 5624 -14787 5636 -14753
rect 5670 -14787 5682 -14753
rect 5624 -14832 5682 -14787
rect 6642 -14277 6700 -14232
rect 6642 -14311 6654 -14277
rect 6688 -14311 6700 -14277
rect 6642 -14345 6700 -14311
rect 6642 -14379 6654 -14345
rect 6688 -14379 6700 -14345
rect 6642 -14413 6700 -14379
rect 6642 -14447 6654 -14413
rect 6688 -14447 6700 -14413
rect 6642 -14481 6700 -14447
rect 6642 -14515 6654 -14481
rect 6688 -14515 6700 -14481
rect 6642 -14549 6700 -14515
rect 6642 -14583 6654 -14549
rect 6688 -14583 6700 -14549
rect 6642 -14617 6700 -14583
rect 6642 -14651 6654 -14617
rect 6688 -14651 6700 -14617
rect 6642 -14685 6700 -14651
rect 6642 -14719 6654 -14685
rect 6688 -14719 6700 -14685
rect 6642 -14753 6700 -14719
rect 6642 -14787 6654 -14753
rect 6688 -14787 6700 -14753
rect 6642 -14832 6700 -14787
rect 7660 -14277 7718 -14232
rect 7660 -14311 7672 -14277
rect 7706 -14311 7718 -14277
rect 7660 -14345 7718 -14311
rect 7660 -14379 7672 -14345
rect 7706 -14379 7718 -14345
rect 7660 -14413 7718 -14379
rect 7660 -14447 7672 -14413
rect 7706 -14447 7718 -14413
rect 7660 -14481 7718 -14447
rect 7660 -14515 7672 -14481
rect 7706 -14515 7718 -14481
rect 7660 -14549 7718 -14515
rect 7660 -14583 7672 -14549
rect 7706 -14583 7718 -14549
rect 7660 -14617 7718 -14583
rect 7660 -14651 7672 -14617
rect 7706 -14651 7718 -14617
rect 7660 -14685 7718 -14651
rect 7660 -14719 7672 -14685
rect 7706 -14719 7718 -14685
rect 7660 -14753 7718 -14719
rect 7660 -14787 7672 -14753
rect 7706 -14787 7718 -14753
rect 7660 -14832 7718 -14787
rect 8678 -14277 8736 -14232
rect 8678 -14311 8690 -14277
rect 8724 -14311 8736 -14277
rect 8678 -14345 8736 -14311
rect 8678 -14379 8690 -14345
rect 8724 -14379 8736 -14345
rect 8678 -14413 8736 -14379
rect 8678 -14447 8690 -14413
rect 8724 -14447 8736 -14413
rect 8678 -14481 8736 -14447
rect 8678 -14515 8690 -14481
rect 8724 -14515 8736 -14481
rect 8678 -14549 8736 -14515
rect 8678 -14583 8690 -14549
rect 8724 -14583 8736 -14549
rect 8678 -14617 8736 -14583
rect 8678 -14651 8690 -14617
rect 8724 -14651 8736 -14617
rect 8678 -14685 8736 -14651
rect 8678 -14719 8690 -14685
rect 8724 -14719 8736 -14685
rect 8678 -14753 8736 -14719
rect 8678 -14787 8690 -14753
rect 8724 -14787 8736 -14753
rect 8678 -14832 8736 -14787
rect 9696 -14277 9754 -14232
rect 9696 -14311 9708 -14277
rect 9742 -14311 9754 -14277
rect 9696 -14345 9754 -14311
rect 9696 -14379 9708 -14345
rect 9742 -14379 9754 -14345
rect 9696 -14413 9754 -14379
rect 9696 -14447 9708 -14413
rect 9742 -14447 9754 -14413
rect 9696 -14481 9754 -14447
rect 9696 -14515 9708 -14481
rect 9742 -14515 9754 -14481
rect 9696 -14549 9754 -14515
rect 9696 -14583 9708 -14549
rect 9742 -14583 9754 -14549
rect 9696 -14617 9754 -14583
rect 9696 -14651 9708 -14617
rect 9742 -14651 9754 -14617
rect 9696 -14685 9754 -14651
rect 9696 -14719 9708 -14685
rect 9742 -14719 9754 -14685
rect 9696 -14753 9754 -14719
rect 9696 -14787 9708 -14753
rect 9742 -14787 9754 -14753
rect 9696 -14832 9754 -14787
rect 10714 -14277 10772 -14232
rect 10714 -14311 10726 -14277
rect 10760 -14311 10772 -14277
rect 10714 -14345 10772 -14311
rect 10714 -14379 10726 -14345
rect 10760 -14379 10772 -14345
rect 10714 -14413 10772 -14379
rect 10714 -14447 10726 -14413
rect 10760 -14447 10772 -14413
rect 10714 -14481 10772 -14447
rect 10714 -14515 10726 -14481
rect 10760 -14515 10772 -14481
rect 10714 -14549 10772 -14515
rect 10714 -14583 10726 -14549
rect 10760 -14583 10772 -14549
rect 10714 -14617 10772 -14583
rect 10714 -14651 10726 -14617
rect 10760 -14651 10772 -14617
rect 10714 -14685 10772 -14651
rect 10714 -14719 10726 -14685
rect 10760 -14719 10772 -14685
rect 10714 -14753 10772 -14719
rect 10714 -14787 10726 -14753
rect 10760 -14787 10772 -14753
rect 10714 -14832 10772 -14787
rect 11732 -14277 11790 -14232
rect 11732 -14311 11744 -14277
rect 11778 -14311 11790 -14277
rect 11732 -14345 11790 -14311
rect 11732 -14379 11744 -14345
rect 11778 -14379 11790 -14345
rect 11732 -14413 11790 -14379
rect 11732 -14447 11744 -14413
rect 11778 -14447 11790 -14413
rect 11732 -14481 11790 -14447
rect 11732 -14515 11744 -14481
rect 11778 -14515 11790 -14481
rect 11732 -14549 11790 -14515
rect 11732 -14583 11744 -14549
rect 11778 -14583 11790 -14549
rect 11732 -14617 11790 -14583
rect 11732 -14651 11744 -14617
rect 11778 -14651 11790 -14617
rect 11732 -14685 11790 -14651
rect 11732 -14719 11744 -14685
rect 11778 -14719 11790 -14685
rect 11732 -14753 11790 -14719
rect 11732 -14787 11744 -14753
rect 11778 -14787 11790 -14753
rect 11732 -14832 11790 -14787
rect 12750 -14277 12808 -14232
rect 12750 -14311 12762 -14277
rect 12796 -14311 12808 -14277
rect 12750 -14345 12808 -14311
rect 12750 -14379 12762 -14345
rect 12796 -14379 12808 -14345
rect 12750 -14413 12808 -14379
rect 12750 -14447 12762 -14413
rect 12796 -14447 12808 -14413
rect 12750 -14481 12808 -14447
rect 12750 -14515 12762 -14481
rect 12796 -14515 12808 -14481
rect 12750 -14549 12808 -14515
rect 12750 -14583 12762 -14549
rect 12796 -14583 12808 -14549
rect 12750 -14617 12808 -14583
rect 12750 -14651 12762 -14617
rect 12796 -14651 12808 -14617
rect 12750 -14685 12808 -14651
rect 12750 -14719 12762 -14685
rect 12796 -14719 12808 -14685
rect 12750 -14753 12808 -14719
rect 12750 -14787 12762 -14753
rect 12796 -14787 12808 -14753
rect 12750 -14832 12808 -14787
rect 13768 -14277 13826 -14232
rect 13768 -14311 13780 -14277
rect 13814 -14311 13826 -14277
rect 13768 -14345 13826 -14311
rect 13768 -14379 13780 -14345
rect 13814 -14379 13826 -14345
rect 13768 -14413 13826 -14379
rect 13768 -14447 13780 -14413
rect 13814 -14447 13826 -14413
rect 13768 -14481 13826 -14447
rect 13768 -14515 13780 -14481
rect 13814 -14515 13826 -14481
rect 13768 -14549 13826 -14515
rect 13768 -14583 13780 -14549
rect 13814 -14583 13826 -14549
rect 13768 -14617 13826 -14583
rect 13768 -14651 13780 -14617
rect 13814 -14651 13826 -14617
rect 13768 -14685 13826 -14651
rect 13768 -14719 13780 -14685
rect 13814 -14719 13826 -14685
rect 13768 -14753 13826 -14719
rect 13768 -14787 13780 -14753
rect 13814 -14787 13826 -14753
rect 13768 -14832 13826 -14787
rect 14786 -14277 14844 -14232
rect 14786 -14311 14798 -14277
rect 14832 -14311 14844 -14277
rect 14786 -14345 14844 -14311
rect 14786 -14379 14798 -14345
rect 14832 -14379 14844 -14345
rect 14786 -14413 14844 -14379
rect 14786 -14447 14798 -14413
rect 14832 -14447 14844 -14413
rect 14786 -14481 14844 -14447
rect 14786 -14515 14798 -14481
rect 14832 -14515 14844 -14481
rect 14786 -14549 14844 -14515
rect 14786 -14583 14798 -14549
rect 14832 -14583 14844 -14549
rect 14786 -14617 14844 -14583
rect 14786 -14651 14798 -14617
rect 14832 -14651 14844 -14617
rect 14786 -14685 14844 -14651
rect 14786 -14719 14798 -14685
rect 14832 -14719 14844 -14685
rect 14786 -14753 14844 -14719
rect 14786 -14787 14798 -14753
rect 14832 -14787 14844 -14753
rect 14786 -14832 14844 -14787
rect 15804 -14277 15862 -14232
rect 15804 -14311 15816 -14277
rect 15850 -14311 15862 -14277
rect 15804 -14345 15862 -14311
rect 15804 -14379 15816 -14345
rect 15850 -14379 15862 -14345
rect 15804 -14413 15862 -14379
rect 15804 -14447 15816 -14413
rect 15850 -14447 15862 -14413
rect 15804 -14481 15862 -14447
rect 15804 -14515 15816 -14481
rect 15850 -14515 15862 -14481
rect 15804 -14549 15862 -14515
rect 15804 -14583 15816 -14549
rect 15850 -14583 15862 -14549
rect 15804 -14617 15862 -14583
rect 15804 -14651 15816 -14617
rect 15850 -14651 15862 -14617
rect 15804 -14685 15862 -14651
rect 15804 -14719 15816 -14685
rect 15850 -14719 15862 -14685
rect 15804 -14753 15862 -14719
rect 15804 -14787 15816 -14753
rect 15850 -14787 15862 -14753
rect 15804 -14832 15862 -14787
rect 16822 -14277 16880 -14232
rect 16822 -14311 16834 -14277
rect 16868 -14311 16880 -14277
rect 16822 -14345 16880 -14311
rect 16822 -14379 16834 -14345
rect 16868 -14379 16880 -14345
rect 16822 -14413 16880 -14379
rect 16822 -14447 16834 -14413
rect 16868 -14447 16880 -14413
rect 16822 -14481 16880 -14447
rect 16822 -14515 16834 -14481
rect 16868 -14515 16880 -14481
rect 16822 -14549 16880 -14515
rect 16822 -14583 16834 -14549
rect 16868 -14583 16880 -14549
rect 16822 -14617 16880 -14583
rect 16822 -14651 16834 -14617
rect 16868 -14651 16880 -14617
rect 16822 -14685 16880 -14651
rect 16822 -14719 16834 -14685
rect 16868 -14719 16880 -14685
rect 16822 -14753 16880 -14719
rect 16822 -14787 16834 -14753
rect 16868 -14787 16880 -14753
rect 16822 -14832 16880 -14787
rect 17840 -14277 17898 -14232
rect 17840 -14311 17852 -14277
rect 17886 -14311 17898 -14277
rect 17840 -14345 17898 -14311
rect 17840 -14379 17852 -14345
rect 17886 -14379 17898 -14345
rect 17840 -14413 17898 -14379
rect 17840 -14447 17852 -14413
rect 17886 -14447 17898 -14413
rect 17840 -14481 17898 -14447
rect 17840 -14515 17852 -14481
rect 17886 -14515 17898 -14481
rect 17840 -14549 17898 -14515
rect 17840 -14583 17852 -14549
rect 17886 -14583 17898 -14549
rect 17840 -14617 17898 -14583
rect 17840 -14651 17852 -14617
rect 17886 -14651 17898 -14617
rect 17840 -14685 17898 -14651
rect 17840 -14719 17852 -14685
rect 17886 -14719 17898 -14685
rect 17840 -14753 17898 -14719
rect 17840 -14787 17852 -14753
rect 17886 -14787 17898 -14753
rect 17840 -14832 17898 -14787
rect 18858 -14277 18916 -14232
rect 18858 -14311 18870 -14277
rect 18904 -14311 18916 -14277
rect 18858 -14345 18916 -14311
rect 18858 -14379 18870 -14345
rect 18904 -14379 18916 -14345
rect 18858 -14413 18916 -14379
rect 18858 -14447 18870 -14413
rect 18904 -14447 18916 -14413
rect 18858 -14481 18916 -14447
rect 18858 -14515 18870 -14481
rect 18904 -14515 18916 -14481
rect 18858 -14549 18916 -14515
rect 18858 -14583 18870 -14549
rect 18904 -14583 18916 -14549
rect 18858 -14617 18916 -14583
rect 18858 -14651 18870 -14617
rect 18904 -14651 18916 -14617
rect 18858 -14685 18916 -14651
rect 18858 -14719 18870 -14685
rect 18904 -14719 18916 -14685
rect 18858 -14753 18916 -14719
rect 18858 -14787 18870 -14753
rect 18904 -14787 18916 -14753
rect 18858 -14832 18916 -14787
rect 19876 -14277 19934 -14232
rect 19876 -14311 19888 -14277
rect 19922 -14311 19934 -14277
rect 19876 -14345 19934 -14311
rect 19876 -14379 19888 -14345
rect 19922 -14379 19934 -14345
rect 19876 -14413 19934 -14379
rect 19876 -14447 19888 -14413
rect 19922 -14447 19934 -14413
rect 19876 -14481 19934 -14447
rect 19876 -14515 19888 -14481
rect 19922 -14515 19934 -14481
rect 19876 -14549 19934 -14515
rect 19876 -14583 19888 -14549
rect 19922 -14583 19934 -14549
rect 19876 -14617 19934 -14583
rect 19876 -14651 19888 -14617
rect 19922 -14651 19934 -14617
rect 19876 -14685 19934 -14651
rect 19876 -14719 19888 -14685
rect 19922 -14719 19934 -14685
rect 19876 -14753 19934 -14719
rect 19876 -14787 19888 -14753
rect 19922 -14787 19934 -14753
rect 19876 -14832 19934 -14787
rect 20894 -14277 20952 -14232
rect 20894 -14311 20906 -14277
rect 20940 -14311 20952 -14277
rect 20894 -14345 20952 -14311
rect 20894 -14379 20906 -14345
rect 20940 -14379 20952 -14345
rect 20894 -14413 20952 -14379
rect 20894 -14447 20906 -14413
rect 20940 -14447 20952 -14413
rect 20894 -14481 20952 -14447
rect 20894 -14515 20906 -14481
rect 20940 -14515 20952 -14481
rect 20894 -14549 20952 -14515
rect 20894 -14583 20906 -14549
rect 20940 -14583 20952 -14549
rect 20894 -14617 20952 -14583
rect 20894 -14651 20906 -14617
rect 20940 -14651 20952 -14617
rect 20894 -14685 20952 -14651
rect 20894 -14719 20906 -14685
rect 20940 -14719 20952 -14685
rect 20894 -14753 20952 -14719
rect 20894 -14787 20906 -14753
rect 20940 -14787 20952 -14753
rect 20894 -14832 20952 -14787
rect 21912 -14277 21970 -14232
rect 21912 -14311 21924 -14277
rect 21958 -14311 21970 -14277
rect 21912 -14345 21970 -14311
rect 21912 -14379 21924 -14345
rect 21958 -14379 21970 -14345
rect 21912 -14413 21970 -14379
rect 21912 -14447 21924 -14413
rect 21958 -14447 21970 -14413
rect 21912 -14481 21970 -14447
rect 21912 -14515 21924 -14481
rect 21958 -14515 21970 -14481
rect 21912 -14549 21970 -14515
rect 21912 -14583 21924 -14549
rect 21958 -14583 21970 -14549
rect 21912 -14617 21970 -14583
rect 21912 -14651 21924 -14617
rect 21958 -14651 21970 -14617
rect 21912 -14685 21970 -14651
rect 21912 -14719 21924 -14685
rect 21958 -14719 21970 -14685
rect 21912 -14753 21970 -14719
rect 21912 -14787 21924 -14753
rect 21958 -14787 21970 -14753
rect 21912 -14832 21970 -14787
rect 22930 -14277 22988 -14232
rect 22930 -14311 22942 -14277
rect 22976 -14311 22988 -14277
rect 22930 -14345 22988 -14311
rect 22930 -14379 22942 -14345
rect 22976 -14379 22988 -14345
rect 22930 -14413 22988 -14379
rect 22930 -14447 22942 -14413
rect 22976 -14447 22988 -14413
rect 22930 -14481 22988 -14447
rect 22930 -14515 22942 -14481
rect 22976 -14515 22988 -14481
rect 22930 -14549 22988 -14515
rect 22930 -14583 22942 -14549
rect 22976 -14583 22988 -14549
rect 22930 -14617 22988 -14583
rect 22930 -14651 22942 -14617
rect 22976 -14651 22988 -14617
rect 22930 -14685 22988 -14651
rect 22930 -14719 22942 -14685
rect 22976 -14719 22988 -14685
rect 22930 -14753 22988 -14719
rect 22930 -14787 22942 -14753
rect 22976 -14787 22988 -14753
rect 22930 -14832 22988 -14787
rect -9196 -15011 -9138 -14966
rect -9196 -15045 -9184 -15011
rect -9150 -15045 -9138 -15011
rect -9196 -15079 -9138 -15045
rect -9196 -15113 -9184 -15079
rect -9150 -15113 -9138 -15079
rect -9196 -15147 -9138 -15113
rect -9196 -15181 -9184 -15147
rect -9150 -15181 -9138 -15147
rect -9196 -15215 -9138 -15181
rect -9196 -15249 -9184 -15215
rect -9150 -15249 -9138 -15215
rect -9196 -15283 -9138 -15249
rect -9196 -15317 -9184 -15283
rect -9150 -15317 -9138 -15283
rect -9196 -15351 -9138 -15317
rect -9196 -15385 -9184 -15351
rect -9150 -15385 -9138 -15351
rect -9196 -15419 -9138 -15385
rect -9196 -15453 -9184 -15419
rect -9150 -15453 -9138 -15419
rect -9196 -15487 -9138 -15453
rect -9196 -15521 -9184 -15487
rect -9150 -15521 -9138 -15487
rect -9196 -15566 -9138 -15521
rect -8178 -15011 -8120 -14966
rect -8178 -15045 -8166 -15011
rect -8132 -15045 -8120 -15011
rect -8178 -15079 -8120 -15045
rect -8178 -15113 -8166 -15079
rect -8132 -15113 -8120 -15079
rect -8178 -15147 -8120 -15113
rect -8178 -15181 -8166 -15147
rect -8132 -15181 -8120 -15147
rect -8178 -15215 -8120 -15181
rect -8178 -15249 -8166 -15215
rect -8132 -15249 -8120 -15215
rect -8178 -15283 -8120 -15249
rect -8178 -15317 -8166 -15283
rect -8132 -15317 -8120 -15283
rect -8178 -15351 -8120 -15317
rect -8178 -15385 -8166 -15351
rect -8132 -15385 -8120 -15351
rect -8178 -15419 -8120 -15385
rect -8178 -15453 -8166 -15419
rect -8132 -15453 -8120 -15419
rect -8178 -15487 -8120 -15453
rect -8178 -15521 -8166 -15487
rect -8132 -15521 -8120 -15487
rect -8178 -15566 -8120 -15521
rect -7160 -15011 -7102 -14966
rect -7160 -15045 -7148 -15011
rect -7114 -15045 -7102 -15011
rect -7160 -15079 -7102 -15045
rect -7160 -15113 -7148 -15079
rect -7114 -15113 -7102 -15079
rect -7160 -15147 -7102 -15113
rect -7160 -15181 -7148 -15147
rect -7114 -15181 -7102 -15147
rect -7160 -15215 -7102 -15181
rect -7160 -15249 -7148 -15215
rect -7114 -15249 -7102 -15215
rect -7160 -15283 -7102 -15249
rect -7160 -15317 -7148 -15283
rect -7114 -15317 -7102 -15283
rect -7160 -15351 -7102 -15317
rect -7160 -15385 -7148 -15351
rect -7114 -15385 -7102 -15351
rect -7160 -15419 -7102 -15385
rect -7160 -15453 -7148 -15419
rect -7114 -15453 -7102 -15419
rect -7160 -15487 -7102 -15453
rect -7160 -15521 -7148 -15487
rect -7114 -15521 -7102 -15487
rect -7160 -15566 -7102 -15521
rect -6142 -15011 -6084 -14966
rect -6142 -15045 -6130 -15011
rect -6096 -15045 -6084 -15011
rect -6142 -15079 -6084 -15045
rect -6142 -15113 -6130 -15079
rect -6096 -15113 -6084 -15079
rect -6142 -15147 -6084 -15113
rect -6142 -15181 -6130 -15147
rect -6096 -15181 -6084 -15147
rect -6142 -15215 -6084 -15181
rect -6142 -15249 -6130 -15215
rect -6096 -15249 -6084 -15215
rect -6142 -15283 -6084 -15249
rect -6142 -15317 -6130 -15283
rect -6096 -15317 -6084 -15283
rect -6142 -15351 -6084 -15317
rect -6142 -15385 -6130 -15351
rect -6096 -15385 -6084 -15351
rect -6142 -15419 -6084 -15385
rect -6142 -15453 -6130 -15419
rect -6096 -15453 -6084 -15419
rect -6142 -15487 -6084 -15453
rect -6142 -15521 -6130 -15487
rect -6096 -15521 -6084 -15487
rect -6142 -15566 -6084 -15521
rect -5124 -15011 -5066 -14966
rect -5124 -15045 -5112 -15011
rect -5078 -15045 -5066 -15011
rect -5124 -15079 -5066 -15045
rect -5124 -15113 -5112 -15079
rect -5078 -15113 -5066 -15079
rect -5124 -15147 -5066 -15113
rect -5124 -15181 -5112 -15147
rect -5078 -15181 -5066 -15147
rect -5124 -15215 -5066 -15181
rect -5124 -15249 -5112 -15215
rect -5078 -15249 -5066 -15215
rect -5124 -15283 -5066 -15249
rect -5124 -15317 -5112 -15283
rect -5078 -15317 -5066 -15283
rect -5124 -15351 -5066 -15317
rect -5124 -15385 -5112 -15351
rect -5078 -15385 -5066 -15351
rect -5124 -15419 -5066 -15385
rect -5124 -15453 -5112 -15419
rect -5078 -15453 -5066 -15419
rect -5124 -15487 -5066 -15453
rect -5124 -15521 -5112 -15487
rect -5078 -15521 -5066 -15487
rect -5124 -15566 -5066 -15521
rect -4106 -15011 -4048 -14966
rect -4106 -15045 -4094 -15011
rect -4060 -15045 -4048 -15011
rect -4106 -15079 -4048 -15045
rect -4106 -15113 -4094 -15079
rect -4060 -15113 -4048 -15079
rect -4106 -15147 -4048 -15113
rect -4106 -15181 -4094 -15147
rect -4060 -15181 -4048 -15147
rect -4106 -15215 -4048 -15181
rect -4106 -15249 -4094 -15215
rect -4060 -15249 -4048 -15215
rect -4106 -15283 -4048 -15249
rect -4106 -15317 -4094 -15283
rect -4060 -15317 -4048 -15283
rect -4106 -15351 -4048 -15317
rect -4106 -15385 -4094 -15351
rect -4060 -15385 -4048 -15351
rect -4106 -15419 -4048 -15385
rect -4106 -15453 -4094 -15419
rect -4060 -15453 -4048 -15419
rect -4106 -15487 -4048 -15453
rect -4106 -15521 -4094 -15487
rect -4060 -15521 -4048 -15487
rect -4106 -15566 -4048 -15521
rect -3088 -15011 -3030 -14966
rect -3088 -15045 -3076 -15011
rect -3042 -15045 -3030 -15011
rect -3088 -15079 -3030 -15045
rect -3088 -15113 -3076 -15079
rect -3042 -15113 -3030 -15079
rect -3088 -15147 -3030 -15113
rect -3088 -15181 -3076 -15147
rect -3042 -15181 -3030 -15147
rect -3088 -15215 -3030 -15181
rect -3088 -15249 -3076 -15215
rect -3042 -15249 -3030 -15215
rect -3088 -15283 -3030 -15249
rect -3088 -15317 -3076 -15283
rect -3042 -15317 -3030 -15283
rect -3088 -15351 -3030 -15317
rect -3088 -15385 -3076 -15351
rect -3042 -15385 -3030 -15351
rect -3088 -15419 -3030 -15385
rect -3088 -15453 -3076 -15419
rect -3042 -15453 -3030 -15419
rect -3088 -15487 -3030 -15453
rect -3088 -15521 -3076 -15487
rect -3042 -15521 -3030 -15487
rect -3088 -15566 -3030 -15521
rect -2070 -15011 -2012 -14966
rect -2070 -15045 -2058 -15011
rect -2024 -15045 -2012 -15011
rect -2070 -15079 -2012 -15045
rect -2070 -15113 -2058 -15079
rect -2024 -15113 -2012 -15079
rect -2070 -15147 -2012 -15113
rect -2070 -15181 -2058 -15147
rect -2024 -15181 -2012 -15147
rect -2070 -15215 -2012 -15181
rect -2070 -15249 -2058 -15215
rect -2024 -15249 -2012 -15215
rect -2070 -15283 -2012 -15249
rect -2070 -15317 -2058 -15283
rect -2024 -15317 -2012 -15283
rect -2070 -15351 -2012 -15317
rect -2070 -15385 -2058 -15351
rect -2024 -15385 -2012 -15351
rect -2070 -15419 -2012 -15385
rect -2070 -15453 -2058 -15419
rect -2024 -15453 -2012 -15419
rect -2070 -15487 -2012 -15453
rect -2070 -15521 -2058 -15487
rect -2024 -15521 -2012 -15487
rect -2070 -15566 -2012 -15521
rect -1052 -15011 -994 -14966
rect -1052 -15045 -1040 -15011
rect -1006 -15045 -994 -15011
rect -1052 -15079 -994 -15045
rect -1052 -15113 -1040 -15079
rect -1006 -15113 -994 -15079
rect -1052 -15147 -994 -15113
rect -1052 -15181 -1040 -15147
rect -1006 -15181 -994 -15147
rect -1052 -15215 -994 -15181
rect -1052 -15249 -1040 -15215
rect -1006 -15249 -994 -15215
rect -1052 -15283 -994 -15249
rect -1052 -15317 -1040 -15283
rect -1006 -15317 -994 -15283
rect -1052 -15351 -994 -15317
rect -1052 -15385 -1040 -15351
rect -1006 -15385 -994 -15351
rect -1052 -15419 -994 -15385
rect -1052 -15453 -1040 -15419
rect -1006 -15453 -994 -15419
rect -1052 -15487 -994 -15453
rect -1052 -15521 -1040 -15487
rect -1006 -15521 -994 -15487
rect -1052 -15566 -994 -15521
rect -34 -15011 24 -14966
rect -34 -15045 -22 -15011
rect 12 -15045 24 -15011
rect -34 -15079 24 -15045
rect -34 -15113 -22 -15079
rect 12 -15113 24 -15079
rect -34 -15147 24 -15113
rect -34 -15181 -22 -15147
rect 12 -15181 24 -15147
rect -34 -15215 24 -15181
rect -34 -15249 -22 -15215
rect 12 -15249 24 -15215
rect -34 -15283 24 -15249
rect -34 -15317 -22 -15283
rect 12 -15317 24 -15283
rect -34 -15351 24 -15317
rect -34 -15385 -22 -15351
rect 12 -15385 24 -15351
rect -34 -15419 24 -15385
rect -34 -15453 -22 -15419
rect 12 -15453 24 -15419
rect -34 -15487 24 -15453
rect -34 -15521 -22 -15487
rect 12 -15521 24 -15487
rect -34 -15566 24 -15521
rect 2570 -15509 2628 -15464
rect 2570 -15543 2582 -15509
rect 2616 -15543 2628 -15509
rect 2570 -15577 2628 -15543
rect 2570 -15611 2582 -15577
rect 2616 -15611 2628 -15577
rect 2570 -15645 2628 -15611
rect 2570 -15679 2582 -15645
rect 2616 -15679 2628 -15645
rect 2570 -15713 2628 -15679
rect 2570 -15747 2582 -15713
rect 2616 -15747 2628 -15713
rect 2570 -15781 2628 -15747
rect -9196 -15829 -9138 -15784
rect -9196 -15863 -9184 -15829
rect -9150 -15863 -9138 -15829
rect -9196 -15897 -9138 -15863
rect -9196 -15931 -9184 -15897
rect -9150 -15931 -9138 -15897
rect -9196 -15965 -9138 -15931
rect -9196 -15999 -9184 -15965
rect -9150 -15999 -9138 -15965
rect -9196 -16033 -9138 -15999
rect -9196 -16067 -9184 -16033
rect -9150 -16067 -9138 -16033
rect -9196 -16101 -9138 -16067
rect -9196 -16135 -9184 -16101
rect -9150 -16135 -9138 -16101
rect -9196 -16169 -9138 -16135
rect -9196 -16203 -9184 -16169
rect -9150 -16203 -9138 -16169
rect -9196 -16237 -9138 -16203
rect -9196 -16271 -9184 -16237
rect -9150 -16271 -9138 -16237
rect -9196 -16305 -9138 -16271
rect -9196 -16339 -9184 -16305
rect -9150 -16339 -9138 -16305
rect -9196 -16384 -9138 -16339
rect -8178 -15829 -8120 -15784
rect -8178 -15863 -8166 -15829
rect -8132 -15863 -8120 -15829
rect -8178 -15897 -8120 -15863
rect -8178 -15931 -8166 -15897
rect -8132 -15931 -8120 -15897
rect -8178 -15965 -8120 -15931
rect -8178 -15999 -8166 -15965
rect -8132 -15999 -8120 -15965
rect -8178 -16033 -8120 -15999
rect -8178 -16067 -8166 -16033
rect -8132 -16067 -8120 -16033
rect -8178 -16101 -8120 -16067
rect -8178 -16135 -8166 -16101
rect -8132 -16135 -8120 -16101
rect -8178 -16169 -8120 -16135
rect -8178 -16203 -8166 -16169
rect -8132 -16203 -8120 -16169
rect -8178 -16237 -8120 -16203
rect -8178 -16271 -8166 -16237
rect -8132 -16271 -8120 -16237
rect -8178 -16305 -8120 -16271
rect -8178 -16339 -8166 -16305
rect -8132 -16339 -8120 -16305
rect -8178 -16384 -8120 -16339
rect -7160 -15829 -7102 -15784
rect -7160 -15863 -7148 -15829
rect -7114 -15863 -7102 -15829
rect -7160 -15897 -7102 -15863
rect -7160 -15931 -7148 -15897
rect -7114 -15931 -7102 -15897
rect -7160 -15965 -7102 -15931
rect -7160 -15999 -7148 -15965
rect -7114 -15999 -7102 -15965
rect -7160 -16033 -7102 -15999
rect -7160 -16067 -7148 -16033
rect -7114 -16067 -7102 -16033
rect -7160 -16101 -7102 -16067
rect -7160 -16135 -7148 -16101
rect -7114 -16135 -7102 -16101
rect -7160 -16169 -7102 -16135
rect -7160 -16203 -7148 -16169
rect -7114 -16203 -7102 -16169
rect -7160 -16237 -7102 -16203
rect -7160 -16271 -7148 -16237
rect -7114 -16271 -7102 -16237
rect -7160 -16305 -7102 -16271
rect -7160 -16339 -7148 -16305
rect -7114 -16339 -7102 -16305
rect -7160 -16384 -7102 -16339
rect -6142 -15829 -6084 -15784
rect -6142 -15863 -6130 -15829
rect -6096 -15863 -6084 -15829
rect -6142 -15897 -6084 -15863
rect -6142 -15931 -6130 -15897
rect -6096 -15931 -6084 -15897
rect -6142 -15965 -6084 -15931
rect -6142 -15999 -6130 -15965
rect -6096 -15999 -6084 -15965
rect -6142 -16033 -6084 -15999
rect -6142 -16067 -6130 -16033
rect -6096 -16067 -6084 -16033
rect -6142 -16101 -6084 -16067
rect -6142 -16135 -6130 -16101
rect -6096 -16135 -6084 -16101
rect -6142 -16169 -6084 -16135
rect -6142 -16203 -6130 -16169
rect -6096 -16203 -6084 -16169
rect -6142 -16237 -6084 -16203
rect -6142 -16271 -6130 -16237
rect -6096 -16271 -6084 -16237
rect -6142 -16305 -6084 -16271
rect -6142 -16339 -6130 -16305
rect -6096 -16339 -6084 -16305
rect -6142 -16384 -6084 -16339
rect -5124 -15829 -5066 -15784
rect -5124 -15863 -5112 -15829
rect -5078 -15863 -5066 -15829
rect -5124 -15897 -5066 -15863
rect -5124 -15931 -5112 -15897
rect -5078 -15931 -5066 -15897
rect -5124 -15965 -5066 -15931
rect -5124 -15999 -5112 -15965
rect -5078 -15999 -5066 -15965
rect -5124 -16033 -5066 -15999
rect -5124 -16067 -5112 -16033
rect -5078 -16067 -5066 -16033
rect -5124 -16101 -5066 -16067
rect -5124 -16135 -5112 -16101
rect -5078 -16135 -5066 -16101
rect -5124 -16169 -5066 -16135
rect -5124 -16203 -5112 -16169
rect -5078 -16203 -5066 -16169
rect -5124 -16237 -5066 -16203
rect -5124 -16271 -5112 -16237
rect -5078 -16271 -5066 -16237
rect -5124 -16305 -5066 -16271
rect -5124 -16339 -5112 -16305
rect -5078 -16339 -5066 -16305
rect -5124 -16384 -5066 -16339
rect -4106 -15829 -4048 -15784
rect -4106 -15863 -4094 -15829
rect -4060 -15863 -4048 -15829
rect -4106 -15897 -4048 -15863
rect -4106 -15931 -4094 -15897
rect -4060 -15931 -4048 -15897
rect -4106 -15965 -4048 -15931
rect -4106 -15999 -4094 -15965
rect -4060 -15999 -4048 -15965
rect -4106 -16033 -4048 -15999
rect -4106 -16067 -4094 -16033
rect -4060 -16067 -4048 -16033
rect -4106 -16101 -4048 -16067
rect -4106 -16135 -4094 -16101
rect -4060 -16135 -4048 -16101
rect -4106 -16169 -4048 -16135
rect -4106 -16203 -4094 -16169
rect -4060 -16203 -4048 -16169
rect -4106 -16237 -4048 -16203
rect -4106 -16271 -4094 -16237
rect -4060 -16271 -4048 -16237
rect -4106 -16305 -4048 -16271
rect -4106 -16339 -4094 -16305
rect -4060 -16339 -4048 -16305
rect -4106 -16384 -4048 -16339
rect -3088 -15829 -3030 -15784
rect -3088 -15863 -3076 -15829
rect -3042 -15863 -3030 -15829
rect -3088 -15897 -3030 -15863
rect -3088 -15931 -3076 -15897
rect -3042 -15931 -3030 -15897
rect -3088 -15965 -3030 -15931
rect -3088 -15999 -3076 -15965
rect -3042 -15999 -3030 -15965
rect -3088 -16033 -3030 -15999
rect -3088 -16067 -3076 -16033
rect -3042 -16067 -3030 -16033
rect -3088 -16101 -3030 -16067
rect -3088 -16135 -3076 -16101
rect -3042 -16135 -3030 -16101
rect -3088 -16169 -3030 -16135
rect -3088 -16203 -3076 -16169
rect -3042 -16203 -3030 -16169
rect -3088 -16237 -3030 -16203
rect -3088 -16271 -3076 -16237
rect -3042 -16271 -3030 -16237
rect -3088 -16305 -3030 -16271
rect -3088 -16339 -3076 -16305
rect -3042 -16339 -3030 -16305
rect -3088 -16384 -3030 -16339
rect -2070 -15829 -2012 -15784
rect -2070 -15863 -2058 -15829
rect -2024 -15863 -2012 -15829
rect -2070 -15897 -2012 -15863
rect -2070 -15931 -2058 -15897
rect -2024 -15931 -2012 -15897
rect -2070 -15965 -2012 -15931
rect -2070 -15999 -2058 -15965
rect -2024 -15999 -2012 -15965
rect -2070 -16033 -2012 -15999
rect -2070 -16067 -2058 -16033
rect -2024 -16067 -2012 -16033
rect -2070 -16101 -2012 -16067
rect -2070 -16135 -2058 -16101
rect -2024 -16135 -2012 -16101
rect -2070 -16169 -2012 -16135
rect -2070 -16203 -2058 -16169
rect -2024 -16203 -2012 -16169
rect -2070 -16237 -2012 -16203
rect -2070 -16271 -2058 -16237
rect -2024 -16271 -2012 -16237
rect -2070 -16305 -2012 -16271
rect -2070 -16339 -2058 -16305
rect -2024 -16339 -2012 -16305
rect -2070 -16384 -2012 -16339
rect -1052 -15829 -994 -15784
rect -1052 -15863 -1040 -15829
rect -1006 -15863 -994 -15829
rect -1052 -15897 -994 -15863
rect -1052 -15931 -1040 -15897
rect -1006 -15931 -994 -15897
rect -1052 -15965 -994 -15931
rect -1052 -15999 -1040 -15965
rect -1006 -15999 -994 -15965
rect -1052 -16033 -994 -15999
rect -1052 -16067 -1040 -16033
rect -1006 -16067 -994 -16033
rect -1052 -16101 -994 -16067
rect -1052 -16135 -1040 -16101
rect -1006 -16135 -994 -16101
rect -1052 -16169 -994 -16135
rect -1052 -16203 -1040 -16169
rect -1006 -16203 -994 -16169
rect -1052 -16237 -994 -16203
rect -1052 -16271 -1040 -16237
rect -1006 -16271 -994 -16237
rect -1052 -16305 -994 -16271
rect -1052 -16339 -1040 -16305
rect -1006 -16339 -994 -16305
rect -1052 -16384 -994 -16339
rect -34 -15829 24 -15784
rect -34 -15863 -22 -15829
rect 12 -15863 24 -15829
rect -34 -15897 24 -15863
rect -34 -15931 -22 -15897
rect 12 -15931 24 -15897
rect -34 -15965 24 -15931
rect -34 -15999 -22 -15965
rect 12 -15999 24 -15965
rect -34 -16033 24 -15999
rect -34 -16067 -22 -16033
rect 12 -16067 24 -16033
rect 2570 -15815 2582 -15781
rect 2616 -15815 2628 -15781
rect 2570 -15849 2628 -15815
rect 2570 -15883 2582 -15849
rect 2616 -15883 2628 -15849
rect 2570 -15917 2628 -15883
rect 2570 -15951 2582 -15917
rect 2616 -15951 2628 -15917
rect 2570 -15985 2628 -15951
rect 2570 -16019 2582 -15985
rect 2616 -16019 2628 -15985
rect 2570 -16064 2628 -16019
rect 3588 -15509 3646 -15464
rect 3588 -15543 3600 -15509
rect 3634 -15543 3646 -15509
rect 3588 -15577 3646 -15543
rect 3588 -15611 3600 -15577
rect 3634 -15611 3646 -15577
rect 3588 -15645 3646 -15611
rect 3588 -15679 3600 -15645
rect 3634 -15679 3646 -15645
rect 3588 -15713 3646 -15679
rect 3588 -15747 3600 -15713
rect 3634 -15747 3646 -15713
rect 3588 -15781 3646 -15747
rect 3588 -15815 3600 -15781
rect 3634 -15815 3646 -15781
rect 3588 -15849 3646 -15815
rect 3588 -15883 3600 -15849
rect 3634 -15883 3646 -15849
rect 3588 -15917 3646 -15883
rect 3588 -15951 3600 -15917
rect 3634 -15951 3646 -15917
rect 3588 -15985 3646 -15951
rect 3588 -16019 3600 -15985
rect 3634 -16019 3646 -15985
rect 3588 -16064 3646 -16019
rect 4606 -15509 4664 -15464
rect 4606 -15543 4618 -15509
rect 4652 -15543 4664 -15509
rect 4606 -15577 4664 -15543
rect 4606 -15611 4618 -15577
rect 4652 -15611 4664 -15577
rect 4606 -15645 4664 -15611
rect 4606 -15679 4618 -15645
rect 4652 -15679 4664 -15645
rect 4606 -15713 4664 -15679
rect 4606 -15747 4618 -15713
rect 4652 -15747 4664 -15713
rect 4606 -15781 4664 -15747
rect 4606 -15815 4618 -15781
rect 4652 -15815 4664 -15781
rect 4606 -15849 4664 -15815
rect 4606 -15883 4618 -15849
rect 4652 -15883 4664 -15849
rect 4606 -15917 4664 -15883
rect 4606 -15951 4618 -15917
rect 4652 -15951 4664 -15917
rect 4606 -15985 4664 -15951
rect 4606 -16019 4618 -15985
rect 4652 -16019 4664 -15985
rect 4606 -16064 4664 -16019
rect 5624 -15509 5682 -15464
rect 5624 -15543 5636 -15509
rect 5670 -15543 5682 -15509
rect 5624 -15577 5682 -15543
rect 5624 -15611 5636 -15577
rect 5670 -15611 5682 -15577
rect 5624 -15645 5682 -15611
rect 5624 -15679 5636 -15645
rect 5670 -15679 5682 -15645
rect 5624 -15713 5682 -15679
rect 5624 -15747 5636 -15713
rect 5670 -15747 5682 -15713
rect 5624 -15781 5682 -15747
rect 5624 -15815 5636 -15781
rect 5670 -15815 5682 -15781
rect 5624 -15849 5682 -15815
rect 5624 -15883 5636 -15849
rect 5670 -15883 5682 -15849
rect 5624 -15917 5682 -15883
rect 5624 -15951 5636 -15917
rect 5670 -15951 5682 -15917
rect 5624 -15985 5682 -15951
rect 5624 -16019 5636 -15985
rect 5670 -16019 5682 -15985
rect 5624 -16064 5682 -16019
rect 6642 -15509 6700 -15464
rect 6642 -15543 6654 -15509
rect 6688 -15543 6700 -15509
rect 6642 -15577 6700 -15543
rect 6642 -15611 6654 -15577
rect 6688 -15611 6700 -15577
rect 6642 -15645 6700 -15611
rect 6642 -15679 6654 -15645
rect 6688 -15679 6700 -15645
rect 6642 -15713 6700 -15679
rect 6642 -15747 6654 -15713
rect 6688 -15747 6700 -15713
rect 6642 -15781 6700 -15747
rect 6642 -15815 6654 -15781
rect 6688 -15815 6700 -15781
rect 6642 -15849 6700 -15815
rect 6642 -15883 6654 -15849
rect 6688 -15883 6700 -15849
rect 6642 -15917 6700 -15883
rect 6642 -15951 6654 -15917
rect 6688 -15951 6700 -15917
rect 6642 -15985 6700 -15951
rect 6642 -16019 6654 -15985
rect 6688 -16019 6700 -15985
rect 6642 -16064 6700 -16019
rect 7660 -15509 7718 -15464
rect 7660 -15543 7672 -15509
rect 7706 -15543 7718 -15509
rect 7660 -15577 7718 -15543
rect 7660 -15611 7672 -15577
rect 7706 -15611 7718 -15577
rect 7660 -15645 7718 -15611
rect 7660 -15679 7672 -15645
rect 7706 -15679 7718 -15645
rect 7660 -15713 7718 -15679
rect 7660 -15747 7672 -15713
rect 7706 -15747 7718 -15713
rect 7660 -15781 7718 -15747
rect 7660 -15815 7672 -15781
rect 7706 -15815 7718 -15781
rect 7660 -15849 7718 -15815
rect 7660 -15883 7672 -15849
rect 7706 -15883 7718 -15849
rect 7660 -15917 7718 -15883
rect 7660 -15951 7672 -15917
rect 7706 -15951 7718 -15917
rect 7660 -15985 7718 -15951
rect 7660 -16019 7672 -15985
rect 7706 -16019 7718 -15985
rect 7660 -16064 7718 -16019
rect 8678 -15509 8736 -15464
rect 8678 -15543 8690 -15509
rect 8724 -15543 8736 -15509
rect 8678 -15577 8736 -15543
rect 8678 -15611 8690 -15577
rect 8724 -15611 8736 -15577
rect 8678 -15645 8736 -15611
rect 8678 -15679 8690 -15645
rect 8724 -15679 8736 -15645
rect 8678 -15713 8736 -15679
rect 8678 -15747 8690 -15713
rect 8724 -15747 8736 -15713
rect 8678 -15781 8736 -15747
rect 8678 -15815 8690 -15781
rect 8724 -15815 8736 -15781
rect 8678 -15849 8736 -15815
rect 8678 -15883 8690 -15849
rect 8724 -15883 8736 -15849
rect 8678 -15917 8736 -15883
rect 8678 -15951 8690 -15917
rect 8724 -15951 8736 -15917
rect 8678 -15985 8736 -15951
rect 8678 -16019 8690 -15985
rect 8724 -16019 8736 -15985
rect 8678 -16064 8736 -16019
rect 9696 -15509 9754 -15464
rect 9696 -15543 9708 -15509
rect 9742 -15543 9754 -15509
rect 9696 -15577 9754 -15543
rect 9696 -15611 9708 -15577
rect 9742 -15611 9754 -15577
rect 9696 -15645 9754 -15611
rect 9696 -15679 9708 -15645
rect 9742 -15679 9754 -15645
rect 9696 -15713 9754 -15679
rect 9696 -15747 9708 -15713
rect 9742 -15747 9754 -15713
rect 9696 -15781 9754 -15747
rect 9696 -15815 9708 -15781
rect 9742 -15815 9754 -15781
rect 9696 -15849 9754 -15815
rect 9696 -15883 9708 -15849
rect 9742 -15883 9754 -15849
rect 9696 -15917 9754 -15883
rect 9696 -15951 9708 -15917
rect 9742 -15951 9754 -15917
rect 9696 -15985 9754 -15951
rect 9696 -16019 9708 -15985
rect 9742 -16019 9754 -15985
rect 9696 -16064 9754 -16019
rect 10714 -15509 10772 -15464
rect 10714 -15543 10726 -15509
rect 10760 -15543 10772 -15509
rect 10714 -15577 10772 -15543
rect 10714 -15611 10726 -15577
rect 10760 -15611 10772 -15577
rect 10714 -15645 10772 -15611
rect 10714 -15679 10726 -15645
rect 10760 -15679 10772 -15645
rect 10714 -15713 10772 -15679
rect 10714 -15747 10726 -15713
rect 10760 -15747 10772 -15713
rect 10714 -15781 10772 -15747
rect 10714 -15815 10726 -15781
rect 10760 -15815 10772 -15781
rect 10714 -15849 10772 -15815
rect 10714 -15883 10726 -15849
rect 10760 -15883 10772 -15849
rect 10714 -15917 10772 -15883
rect 10714 -15951 10726 -15917
rect 10760 -15951 10772 -15917
rect 10714 -15985 10772 -15951
rect 10714 -16019 10726 -15985
rect 10760 -16019 10772 -15985
rect 10714 -16064 10772 -16019
rect 11732 -15509 11790 -15464
rect 11732 -15543 11744 -15509
rect 11778 -15543 11790 -15509
rect 11732 -15577 11790 -15543
rect 11732 -15611 11744 -15577
rect 11778 -15611 11790 -15577
rect 11732 -15645 11790 -15611
rect 11732 -15679 11744 -15645
rect 11778 -15679 11790 -15645
rect 11732 -15713 11790 -15679
rect 11732 -15747 11744 -15713
rect 11778 -15747 11790 -15713
rect 11732 -15781 11790 -15747
rect 11732 -15815 11744 -15781
rect 11778 -15815 11790 -15781
rect 11732 -15849 11790 -15815
rect 11732 -15883 11744 -15849
rect 11778 -15883 11790 -15849
rect 11732 -15917 11790 -15883
rect 11732 -15951 11744 -15917
rect 11778 -15951 11790 -15917
rect 11732 -15985 11790 -15951
rect 11732 -16019 11744 -15985
rect 11778 -16019 11790 -15985
rect 11732 -16064 11790 -16019
rect 12750 -15509 12808 -15464
rect 12750 -15543 12762 -15509
rect 12796 -15543 12808 -15509
rect 12750 -15577 12808 -15543
rect 12750 -15611 12762 -15577
rect 12796 -15611 12808 -15577
rect 12750 -15645 12808 -15611
rect 12750 -15679 12762 -15645
rect 12796 -15679 12808 -15645
rect 12750 -15713 12808 -15679
rect 12750 -15747 12762 -15713
rect 12796 -15747 12808 -15713
rect 12750 -15781 12808 -15747
rect 12750 -15815 12762 -15781
rect 12796 -15815 12808 -15781
rect 12750 -15849 12808 -15815
rect 12750 -15883 12762 -15849
rect 12796 -15883 12808 -15849
rect 12750 -15917 12808 -15883
rect 12750 -15951 12762 -15917
rect 12796 -15951 12808 -15917
rect 12750 -15985 12808 -15951
rect 12750 -16019 12762 -15985
rect 12796 -16019 12808 -15985
rect 12750 -16064 12808 -16019
rect 13768 -15509 13826 -15464
rect 13768 -15543 13780 -15509
rect 13814 -15543 13826 -15509
rect 13768 -15577 13826 -15543
rect 13768 -15611 13780 -15577
rect 13814 -15611 13826 -15577
rect 13768 -15645 13826 -15611
rect 13768 -15679 13780 -15645
rect 13814 -15679 13826 -15645
rect 13768 -15713 13826 -15679
rect 13768 -15747 13780 -15713
rect 13814 -15747 13826 -15713
rect 13768 -15781 13826 -15747
rect 13768 -15815 13780 -15781
rect 13814 -15815 13826 -15781
rect 13768 -15849 13826 -15815
rect 13768 -15883 13780 -15849
rect 13814 -15883 13826 -15849
rect 13768 -15917 13826 -15883
rect 13768 -15951 13780 -15917
rect 13814 -15951 13826 -15917
rect 13768 -15985 13826 -15951
rect 13768 -16019 13780 -15985
rect 13814 -16019 13826 -15985
rect 13768 -16064 13826 -16019
rect 14786 -15509 14844 -15464
rect 14786 -15543 14798 -15509
rect 14832 -15543 14844 -15509
rect 14786 -15577 14844 -15543
rect 14786 -15611 14798 -15577
rect 14832 -15611 14844 -15577
rect 14786 -15645 14844 -15611
rect 14786 -15679 14798 -15645
rect 14832 -15679 14844 -15645
rect 14786 -15713 14844 -15679
rect 14786 -15747 14798 -15713
rect 14832 -15747 14844 -15713
rect 14786 -15781 14844 -15747
rect 14786 -15815 14798 -15781
rect 14832 -15815 14844 -15781
rect 14786 -15849 14844 -15815
rect 14786 -15883 14798 -15849
rect 14832 -15883 14844 -15849
rect 14786 -15917 14844 -15883
rect 14786 -15951 14798 -15917
rect 14832 -15951 14844 -15917
rect 14786 -15985 14844 -15951
rect 14786 -16019 14798 -15985
rect 14832 -16019 14844 -15985
rect 14786 -16064 14844 -16019
rect 15804 -15509 15862 -15464
rect 15804 -15543 15816 -15509
rect 15850 -15543 15862 -15509
rect 15804 -15577 15862 -15543
rect 15804 -15611 15816 -15577
rect 15850 -15611 15862 -15577
rect 15804 -15645 15862 -15611
rect 15804 -15679 15816 -15645
rect 15850 -15679 15862 -15645
rect 15804 -15713 15862 -15679
rect 15804 -15747 15816 -15713
rect 15850 -15747 15862 -15713
rect 15804 -15781 15862 -15747
rect 15804 -15815 15816 -15781
rect 15850 -15815 15862 -15781
rect 15804 -15849 15862 -15815
rect 15804 -15883 15816 -15849
rect 15850 -15883 15862 -15849
rect 15804 -15917 15862 -15883
rect 15804 -15951 15816 -15917
rect 15850 -15951 15862 -15917
rect 15804 -15985 15862 -15951
rect 15804 -16019 15816 -15985
rect 15850 -16019 15862 -15985
rect 15804 -16064 15862 -16019
rect 16822 -15509 16880 -15464
rect 16822 -15543 16834 -15509
rect 16868 -15543 16880 -15509
rect 16822 -15577 16880 -15543
rect 16822 -15611 16834 -15577
rect 16868 -15611 16880 -15577
rect 16822 -15645 16880 -15611
rect 16822 -15679 16834 -15645
rect 16868 -15679 16880 -15645
rect 16822 -15713 16880 -15679
rect 16822 -15747 16834 -15713
rect 16868 -15747 16880 -15713
rect 16822 -15781 16880 -15747
rect 16822 -15815 16834 -15781
rect 16868 -15815 16880 -15781
rect 16822 -15849 16880 -15815
rect 16822 -15883 16834 -15849
rect 16868 -15883 16880 -15849
rect 16822 -15917 16880 -15883
rect 16822 -15951 16834 -15917
rect 16868 -15951 16880 -15917
rect 16822 -15985 16880 -15951
rect 16822 -16019 16834 -15985
rect 16868 -16019 16880 -15985
rect 16822 -16064 16880 -16019
rect 17840 -15509 17898 -15464
rect 17840 -15543 17852 -15509
rect 17886 -15543 17898 -15509
rect 17840 -15577 17898 -15543
rect 17840 -15611 17852 -15577
rect 17886 -15611 17898 -15577
rect 17840 -15645 17898 -15611
rect 17840 -15679 17852 -15645
rect 17886 -15679 17898 -15645
rect 17840 -15713 17898 -15679
rect 17840 -15747 17852 -15713
rect 17886 -15747 17898 -15713
rect 17840 -15781 17898 -15747
rect 17840 -15815 17852 -15781
rect 17886 -15815 17898 -15781
rect 17840 -15849 17898 -15815
rect 17840 -15883 17852 -15849
rect 17886 -15883 17898 -15849
rect 17840 -15917 17898 -15883
rect 17840 -15951 17852 -15917
rect 17886 -15951 17898 -15917
rect 17840 -15985 17898 -15951
rect 17840 -16019 17852 -15985
rect 17886 -16019 17898 -15985
rect 17840 -16064 17898 -16019
rect 18858 -15509 18916 -15464
rect 18858 -15543 18870 -15509
rect 18904 -15543 18916 -15509
rect 18858 -15577 18916 -15543
rect 18858 -15611 18870 -15577
rect 18904 -15611 18916 -15577
rect 18858 -15645 18916 -15611
rect 18858 -15679 18870 -15645
rect 18904 -15679 18916 -15645
rect 18858 -15713 18916 -15679
rect 18858 -15747 18870 -15713
rect 18904 -15747 18916 -15713
rect 18858 -15781 18916 -15747
rect 18858 -15815 18870 -15781
rect 18904 -15815 18916 -15781
rect 18858 -15849 18916 -15815
rect 18858 -15883 18870 -15849
rect 18904 -15883 18916 -15849
rect 18858 -15917 18916 -15883
rect 18858 -15951 18870 -15917
rect 18904 -15951 18916 -15917
rect 18858 -15985 18916 -15951
rect 18858 -16019 18870 -15985
rect 18904 -16019 18916 -15985
rect 18858 -16064 18916 -16019
rect 19876 -15509 19934 -15464
rect 19876 -15543 19888 -15509
rect 19922 -15543 19934 -15509
rect 19876 -15577 19934 -15543
rect 19876 -15611 19888 -15577
rect 19922 -15611 19934 -15577
rect 19876 -15645 19934 -15611
rect 19876 -15679 19888 -15645
rect 19922 -15679 19934 -15645
rect 19876 -15713 19934 -15679
rect 19876 -15747 19888 -15713
rect 19922 -15747 19934 -15713
rect 19876 -15781 19934 -15747
rect 19876 -15815 19888 -15781
rect 19922 -15815 19934 -15781
rect 19876 -15849 19934 -15815
rect 19876 -15883 19888 -15849
rect 19922 -15883 19934 -15849
rect 19876 -15917 19934 -15883
rect 19876 -15951 19888 -15917
rect 19922 -15951 19934 -15917
rect 19876 -15985 19934 -15951
rect 19876 -16019 19888 -15985
rect 19922 -16019 19934 -15985
rect 19876 -16064 19934 -16019
rect 20894 -15509 20952 -15464
rect 20894 -15543 20906 -15509
rect 20940 -15543 20952 -15509
rect 20894 -15577 20952 -15543
rect 20894 -15611 20906 -15577
rect 20940 -15611 20952 -15577
rect 20894 -15645 20952 -15611
rect 20894 -15679 20906 -15645
rect 20940 -15679 20952 -15645
rect 20894 -15713 20952 -15679
rect 20894 -15747 20906 -15713
rect 20940 -15747 20952 -15713
rect 20894 -15781 20952 -15747
rect 20894 -15815 20906 -15781
rect 20940 -15815 20952 -15781
rect 20894 -15849 20952 -15815
rect 20894 -15883 20906 -15849
rect 20940 -15883 20952 -15849
rect 20894 -15917 20952 -15883
rect 20894 -15951 20906 -15917
rect 20940 -15951 20952 -15917
rect 20894 -15985 20952 -15951
rect 20894 -16019 20906 -15985
rect 20940 -16019 20952 -15985
rect 20894 -16064 20952 -16019
rect 21912 -15509 21970 -15464
rect 21912 -15543 21924 -15509
rect 21958 -15543 21970 -15509
rect 21912 -15577 21970 -15543
rect 21912 -15611 21924 -15577
rect 21958 -15611 21970 -15577
rect 21912 -15645 21970 -15611
rect 21912 -15679 21924 -15645
rect 21958 -15679 21970 -15645
rect 21912 -15713 21970 -15679
rect 21912 -15747 21924 -15713
rect 21958 -15747 21970 -15713
rect 21912 -15781 21970 -15747
rect 21912 -15815 21924 -15781
rect 21958 -15815 21970 -15781
rect 21912 -15849 21970 -15815
rect 21912 -15883 21924 -15849
rect 21958 -15883 21970 -15849
rect 21912 -15917 21970 -15883
rect 21912 -15951 21924 -15917
rect 21958 -15951 21970 -15917
rect 21912 -15985 21970 -15951
rect 21912 -16019 21924 -15985
rect 21958 -16019 21970 -15985
rect 21912 -16064 21970 -16019
rect 22930 -15509 22988 -15464
rect 22930 -15543 22942 -15509
rect 22976 -15543 22988 -15509
rect 22930 -15577 22988 -15543
rect 22930 -15611 22942 -15577
rect 22976 -15611 22988 -15577
rect 22930 -15645 22988 -15611
rect 22930 -15679 22942 -15645
rect 22976 -15679 22988 -15645
rect 22930 -15713 22988 -15679
rect 22930 -15747 22942 -15713
rect 22976 -15747 22988 -15713
rect 22930 -15781 22988 -15747
rect 22930 -15815 22942 -15781
rect 22976 -15815 22988 -15781
rect 22930 -15849 22988 -15815
rect 22930 -15883 22942 -15849
rect 22976 -15883 22988 -15849
rect 22930 -15917 22988 -15883
rect 22930 -15951 22942 -15917
rect 22976 -15951 22988 -15917
rect 22930 -15985 22988 -15951
rect 22930 -16019 22942 -15985
rect 22976 -16019 22988 -15985
rect 22930 -16064 22988 -16019
rect -34 -16101 24 -16067
rect -34 -16135 -22 -16101
rect 12 -16135 24 -16101
rect -34 -16169 24 -16135
rect -34 -16203 -22 -16169
rect 12 -16203 24 -16169
rect -34 -16237 24 -16203
rect -34 -16271 -22 -16237
rect 12 -16271 24 -16237
rect -34 -16305 24 -16271
rect -34 -16339 -22 -16305
rect 12 -16339 24 -16305
rect -34 -16384 24 -16339
rect -9196 -16647 -9138 -16602
rect -9196 -16681 -9184 -16647
rect -9150 -16681 -9138 -16647
rect -9196 -16715 -9138 -16681
rect -9196 -16749 -9184 -16715
rect -9150 -16749 -9138 -16715
rect -9196 -16783 -9138 -16749
rect -9196 -16817 -9184 -16783
rect -9150 -16817 -9138 -16783
rect -9196 -16851 -9138 -16817
rect -9196 -16885 -9184 -16851
rect -9150 -16885 -9138 -16851
rect -9196 -16919 -9138 -16885
rect -9196 -16953 -9184 -16919
rect -9150 -16953 -9138 -16919
rect -9196 -16987 -9138 -16953
rect -9196 -17021 -9184 -16987
rect -9150 -17021 -9138 -16987
rect -9196 -17055 -9138 -17021
rect -9196 -17089 -9184 -17055
rect -9150 -17089 -9138 -17055
rect -9196 -17123 -9138 -17089
rect -9196 -17157 -9184 -17123
rect -9150 -17157 -9138 -17123
rect -9196 -17202 -9138 -17157
rect -8178 -16647 -8120 -16602
rect -8178 -16681 -8166 -16647
rect -8132 -16681 -8120 -16647
rect -8178 -16715 -8120 -16681
rect -8178 -16749 -8166 -16715
rect -8132 -16749 -8120 -16715
rect -8178 -16783 -8120 -16749
rect -8178 -16817 -8166 -16783
rect -8132 -16817 -8120 -16783
rect -8178 -16851 -8120 -16817
rect -8178 -16885 -8166 -16851
rect -8132 -16885 -8120 -16851
rect -8178 -16919 -8120 -16885
rect -8178 -16953 -8166 -16919
rect -8132 -16953 -8120 -16919
rect -8178 -16987 -8120 -16953
rect -8178 -17021 -8166 -16987
rect -8132 -17021 -8120 -16987
rect -8178 -17055 -8120 -17021
rect -8178 -17089 -8166 -17055
rect -8132 -17089 -8120 -17055
rect -8178 -17123 -8120 -17089
rect -8178 -17157 -8166 -17123
rect -8132 -17157 -8120 -17123
rect -8178 -17202 -8120 -17157
rect -7160 -16647 -7102 -16602
rect -7160 -16681 -7148 -16647
rect -7114 -16681 -7102 -16647
rect -7160 -16715 -7102 -16681
rect -7160 -16749 -7148 -16715
rect -7114 -16749 -7102 -16715
rect -7160 -16783 -7102 -16749
rect -7160 -16817 -7148 -16783
rect -7114 -16817 -7102 -16783
rect -7160 -16851 -7102 -16817
rect -7160 -16885 -7148 -16851
rect -7114 -16885 -7102 -16851
rect -7160 -16919 -7102 -16885
rect -7160 -16953 -7148 -16919
rect -7114 -16953 -7102 -16919
rect -7160 -16987 -7102 -16953
rect -7160 -17021 -7148 -16987
rect -7114 -17021 -7102 -16987
rect -7160 -17055 -7102 -17021
rect -7160 -17089 -7148 -17055
rect -7114 -17089 -7102 -17055
rect -7160 -17123 -7102 -17089
rect -7160 -17157 -7148 -17123
rect -7114 -17157 -7102 -17123
rect -7160 -17202 -7102 -17157
rect -6142 -16647 -6084 -16602
rect -6142 -16681 -6130 -16647
rect -6096 -16681 -6084 -16647
rect -6142 -16715 -6084 -16681
rect -6142 -16749 -6130 -16715
rect -6096 -16749 -6084 -16715
rect -6142 -16783 -6084 -16749
rect -6142 -16817 -6130 -16783
rect -6096 -16817 -6084 -16783
rect -6142 -16851 -6084 -16817
rect -6142 -16885 -6130 -16851
rect -6096 -16885 -6084 -16851
rect -6142 -16919 -6084 -16885
rect -6142 -16953 -6130 -16919
rect -6096 -16953 -6084 -16919
rect -6142 -16987 -6084 -16953
rect -6142 -17021 -6130 -16987
rect -6096 -17021 -6084 -16987
rect -6142 -17055 -6084 -17021
rect -6142 -17089 -6130 -17055
rect -6096 -17089 -6084 -17055
rect -6142 -17123 -6084 -17089
rect -6142 -17157 -6130 -17123
rect -6096 -17157 -6084 -17123
rect -6142 -17202 -6084 -17157
rect -5124 -16647 -5066 -16602
rect -5124 -16681 -5112 -16647
rect -5078 -16681 -5066 -16647
rect -5124 -16715 -5066 -16681
rect -5124 -16749 -5112 -16715
rect -5078 -16749 -5066 -16715
rect -5124 -16783 -5066 -16749
rect -5124 -16817 -5112 -16783
rect -5078 -16817 -5066 -16783
rect -5124 -16851 -5066 -16817
rect -5124 -16885 -5112 -16851
rect -5078 -16885 -5066 -16851
rect -5124 -16919 -5066 -16885
rect -5124 -16953 -5112 -16919
rect -5078 -16953 -5066 -16919
rect -5124 -16987 -5066 -16953
rect -5124 -17021 -5112 -16987
rect -5078 -17021 -5066 -16987
rect -5124 -17055 -5066 -17021
rect -5124 -17089 -5112 -17055
rect -5078 -17089 -5066 -17055
rect -5124 -17123 -5066 -17089
rect -5124 -17157 -5112 -17123
rect -5078 -17157 -5066 -17123
rect -5124 -17202 -5066 -17157
rect -4106 -16647 -4048 -16602
rect -4106 -16681 -4094 -16647
rect -4060 -16681 -4048 -16647
rect -4106 -16715 -4048 -16681
rect -4106 -16749 -4094 -16715
rect -4060 -16749 -4048 -16715
rect -4106 -16783 -4048 -16749
rect -4106 -16817 -4094 -16783
rect -4060 -16817 -4048 -16783
rect -4106 -16851 -4048 -16817
rect -4106 -16885 -4094 -16851
rect -4060 -16885 -4048 -16851
rect -4106 -16919 -4048 -16885
rect -4106 -16953 -4094 -16919
rect -4060 -16953 -4048 -16919
rect -4106 -16987 -4048 -16953
rect -4106 -17021 -4094 -16987
rect -4060 -17021 -4048 -16987
rect -4106 -17055 -4048 -17021
rect -4106 -17089 -4094 -17055
rect -4060 -17089 -4048 -17055
rect -4106 -17123 -4048 -17089
rect -4106 -17157 -4094 -17123
rect -4060 -17157 -4048 -17123
rect -4106 -17202 -4048 -17157
rect -3088 -16647 -3030 -16602
rect -3088 -16681 -3076 -16647
rect -3042 -16681 -3030 -16647
rect -3088 -16715 -3030 -16681
rect -3088 -16749 -3076 -16715
rect -3042 -16749 -3030 -16715
rect -3088 -16783 -3030 -16749
rect -3088 -16817 -3076 -16783
rect -3042 -16817 -3030 -16783
rect -3088 -16851 -3030 -16817
rect -3088 -16885 -3076 -16851
rect -3042 -16885 -3030 -16851
rect -3088 -16919 -3030 -16885
rect -3088 -16953 -3076 -16919
rect -3042 -16953 -3030 -16919
rect -3088 -16987 -3030 -16953
rect -3088 -17021 -3076 -16987
rect -3042 -17021 -3030 -16987
rect -3088 -17055 -3030 -17021
rect -3088 -17089 -3076 -17055
rect -3042 -17089 -3030 -17055
rect -3088 -17123 -3030 -17089
rect -3088 -17157 -3076 -17123
rect -3042 -17157 -3030 -17123
rect -3088 -17202 -3030 -17157
rect -2070 -16647 -2012 -16602
rect -2070 -16681 -2058 -16647
rect -2024 -16681 -2012 -16647
rect -2070 -16715 -2012 -16681
rect -2070 -16749 -2058 -16715
rect -2024 -16749 -2012 -16715
rect -2070 -16783 -2012 -16749
rect -2070 -16817 -2058 -16783
rect -2024 -16817 -2012 -16783
rect -2070 -16851 -2012 -16817
rect -2070 -16885 -2058 -16851
rect -2024 -16885 -2012 -16851
rect -2070 -16919 -2012 -16885
rect -2070 -16953 -2058 -16919
rect -2024 -16953 -2012 -16919
rect -2070 -16987 -2012 -16953
rect -2070 -17021 -2058 -16987
rect -2024 -17021 -2012 -16987
rect -2070 -17055 -2012 -17021
rect -2070 -17089 -2058 -17055
rect -2024 -17089 -2012 -17055
rect -2070 -17123 -2012 -17089
rect -2070 -17157 -2058 -17123
rect -2024 -17157 -2012 -17123
rect -2070 -17202 -2012 -17157
rect -1052 -16647 -994 -16602
rect -1052 -16681 -1040 -16647
rect -1006 -16681 -994 -16647
rect -1052 -16715 -994 -16681
rect -1052 -16749 -1040 -16715
rect -1006 -16749 -994 -16715
rect -1052 -16783 -994 -16749
rect -1052 -16817 -1040 -16783
rect -1006 -16817 -994 -16783
rect -1052 -16851 -994 -16817
rect -1052 -16885 -1040 -16851
rect -1006 -16885 -994 -16851
rect -1052 -16919 -994 -16885
rect -1052 -16953 -1040 -16919
rect -1006 -16953 -994 -16919
rect -1052 -16987 -994 -16953
rect -1052 -17021 -1040 -16987
rect -1006 -17021 -994 -16987
rect -1052 -17055 -994 -17021
rect -1052 -17089 -1040 -17055
rect -1006 -17089 -994 -17055
rect -1052 -17123 -994 -17089
rect -1052 -17157 -1040 -17123
rect -1006 -17157 -994 -17123
rect -1052 -17202 -994 -17157
rect -34 -16647 24 -16602
rect -34 -16681 -22 -16647
rect 12 -16681 24 -16647
rect -34 -16715 24 -16681
rect -34 -16749 -22 -16715
rect 12 -16749 24 -16715
rect -34 -16783 24 -16749
rect -34 -16817 -22 -16783
rect 12 -16817 24 -16783
rect -34 -16851 24 -16817
rect -34 -16885 -22 -16851
rect 12 -16885 24 -16851
rect -34 -16919 24 -16885
rect -34 -16953 -22 -16919
rect 12 -16953 24 -16919
rect -34 -16987 24 -16953
rect -34 -17021 -22 -16987
rect 12 -17021 24 -16987
rect -34 -17055 24 -17021
rect -34 -17089 -22 -17055
rect 12 -17089 24 -17055
rect -34 -17123 24 -17089
rect -34 -17157 -22 -17123
rect 12 -17157 24 -17123
rect -34 -17202 24 -17157
rect 2568 -16743 2626 -16698
rect 2568 -16777 2580 -16743
rect 2614 -16777 2626 -16743
rect 2568 -16811 2626 -16777
rect 2568 -16845 2580 -16811
rect 2614 -16845 2626 -16811
rect 2568 -16879 2626 -16845
rect 2568 -16913 2580 -16879
rect 2614 -16913 2626 -16879
rect 2568 -16947 2626 -16913
rect 2568 -16981 2580 -16947
rect 2614 -16981 2626 -16947
rect 2568 -17015 2626 -16981
rect 2568 -17049 2580 -17015
rect 2614 -17049 2626 -17015
rect 2568 -17083 2626 -17049
rect 2568 -17117 2580 -17083
rect 2614 -17117 2626 -17083
rect 2568 -17151 2626 -17117
rect 2568 -17185 2580 -17151
rect 2614 -17185 2626 -17151
rect 2568 -17219 2626 -17185
rect 2568 -17253 2580 -17219
rect 2614 -17253 2626 -17219
rect 2568 -17298 2626 -17253
rect 3586 -16743 3644 -16698
rect 3586 -16777 3598 -16743
rect 3632 -16777 3644 -16743
rect 3586 -16811 3644 -16777
rect 3586 -16845 3598 -16811
rect 3632 -16845 3644 -16811
rect 3586 -16879 3644 -16845
rect 3586 -16913 3598 -16879
rect 3632 -16913 3644 -16879
rect 3586 -16947 3644 -16913
rect 3586 -16981 3598 -16947
rect 3632 -16981 3644 -16947
rect 3586 -17015 3644 -16981
rect 3586 -17049 3598 -17015
rect 3632 -17049 3644 -17015
rect 3586 -17083 3644 -17049
rect 3586 -17117 3598 -17083
rect 3632 -17117 3644 -17083
rect 3586 -17151 3644 -17117
rect 3586 -17185 3598 -17151
rect 3632 -17185 3644 -17151
rect 3586 -17219 3644 -17185
rect 3586 -17253 3598 -17219
rect 3632 -17253 3644 -17219
rect 3586 -17298 3644 -17253
rect 4604 -16743 4662 -16698
rect 4604 -16777 4616 -16743
rect 4650 -16777 4662 -16743
rect 4604 -16811 4662 -16777
rect 4604 -16845 4616 -16811
rect 4650 -16845 4662 -16811
rect 4604 -16879 4662 -16845
rect 4604 -16913 4616 -16879
rect 4650 -16913 4662 -16879
rect 4604 -16947 4662 -16913
rect 4604 -16981 4616 -16947
rect 4650 -16981 4662 -16947
rect 4604 -17015 4662 -16981
rect 4604 -17049 4616 -17015
rect 4650 -17049 4662 -17015
rect 4604 -17083 4662 -17049
rect 4604 -17117 4616 -17083
rect 4650 -17117 4662 -17083
rect 4604 -17151 4662 -17117
rect 4604 -17185 4616 -17151
rect 4650 -17185 4662 -17151
rect 4604 -17219 4662 -17185
rect 4604 -17253 4616 -17219
rect 4650 -17253 4662 -17219
rect 4604 -17298 4662 -17253
rect 5622 -16743 5680 -16698
rect 5622 -16777 5634 -16743
rect 5668 -16777 5680 -16743
rect 5622 -16811 5680 -16777
rect 5622 -16845 5634 -16811
rect 5668 -16845 5680 -16811
rect 5622 -16879 5680 -16845
rect 5622 -16913 5634 -16879
rect 5668 -16913 5680 -16879
rect 5622 -16947 5680 -16913
rect 5622 -16981 5634 -16947
rect 5668 -16981 5680 -16947
rect 5622 -17015 5680 -16981
rect 5622 -17049 5634 -17015
rect 5668 -17049 5680 -17015
rect 5622 -17083 5680 -17049
rect 5622 -17117 5634 -17083
rect 5668 -17117 5680 -17083
rect 5622 -17151 5680 -17117
rect 5622 -17185 5634 -17151
rect 5668 -17185 5680 -17151
rect 5622 -17219 5680 -17185
rect 5622 -17253 5634 -17219
rect 5668 -17253 5680 -17219
rect 5622 -17298 5680 -17253
rect 6640 -16743 6698 -16698
rect 6640 -16777 6652 -16743
rect 6686 -16777 6698 -16743
rect 6640 -16811 6698 -16777
rect 6640 -16845 6652 -16811
rect 6686 -16845 6698 -16811
rect 6640 -16879 6698 -16845
rect 6640 -16913 6652 -16879
rect 6686 -16913 6698 -16879
rect 6640 -16947 6698 -16913
rect 6640 -16981 6652 -16947
rect 6686 -16981 6698 -16947
rect 6640 -17015 6698 -16981
rect 6640 -17049 6652 -17015
rect 6686 -17049 6698 -17015
rect 6640 -17083 6698 -17049
rect 6640 -17117 6652 -17083
rect 6686 -17117 6698 -17083
rect 6640 -17151 6698 -17117
rect 6640 -17185 6652 -17151
rect 6686 -17185 6698 -17151
rect 6640 -17219 6698 -17185
rect 6640 -17253 6652 -17219
rect 6686 -17253 6698 -17219
rect 6640 -17298 6698 -17253
rect 7658 -16743 7716 -16698
rect 7658 -16777 7670 -16743
rect 7704 -16777 7716 -16743
rect 7658 -16811 7716 -16777
rect 7658 -16845 7670 -16811
rect 7704 -16845 7716 -16811
rect 7658 -16879 7716 -16845
rect 7658 -16913 7670 -16879
rect 7704 -16913 7716 -16879
rect 7658 -16947 7716 -16913
rect 7658 -16981 7670 -16947
rect 7704 -16981 7716 -16947
rect 7658 -17015 7716 -16981
rect 7658 -17049 7670 -17015
rect 7704 -17049 7716 -17015
rect 7658 -17083 7716 -17049
rect 7658 -17117 7670 -17083
rect 7704 -17117 7716 -17083
rect 7658 -17151 7716 -17117
rect 7658 -17185 7670 -17151
rect 7704 -17185 7716 -17151
rect 7658 -17219 7716 -17185
rect 7658 -17253 7670 -17219
rect 7704 -17253 7716 -17219
rect 7658 -17298 7716 -17253
rect 8676 -16743 8734 -16698
rect 8676 -16777 8688 -16743
rect 8722 -16777 8734 -16743
rect 8676 -16811 8734 -16777
rect 8676 -16845 8688 -16811
rect 8722 -16845 8734 -16811
rect 8676 -16879 8734 -16845
rect 8676 -16913 8688 -16879
rect 8722 -16913 8734 -16879
rect 8676 -16947 8734 -16913
rect 8676 -16981 8688 -16947
rect 8722 -16981 8734 -16947
rect 8676 -17015 8734 -16981
rect 8676 -17049 8688 -17015
rect 8722 -17049 8734 -17015
rect 8676 -17083 8734 -17049
rect 8676 -17117 8688 -17083
rect 8722 -17117 8734 -17083
rect 8676 -17151 8734 -17117
rect 8676 -17185 8688 -17151
rect 8722 -17185 8734 -17151
rect 8676 -17219 8734 -17185
rect 8676 -17253 8688 -17219
rect 8722 -17253 8734 -17219
rect 8676 -17298 8734 -17253
rect 9694 -16743 9752 -16698
rect 9694 -16777 9706 -16743
rect 9740 -16777 9752 -16743
rect 9694 -16811 9752 -16777
rect 9694 -16845 9706 -16811
rect 9740 -16845 9752 -16811
rect 9694 -16879 9752 -16845
rect 9694 -16913 9706 -16879
rect 9740 -16913 9752 -16879
rect 9694 -16947 9752 -16913
rect 9694 -16981 9706 -16947
rect 9740 -16981 9752 -16947
rect 9694 -17015 9752 -16981
rect 9694 -17049 9706 -17015
rect 9740 -17049 9752 -17015
rect 9694 -17083 9752 -17049
rect 9694 -17117 9706 -17083
rect 9740 -17117 9752 -17083
rect 9694 -17151 9752 -17117
rect 9694 -17185 9706 -17151
rect 9740 -17185 9752 -17151
rect 9694 -17219 9752 -17185
rect 9694 -17253 9706 -17219
rect 9740 -17253 9752 -17219
rect 9694 -17298 9752 -17253
rect 10712 -16743 10770 -16698
rect 10712 -16777 10724 -16743
rect 10758 -16777 10770 -16743
rect 10712 -16811 10770 -16777
rect 10712 -16845 10724 -16811
rect 10758 -16845 10770 -16811
rect 10712 -16879 10770 -16845
rect 10712 -16913 10724 -16879
rect 10758 -16913 10770 -16879
rect 10712 -16947 10770 -16913
rect 10712 -16981 10724 -16947
rect 10758 -16981 10770 -16947
rect 10712 -17015 10770 -16981
rect 10712 -17049 10724 -17015
rect 10758 -17049 10770 -17015
rect 10712 -17083 10770 -17049
rect 10712 -17117 10724 -17083
rect 10758 -17117 10770 -17083
rect 10712 -17151 10770 -17117
rect 10712 -17185 10724 -17151
rect 10758 -17185 10770 -17151
rect 10712 -17219 10770 -17185
rect 10712 -17253 10724 -17219
rect 10758 -17253 10770 -17219
rect 10712 -17298 10770 -17253
rect 11730 -16743 11788 -16698
rect 11730 -16777 11742 -16743
rect 11776 -16777 11788 -16743
rect 11730 -16811 11788 -16777
rect 11730 -16845 11742 -16811
rect 11776 -16845 11788 -16811
rect 11730 -16879 11788 -16845
rect 11730 -16913 11742 -16879
rect 11776 -16913 11788 -16879
rect 11730 -16947 11788 -16913
rect 11730 -16981 11742 -16947
rect 11776 -16981 11788 -16947
rect 11730 -17015 11788 -16981
rect 11730 -17049 11742 -17015
rect 11776 -17049 11788 -17015
rect 11730 -17083 11788 -17049
rect 11730 -17117 11742 -17083
rect 11776 -17117 11788 -17083
rect 11730 -17151 11788 -17117
rect 11730 -17185 11742 -17151
rect 11776 -17185 11788 -17151
rect 11730 -17219 11788 -17185
rect 11730 -17253 11742 -17219
rect 11776 -17253 11788 -17219
rect 11730 -17298 11788 -17253
rect 12748 -16743 12806 -16698
rect 12748 -16777 12760 -16743
rect 12794 -16777 12806 -16743
rect 12748 -16811 12806 -16777
rect 12748 -16845 12760 -16811
rect 12794 -16845 12806 -16811
rect 12748 -16879 12806 -16845
rect 12748 -16913 12760 -16879
rect 12794 -16913 12806 -16879
rect 12748 -16947 12806 -16913
rect 12748 -16981 12760 -16947
rect 12794 -16981 12806 -16947
rect 12748 -17015 12806 -16981
rect 12748 -17049 12760 -17015
rect 12794 -17049 12806 -17015
rect 12748 -17083 12806 -17049
rect 12748 -17117 12760 -17083
rect 12794 -17117 12806 -17083
rect 12748 -17151 12806 -17117
rect 12748 -17185 12760 -17151
rect 12794 -17185 12806 -17151
rect 12748 -17219 12806 -17185
rect 12748 -17253 12760 -17219
rect 12794 -17253 12806 -17219
rect 12748 -17298 12806 -17253
rect 13766 -16743 13824 -16698
rect 13766 -16777 13778 -16743
rect 13812 -16777 13824 -16743
rect 13766 -16811 13824 -16777
rect 13766 -16845 13778 -16811
rect 13812 -16845 13824 -16811
rect 13766 -16879 13824 -16845
rect 13766 -16913 13778 -16879
rect 13812 -16913 13824 -16879
rect 13766 -16947 13824 -16913
rect 13766 -16981 13778 -16947
rect 13812 -16981 13824 -16947
rect 13766 -17015 13824 -16981
rect 13766 -17049 13778 -17015
rect 13812 -17049 13824 -17015
rect 13766 -17083 13824 -17049
rect 13766 -17117 13778 -17083
rect 13812 -17117 13824 -17083
rect 13766 -17151 13824 -17117
rect 13766 -17185 13778 -17151
rect 13812 -17185 13824 -17151
rect 13766 -17219 13824 -17185
rect 13766 -17253 13778 -17219
rect 13812 -17253 13824 -17219
rect 13766 -17298 13824 -17253
rect 14784 -16743 14842 -16698
rect 14784 -16777 14796 -16743
rect 14830 -16777 14842 -16743
rect 14784 -16811 14842 -16777
rect 14784 -16845 14796 -16811
rect 14830 -16845 14842 -16811
rect 14784 -16879 14842 -16845
rect 14784 -16913 14796 -16879
rect 14830 -16913 14842 -16879
rect 14784 -16947 14842 -16913
rect 14784 -16981 14796 -16947
rect 14830 -16981 14842 -16947
rect 14784 -17015 14842 -16981
rect 14784 -17049 14796 -17015
rect 14830 -17049 14842 -17015
rect 14784 -17083 14842 -17049
rect 14784 -17117 14796 -17083
rect 14830 -17117 14842 -17083
rect 14784 -17151 14842 -17117
rect 14784 -17185 14796 -17151
rect 14830 -17185 14842 -17151
rect 14784 -17219 14842 -17185
rect 14784 -17253 14796 -17219
rect 14830 -17253 14842 -17219
rect 14784 -17298 14842 -17253
rect 15802 -16743 15860 -16698
rect 15802 -16777 15814 -16743
rect 15848 -16777 15860 -16743
rect 15802 -16811 15860 -16777
rect 15802 -16845 15814 -16811
rect 15848 -16845 15860 -16811
rect 15802 -16879 15860 -16845
rect 15802 -16913 15814 -16879
rect 15848 -16913 15860 -16879
rect 15802 -16947 15860 -16913
rect 15802 -16981 15814 -16947
rect 15848 -16981 15860 -16947
rect 15802 -17015 15860 -16981
rect 15802 -17049 15814 -17015
rect 15848 -17049 15860 -17015
rect 15802 -17083 15860 -17049
rect 15802 -17117 15814 -17083
rect 15848 -17117 15860 -17083
rect 15802 -17151 15860 -17117
rect 15802 -17185 15814 -17151
rect 15848 -17185 15860 -17151
rect 15802 -17219 15860 -17185
rect 15802 -17253 15814 -17219
rect 15848 -17253 15860 -17219
rect 15802 -17298 15860 -17253
rect 16820 -16743 16878 -16698
rect 16820 -16777 16832 -16743
rect 16866 -16777 16878 -16743
rect 16820 -16811 16878 -16777
rect 16820 -16845 16832 -16811
rect 16866 -16845 16878 -16811
rect 16820 -16879 16878 -16845
rect 16820 -16913 16832 -16879
rect 16866 -16913 16878 -16879
rect 16820 -16947 16878 -16913
rect 16820 -16981 16832 -16947
rect 16866 -16981 16878 -16947
rect 16820 -17015 16878 -16981
rect 16820 -17049 16832 -17015
rect 16866 -17049 16878 -17015
rect 16820 -17083 16878 -17049
rect 16820 -17117 16832 -17083
rect 16866 -17117 16878 -17083
rect 16820 -17151 16878 -17117
rect 16820 -17185 16832 -17151
rect 16866 -17185 16878 -17151
rect 16820 -17219 16878 -17185
rect 16820 -17253 16832 -17219
rect 16866 -17253 16878 -17219
rect 16820 -17298 16878 -17253
rect 17838 -16743 17896 -16698
rect 17838 -16777 17850 -16743
rect 17884 -16777 17896 -16743
rect 17838 -16811 17896 -16777
rect 17838 -16845 17850 -16811
rect 17884 -16845 17896 -16811
rect 17838 -16879 17896 -16845
rect 17838 -16913 17850 -16879
rect 17884 -16913 17896 -16879
rect 17838 -16947 17896 -16913
rect 17838 -16981 17850 -16947
rect 17884 -16981 17896 -16947
rect 17838 -17015 17896 -16981
rect 17838 -17049 17850 -17015
rect 17884 -17049 17896 -17015
rect 17838 -17083 17896 -17049
rect 17838 -17117 17850 -17083
rect 17884 -17117 17896 -17083
rect 17838 -17151 17896 -17117
rect 17838 -17185 17850 -17151
rect 17884 -17185 17896 -17151
rect 17838 -17219 17896 -17185
rect 17838 -17253 17850 -17219
rect 17884 -17253 17896 -17219
rect 17838 -17298 17896 -17253
rect 18856 -16743 18914 -16698
rect 18856 -16777 18868 -16743
rect 18902 -16777 18914 -16743
rect 18856 -16811 18914 -16777
rect 18856 -16845 18868 -16811
rect 18902 -16845 18914 -16811
rect 18856 -16879 18914 -16845
rect 18856 -16913 18868 -16879
rect 18902 -16913 18914 -16879
rect 18856 -16947 18914 -16913
rect 18856 -16981 18868 -16947
rect 18902 -16981 18914 -16947
rect 18856 -17015 18914 -16981
rect 18856 -17049 18868 -17015
rect 18902 -17049 18914 -17015
rect 18856 -17083 18914 -17049
rect 18856 -17117 18868 -17083
rect 18902 -17117 18914 -17083
rect 18856 -17151 18914 -17117
rect 18856 -17185 18868 -17151
rect 18902 -17185 18914 -17151
rect 18856 -17219 18914 -17185
rect 18856 -17253 18868 -17219
rect 18902 -17253 18914 -17219
rect 18856 -17298 18914 -17253
rect 19874 -16743 19932 -16698
rect 19874 -16777 19886 -16743
rect 19920 -16777 19932 -16743
rect 19874 -16811 19932 -16777
rect 19874 -16845 19886 -16811
rect 19920 -16845 19932 -16811
rect 19874 -16879 19932 -16845
rect 19874 -16913 19886 -16879
rect 19920 -16913 19932 -16879
rect 19874 -16947 19932 -16913
rect 19874 -16981 19886 -16947
rect 19920 -16981 19932 -16947
rect 19874 -17015 19932 -16981
rect 19874 -17049 19886 -17015
rect 19920 -17049 19932 -17015
rect 19874 -17083 19932 -17049
rect 19874 -17117 19886 -17083
rect 19920 -17117 19932 -17083
rect 19874 -17151 19932 -17117
rect 19874 -17185 19886 -17151
rect 19920 -17185 19932 -17151
rect 19874 -17219 19932 -17185
rect 19874 -17253 19886 -17219
rect 19920 -17253 19932 -17219
rect 19874 -17298 19932 -17253
rect 20892 -16743 20950 -16698
rect 20892 -16777 20904 -16743
rect 20938 -16777 20950 -16743
rect 20892 -16811 20950 -16777
rect 20892 -16845 20904 -16811
rect 20938 -16845 20950 -16811
rect 20892 -16879 20950 -16845
rect 20892 -16913 20904 -16879
rect 20938 -16913 20950 -16879
rect 20892 -16947 20950 -16913
rect 20892 -16981 20904 -16947
rect 20938 -16981 20950 -16947
rect 20892 -17015 20950 -16981
rect 20892 -17049 20904 -17015
rect 20938 -17049 20950 -17015
rect 20892 -17083 20950 -17049
rect 20892 -17117 20904 -17083
rect 20938 -17117 20950 -17083
rect 20892 -17151 20950 -17117
rect 20892 -17185 20904 -17151
rect 20938 -17185 20950 -17151
rect 20892 -17219 20950 -17185
rect 20892 -17253 20904 -17219
rect 20938 -17253 20950 -17219
rect 20892 -17298 20950 -17253
rect 21910 -16743 21968 -16698
rect 21910 -16777 21922 -16743
rect 21956 -16777 21968 -16743
rect 21910 -16811 21968 -16777
rect 21910 -16845 21922 -16811
rect 21956 -16845 21968 -16811
rect 21910 -16879 21968 -16845
rect 21910 -16913 21922 -16879
rect 21956 -16913 21968 -16879
rect 21910 -16947 21968 -16913
rect 21910 -16981 21922 -16947
rect 21956 -16981 21968 -16947
rect 21910 -17015 21968 -16981
rect 21910 -17049 21922 -17015
rect 21956 -17049 21968 -17015
rect 21910 -17083 21968 -17049
rect 21910 -17117 21922 -17083
rect 21956 -17117 21968 -17083
rect 21910 -17151 21968 -17117
rect 21910 -17185 21922 -17151
rect 21956 -17185 21968 -17151
rect 21910 -17219 21968 -17185
rect 21910 -17253 21922 -17219
rect 21956 -17253 21968 -17219
rect 21910 -17298 21968 -17253
rect 22928 -16743 22986 -16698
rect 22928 -16777 22940 -16743
rect 22974 -16777 22986 -16743
rect 22928 -16811 22986 -16777
rect 22928 -16845 22940 -16811
rect 22974 -16845 22986 -16811
rect 22928 -16879 22986 -16845
rect 22928 -16913 22940 -16879
rect 22974 -16913 22986 -16879
rect 22928 -16947 22986 -16913
rect 22928 -16981 22940 -16947
rect 22974 -16981 22986 -16947
rect 22928 -17015 22986 -16981
rect 22928 -17049 22940 -17015
rect 22974 -17049 22986 -17015
rect 22928 -17083 22986 -17049
rect 22928 -17117 22940 -17083
rect 22974 -17117 22986 -17083
rect 22928 -17151 22986 -17117
rect 22928 -17185 22940 -17151
rect 22974 -17185 22986 -17151
rect 22928 -17219 22986 -17185
rect 22928 -17253 22940 -17219
rect 22974 -17253 22986 -17219
rect 22928 -17298 22986 -17253
rect -9196 -17465 -9138 -17420
rect -9196 -17499 -9184 -17465
rect -9150 -17499 -9138 -17465
rect -9196 -17533 -9138 -17499
rect -9196 -17567 -9184 -17533
rect -9150 -17567 -9138 -17533
rect -9196 -17601 -9138 -17567
rect -9196 -17635 -9184 -17601
rect -9150 -17635 -9138 -17601
rect -9196 -17669 -9138 -17635
rect -9196 -17703 -9184 -17669
rect -9150 -17703 -9138 -17669
rect -9196 -17737 -9138 -17703
rect -9196 -17771 -9184 -17737
rect -9150 -17771 -9138 -17737
rect -9196 -17805 -9138 -17771
rect -9196 -17839 -9184 -17805
rect -9150 -17839 -9138 -17805
rect -9196 -17873 -9138 -17839
rect -9196 -17907 -9184 -17873
rect -9150 -17907 -9138 -17873
rect -9196 -17941 -9138 -17907
rect -9196 -17975 -9184 -17941
rect -9150 -17975 -9138 -17941
rect -9196 -18020 -9138 -17975
rect -8178 -17465 -8120 -17420
rect -8178 -17499 -8166 -17465
rect -8132 -17499 -8120 -17465
rect -8178 -17533 -8120 -17499
rect -8178 -17567 -8166 -17533
rect -8132 -17567 -8120 -17533
rect -8178 -17601 -8120 -17567
rect -8178 -17635 -8166 -17601
rect -8132 -17635 -8120 -17601
rect -8178 -17669 -8120 -17635
rect -8178 -17703 -8166 -17669
rect -8132 -17703 -8120 -17669
rect -8178 -17737 -8120 -17703
rect -8178 -17771 -8166 -17737
rect -8132 -17771 -8120 -17737
rect -8178 -17805 -8120 -17771
rect -8178 -17839 -8166 -17805
rect -8132 -17839 -8120 -17805
rect -8178 -17873 -8120 -17839
rect -8178 -17907 -8166 -17873
rect -8132 -17907 -8120 -17873
rect -8178 -17941 -8120 -17907
rect -8178 -17975 -8166 -17941
rect -8132 -17975 -8120 -17941
rect -8178 -18020 -8120 -17975
rect -7160 -17465 -7102 -17420
rect -7160 -17499 -7148 -17465
rect -7114 -17499 -7102 -17465
rect -7160 -17533 -7102 -17499
rect -7160 -17567 -7148 -17533
rect -7114 -17567 -7102 -17533
rect -7160 -17601 -7102 -17567
rect -7160 -17635 -7148 -17601
rect -7114 -17635 -7102 -17601
rect -7160 -17669 -7102 -17635
rect -7160 -17703 -7148 -17669
rect -7114 -17703 -7102 -17669
rect -7160 -17737 -7102 -17703
rect -7160 -17771 -7148 -17737
rect -7114 -17771 -7102 -17737
rect -7160 -17805 -7102 -17771
rect -7160 -17839 -7148 -17805
rect -7114 -17839 -7102 -17805
rect -7160 -17873 -7102 -17839
rect -7160 -17907 -7148 -17873
rect -7114 -17907 -7102 -17873
rect -7160 -17941 -7102 -17907
rect -7160 -17975 -7148 -17941
rect -7114 -17975 -7102 -17941
rect -7160 -18020 -7102 -17975
rect -6142 -17465 -6084 -17420
rect -6142 -17499 -6130 -17465
rect -6096 -17499 -6084 -17465
rect -6142 -17533 -6084 -17499
rect -6142 -17567 -6130 -17533
rect -6096 -17567 -6084 -17533
rect -6142 -17601 -6084 -17567
rect -6142 -17635 -6130 -17601
rect -6096 -17635 -6084 -17601
rect -6142 -17669 -6084 -17635
rect -6142 -17703 -6130 -17669
rect -6096 -17703 -6084 -17669
rect -6142 -17737 -6084 -17703
rect -6142 -17771 -6130 -17737
rect -6096 -17771 -6084 -17737
rect -6142 -17805 -6084 -17771
rect -6142 -17839 -6130 -17805
rect -6096 -17839 -6084 -17805
rect -6142 -17873 -6084 -17839
rect -6142 -17907 -6130 -17873
rect -6096 -17907 -6084 -17873
rect -6142 -17941 -6084 -17907
rect -6142 -17975 -6130 -17941
rect -6096 -17975 -6084 -17941
rect -6142 -18020 -6084 -17975
rect -5124 -17465 -5066 -17420
rect -5124 -17499 -5112 -17465
rect -5078 -17499 -5066 -17465
rect -5124 -17533 -5066 -17499
rect -5124 -17567 -5112 -17533
rect -5078 -17567 -5066 -17533
rect -5124 -17601 -5066 -17567
rect -5124 -17635 -5112 -17601
rect -5078 -17635 -5066 -17601
rect -5124 -17669 -5066 -17635
rect -5124 -17703 -5112 -17669
rect -5078 -17703 -5066 -17669
rect -5124 -17737 -5066 -17703
rect -5124 -17771 -5112 -17737
rect -5078 -17771 -5066 -17737
rect -5124 -17805 -5066 -17771
rect -5124 -17839 -5112 -17805
rect -5078 -17839 -5066 -17805
rect -5124 -17873 -5066 -17839
rect -5124 -17907 -5112 -17873
rect -5078 -17907 -5066 -17873
rect -5124 -17941 -5066 -17907
rect -5124 -17975 -5112 -17941
rect -5078 -17975 -5066 -17941
rect -5124 -18020 -5066 -17975
rect -4106 -17465 -4048 -17420
rect -4106 -17499 -4094 -17465
rect -4060 -17499 -4048 -17465
rect -4106 -17533 -4048 -17499
rect -4106 -17567 -4094 -17533
rect -4060 -17567 -4048 -17533
rect -4106 -17601 -4048 -17567
rect -4106 -17635 -4094 -17601
rect -4060 -17635 -4048 -17601
rect -4106 -17669 -4048 -17635
rect -4106 -17703 -4094 -17669
rect -4060 -17703 -4048 -17669
rect -4106 -17737 -4048 -17703
rect -4106 -17771 -4094 -17737
rect -4060 -17771 -4048 -17737
rect -4106 -17805 -4048 -17771
rect -4106 -17839 -4094 -17805
rect -4060 -17839 -4048 -17805
rect -4106 -17873 -4048 -17839
rect -4106 -17907 -4094 -17873
rect -4060 -17907 -4048 -17873
rect -4106 -17941 -4048 -17907
rect -4106 -17975 -4094 -17941
rect -4060 -17975 -4048 -17941
rect -4106 -18020 -4048 -17975
rect -3088 -17465 -3030 -17420
rect -3088 -17499 -3076 -17465
rect -3042 -17499 -3030 -17465
rect -3088 -17533 -3030 -17499
rect -3088 -17567 -3076 -17533
rect -3042 -17567 -3030 -17533
rect -3088 -17601 -3030 -17567
rect -3088 -17635 -3076 -17601
rect -3042 -17635 -3030 -17601
rect -3088 -17669 -3030 -17635
rect -3088 -17703 -3076 -17669
rect -3042 -17703 -3030 -17669
rect -3088 -17737 -3030 -17703
rect -3088 -17771 -3076 -17737
rect -3042 -17771 -3030 -17737
rect -3088 -17805 -3030 -17771
rect -3088 -17839 -3076 -17805
rect -3042 -17839 -3030 -17805
rect -3088 -17873 -3030 -17839
rect -3088 -17907 -3076 -17873
rect -3042 -17907 -3030 -17873
rect -3088 -17941 -3030 -17907
rect -3088 -17975 -3076 -17941
rect -3042 -17975 -3030 -17941
rect -3088 -18020 -3030 -17975
rect -2070 -17465 -2012 -17420
rect -2070 -17499 -2058 -17465
rect -2024 -17499 -2012 -17465
rect -2070 -17533 -2012 -17499
rect -2070 -17567 -2058 -17533
rect -2024 -17567 -2012 -17533
rect -2070 -17601 -2012 -17567
rect -2070 -17635 -2058 -17601
rect -2024 -17635 -2012 -17601
rect -2070 -17669 -2012 -17635
rect -2070 -17703 -2058 -17669
rect -2024 -17703 -2012 -17669
rect -2070 -17737 -2012 -17703
rect -2070 -17771 -2058 -17737
rect -2024 -17771 -2012 -17737
rect -2070 -17805 -2012 -17771
rect -2070 -17839 -2058 -17805
rect -2024 -17839 -2012 -17805
rect -2070 -17873 -2012 -17839
rect -2070 -17907 -2058 -17873
rect -2024 -17907 -2012 -17873
rect -2070 -17941 -2012 -17907
rect -2070 -17975 -2058 -17941
rect -2024 -17975 -2012 -17941
rect -2070 -18020 -2012 -17975
rect -1052 -17465 -994 -17420
rect -1052 -17499 -1040 -17465
rect -1006 -17499 -994 -17465
rect -1052 -17533 -994 -17499
rect -1052 -17567 -1040 -17533
rect -1006 -17567 -994 -17533
rect -1052 -17601 -994 -17567
rect -1052 -17635 -1040 -17601
rect -1006 -17635 -994 -17601
rect -1052 -17669 -994 -17635
rect -1052 -17703 -1040 -17669
rect -1006 -17703 -994 -17669
rect -1052 -17737 -994 -17703
rect -1052 -17771 -1040 -17737
rect -1006 -17771 -994 -17737
rect -1052 -17805 -994 -17771
rect -1052 -17839 -1040 -17805
rect -1006 -17839 -994 -17805
rect -1052 -17873 -994 -17839
rect -1052 -17907 -1040 -17873
rect -1006 -17907 -994 -17873
rect -1052 -17941 -994 -17907
rect -1052 -17975 -1040 -17941
rect -1006 -17975 -994 -17941
rect -1052 -18020 -994 -17975
rect -34 -17465 24 -17420
rect -34 -17499 -22 -17465
rect 12 -17499 24 -17465
rect -34 -17533 24 -17499
rect -34 -17567 -22 -17533
rect 12 -17567 24 -17533
rect -34 -17601 24 -17567
rect -34 -17635 -22 -17601
rect 12 -17635 24 -17601
rect -34 -17669 24 -17635
rect -34 -17703 -22 -17669
rect 12 -17703 24 -17669
rect -34 -17737 24 -17703
rect -34 -17771 -22 -17737
rect 12 -17771 24 -17737
rect -34 -17805 24 -17771
rect -34 -17839 -22 -17805
rect 12 -17839 24 -17805
rect -34 -17873 24 -17839
rect -34 -17907 -22 -17873
rect 12 -17907 24 -17873
rect -34 -17941 24 -17907
rect -34 -17975 -22 -17941
rect 12 -17975 24 -17941
rect -34 -18020 24 -17975
rect 2568 -17977 2626 -17932
rect 2568 -18011 2580 -17977
rect 2614 -18011 2626 -17977
rect 2568 -18045 2626 -18011
rect 2568 -18079 2580 -18045
rect 2614 -18079 2626 -18045
rect 2568 -18113 2626 -18079
rect 2568 -18147 2580 -18113
rect 2614 -18147 2626 -18113
rect 2568 -18181 2626 -18147
rect 2568 -18215 2580 -18181
rect 2614 -18215 2626 -18181
rect -9196 -18283 -9138 -18238
rect -9196 -18317 -9184 -18283
rect -9150 -18317 -9138 -18283
rect -9196 -18351 -9138 -18317
rect -9196 -18385 -9184 -18351
rect -9150 -18385 -9138 -18351
rect -9196 -18419 -9138 -18385
rect -9196 -18453 -9184 -18419
rect -9150 -18453 -9138 -18419
rect -9196 -18487 -9138 -18453
rect -9196 -18521 -9184 -18487
rect -9150 -18521 -9138 -18487
rect -9196 -18555 -9138 -18521
rect -9196 -18589 -9184 -18555
rect -9150 -18589 -9138 -18555
rect -9196 -18623 -9138 -18589
rect -9196 -18657 -9184 -18623
rect -9150 -18657 -9138 -18623
rect -9196 -18691 -9138 -18657
rect -9196 -18725 -9184 -18691
rect -9150 -18725 -9138 -18691
rect -9196 -18759 -9138 -18725
rect -9196 -18793 -9184 -18759
rect -9150 -18793 -9138 -18759
rect -9196 -18838 -9138 -18793
rect -8178 -18283 -8120 -18238
rect -8178 -18317 -8166 -18283
rect -8132 -18317 -8120 -18283
rect -8178 -18351 -8120 -18317
rect -8178 -18385 -8166 -18351
rect -8132 -18385 -8120 -18351
rect -8178 -18419 -8120 -18385
rect -8178 -18453 -8166 -18419
rect -8132 -18453 -8120 -18419
rect -8178 -18487 -8120 -18453
rect -8178 -18521 -8166 -18487
rect -8132 -18521 -8120 -18487
rect -8178 -18555 -8120 -18521
rect -8178 -18589 -8166 -18555
rect -8132 -18589 -8120 -18555
rect -8178 -18623 -8120 -18589
rect -8178 -18657 -8166 -18623
rect -8132 -18657 -8120 -18623
rect -8178 -18691 -8120 -18657
rect -8178 -18725 -8166 -18691
rect -8132 -18725 -8120 -18691
rect -8178 -18759 -8120 -18725
rect -8178 -18793 -8166 -18759
rect -8132 -18793 -8120 -18759
rect -8178 -18838 -8120 -18793
rect -7160 -18283 -7102 -18238
rect -7160 -18317 -7148 -18283
rect -7114 -18317 -7102 -18283
rect -7160 -18351 -7102 -18317
rect -7160 -18385 -7148 -18351
rect -7114 -18385 -7102 -18351
rect -7160 -18419 -7102 -18385
rect -7160 -18453 -7148 -18419
rect -7114 -18453 -7102 -18419
rect -7160 -18487 -7102 -18453
rect -7160 -18521 -7148 -18487
rect -7114 -18521 -7102 -18487
rect -7160 -18555 -7102 -18521
rect -7160 -18589 -7148 -18555
rect -7114 -18589 -7102 -18555
rect -7160 -18623 -7102 -18589
rect -7160 -18657 -7148 -18623
rect -7114 -18657 -7102 -18623
rect -7160 -18691 -7102 -18657
rect -7160 -18725 -7148 -18691
rect -7114 -18725 -7102 -18691
rect -7160 -18759 -7102 -18725
rect -7160 -18793 -7148 -18759
rect -7114 -18793 -7102 -18759
rect -7160 -18838 -7102 -18793
rect -6142 -18283 -6084 -18238
rect -6142 -18317 -6130 -18283
rect -6096 -18317 -6084 -18283
rect -6142 -18351 -6084 -18317
rect -6142 -18385 -6130 -18351
rect -6096 -18385 -6084 -18351
rect -6142 -18419 -6084 -18385
rect -6142 -18453 -6130 -18419
rect -6096 -18453 -6084 -18419
rect -6142 -18487 -6084 -18453
rect -6142 -18521 -6130 -18487
rect -6096 -18521 -6084 -18487
rect -6142 -18555 -6084 -18521
rect -6142 -18589 -6130 -18555
rect -6096 -18589 -6084 -18555
rect -6142 -18623 -6084 -18589
rect -6142 -18657 -6130 -18623
rect -6096 -18657 -6084 -18623
rect -6142 -18691 -6084 -18657
rect -6142 -18725 -6130 -18691
rect -6096 -18725 -6084 -18691
rect -6142 -18759 -6084 -18725
rect -6142 -18793 -6130 -18759
rect -6096 -18793 -6084 -18759
rect -6142 -18838 -6084 -18793
rect -5124 -18283 -5066 -18238
rect -5124 -18317 -5112 -18283
rect -5078 -18317 -5066 -18283
rect -5124 -18351 -5066 -18317
rect -5124 -18385 -5112 -18351
rect -5078 -18385 -5066 -18351
rect -5124 -18419 -5066 -18385
rect -5124 -18453 -5112 -18419
rect -5078 -18453 -5066 -18419
rect -5124 -18487 -5066 -18453
rect -5124 -18521 -5112 -18487
rect -5078 -18521 -5066 -18487
rect -5124 -18555 -5066 -18521
rect -5124 -18589 -5112 -18555
rect -5078 -18589 -5066 -18555
rect -5124 -18623 -5066 -18589
rect -5124 -18657 -5112 -18623
rect -5078 -18657 -5066 -18623
rect -5124 -18691 -5066 -18657
rect -5124 -18725 -5112 -18691
rect -5078 -18725 -5066 -18691
rect -5124 -18759 -5066 -18725
rect -5124 -18793 -5112 -18759
rect -5078 -18793 -5066 -18759
rect -5124 -18838 -5066 -18793
rect -4106 -18283 -4048 -18238
rect -4106 -18317 -4094 -18283
rect -4060 -18317 -4048 -18283
rect -4106 -18351 -4048 -18317
rect -4106 -18385 -4094 -18351
rect -4060 -18385 -4048 -18351
rect -4106 -18419 -4048 -18385
rect -4106 -18453 -4094 -18419
rect -4060 -18453 -4048 -18419
rect -4106 -18487 -4048 -18453
rect -4106 -18521 -4094 -18487
rect -4060 -18521 -4048 -18487
rect -4106 -18555 -4048 -18521
rect -4106 -18589 -4094 -18555
rect -4060 -18589 -4048 -18555
rect -4106 -18623 -4048 -18589
rect -4106 -18657 -4094 -18623
rect -4060 -18657 -4048 -18623
rect -4106 -18691 -4048 -18657
rect -4106 -18725 -4094 -18691
rect -4060 -18725 -4048 -18691
rect -4106 -18759 -4048 -18725
rect -4106 -18793 -4094 -18759
rect -4060 -18793 -4048 -18759
rect -4106 -18838 -4048 -18793
rect -3088 -18283 -3030 -18238
rect -3088 -18317 -3076 -18283
rect -3042 -18317 -3030 -18283
rect -3088 -18351 -3030 -18317
rect -3088 -18385 -3076 -18351
rect -3042 -18385 -3030 -18351
rect -3088 -18419 -3030 -18385
rect -3088 -18453 -3076 -18419
rect -3042 -18453 -3030 -18419
rect -3088 -18487 -3030 -18453
rect -3088 -18521 -3076 -18487
rect -3042 -18521 -3030 -18487
rect -3088 -18555 -3030 -18521
rect -3088 -18589 -3076 -18555
rect -3042 -18589 -3030 -18555
rect -3088 -18623 -3030 -18589
rect -3088 -18657 -3076 -18623
rect -3042 -18657 -3030 -18623
rect -3088 -18691 -3030 -18657
rect -3088 -18725 -3076 -18691
rect -3042 -18725 -3030 -18691
rect -3088 -18759 -3030 -18725
rect -3088 -18793 -3076 -18759
rect -3042 -18793 -3030 -18759
rect -3088 -18838 -3030 -18793
rect -2070 -18283 -2012 -18238
rect -2070 -18317 -2058 -18283
rect -2024 -18317 -2012 -18283
rect -2070 -18351 -2012 -18317
rect -2070 -18385 -2058 -18351
rect -2024 -18385 -2012 -18351
rect -2070 -18419 -2012 -18385
rect -2070 -18453 -2058 -18419
rect -2024 -18453 -2012 -18419
rect -2070 -18487 -2012 -18453
rect -2070 -18521 -2058 -18487
rect -2024 -18521 -2012 -18487
rect -2070 -18555 -2012 -18521
rect -2070 -18589 -2058 -18555
rect -2024 -18589 -2012 -18555
rect -2070 -18623 -2012 -18589
rect -2070 -18657 -2058 -18623
rect -2024 -18657 -2012 -18623
rect -2070 -18691 -2012 -18657
rect -2070 -18725 -2058 -18691
rect -2024 -18725 -2012 -18691
rect -2070 -18759 -2012 -18725
rect -2070 -18793 -2058 -18759
rect -2024 -18793 -2012 -18759
rect -2070 -18838 -2012 -18793
rect -1052 -18283 -994 -18238
rect -1052 -18317 -1040 -18283
rect -1006 -18317 -994 -18283
rect -1052 -18351 -994 -18317
rect -1052 -18385 -1040 -18351
rect -1006 -18385 -994 -18351
rect -1052 -18419 -994 -18385
rect -1052 -18453 -1040 -18419
rect -1006 -18453 -994 -18419
rect -1052 -18487 -994 -18453
rect -1052 -18521 -1040 -18487
rect -1006 -18521 -994 -18487
rect -1052 -18555 -994 -18521
rect -1052 -18589 -1040 -18555
rect -1006 -18589 -994 -18555
rect -1052 -18623 -994 -18589
rect -1052 -18657 -1040 -18623
rect -1006 -18657 -994 -18623
rect -1052 -18691 -994 -18657
rect -1052 -18725 -1040 -18691
rect -1006 -18725 -994 -18691
rect -1052 -18759 -994 -18725
rect -1052 -18793 -1040 -18759
rect -1006 -18793 -994 -18759
rect -1052 -18838 -994 -18793
rect -34 -18283 24 -18238
rect -34 -18317 -22 -18283
rect 12 -18317 24 -18283
rect -34 -18351 24 -18317
rect -34 -18385 -22 -18351
rect 12 -18385 24 -18351
rect -34 -18419 24 -18385
rect -34 -18453 -22 -18419
rect 12 -18453 24 -18419
rect -34 -18487 24 -18453
rect -34 -18521 -22 -18487
rect 12 -18521 24 -18487
rect -34 -18555 24 -18521
rect 2568 -18249 2626 -18215
rect 2568 -18283 2580 -18249
rect 2614 -18283 2626 -18249
rect 2568 -18317 2626 -18283
rect 2568 -18351 2580 -18317
rect 2614 -18351 2626 -18317
rect 2568 -18385 2626 -18351
rect 2568 -18419 2580 -18385
rect 2614 -18419 2626 -18385
rect 2568 -18453 2626 -18419
rect 2568 -18487 2580 -18453
rect 2614 -18487 2626 -18453
rect 2568 -18532 2626 -18487
rect 3586 -17977 3644 -17932
rect 3586 -18011 3598 -17977
rect 3632 -18011 3644 -17977
rect 3586 -18045 3644 -18011
rect 3586 -18079 3598 -18045
rect 3632 -18079 3644 -18045
rect 3586 -18113 3644 -18079
rect 3586 -18147 3598 -18113
rect 3632 -18147 3644 -18113
rect 3586 -18181 3644 -18147
rect 3586 -18215 3598 -18181
rect 3632 -18215 3644 -18181
rect 3586 -18249 3644 -18215
rect 3586 -18283 3598 -18249
rect 3632 -18283 3644 -18249
rect 3586 -18317 3644 -18283
rect 3586 -18351 3598 -18317
rect 3632 -18351 3644 -18317
rect 3586 -18385 3644 -18351
rect 3586 -18419 3598 -18385
rect 3632 -18419 3644 -18385
rect 3586 -18453 3644 -18419
rect 3586 -18487 3598 -18453
rect 3632 -18487 3644 -18453
rect 3586 -18532 3644 -18487
rect 4604 -17977 4662 -17932
rect 4604 -18011 4616 -17977
rect 4650 -18011 4662 -17977
rect 4604 -18045 4662 -18011
rect 4604 -18079 4616 -18045
rect 4650 -18079 4662 -18045
rect 4604 -18113 4662 -18079
rect 4604 -18147 4616 -18113
rect 4650 -18147 4662 -18113
rect 4604 -18181 4662 -18147
rect 4604 -18215 4616 -18181
rect 4650 -18215 4662 -18181
rect 4604 -18249 4662 -18215
rect 4604 -18283 4616 -18249
rect 4650 -18283 4662 -18249
rect 4604 -18317 4662 -18283
rect 4604 -18351 4616 -18317
rect 4650 -18351 4662 -18317
rect 4604 -18385 4662 -18351
rect 4604 -18419 4616 -18385
rect 4650 -18419 4662 -18385
rect 4604 -18453 4662 -18419
rect 4604 -18487 4616 -18453
rect 4650 -18487 4662 -18453
rect 4604 -18532 4662 -18487
rect 5622 -17977 5680 -17932
rect 5622 -18011 5634 -17977
rect 5668 -18011 5680 -17977
rect 5622 -18045 5680 -18011
rect 5622 -18079 5634 -18045
rect 5668 -18079 5680 -18045
rect 5622 -18113 5680 -18079
rect 5622 -18147 5634 -18113
rect 5668 -18147 5680 -18113
rect 5622 -18181 5680 -18147
rect 5622 -18215 5634 -18181
rect 5668 -18215 5680 -18181
rect 5622 -18249 5680 -18215
rect 5622 -18283 5634 -18249
rect 5668 -18283 5680 -18249
rect 5622 -18317 5680 -18283
rect 5622 -18351 5634 -18317
rect 5668 -18351 5680 -18317
rect 5622 -18385 5680 -18351
rect 5622 -18419 5634 -18385
rect 5668 -18419 5680 -18385
rect 5622 -18453 5680 -18419
rect 5622 -18487 5634 -18453
rect 5668 -18487 5680 -18453
rect 5622 -18532 5680 -18487
rect 6640 -17977 6698 -17932
rect 6640 -18011 6652 -17977
rect 6686 -18011 6698 -17977
rect 6640 -18045 6698 -18011
rect 6640 -18079 6652 -18045
rect 6686 -18079 6698 -18045
rect 6640 -18113 6698 -18079
rect 6640 -18147 6652 -18113
rect 6686 -18147 6698 -18113
rect 6640 -18181 6698 -18147
rect 6640 -18215 6652 -18181
rect 6686 -18215 6698 -18181
rect 6640 -18249 6698 -18215
rect 6640 -18283 6652 -18249
rect 6686 -18283 6698 -18249
rect 6640 -18317 6698 -18283
rect 6640 -18351 6652 -18317
rect 6686 -18351 6698 -18317
rect 6640 -18385 6698 -18351
rect 6640 -18419 6652 -18385
rect 6686 -18419 6698 -18385
rect 6640 -18453 6698 -18419
rect 6640 -18487 6652 -18453
rect 6686 -18487 6698 -18453
rect 6640 -18532 6698 -18487
rect 7658 -17977 7716 -17932
rect 7658 -18011 7670 -17977
rect 7704 -18011 7716 -17977
rect 7658 -18045 7716 -18011
rect 7658 -18079 7670 -18045
rect 7704 -18079 7716 -18045
rect 7658 -18113 7716 -18079
rect 7658 -18147 7670 -18113
rect 7704 -18147 7716 -18113
rect 7658 -18181 7716 -18147
rect 7658 -18215 7670 -18181
rect 7704 -18215 7716 -18181
rect 7658 -18249 7716 -18215
rect 7658 -18283 7670 -18249
rect 7704 -18283 7716 -18249
rect 7658 -18317 7716 -18283
rect 7658 -18351 7670 -18317
rect 7704 -18351 7716 -18317
rect 7658 -18385 7716 -18351
rect 7658 -18419 7670 -18385
rect 7704 -18419 7716 -18385
rect 7658 -18453 7716 -18419
rect 7658 -18487 7670 -18453
rect 7704 -18487 7716 -18453
rect 7658 -18532 7716 -18487
rect 8676 -17977 8734 -17932
rect 8676 -18011 8688 -17977
rect 8722 -18011 8734 -17977
rect 8676 -18045 8734 -18011
rect 8676 -18079 8688 -18045
rect 8722 -18079 8734 -18045
rect 8676 -18113 8734 -18079
rect 8676 -18147 8688 -18113
rect 8722 -18147 8734 -18113
rect 8676 -18181 8734 -18147
rect 8676 -18215 8688 -18181
rect 8722 -18215 8734 -18181
rect 8676 -18249 8734 -18215
rect 8676 -18283 8688 -18249
rect 8722 -18283 8734 -18249
rect 8676 -18317 8734 -18283
rect 8676 -18351 8688 -18317
rect 8722 -18351 8734 -18317
rect 8676 -18385 8734 -18351
rect 8676 -18419 8688 -18385
rect 8722 -18419 8734 -18385
rect 8676 -18453 8734 -18419
rect 8676 -18487 8688 -18453
rect 8722 -18487 8734 -18453
rect 8676 -18532 8734 -18487
rect 9694 -17977 9752 -17932
rect 9694 -18011 9706 -17977
rect 9740 -18011 9752 -17977
rect 9694 -18045 9752 -18011
rect 9694 -18079 9706 -18045
rect 9740 -18079 9752 -18045
rect 9694 -18113 9752 -18079
rect 9694 -18147 9706 -18113
rect 9740 -18147 9752 -18113
rect 9694 -18181 9752 -18147
rect 9694 -18215 9706 -18181
rect 9740 -18215 9752 -18181
rect 9694 -18249 9752 -18215
rect 9694 -18283 9706 -18249
rect 9740 -18283 9752 -18249
rect 9694 -18317 9752 -18283
rect 9694 -18351 9706 -18317
rect 9740 -18351 9752 -18317
rect 9694 -18385 9752 -18351
rect 9694 -18419 9706 -18385
rect 9740 -18419 9752 -18385
rect 9694 -18453 9752 -18419
rect 9694 -18487 9706 -18453
rect 9740 -18487 9752 -18453
rect 9694 -18532 9752 -18487
rect 10712 -17977 10770 -17932
rect 10712 -18011 10724 -17977
rect 10758 -18011 10770 -17977
rect 10712 -18045 10770 -18011
rect 10712 -18079 10724 -18045
rect 10758 -18079 10770 -18045
rect 10712 -18113 10770 -18079
rect 10712 -18147 10724 -18113
rect 10758 -18147 10770 -18113
rect 10712 -18181 10770 -18147
rect 10712 -18215 10724 -18181
rect 10758 -18215 10770 -18181
rect 10712 -18249 10770 -18215
rect 10712 -18283 10724 -18249
rect 10758 -18283 10770 -18249
rect 10712 -18317 10770 -18283
rect 10712 -18351 10724 -18317
rect 10758 -18351 10770 -18317
rect 10712 -18385 10770 -18351
rect 10712 -18419 10724 -18385
rect 10758 -18419 10770 -18385
rect 10712 -18453 10770 -18419
rect 10712 -18487 10724 -18453
rect 10758 -18487 10770 -18453
rect 10712 -18532 10770 -18487
rect 11730 -17977 11788 -17932
rect 11730 -18011 11742 -17977
rect 11776 -18011 11788 -17977
rect 11730 -18045 11788 -18011
rect 11730 -18079 11742 -18045
rect 11776 -18079 11788 -18045
rect 11730 -18113 11788 -18079
rect 11730 -18147 11742 -18113
rect 11776 -18147 11788 -18113
rect 11730 -18181 11788 -18147
rect 11730 -18215 11742 -18181
rect 11776 -18215 11788 -18181
rect 11730 -18249 11788 -18215
rect 11730 -18283 11742 -18249
rect 11776 -18283 11788 -18249
rect 11730 -18317 11788 -18283
rect 11730 -18351 11742 -18317
rect 11776 -18351 11788 -18317
rect 11730 -18385 11788 -18351
rect 11730 -18419 11742 -18385
rect 11776 -18419 11788 -18385
rect 11730 -18453 11788 -18419
rect 11730 -18487 11742 -18453
rect 11776 -18487 11788 -18453
rect 11730 -18532 11788 -18487
rect 12748 -17977 12806 -17932
rect 12748 -18011 12760 -17977
rect 12794 -18011 12806 -17977
rect 12748 -18045 12806 -18011
rect 12748 -18079 12760 -18045
rect 12794 -18079 12806 -18045
rect 12748 -18113 12806 -18079
rect 12748 -18147 12760 -18113
rect 12794 -18147 12806 -18113
rect 12748 -18181 12806 -18147
rect 12748 -18215 12760 -18181
rect 12794 -18215 12806 -18181
rect 12748 -18249 12806 -18215
rect 12748 -18283 12760 -18249
rect 12794 -18283 12806 -18249
rect 12748 -18317 12806 -18283
rect 12748 -18351 12760 -18317
rect 12794 -18351 12806 -18317
rect 12748 -18385 12806 -18351
rect 12748 -18419 12760 -18385
rect 12794 -18419 12806 -18385
rect 12748 -18453 12806 -18419
rect 12748 -18487 12760 -18453
rect 12794 -18487 12806 -18453
rect 12748 -18532 12806 -18487
rect 13766 -17977 13824 -17932
rect 13766 -18011 13778 -17977
rect 13812 -18011 13824 -17977
rect 13766 -18045 13824 -18011
rect 13766 -18079 13778 -18045
rect 13812 -18079 13824 -18045
rect 13766 -18113 13824 -18079
rect 13766 -18147 13778 -18113
rect 13812 -18147 13824 -18113
rect 13766 -18181 13824 -18147
rect 13766 -18215 13778 -18181
rect 13812 -18215 13824 -18181
rect 13766 -18249 13824 -18215
rect 13766 -18283 13778 -18249
rect 13812 -18283 13824 -18249
rect 13766 -18317 13824 -18283
rect 13766 -18351 13778 -18317
rect 13812 -18351 13824 -18317
rect 13766 -18385 13824 -18351
rect 13766 -18419 13778 -18385
rect 13812 -18419 13824 -18385
rect 13766 -18453 13824 -18419
rect 13766 -18487 13778 -18453
rect 13812 -18487 13824 -18453
rect 13766 -18532 13824 -18487
rect 14784 -17977 14842 -17932
rect 14784 -18011 14796 -17977
rect 14830 -18011 14842 -17977
rect 14784 -18045 14842 -18011
rect 14784 -18079 14796 -18045
rect 14830 -18079 14842 -18045
rect 14784 -18113 14842 -18079
rect 14784 -18147 14796 -18113
rect 14830 -18147 14842 -18113
rect 14784 -18181 14842 -18147
rect 14784 -18215 14796 -18181
rect 14830 -18215 14842 -18181
rect 14784 -18249 14842 -18215
rect 14784 -18283 14796 -18249
rect 14830 -18283 14842 -18249
rect 14784 -18317 14842 -18283
rect 14784 -18351 14796 -18317
rect 14830 -18351 14842 -18317
rect 14784 -18385 14842 -18351
rect 14784 -18419 14796 -18385
rect 14830 -18419 14842 -18385
rect 14784 -18453 14842 -18419
rect 14784 -18487 14796 -18453
rect 14830 -18487 14842 -18453
rect 14784 -18532 14842 -18487
rect 15802 -17977 15860 -17932
rect 15802 -18011 15814 -17977
rect 15848 -18011 15860 -17977
rect 15802 -18045 15860 -18011
rect 15802 -18079 15814 -18045
rect 15848 -18079 15860 -18045
rect 15802 -18113 15860 -18079
rect 15802 -18147 15814 -18113
rect 15848 -18147 15860 -18113
rect 15802 -18181 15860 -18147
rect 15802 -18215 15814 -18181
rect 15848 -18215 15860 -18181
rect 15802 -18249 15860 -18215
rect 15802 -18283 15814 -18249
rect 15848 -18283 15860 -18249
rect 15802 -18317 15860 -18283
rect 15802 -18351 15814 -18317
rect 15848 -18351 15860 -18317
rect 15802 -18385 15860 -18351
rect 15802 -18419 15814 -18385
rect 15848 -18419 15860 -18385
rect 15802 -18453 15860 -18419
rect 15802 -18487 15814 -18453
rect 15848 -18487 15860 -18453
rect 15802 -18532 15860 -18487
rect 16820 -17977 16878 -17932
rect 16820 -18011 16832 -17977
rect 16866 -18011 16878 -17977
rect 16820 -18045 16878 -18011
rect 16820 -18079 16832 -18045
rect 16866 -18079 16878 -18045
rect 16820 -18113 16878 -18079
rect 16820 -18147 16832 -18113
rect 16866 -18147 16878 -18113
rect 16820 -18181 16878 -18147
rect 16820 -18215 16832 -18181
rect 16866 -18215 16878 -18181
rect 16820 -18249 16878 -18215
rect 16820 -18283 16832 -18249
rect 16866 -18283 16878 -18249
rect 16820 -18317 16878 -18283
rect 16820 -18351 16832 -18317
rect 16866 -18351 16878 -18317
rect 16820 -18385 16878 -18351
rect 16820 -18419 16832 -18385
rect 16866 -18419 16878 -18385
rect 16820 -18453 16878 -18419
rect 16820 -18487 16832 -18453
rect 16866 -18487 16878 -18453
rect 16820 -18532 16878 -18487
rect 17838 -17977 17896 -17932
rect 17838 -18011 17850 -17977
rect 17884 -18011 17896 -17977
rect 17838 -18045 17896 -18011
rect 17838 -18079 17850 -18045
rect 17884 -18079 17896 -18045
rect 17838 -18113 17896 -18079
rect 17838 -18147 17850 -18113
rect 17884 -18147 17896 -18113
rect 17838 -18181 17896 -18147
rect 17838 -18215 17850 -18181
rect 17884 -18215 17896 -18181
rect 17838 -18249 17896 -18215
rect 17838 -18283 17850 -18249
rect 17884 -18283 17896 -18249
rect 17838 -18317 17896 -18283
rect 17838 -18351 17850 -18317
rect 17884 -18351 17896 -18317
rect 17838 -18385 17896 -18351
rect 17838 -18419 17850 -18385
rect 17884 -18419 17896 -18385
rect 17838 -18453 17896 -18419
rect 17838 -18487 17850 -18453
rect 17884 -18487 17896 -18453
rect 17838 -18532 17896 -18487
rect 18856 -17977 18914 -17932
rect 18856 -18011 18868 -17977
rect 18902 -18011 18914 -17977
rect 18856 -18045 18914 -18011
rect 18856 -18079 18868 -18045
rect 18902 -18079 18914 -18045
rect 18856 -18113 18914 -18079
rect 18856 -18147 18868 -18113
rect 18902 -18147 18914 -18113
rect 18856 -18181 18914 -18147
rect 18856 -18215 18868 -18181
rect 18902 -18215 18914 -18181
rect 18856 -18249 18914 -18215
rect 18856 -18283 18868 -18249
rect 18902 -18283 18914 -18249
rect 18856 -18317 18914 -18283
rect 18856 -18351 18868 -18317
rect 18902 -18351 18914 -18317
rect 18856 -18385 18914 -18351
rect 18856 -18419 18868 -18385
rect 18902 -18419 18914 -18385
rect 18856 -18453 18914 -18419
rect 18856 -18487 18868 -18453
rect 18902 -18487 18914 -18453
rect 18856 -18532 18914 -18487
rect 19874 -17977 19932 -17932
rect 19874 -18011 19886 -17977
rect 19920 -18011 19932 -17977
rect 19874 -18045 19932 -18011
rect 19874 -18079 19886 -18045
rect 19920 -18079 19932 -18045
rect 19874 -18113 19932 -18079
rect 19874 -18147 19886 -18113
rect 19920 -18147 19932 -18113
rect 19874 -18181 19932 -18147
rect 19874 -18215 19886 -18181
rect 19920 -18215 19932 -18181
rect 19874 -18249 19932 -18215
rect 19874 -18283 19886 -18249
rect 19920 -18283 19932 -18249
rect 19874 -18317 19932 -18283
rect 19874 -18351 19886 -18317
rect 19920 -18351 19932 -18317
rect 19874 -18385 19932 -18351
rect 19874 -18419 19886 -18385
rect 19920 -18419 19932 -18385
rect 19874 -18453 19932 -18419
rect 19874 -18487 19886 -18453
rect 19920 -18487 19932 -18453
rect 19874 -18532 19932 -18487
rect 20892 -17977 20950 -17932
rect 20892 -18011 20904 -17977
rect 20938 -18011 20950 -17977
rect 20892 -18045 20950 -18011
rect 20892 -18079 20904 -18045
rect 20938 -18079 20950 -18045
rect 20892 -18113 20950 -18079
rect 20892 -18147 20904 -18113
rect 20938 -18147 20950 -18113
rect 20892 -18181 20950 -18147
rect 20892 -18215 20904 -18181
rect 20938 -18215 20950 -18181
rect 20892 -18249 20950 -18215
rect 20892 -18283 20904 -18249
rect 20938 -18283 20950 -18249
rect 20892 -18317 20950 -18283
rect 20892 -18351 20904 -18317
rect 20938 -18351 20950 -18317
rect 20892 -18385 20950 -18351
rect 20892 -18419 20904 -18385
rect 20938 -18419 20950 -18385
rect 20892 -18453 20950 -18419
rect 20892 -18487 20904 -18453
rect 20938 -18487 20950 -18453
rect 20892 -18532 20950 -18487
rect 21910 -17977 21968 -17932
rect 21910 -18011 21922 -17977
rect 21956 -18011 21968 -17977
rect 21910 -18045 21968 -18011
rect 21910 -18079 21922 -18045
rect 21956 -18079 21968 -18045
rect 21910 -18113 21968 -18079
rect 21910 -18147 21922 -18113
rect 21956 -18147 21968 -18113
rect 21910 -18181 21968 -18147
rect 21910 -18215 21922 -18181
rect 21956 -18215 21968 -18181
rect 21910 -18249 21968 -18215
rect 21910 -18283 21922 -18249
rect 21956 -18283 21968 -18249
rect 21910 -18317 21968 -18283
rect 21910 -18351 21922 -18317
rect 21956 -18351 21968 -18317
rect 21910 -18385 21968 -18351
rect 21910 -18419 21922 -18385
rect 21956 -18419 21968 -18385
rect 21910 -18453 21968 -18419
rect 21910 -18487 21922 -18453
rect 21956 -18487 21968 -18453
rect 21910 -18532 21968 -18487
rect 22928 -17977 22986 -17932
rect 22928 -18011 22940 -17977
rect 22974 -18011 22986 -17977
rect 22928 -18045 22986 -18011
rect 22928 -18079 22940 -18045
rect 22974 -18079 22986 -18045
rect 22928 -18113 22986 -18079
rect 22928 -18147 22940 -18113
rect 22974 -18147 22986 -18113
rect 22928 -18181 22986 -18147
rect 22928 -18215 22940 -18181
rect 22974 -18215 22986 -18181
rect 22928 -18249 22986 -18215
rect 22928 -18283 22940 -18249
rect 22974 -18283 22986 -18249
rect 22928 -18317 22986 -18283
rect 22928 -18351 22940 -18317
rect 22974 -18351 22986 -18317
rect 22928 -18385 22986 -18351
rect 22928 -18419 22940 -18385
rect 22974 -18419 22986 -18385
rect 22928 -18453 22986 -18419
rect 22928 -18487 22940 -18453
rect 22974 -18487 22986 -18453
rect 22928 -18532 22986 -18487
rect -34 -18589 -22 -18555
rect 12 -18589 24 -18555
rect -34 -18623 24 -18589
rect -34 -18657 -22 -18623
rect 12 -18657 24 -18623
rect -34 -18691 24 -18657
rect -34 -18725 -22 -18691
rect 12 -18725 24 -18691
rect -34 -18759 24 -18725
rect -34 -18793 -22 -18759
rect 12 -18793 24 -18759
rect -34 -18838 24 -18793
rect 2568 -19209 2626 -19164
rect 2568 -19243 2580 -19209
rect 2614 -19243 2626 -19209
rect 2568 -19277 2626 -19243
rect 2568 -19311 2580 -19277
rect 2614 -19311 2626 -19277
rect 2568 -19345 2626 -19311
rect 2568 -19379 2580 -19345
rect 2614 -19379 2626 -19345
rect 2568 -19413 2626 -19379
rect 2568 -19447 2580 -19413
rect 2614 -19447 2626 -19413
rect 2568 -19481 2626 -19447
rect 2568 -19515 2580 -19481
rect 2614 -19515 2626 -19481
rect 2568 -19549 2626 -19515
rect 2568 -19583 2580 -19549
rect 2614 -19583 2626 -19549
rect 2568 -19617 2626 -19583
rect 2568 -19651 2580 -19617
rect 2614 -19651 2626 -19617
rect 2568 -19685 2626 -19651
rect 2568 -19719 2580 -19685
rect 2614 -19719 2626 -19685
rect 2568 -19764 2626 -19719
rect 3586 -19209 3644 -19164
rect 3586 -19243 3598 -19209
rect 3632 -19243 3644 -19209
rect 3586 -19277 3644 -19243
rect 3586 -19311 3598 -19277
rect 3632 -19311 3644 -19277
rect 3586 -19345 3644 -19311
rect 3586 -19379 3598 -19345
rect 3632 -19379 3644 -19345
rect 3586 -19413 3644 -19379
rect 3586 -19447 3598 -19413
rect 3632 -19447 3644 -19413
rect 3586 -19481 3644 -19447
rect 3586 -19515 3598 -19481
rect 3632 -19515 3644 -19481
rect 3586 -19549 3644 -19515
rect 3586 -19583 3598 -19549
rect 3632 -19583 3644 -19549
rect 3586 -19617 3644 -19583
rect 3586 -19651 3598 -19617
rect 3632 -19651 3644 -19617
rect 3586 -19685 3644 -19651
rect 3586 -19719 3598 -19685
rect 3632 -19719 3644 -19685
rect 3586 -19764 3644 -19719
rect 4604 -19209 4662 -19164
rect 4604 -19243 4616 -19209
rect 4650 -19243 4662 -19209
rect 4604 -19277 4662 -19243
rect 4604 -19311 4616 -19277
rect 4650 -19311 4662 -19277
rect 4604 -19345 4662 -19311
rect 4604 -19379 4616 -19345
rect 4650 -19379 4662 -19345
rect 4604 -19413 4662 -19379
rect 4604 -19447 4616 -19413
rect 4650 -19447 4662 -19413
rect 4604 -19481 4662 -19447
rect 4604 -19515 4616 -19481
rect 4650 -19515 4662 -19481
rect 4604 -19549 4662 -19515
rect 4604 -19583 4616 -19549
rect 4650 -19583 4662 -19549
rect 4604 -19617 4662 -19583
rect 4604 -19651 4616 -19617
rect 4650 -19651 4662 -19617
rect 4604 -19685 4662 -19651
rect 4604 -19719 4616 -19685
rect 4650 -19719 4662 -19685
rect 4604 -19764 4662 -19719
rect 5622 -19209 5680 -19164
rect 5622 -19243 5634 -19209
rect 5668 -19243 5680 -19209
rect 5622 -19277 5680 -19243
rect 5622 -19311 5634 -19277
rect 5668 -19311 5680 -19277
rect 5622 -19345 5680 -19311
rect 5622 -19379 5634 -19345
rect 5668 -19379 5680 -19345
rect 5622 -19413 5680 -19379
rect 5622 -19447 5634 -19413
rect 5668 -19447 5680 -19413
rect 5622 -19481 5680 -19447
rect 5622 -19515 5634 -19481
rect 5668 -19515 5680 -19481
rect 5622 -19549 5680 -19515
rect 5622 -19583 5634 -19549
rect 5668 -19583 5680 -19549
rect 5622 -19617 5680 -19583
rect 5622 -19651 5634 -19617
rect 5668 -19651 5680 -19617
rect 5622 -19685 5680 -19651
rect 5622 -19719 5634 -19685
rect 5668 -19719 5680 -19685
rect 5622 -19764 5680 -19719
rect 6640 -19209 6698 -19164
rect 6640 -19243 6652 -19209
rect 6686 -19243 6698 -19209
rect 6640 -19277 6698 -19243
rect 6640 -19311 6652 -19277
rect 6686 -19311 6698 -19277
rect 6640 -19345 6698 -19311
rect 6640 -19379 6652 -19345
rect 6686 -19379 6698 -19345
rect 6640 -19413 6698 -19379
rect 6640 -19447 6652 -19413
rect 6686 -19447 6698 -19413
rect 6640 -19481 6698 -19447
rect 6640 -19515 6652 -19481
rect 6686 -19515 6698 -19481
rect 6640 -19549 6698 -19515
rect 6640 -19583 6652 -19549
rect 6686 -19583 6698 -19549
rect 6640 -19617 6698 -19583
rect 6640 -19651 6652 -19617
rect 6686 -19651 6698 -19617
rect 6640 -19685 6698 -19651
rect 6640 -19719 6652 -19685
rect 6686 -19719 6698 -19685
rect 6640 -19764 6698 -19719
rect 7658 -19209 7716 -19164
rect 7658 -19243 7670 -19209
rect 7704 -19243 7716 -19209
rect 7658 -19277 7716 -19243
rect 7658 -19311 7670 -19277
rect 7704 -19311 7716 -19277
rect 7658 -19345 7716 -19311
rect 7658 -19379 7670 -19345
rect 7704 -19379 7716 -19345
rect 7658 -19413 7716 -19379
rect 7658 -19447 7670 -19413
rect 7704 -19447 7716 -19413
rect 7658 -19481 7716 -19447
rect 7658 -19515 7670 -19481
rect 7704 -19515 7716 -19481
rect 7658 -19549 7716 -19515
rect 7658 -19583 7670 -19549
rect 7704 -19583 7716 -19549
rect 7658 -19617 7716 -19583
rect 7658 -19651 7670 -19617
rect 7704 -19651 7716 -19617
rect 7658 -19685 7716 -19651
rect 7658 -19719 7670 -19685
rect 7704 -19719 7716 -19685
rect 7658 -19764 7716 -19719
rect 8676 -19209 8734 -19164
rect 8676 -19243 8688 -19209
rect 8722 -19243 8734 -19209
rect 8676 -19277 8734 -19243
rect 8676 -19311 8688 -19277
rect 8722 -19311 8734 -19277
rect 8676 -19345 8734 -19311
rect 8676 -19379 8688 -19345
rect 8722 -19379 8734 -19345
rect 8676 -19413 8734 -19379
rect 8676 -19447 8688 -19413
rect 8722 -19447 8734 -19413
rect 8676 -19481 8734 -19447
rect 8676 -19515 8688 -19481
rect 8722 -19515 8734 -19481
rect 8676 -19549 8734 -19515
rect 8676 -19583 8688 -19549
rect 8722 -19583 8734 -19549
rect 8676 -19617 8734 -19583
rect 8676 -19651 8688 -19617
rect 8722 -19651 8734 -19617
rect 8676 -19685 8734 -19651
rect 8676 -19719 8688 -19685
rect 8722 -19719 8734 -19685
rect 8676 -19764 8734 -19719
rect 9694 -19209 9752 -19164
rect 9694 -19243 9706 -19209
rect 9740 -19243 9752 -19209
rect 9694 -19277 9752 -19243
rect 9694 -19311 9706 -19277
rect 9740 -19311 9752 -19277
rect 9694 -19345 9752 -19311
rect 9694 -19379 9706 -19345
rect 9740 -19379 9752 -19345
rect 9694 -19413 9752 -19379
rect 9694 -19447 9706 -19413
rect 9740 -19447 9752 -19413
rect 9694 -19481 9752 -19447
rect 9694 -19515 9706 -19481
rect 9740 -19515 9752 -19481
rect 9694 -19549 9752 -19515
rect 9694 -19583 9706 -19549
rect 9740 -19583 9752 -19549
rect 9694 -19617 9752 -19583
rect 9694 -19651 9706 -19617
rect 9740 -19651 9752 -19617
rect 9694 -19685 9752 -19651
rect 9694 -19719 9706 -19685
rect 9740 -19719 9752 -19685
rect 9694 -19764 9752 -19719
rect 10712 -19209 10770 -19164
rect 10712 -19243 10724 -19209
rect 10758 -19243 10770 -19209
rect 10712 -19277 10770 -19243
rect 10712 -19311 10724 -19277
rect 10758 -19311 10770 -19277
rect 10712 -19345 10770 -19311
rect 10712 -19379 10724 -19345
rect 10758 -19379 10770 -19345
rect 10712 -19413 10770 -19379
rect 10712 -19447 10724 -19413
rect 10758 -19447 10770 -19413
rect 10712 -19481 10770 -19447
rect 10712 -19515 10724 -19481
rect 10758 -19515 10770 -19481
rect 10712 -19549 10770 -19515
rect 10712 -19583 10724 -19549
rect 10758 -19583 10770 -19549
rect 10712 -19617 10770 -19583
rect 10712 -19651 10724 -19617
rect 10758 -19651 10770 -19617
rect 10712 -19685 10770 -19651
rect 10712 -19719 10724 -19685
rect 10758 -19719 10770 -19685
rect 10712 -19764 10770 -19719
rect 11730 -19209 11788 -19164
rect 11730 -19243 11742 -19209
rect 11776 -19243 11788 -19209
rect 11730 -19277 11788 -19243
rect 11730 -19311 11742 -19277
rect 11776 -19311 11788 -19277
rect 11730 -19345 11788 -19311
rect 11730 -19379 11742 -19345
rect 11776 -19379 11788 -19345
rect 11730 -19413 11788 -19379
rect 11730 -19447 11742 -19413
rect 11776 -19447 11788 -19413
rect 11730 -19481 11788 -19447
rect 11730 -19515 11742 -19481
rect 11776 -19515 11788 -19481
rect 11730 -19549 11788 -19515
rect 11730 -19583 11742 -19549
rect 11776 -19583 11788 -19549
rect 11730 -19617 11788 -19583
rect 11730 -19651 11742 -19617
rect 11776 -19651 11788 -19617
rect 11730 -19685 11788 -19651
rect 11730 -19719 11742 -19685
rect 11776 -19719 11788 -19685
rect 11730 -19764 11788 -19719
rect 12748 -19209 12806 -19164
rect 12748 -19243 12760 -19209
rect 12794 -19243 12806 -19209
rect 12748 -19277 12806 -19243
rect 12748 -19311 12760 -19277
rect 12794 -19311 12806 -19277
rect 12748 -19345 12806 -19311
rect 12748 -19379 12760 -19345
rect 12794 -19379 12806 -19345
rect 12748 -19413 12806 -19379
rect 12748 -19447 12760 -19413
rect 12794 -19447 12806 -19413
rect 12748 -19481 12806 -19447
rect 12748 -19515 12760 -19481
rect 12794 -19515 12806 -19481
rect 12748 -19549 12806 -19515
rect 12748 -19583 12760 -19549
rect 12794 -19583 12806 -19549
rect 12748 -19617 12806 -19583
rect 12748 -19651 12760 -19617
rect 12794 -19651 12806 -19617
rect 12748 -19685 12806 -19651
rect 12748 -19719 12760 -19685
rect 12794 -19719 12806 -19685
rect 12748 -19764 12806 -19719
rect 13766 -19209 13824 -19164
rect 13766 -19243 13778 -19209
rect 13812 -19243 13824 -19209
rect 13766 -19277 13824 -19243
rect 13766 -19311 13778 -19277
rect 13812 -19311 13824 -19277
rect 13766 -19345 13824 -19311
rect 13766 -19379 13778 -19345
rect 13812 -19379 13824 -19345
rect 13766 -19413 13824 -19379
rect 13766 -19447 13778 -19413
rect 13812 -19447 13824 -19413
rect 13766 -19481 13824 -19447
rect 13766 -19515 13778 -19481
rect 13812 -19515 13824 -19481
rect 13766 -19549 13824 -19515
rect 13766 -19583 13778 -19549
rect 13812 -19583 13824 -19549
rect 13766 -19617 13824 -19583
rect 13766 -19651 13778 -19617
rect 13812 -19651 13824 -19617
rect 13766 -19685 13824 -19651
rect 13766 -19719 13778 -19685
rect 13812 -19719 13824 -19685
rect 13766 -19764 13824 -19719
rect 14784 -19209 14842 -19164
rect 14784 -19243 14796 -19209
rect 14830 -19243 14842 -19209
rect 14784 -19277 14842 -19243
rect 14784 -19311 14796 -19277
rect 14830 -19311 14842 -19277
rect 14784 -19345 14842 -19311
rect 14784 -19379 14796 -19345
rect 14830 -19379 14842 -19345
rect 14784 -19413 14842 -19379
rect 14784 -19447 14796 -19413
rect 14830 -19447 14842 -19413
rect 14784 -19481 14842 -19447
rect 14784 -19515 14796 -19481
rect 14830 -19515 14842 -19481
rect 14784 -19549 14842 -19515
rect 14784 -19583 14796 -19549
rect 14830 -19583 14842 -19549
rect 14784 -19617 14842 -19583
rect 14784 -19651 14796 -19617
rect 14830 -19651 14842 -19617
rect 14784 -19685 14842 -19651
rect 14784 -19719 14796 -19685
rect 14830 -19719 14842 -19685
rect 14784 -19764 14842 -19719
rect 15802 -19209 15860 -19164
rect 15802 -19243 15814 -19209
rect 15848 -19243 15860 -19209
rect 15802 -19277 15860 -19243
rect 15802 -19311 15814 -19277
rect 15848 -19311 15860 -19277
rect 15802 -19345 15860 -19311
rect 15802 -19379 15814 -19345
rect 15848 -19379 15860 -19345
rect 15802 -19413 15860 -19379
rect 15802 -19447 15814 -19413
rect 15848 -19447 15860 -19413
rect 15802 -19481 15860 -19447
rect 15802 -19515 15814 -19481
rect 15848 -19515 15860 -19481
rect 15802 -19549 15860 -19515
rect 15802 -19583 15814 -19549
rect 15848 -19583 15860 -19549
rect 15802 -19617 15860 -19583
rect 15802 -19651 15814 -19617
rect 15848 -19651 15860 -19617
rect 15802 -19685 15860 -19651
rect 15802 -19719 15814 -19685
rect 15848 -19719 15860 -19685
rect 15802 -19764 15860 -19719
rect 16820 -19209 16878 -19164
rect 16820 -19243 16832 -19209
rect 16866 -19243 16878 -19209
rect 16820 -19277 16878 -19243
rect 16820 -19311 16832 -19277
rect 16866 -19311 16878 -19277
rect 16820 -19345 16878 -19311
rect 16820 -19379 16832 -19345
rect 16866 -19379 16878 -19345
rect 16820 -19413 16878 -19379
rect 16820 -19447 16832 -19413
rect 16866 -19447 16878 -19413
rect 16820 -19481 16878 -19447
rect 16820 -19515 16832 -19481
rect 16866 -19515 16878 -19481
rect 16820 -19549 16878 -19515
rect 16820 -19583 16832 -19549
rect 16866 -19583 16878 -19549
rect 16820 -19617 16878 -19583
rect 16820 -19651 16832 -19617
rect 16866 -19651 16878 -19617
rect 16820 -19685 16878 -19651
rect 16820 -19719 16832 -19685
rect 16866 -19719 16878 -19685
rect 16820 -19764 16878 -19719
rect 17838 -19209 17896 -19164
rect 17838 -19243 17850 -19209
rect 17884 -19243 17896 -19209
rect 17838 -19277 17896 -19243
rect 17838 -19311 17850 -19277
rect 17884 -19311 17896 -19277
rect 17838 -19345 17896 -19311
rect 17838 -19379 17850 -19345
rect 17884 -19379 17896 -19345
rect 17838 -19413 17896 -19379
rect 17838 -19447 17850 -19413
rect 17884 -19447 17896 -19413
rect 17838 -19481 17896 -19447
rect 17838 -19515 17850 -19481
rect 17884 -19515 17896 -19481
rect 17838 -19549 17896 -19515
rect 17838 -19583 17850 -19549
rect 17884 -19583 17896 -19549
rect 17838 -19617 17896 -19583
rect 17838 -19651 17850 -19617
rect 17884 -19651 17896 -19617
rect 17838 -19685 17896 -19651
rect 17838 -19719 17850 -19685
rect 17884 -19719 17896 -19685
rect 17838 -19764 17896 -19719
rect 18856 -19209 18914 -19164
rect 18856 -19243 18868 -19209
rect 18902 -19243 18914 -19209
rect 18856 -19277 18914 -19243
rect 18856 -19311 18868 -19277
rect 18902 -19311 18914 -19277
rect 18856 -19345 18914 -19311
rect 18856 -19379 18868 -19345
rect 18902 -19379 18914 -19345
rect 18856 -19413 18914 -19379
rect 18856 -19447 18868 -19413
rect 18902 -19447 18914 -19413
rect 18856 -19481 18914 -19447
rect 18856 -19515 18868 -19481
rect 18902 -19515 18914 -19481
rect 18856 -19549 18914 -19515
rect 18856 -19583 18868 -19549
rect 18902 -19583 18914 -19549
rect 18856 -19617 18914 -19583
rect 18856 -19651 18868 -19617
rect 18902 -19651 18914 -19617
rect 18856 -19685 18914 -19651
rect 18856 -19719 18868 -19685
rect 18902 -19719 18914 -19685
rect 18856 -19764 18914 -19719
rect 19874 -19209 19932 -19164
rect 19874 -19243 19886 -19209
rect 19920 -19243 19932 -19209
rect 19874 -19277 19932 -19243
rect 19874 -19311 19886 -19277
rect 19920 -19311 19932 -19277
rect 19874 -19345 19932 -19311
rect 19874 -19379 19886 -19345
rect 19920 -19379 19932 -19345
rect 19874 -19413 19932 -19379
rect 19874 -19447 19886 -19413
rect 19920 -19447 19932 -19413
rect 19874 -19481 19932 -19447
rect 19874 -19515 19886 -19481
rect 19920 -19515 19932 -19481
rect 19874 -19549 19932 -19515
rect 19874 -19583 19886 -19549
rect 19920 -19583 19932 -19549
rect 19874 -19617 19932 -19583
rect 19874 -19651 19886 -19617
rect 19920 -19651 19932 -19617
rect 19874 -19685 19932 -19651
rect 19874 -19719 19886 -19685
rect 19920 -19719 19932 -19685
rect 19874 -19764 19932 -19719
rect 20892 -19209 20950 -19164
rect 20892 -19243 20904 -19209
rect 20938 -19243 20950 -19209
rect 20892 -19277 20950 -19243
rect 20892 -19311 20904 -19277
rect 20938 -19311 20950 -19277
rect 20892 -19345 20950 -19311
rect 20892 -19379 20904 -19345
rect 20938 -19379 20950 -19345
rect 20892 -19413 20950 -19379
rect 20892 -19447 20904 -19413
rect 20938 -19447 20950 -19413
rect 20892 -19481 20950 -19447
rect 20892 -19515 20904 -19481
rect 20938 -19515 20950 -19481
rect 20892 -19549 20950 -19515
rect 20892 -19583 20904 -19549
rect 20938 -19583 20950 -19549
rect 20892 -19617 20950 -19583
rect 20892 -19651 20904 -19617
rect 20938 -19651 20950 -19617
rect 20892 -19685 20950 -19651
rect 20892 -19719 20904 -19685
rect 20938 -19719 20950 -19685
rect 20892 -19764 20950 -19719
rect 21910 -19209 21968 -19164
rect 21910 -19243 21922 -19209
rect 21956 -19243 21968 -19209
rect 21910 -19277 21968 -19243
rect 21910 -19311 21922 -19277
rect 21956 -19311 21968 -19277
rect 21910 -19345 21968 -19311
rect 21910 -19379 21922 -19345
rect 21956 -19379 21968 -19345
rect 21910 -19413 21968 -19379
rect 21910 -19447 21922 -19413
rect 21956 -19447 21968 -19413
rect 21910 -19481 21968 -19447
rect 21910 -19515 21922 -19481
rect 21956 -19515 21968 -19481
rect 21910 -19549 21968 -19515
rect 21910 -19583 21922 -19549
rect 21956 -19583 21968 -19549
rect 21910 -19617 21968 -19583
rect 21910 -19651 21922 -19617
rect 21956 -19651 21968 -19617
rect 21910 -19685 21968 -19651
rect 21910 -19719 21922 -19685
rect 21956 -19719 21968 -19685
rect 21910 -19764 21968 -19719
rect 22928 -19209 22986 -19164
rect 22928 -19243 22940 -19209
rect 22974 -19243 22986 -19209
rect 22928 -19277 22986 -19243
rect 22928 -19311 22940 -19277
rect 22974 -19311 22986 -19277
rect 22928 -19345 22986 -19311
rect 22928 -19379 22940 -19345
rect 22974 -19379 22986 -19345
rect 22928 -19413 22986 -19379
rect 22928 -19447 22940 -19413
rect 22974 -19447 22986 -19413
rect 22928 -19481 22986 -19447
rect 22928 -19515 22940 -19481
rect 22974 -19515 22986 -19481
rect 22928 -19549 22986 -19515
rect 22928 -19583 22940 -19549
rect 22974 -19583 22986 -19549
rect 22928 -19617 22986 -19583
rect 22928 -19651 22940 -19617
rect 22974 -19651 22986 -19617
rect 22928 -19685 22986 -19651
rect 22928 -19719 22940 -19685
rect 22974 -19719 22986 -19685
rect 22928 -19764 22986 -19719
rect 2568 -20443 2626 -20398
rect 2568 -20477 2580 -20443
rect 2614 -20477 2626 -20443
rect 2568 -20511 2626 -20477
rect 2568 -20545 2580 -20511
rect 2614 -20545 2626 -20511
rect 2568 -20579 2626 -20545
rect 2568 -20613 2580 -20579
rect 2614 -20613 2626 -20579
rect 2568 -20647 2626 -20613
rect 2568 -20681 2580 -20647
rect 2614 -20681 2626 -20647
rect 2568 -20715 2626 -20681
rect 2568 -20749 2580 -20715
rect 2614 -20749 2626 -20715
rect 2568 -20783 2626 -20749
rect 2568 -20817 2580 -20783
rect 2614 -20817 2626 -20783
rect 2568 -20851 2626 -20817
rect 2568 -20885 2580 -20851
rect 2614 -20885 2626 -20851
rect 2568 -20919 2626 -20885
rect 2568 -20953 2580 -20919
rect 2614 -20953 2626 -20919
rect 2568 -20998 2626 -20953
rect 3586 -20443 3644 -20398
rect 3586 -20477 3598 -20443
rect 3632 -20477 3644 -20443
rect 3586 -20511 3644 -20477
rect 3586 -20545 3598 -20511
rect 3632 -20545 3644 -20511
rect 3586 -20579 3644 -20545
rect 3586 -20613 3598 -20579
rect 3632 -20613 3644 -20579
rect 3586 -20647 3644 -20613
rect 3586 -20681 3598 -20647
rect 3632 -20681 3644 -20647
rect 3586 -20715 3644 -20681
rect 3586 -20749 3598 -20715
rect 3632 -20749 3644 -20715
rect 3586 -20783 3644 -20749
rect 3586 -20817 3598 -20783
rect 3632 -20817 3644 -20783
rect 3586 -20851 3644 -20817
rect 3586 -20885 3598 -20851
rect 3632 -20885 3644 -20851
rect 3586 -20919 3644 -20885
rect 3586 -20953 3598 -20919
rect 3632 -20953 3644 -20919
rect 3586 -20998 3644 -20953
rect 4604 -20443 4662 -20398
rect 4604 -20477 4616 -20443
rect 4650 -20477 4662 -20443
rect 4604 -20511 4662 -20477
rect 4604 -20545 4616 -20511
rect 4650 -20545 4662 -20511
rect 4604 -20579 4662 -20545
rect 4604 -20613 4616 -20579
rect 4650 -20613 4662 -20579
rect 4604 -20647 4662 -20613
rect 4604 -20681 4616 -20647
rect 4650 -20681 4662 -20647
rect 4604 -20715 4662 -20681
rect 4604 -20749 4616 -20715
rect 4650 -20749 4662 -20715
rect 4604 -20783 4662 -20749
rect 4604 -20817 4616 -20783
rect 4650 -20817 4662 -20783
rect 4604 -20851 4662 -20817
rect 4604 -20885 4616 -20851
rect 4650 -20885 4662 -20851
rect 4604 -20919 4662 -20885
rect 4604 -20953 4616 -20919
rect 4650 -20953 4662 -20919
rect 4604 -20998 4662 -20953
rect 5622 -20443 5680 -20398
rect 5622 -20477 5634 -20443
rect 5668 -20477 5680 -20443
rect 5622 -20511 5680 -20477
rect 5622 -20545 5634 -20511
rect 5668 -20545 5680 -20511
rect 5622 -20579 5680 -20545
rect 5622 -20613 5634 -20579
rect 5668 -20613 5680 -20579
rect 5622 -20647 5680 -20613
rect 5622 -20681 5634 -20647
rect 5668 -20681 5680 -20647
rect 5622 -20715 5680 -20681
rect 5622 -20749 5634 -20715
rect 5668 -20749 5680 -20715
rect 5622 -20783 5680 -20749
rect 5622 -20817 5634 -20783
rect 5668 -20817 5680 -20783
rect 5622 -20851 5680 -20817
rect 5622 -20885 5634 -20851
rect 5668 -20885 5680 -20851
rect 5622 -20919 5680 -20885
rect 5622 -20953 5634 -20919
rect 5668 -20953 5680 -20919
rect 5622 -20998 5680 -20953
rect 6640 -20443 6698 -20398
rect 6640 -20477 6652 -20443
rect 6686 -20477 6698 -20443
rect 6640 -20511 6698 -20477
rect 6640 -20545 6652 -20511
rect 6686 -20545 6698 -20511
rect 6640 -20579 6698 -20545
rect 6640 -20613 6652 -20579
rect 6686 -20613 6698 -20579
rect 6640 -20647 6698 -20613
rect 6640 -20681 6652 -20647
rect 6686 -20681 6698 -20647
rect 6640 -20715 6698 -20681
rect 6640 -20749 6652 -20715
rect 6686 -20749 6698 -20715
rect 6640 -20783 6698 -20749
rect 6640 -20817 6652 -20783
rect 6686 -20817 6698 -20783
rect 6640 -20851 6698 -20817
rect 6640 -20885 6652 -20851
rect 6686 -20885 6698 -20851
rect 6640 -20919 6698 -20885
rect 6640 -20953 6652 -20919
rect 6686 -20953 6698 -20919
rect 6640 -20998 6698 -20953
rect 7658 -20443 7716 -20398
rect 7658 -20477 7670 -20443
rect 7704 -20477 7716 -20443
rect 7658 -20511 7716 -20477
rect 7658 -20545 7670 -20511
rect 7704 -20545 7716 -20511
rect 7658 -20579 7716 -20545
rect 7658 -20613 7670 -20579
rect 7704 -20613 7716 -20579
rect 7658 -20647 7716 -20613
rect 7658 -20681 7670 -20647
rect 7704 -20681 7716 -20647
rect 7658 -20715 7716 -20681
rect 7658 -20749 7670 -20715
rect 7704 -20749 7716 -20715
rect 7658 -20783 7716 -20749
rect 7658 -20817 7670 -20783
rect 7704 -20817 7716 -20783
rect 7658 -20851 7716 -20817
rect 7658 -20885 7670 -20851
rect 7704 -20885 7716 -20851
rect 7658 -20919 7716 -20885
rect 7658 -20953 7670 -20919
rect 7704 -20953 7716 -20919
rect 7658 -20998 7716 -20953
rect 8676 -20443 8734 -20398
rect 8676 -20477 8688 -20443
rect 8722 -20477 8734 -20443
rect 8676 -20511 8734 -20477
rect 8676 -20545 8688 -20511
rect 8722 -20545 8734 -20511
rect 8676 -20579 8734 -20545
rect 8676 -20613 8688 -20579
rect 8722 -20613 8734 -20579
rect 8676 -20647 8734 -20613
rect 8676 -20681 8688 -20647
rect 8722 -20681 8734 -20647
rect 8676 -20715 8734 -20681
rect 8676 -20749 8688 -20715
rect 8722 -20749 8734 -20715
rect 8676 -20783 8734 -20749
rect 8676 -20817 8688 -20783
rect 8722 -20817 8734 -20783
rect 8676 -20851 8734 -20817
rect 8676 -20885 8688 -20851
rect 8722 -20885 8734 -20851
rect 8676 -20919 8734 -20885
rect 8676 -20953 8688 -20919
rect 8722 -20953 8734 -20919
rect 8676 -20998 8734 -20953
rect 9694 -20443 9752 -20398
rect 9694 -20477 9706 -20443
rect 9740 -20477 9752 -20443
rect 9694 -20511 9752 -20477
rect 9694 -20545 9706 -20511
rect 9740 -20545 9752 -20511
rect 9694 -20579 9752 -20545
rect 9694 -20613 9706 -20579
rect 9740 -20613 9752 -20579
rect 9694 -20647 9752 -20613
rect 9694 -20681 9706 -20647
rect 9740 -20681 9752 -20647
rect 9694 -20715 9752 -20681
rect 9694 -20749 9706 -20715
rect 9740 -20749 9752 -20715
rect 9694 -20783 9752 -20749
rect 9694 -20817 9706 -20783
rect 9740 -20817 9752 -20783
rect 9694 -20851 9752 -20817
rect 9694 -20885 9706 -20851
rect 9740 -20885 9752 -20851
rect 9694 -20919 9752 -20885
rect 9694 -20953 9706 -20919
rect 9740 -20953 9752 -20919
rect 9694 -20998 9752 -20953
rect 10712 -20443 10770 -20398
rect 10712 -20477 10724 -20443
rect 10758 -20477 10770 -20443
rect 10712 -20511 10770 -20477
rect 10712 -20545 10724 -20511
rect 10758 -20545 10770 -20511
rect 10712 -20579 10770 -20545
rect 10712 -20613 10724 -20579
rect 10758 -20613 10770 -20579
rect 10712 -20647 10770 -20613
rect 10712 -20681 10724 -20647
rect 10758 -20681 10770 -20647
rect 10712 -20715 10770 -20681
rect 10712 -20749 10724 -20715
rect 10758 -20749 10770 -20715
rect 10712 -20783 10770 -20749
rect 10712 -20817 10724 -20783
rect 10758 -20817 10770 -20783
rect 10712 -20851 10770 -20817
rect 10712 -20885 10724 -20851
rect 10758 -20885 10770 -20851
rect 10712 -20919 10770 -20885
rect 10712 -20953 10724 -20919
rect 10758 -20953 10770 -20919
rect 10712 -20998 10770 -20953
rect 11730 -20443 11788 -20398
rect 11730 -20477 11742 -20443
rect 11776 -20477 11788 -20443
rect 11730 -20511 11788 -20477
rect 11730 -20545 11742 -20511
rect 11776 -20545 11788 -20511
rect 11730 -20579 11788 -20545
rect 11730 -20613 11742 -20579
rect 11776 -20613 11788 -20579
rect 11730 -20647 11788 -20613
rect 11730 -20681 11742 -20647
rect 11776 -20681 11788 -20647
rect 11730 -20715 11788 -20681
rect 11730 -20749 11742 -20715
rect 11776 -20749 11788 -20715
rect 11730 -20783 11788 -20749
rect 11730 -20817 11742 -20783
rect 11776 -20817 11788 -20783
rect 11730 -20851 11788 -20817
rect 11730 -20885 11742 -20851
rect 11776 -20885 11788 -20851
rect 11730 -20919 11788 -20885
rect 11730 -20953 11742 -20919
rect 11776 -20953 11788 -20919
rect 11730 -20998 11788 -20953
rect 12748 -20443 12806 -20398
rect 12748 -20477 12760 -20443
rect 12794 -20477 12806 -20443
rect 12748 -20511 12806 -20477
rect 12748 -20545 12760 -20511
rect 12794 -20545 12806 -20511
rect 12748 -20579 12806 -20545
rect 12748 -20613 12760 -20579
rect 12794 -20613 12806 -20579
rect 12748 -20647 12806 -20613
rect 12748 -20681 12760 -20647
rect 12794 -20681 12806 -20647
rect 12748 -20715 12806 -20681
rect 12748 -20749 12760 -20715
rect 12794 -20749 12806 -20715
rect 12748 -20783 12806 -20749
rect 12748 -20817 12760 -20783
rect 12794 -20817 12806 -20783
rect 12748 -20851 12806 -20817
rect 12748 -20885 12760 -20851
rect 12794 -20885 12806 -20851
rect 12748 -20919 12806 -20885
rect 12748 -20953 12760 -20919
rect 12794 -20953 12806 -20919
rect 12748 -20998 12806 -20953
rect 13766 -20443 13824 -20398
rect 13766 -20477 13778 -20443
rect 13812 -20477 13824 -20443
rect 13766 -20511 13824 -20477
rect 13766 -20545 13778 -20511
rect 13812 -20545 13824 -20511
rect 13766 -20579 13824 -20545
rect 13766 -20613 13778 -20579
rect 13812 -20613 13824 -20579
rect 13766 -20647 13824 -20613
rect 13766 -20681 13778 -20647
rect 13812 -20681 13824 -20647
rect 13766 -20715 13824 -20681
rect 13766 -20749 13778 -20715
rect 13812 -20749 13824 -20715
rect 13766 -20783 13824 -20749
rect 13766 -20817 13778 -20783
rect 13812 -20817 13824 -20783
rect 13766 -20851 13824 -20817
rect 13766 -20885 13778 -20851
rect 13812 -20885 13824 -20851
rect 13766 -20919 13824 -20885
rect 13766 -20953 13778 -20919
rect 13812 -20953 13824 -20919
rect 13766 -20998 13824 -20953
rect 14784 -20443 14842 -20398
rect 14784 -20477 14796 -20443
rect 14830 -20477 14842 -20443
rect 14784 -20511 14842 -20477
rect 14784 -20545 14796 -20511
rect 14830 -20545 14842 -20511
rect 14784 -20579 14842 -20545
rect 14784 -20613 14796 -20579
rect 14830 -20613 14842 -20579
rect 14784 -20647 14842 -20613
rect 14784 -20681 14796 -20647
rect 14830 -20681 14842 -20647
rect 14784 -20715 14842 -20681
rect 14784 -20749 14796 -20715
rect 14830 -20749 14842 -20715
rect 14784 -20783 14842 -20749
rect 14784 -20817 14796 -20783
rect 14830 -20817 14842 -20783
rect 14784 -20851 14842 -20817
rect 14784 -20885 14796 -20851
rect 14830 -20885 14842 -20851
rect 14784 -20919 14842 -20885
rect 14784 -20953 14796 -20919
rect 14830 -20953 14842 -20919
rect 14784 -20998 14842 -20953
rect 15802 -20443 15860 -20398
rect 15802 -20477 15814 -20443
rect 15848 -20477 15860 -20443
rect 15802 -20511 15860 -20477
rect 15802 -20545 15814 -20511
rect 15848 -20545 15860 -20511
rect 15802 -20579 15860 -20545
rect 15802 -20613 15814 -20579
rect 15848 -20613 15860 -20579
rect 15802 -20647 15860 -20613
rect 15802 -20681 15814 -20647
rect 15848 -20681 15860 -20647
rect 15802 -20715 15860 -20681
rect 15802 -20749 15814 -20715
rect 15848 -20749 15860 -20715
rect 15802 -20783 15860 -20749
rect 15802 -20817 15814 -20783
rect 15848 -20817 15860 -20783
rect 15802 -20851 15860 -20817
rect 15802 -20885 15814 -20851
rect 15848 -20885 15860 -20851
rect 15802 -20919 15860 -20885
rect 15802 -20953 15814 -20919
rect 15848 -20953 15860 -20919
rect 15802 -20998 15860 -20953
rect 16820 -20443 16878 -20398
rect 16820 -20477 16832 -20443
rect 16866 -20477 16878 -20443
rect 16820 -20511 16878 -20477
rect 16820 -20545 16832 -20511
rect 16866 -20545 16878 -20511
rect 16820 -20579 16878 -20545
rect 16820 -20613 16832 -20579
rect 16866 -20613 16878 -20579
rect 16820 -20647 16878 -20613
rect 16820 -20681 16832 -20647
rect 16866 -20681 16878 -20647
rect 16820 -20715 16878 -20681
rect 16820 -20749 16832 -20715
rect 16866 -20749 16878 -20715
rect 16820 -20783 16878 -20749
rect 16820 -20817 16832 -20783
rect 16866 -20817 16878 -20783
rect 16820 -20851 16878 -20817
rect 16820 -20885 16832 -20851
rect 16866 -20885 16878 -20851
rect 16820 -20919 16878 -20885
rect 16820 -20953 16832 -20919
rect 16866 -20953 16878 -20919
rect 16820 -20998 16878 -20953
rect 17838 -20443 17896 -20398
rect 17838 -20477 17850 -20443
rect 17884 -20477 17896 -20443
rect 17838 -20511 17896 -20477
rect 17838 -20545 17850 -20511
rect 17884 -20545 17896 -20511
rect 17838 -20579 17896 -20545
rect 17838 -20613 17850 -20579
rect 17884 -20613 17896 -20579
rect 17838 -20647 17896 -20613
rect 17838 -20681 17850 -20647
rect 17884 -20681 17896 -20647
rect 17838 -20715 17896 -20681
rect 17838 -20749 17850 -20715
rect 17884 -20749 17896 -20715
rect 17838 -20783 17896 -20749
rect 17838 -20817 17850 -20783
rect 17884 -20817 17896 -20783
rect 17838 -20851 17896 -20817
rect 17838 -20885 17850 -20851
rect 17884 -20885 17896 -20851
rect 17838 -20919 17896 -20885
rect 17838 -20953 17850 -20919
rect 17884 -20953 17896 -20919
rect 17838 -20998 17896 -20953
rect 18856 -20443 18914 -20398
rect 18856 -20477 18868 -20443
rect 18902 -20477 18914 -20443
rect 18856 -20511 18914 -20477
rect 18856 -20545 18868 -20511
rect 18902 -20545 18914 -20511
rect 18856 -20579 18914 -20545
rect 18856 -20613 18868 -20579
rect 18902 -20613 18914 -20579
rect 18856 -20647 18914 -20613
rect 18856 -20681 18868 -20647
rect 18902 -20681 18914 -20647
rect 18856 -20715 18914 -20681
rect 18856 -20749 18868 -20715
rect 18902 -20749 18914 -20715
rect 18856 -20783 18914 -20749
rect 18856 -20817 18868 -20783
rect 18902 -20817 18914 -20783
rect 18856 -20851 18914 -20817
rect 18856 -20885 18868 -20851
rect 18902 -20885 18914 -20851
rect 18856 -20919 18914 -20885
rect 18856 -20953 18868 -20919
rect 18902 -20953 18914 -20919
rect 18856 -20998 18914 -20953
rect 19874 -20443 19932 -20398
rect 19874 -20477 19886 -20443
rect 19920 -20477 19932 -20443
rect 19874 -20511 19932 -20477
rect 19874 -20545 19886 -20511
rect 19920 -20545 19932 -20511
rect 19874 -20579 19932 -20545
rect 19874 -20613 19886 -20579
rect 19920 -20613 19932 -20579
rect 19874 -20647 19932 -20613
rect 19874 -20681 19886 -20647
rect 19920 -20681 19932 -20647
rect 19874 -20715 19932 -20681
rect 19874 -20749 19886 -20715
rect 19920 -20749 19932 -20715
rect 19874 -20783 19932 -20749
rect 19874 -20817 19886 -20783
rect 19920 -20817 19932 -20783
rect 19874 -20851 19932 -20817
rect 19874 -20885 19886 -20851
rect 19920 -20885 19932 -20851
rect 19874 -20919 19932 -20885
rect 19874 -20953 19886 -20919
rect 19920 -20953 19932 -20919
rect 19874 -20998 19932 -20953
rect 20892 -20443 20950 -20398
rect 20892 -20477 20904 -20443
rect 20938 -20477 20950 -20443
rect 20892 -20511 20950 -20477
rect 20892 -20545 20904 -20511
rect 20938 -20545 20950 -20511
rect 20892 -20579 20950 -20545
rect 20892 -20613 20904 -20579
rect 20938 -20613 20950 -20579
rect 20892 -20647 20950 -20613
rect 20892 -20681 20904 -20647
rect 20938 -20681 20950 -20647
rect 20892 -20715 20950 -20681
rect 20892 -20749 20904 -20715
rect 20938 -20749 20950 -20715
rect 20892 -20783 20950 -20749
rect 20892 -20817 20904 -20783
rect 20938 -20817 20950 -20783
rect 20892 -20851 20950 -20817
rect 20892 -20885 20904 -20851
rect 20938 -20885 20950 -20851
rect 20892 -20919 20950 -20885
rect 20892 -20953 20904 -20919
rect 20938 -20953 20950 -20919
rect 20892 -20998 20950 -20953
rect 21910 -20443 21968 -20398
rect 21910 -20477 21922 -20443
rect 21956 -20477 21968 -20443
rect 21910 -20511 21968 -20477
rect 21910 -20545 21922 -20511
rect 21956 -20545 21968 -20511
rect 21910 -20579 21968 -20545
rect 21910 -20613 21922 -20579
rect 21956 -20613 21968 -20579
rect 21910 -20647 21968 -20613
rect 21910 -20681 21922 -20647
rect 21956 -20681 21968 -20647
rect 21910 -20715 21968 -20681
rect 21910 -20749 21922 -20715
rect 21956 -20749 21968 -20715
rect 21910 -20783 21968 -20749
rect 21910 -20817 21922 -20783
rect 21956 -20817 21968 -20783
rect 21910 -20851 21968 -20817
rect 21910 -20885 21922 -20851
rect 21956 -20885 21968 -20851
rect 21910 -20919 21968 -20885
rect 21910 -20953 21922 -20919
rect 21956 -20953 21968 -20919
rect 21910 -20998 21968 -20953
rect 22928 -20443 22986 -20398
rect 22928 -20477 22940 -20443
rect 22974 -20477 22986 -20443
rect 22928 -20511 22986 -20477
rect 22928 -20545 22940 -20511
rect 22974 -20545 22986 -20511
rect 22928 -20579 22986 -20545
rect 22928 -20613 22940 -20579
rect 22974 -20613 22986 -20579
rect 22928 -20647 22986 -20613
rect 22928 -20681 22940 -20647
rect 22974 -20681 22986 -20647
rect 22928 -20715 22986 -20681
rect 22928 -20749 22940 -20715
rect 22974 -20749 22986 -20715
rect 22928 -20783 22986 -20749
rect 22928 -20817 22940 -20783
rect 22974 -20817 22986 -20783
rect 22928 -20851 22986 -20817
rect 22928 -20885 22940 -20851
rect 22974 -20885 22986 -20851
rect 22928 -20919 22986 -20885
rect 22928 -20953 22940 -20919
rect 22974 -20953 22986 -20919
rect 22928 -20998 22986 -20953
rect 2568 -21677 2626 -21632
rect 2568 -21711 2580 -21677
rect 2614 -21711 2626 -21677
rect 2568 -21745 2626 -21711
rect 2568 -21779 2580 -21745
rect 2614 -21779 2626 -21745
rect 2568 -21813 2626 -21779
rect 2568 -21847 2580 -21813
rect 2614 -21847 2626 -21813
rect 2568 -21881 2626 -21847
rect 2568 -21915 2580 -21881
rect 2614 -21915 2626 -21881
rect 2568 -21949 2626 -21915
rect 2568 -21983 2580 -21949
rect 2614 -21983 2626 -21949
rect 2568 -22017 2626 -21983
rect 2568 -22051 2580 -22017
rect 2614 -22051 2626 -22017
rect 2568 -22085 2626 -22051
rect 2568 -22119 2580 -22085
rect 2614 -22119 2626 -22085
rect 2568 -22153 2626 -22119
rect 2568 -22187 2580 -22153
rect 2614 -22187 2626 -22153
rect 2568 -22232 2626 -22187
rect 3586 -21677 3644 -21632
rect 3586 -21711 3598 -21677
rect 3632 -21711 3644 -21677
rect 3586 -21745 3644 -21711
rect 3586 -21779 3598 -21745
rect 3632 -21779 3644 -21745
rect 3586 -21813 3644 -21779
rect 3586 -21847 3598 -21813
rect 3632 -21847 3644 -21813
rect 3586 -21881 3644 -21847
rect 3586 -21915 3598 -21881
rect 3632 -21915 3644 -21881
rect 3586 -21949 3644 -21915
rect 3586 -21983 3598 -21949
rect 3632 -21983 3644 -21949
rect 3586 -22017 3644 -21983
rect 3586 -22051 3598 -22017
rect 3632 -22051 3644 -22017
rect 3586 -22085 3644 -22051
rect 3586 -22119 3598 -22085
rect 3632 -22119 3644 -22085
rect 3586 -22153 3644 -22119
rect 3586 -22187 3598 -22153
rect 3632 -22187 3644 -22153
rect 3586 -22232 3644 -22187
rect 4604 -21677 4662 -21632
rect 4604 -21711 4616 -21677
rect 4650 -21711 4662 -21677
rect 4604 -21745 4662 -21711
rect 4604 -21779 4616 -21745
rect 4650 -21779 4662 -21745
rect 4604 -21813 4662 -21779
rect 4604 -21847 4616 -21813
rect 4650 -21847 4662 -21813
rect 4604 -21881 4662 -21847
rect 4604 -21915 4616 -21881
rect 4650 -21915 4662 -21881
rect 4604 -21949 4662 -21915
rect 4604 -21983 4616 -21949
rect 4650 -21983 4662 -21949
rect 4604 -22017 4662 -21983
rect 4604 -22051 4616 -22017
rect 4650 -22051 4662 -22017
rect 4604 -22085 4662 -22051
rect 4604 -22119 4616 -22085
rect 4650 -22119 4662 -22085
rect 4604 -22153 4662 -22119
rect 4604 -22187 4616 -22153
rect 4650 -22187 4662 -22153
rect 4604 -22232 4662 -22187
rect 5622 -21677 5680 -21632
rect 5622 -21711 5634 -21677
rect 5668 -21711 5680 -21677
rect 5622 -21745 5680 -21711
rect 5622 -21779 5634 -21745
rect 5668 -21779 5680 -21745
rect 5622 -21813 5680 -21779
rect 5622 -21847 5634 -21813
rect 5668 -21847 5680 -21813
rect 5622 -21881 5680 -21847
rect 5622 -21915 5634 -21881
rect 5668 -21915 5680 -21881
rect 5622 -21949 5680 -21915
rect 5622 -21983 5634 -21949
rect 5668 -21983 5680 -21949
rect 5622 -22017 5680 -21983
rect 5622 -22051 5634 -22017
rect 5668 -22051 5680 -22017
rect 5622 -22085 5680 -22051
rect 5622 -22119 5634 -22085
rect 5668 -22119 5680 -22085
rect 5622 -22153 5680 -22119
rect 5622 -22187 5634 -22153
rect 5668 -22187 5680 -22153
rect 5622 -22232 5680 -22187
rect 6640 -21677 6698 -21632
rect 6640 -21711 6652 -21677
rect 6686 -21711 6698 -21677
rect 6640 -21745 6698 -21711
rect 6640 -21779 6652 -21745
rect 6686 -21779 6698 -21745
rect 6640 -21813 6698 -21779
rect 6640 -21847 6652 -21813
rect 6686 -21847 6698 -21813
rect 6640 -21881 6698 -21847
rect 6640 -21915 6652 -21881
rect 6686 -21915 6698 -21881
rect 6640 -21949 6698 -21915
rect 6640 -21983 6652 -21949
rect 6686 -21983 6698 -21949
rect 6640 -22017 6698 -21983
rect 6640 -22051 6652 -22017
rect 6686 -22051 6698 -22017
rect 6640 -22085 6698 -22051
rect 6640 -22119 6652 -22085
rect 6686 -22119 6698 -22085
rect 6640 -22153 6698 -22119
rect 6640 -22187 6652 -22153
rect 6686 -22187 6698 -22153
rect 6640 -22232 6698 -22187
rect 7658 -21677 7716 -21632
rect 7658 -21711 7670 -21677
rect 7704 -21711 7716 -21677
rect 7658 -21745 7716 -21711
rect 7658 -21779 7670 -21745
rect 7704 -21779 7716 -21745
rect 7658 -21813 7716 -21779
rect 7658 -21847 7670 -21813
rect 7704 -21847 7716 -21813
rect 7658 -21881 7716 -21847
rect 7658 -21915 7670 -21881
rect 7704 -21915 7716 -21881
rect 7658 -21949 7716 -21915
rect 7658 -21983 7670 -21949
rect 7704 -21983 7716 -21949
rect 7658 -22017 7716 -21983
rect 7658 -22051 7670 -22017
rect 7704 -22051 7716 -22017
rect 7658 -22085 7716 -22051
rect 7658 -22119 7670 -22085
rect 7704 -22119 7716 -22085
rect 7658 -22153 7716 -22119
rect 7658 -22187 7670 -22153
rect 7704 -22187 7716 -22153
rect 7658 -22232 7716 -22187
rect 8676 -21677 8734 -21632
rect 8676 -21711 8688 -21677
rect 8722 -21711 8734 -21677
rect 8676 -21745 8734 -21711
rect 8676 -21779 8688 -21745
rect 8722 -21779 8734 -21745
rect 8676 -21813 8734 -21779
rect 8676 -21847 8688 -21813
rect 8722 -21847 8734 -21813
rect 8676 -21881 8734 -21847
rect 8676 -21915 8688 -21881
rect 8722 -21915 8734 -21881
rect 8676 -21949 8734 -21915
rect 8676 -21983 8688 -21949
rect 8722 -21983 8734 -21949
rect 8676 -22017 8734 -21983
rect 8676 -22051 8688 -22017
rect 8722 -22051 8734 -22017
rect 8676 -22085 8734 -22051
rect 8676 -22119 8688 -22085
rect 8722 -22119 8734 -22085
rect 8676 -22153 8734 -22119
rect 8676 -22187 8688 -22153
rect 8722 -22187 8734 -22153
rect 8676 -22232 8734 -22187
rect 9694 -21677 9752 -21632
rect 9694 -21711 9706 -21677
rect 9740 -21711 9752 -21677
rect 9694 -21745 9752 -21711
rect 9694 -21779 9706 -21745
rect 9740 -21779 9752 -21745
rect 9694 -21813 9752 -21779
rect 9694 -21847 9706 -21813
rect 9740 -21847 9752 -21813
rect 9694 -21881 9752 -21847
rect 9694 -21915 9706 -21881
rect 9740 -21915 9752 -21881
rect 9694 -21949 9752 -21915
rect 9694 -21983 9706 -21949
rect 9740 -21983 9752 -21949
rect 9694 -22017 9752 -21983
rect 9694 -22051 9706 -22017
rect 9740 -22051 9752 -22017
rect 9694 -22085 9752 -22051
rect 9694 -22119 9706 -22085
rect 9740 -22119 9752 -22085
rect 9694 -22153 9752 -22119
rect 9694 -22187 9706 -22153
rect 9740 -22187 9752 -22153
rect 9694 -22232 9752 -22187
rect 10712 -21677 10770 -21632
rect 10712 -21711 10724 -21677
rect 10758 -21711 10770 -21677
rect 10712 -21745 10770 -21711
rect 10712 -21779 10724 -21745
rect 10758 -21779 10770 -21745
rect 10712 -21813 10770 -21779
rect 10712 -21847 10724 -21813
rect 10758 -21847 10770 -21813
rect 10712 -21881 10770 -21847
rect 10712 -21915 10724 -21881
rect 10758 -21915 10770 -21881
rect 10712 -21949 10770 -21915
rect 10712 -21983 10724 -21949
rect 10758 -21983 10770 -21949
rect 10712 -22017 10770 -21983
rect 10712 -22051 10724 -22017
rect 10758 -22051 10770 -22017
rect 10712 -22085 10770 -22051
rect 10712 -22119 10724 -22085
rect 10758 -22119 10770 -22085
rect 10712 -22153 10770 -22119
rect 10712 -22187 10724 -22153
rect 10758 -22187 10770 -22153
rect 10712 -22232 10770 -22187
rect 11730 -21677 11788 -21632
rect 11730 -21711 11742 -21677
rect 11776 -21711 11788 -21677
rect 11730 -21745 11788 -21711
rect 11730 -21779 11742 -21745
rect 11776 -21779 11788 -21745
rect 11730 -21813 11788 -21779
rect 11730 -21847 11742 -21813
rect 11776 -21847 11788 -21813
rect 11730 -21881 11788 -21847
rect 11730 -21915 11742 -21881
rect 11776 -21915 11788 -21881
rect 11730 -21949 11788 -21915
rect 11730 -21983 11742 -21949
rect 11776 -21983 11788 -21949
rect 11730 -22017 11788 -21983
rect 11730 -22051 11742 -22017
rect 11776 -22051 11788 -22017
rect 11730 -22085 11788 -22051
rect 11730 -22119 11742 -22085
rect 11776 -22119 11788 -22085
rect 11730 -22153 11788 -22119
rect 11730 -22187 11742 -22153
rect 11776 -22187 11788 -22153
rect 11730 -22232 11788 -22187
rect 12748 -21677 12806 -21632
rect 12748 -21711 12760 -21677
rect 12794 -21711 12806 -21677
rect 12748 -21745 12806 -21711
rect 12748 -21779 12760 -21745
rect 12794 -21779 12806 -21745
rect 12748 -21813 12806 -21779
rect 12748 -21847 12760 -21813
rect 12794 -21847 12806 -21813
rect 12748 -21881 12806 -21847
rect 12748 -21915 12760 -21881
rect 12794 -21915 12806 -21881
rect 12748 -21949 12806 -21915
rect 12748 -21983 12760 -21949
rect 12794 -21983 12806 -21949
rect 12748 -22017 12806 -21983
rect 12748 -22051 12760 -22017
rect 12794 -22051 12806 -22017
rect 12748 -22085 12806 -22051
rect 12748 -22119 12760 -22085
rect 12794 -22119 12806 -22085
rect 12748 -22153 12806 -22119
rect 12748 -22187 12760 -22153
rect 12794 -22187 12806 -22153
rect 12748 -22232 12806 -22187
rect 13766 -21677 13824 -21632
rect 13766 -21711 13778 -21677
rect 13812 -21711 13824 -21677
rect 13766 -21745 13824 -21711
rect 13766 -21779 13778 -21745
rect 13812 -21779 13824 -21745
rect 13766 -21813 13824 -21779
rect 13766 -21847 13778 -21813
rect 13812 -21847 13824 -21813
rect 13766 -21881 13824 -21847
rect 13766 -21915 13778 -21881
rect 13812 -21915 13824 -21881
rect 13766 -21949 13824 -21915
rect 13766 -21983 13778 -21949
rect 13812 -21983 13824 -21949
rect 13766 -22017 13824 -21983
rect 13766 -22051 13778 -22017
rect 13812 -22051 13824 -22017
rect 13766 -22085 13824 -22051
rect 13766 -22119 13778 -22085
rect 13812 -22119 13824 -22085
rect 13766 -22153 13824 -22119
rect 13766 -22187 13778 -22153
rect 13812 -22187 13824 -22153
rect 13766 -22232 13824 -22187
rect 14784 -21677 14842 -21632
rect 14784 -21711 14796 -21677
rect 14830 -21711 14842 -21677
rect 14784 -21745 14842 -21711
rect 14784 -21779 14796 -21745
rect 14830 -21779 14842 -21745
rect 14784 -21813 14842 -21779
rect 14784 -21847 14796 -21813
rect 14830 -21847 14842 -21813
rect 14784 -21881 14842 -21847
rect 14784 -21915 14796 -21881
rect 14830 -21915 14842 -21881
rect 14784 -21949 14842 -21915
rect 14784 -21983 14796 -21949
rect 14830 -21983 14842 -21949
rect 14784 -22017 14842 -21983
rect 14784 -22051 14796 -22017
rect 14830 -22051 14842 -22017
rect 14784 -22085 14842 -22051
rect 14784 -22119 14796 -22085
rect 14830 -22119 14842 -22085
rect 14784 -22153 14842 -22119
rect 14784 -22187 14796 -22153
rect 14830 -22187 14842 -22153
rect 14784 -22232 14842 -22187
rect 15802 -21677 15860 -21632
rect 15802 -21711 15814 -21677
rect 15848 -21711 15860 -21677
rect 15802 -21745 15860 -21711
rect 15802 -21779 15814 -21745
rect 15848 -21779 15860 -21745
rect 15802 -21813 15860 -21779
rect 15802 -21847 15814 -21813
rect 15848 -21847 15860 -21813
rect 15802 -21881 15860 -21847
rect 15802 -21915 15814 -21881
rect 15848 -21915 15860 -21881
rect 15802 -21949 15860 -21915
rect 15802 -21983 15814 -21949
rect 15848 -21983 15860 -21949
rect 15802 -22017 15860 -21983
rect 15802 -22051 15814 -22017
rect 15848 -22051 15860 -22017
rect 15802 -22085 15860 -22051
rect 15802 -22119 15814 -22085
rect 15848 -22119 15860 -22085
rect 15802 -22153 15860 -22119
rect 15802 -22187 15814 -22153
rect 15848 -22187 15860 -22153
rect 15802 -22232 15860 -22187
rect 16820 -21677 16878 -21632
rect 16820 -21711 16832 -21677
rect 16866 -21711 16878 -21677
rect 16820 -21745 16878 -21711
rect 16820 -21779 16832 -21745
rect 16866 -21779 16878 -21745
rect 16820 -21813 16878 -21779
rect 16820 -21847 16832 -21813
rect 16866 -21847 16878 -21813
rect 16820 -21881 16878 -21847
rect 16820 -21915 16832 -21881
rect 16866 -21915 16878 -21881
rect 16820 -21949 16878 -21915
rect 16820 -21983 16832 -21949
rect 16866 -21983 16878 -21949
rect 16820 -22017 16878 -21983
rect 16820 -22051 16832 -22017
rect 16866 -22051 16878 -22017
rect 16820 -22085 16878 -22051
rect 16820 -22119 16832 -22085
rect 16866 -22119 16878 -22085
rect 16820 -22153 16878 -22119
rect 16820 -22187 16832 -22153
rect 16866 -22187 16878 -22153
rect 16820 -22232 16878 -22187
rect 17838 -21677 17896 -21632
rect 17838 -21711 17850 -21677
rect 17884 -21711 17896 -21677
rect 17838 -21745 17896 -21711
rect 17838 -21779 17850 -21745
rect 17884 -21779 17896 -21745
rect 17838 -21813 17896 -21779
rect 17838 -21847 17850 -21813
rect 17884 -21847 17896 -21813
rect 17838 -21881 17896 -21847
rect 17838 -21915 17850 -21881
rect 17884 -21915 17896 -21881
rect 17838 -21949 17896 -21915
rect 17838 -21983 17850 -21949
rect 17884 -21983 17896 -21949
rect 17838 -22017 17896 -21983
rect 17838 -22051 17850 -22017
rect 17884 -22051 17896 -22017
rect 17838 -22085 17896 -22051
rect 17838 -22119 17850 -22085
rect 17884 -22119 17896 -22085
rect 17838 -22153 17896 -22119
rect 17838 -22187 17850 -22153
rect 17884 -22187 17896 -22153
rect 17838 -22232 17896 -22187
rect 18856 -21677 18914 -21632
rect 18856 -21711 18868 -21677
rect 18902 -21711 18914 -21677
rect 18856 -21745 18914 -21711
rect 18856 -21779 18868 -21745
rect 18902 -21779 18914 -21745
rect 18856 -21813 18914 -21779
rect 18856 -21847 18868 -21813
rect 18902 -21847 18914 -21813
rect 18856 -21881 18914 -21847
rect 18856 -21915 18868 -21881
rect 18902 -21915 18914 -21881
rect 18856 -21949 18914 -21915
rect 18856 -21983 18868 -21949
rect 18902 -21983 18914 -21949
rect 18856 -22017 18914 -21983
rect 18856 -22051 18868 -22017
rect 18902 -22051 18914 -22017
rect 18856 -22085 18914 -22051
rect 18856 -22119 18868 -22085
rect 18902 -22119 18914 -22085
rect 18856 -22153 18914 -22119
rect 18856 -22187 18868 -22153
rect 18902 -22187 18914 -22153
rect 18856 -22232 18914 -22187
rect 19874 -21677 19932 -21632
rect 19874 -21711 19886 -21677
rect 19920 -21711 19932 -21677
rect 19874 -21745 19932 -21711
rect 19874 -21779 19886 -21745
rect 19920 -21779 19932 -21745
rect 19874 -21813 19932 -21779
rect 19874 -21847 19886 -21813
rect 19920 -21847 19932 -21813
rect 19874 -21881 19932 -21847
rect 19874 -21915 19886 -21881
rect 19920 -21915 19932 -21881
rect 19874 -21949 19932 -21915
rect 19874 -21983 19886 -21949
rect 19920 -21983 19932 -21949
rect 19874 -22017 19932 -21983
rect 19874 -22051 19886 -22017
rect 19920 -22051 19932 -22017
rect 19874 -22085 19932 -22051
rect 19874 -22119 19886 -22085
rect 19920 -22119 19932 -22085
rect 19874 -22153 19932 -22119
rect 19874 -22187 19886 -22153
rect 19920 -22187 19932 -22153
rect 19874 -22232 19932 -22187
rect 20892 -21677 20950 -21632
rect 20892 -21711 20904 -21677
rect 20938 -21711 20950 -21677
rect 20892 -21745 20950 -21711
rect 20892 -21779 20904 -21745
rect 20938 -21779 20950 -21745
rect 20892 -21813 20950 -21779
rect 20892 -21847 20904 -21813
rect 20938 -21847 20950 -21813
rect 20892 -21881 20950 -21847
rect 20892 -21915 20904 -21881
rect 20938 -21915 20950 -21881
rect 20892 -21949 20950 -21915
rect 20892 -21983 20904 -21949
rect 20938 -21983 20950 -21949
rect 20892 -22017 20950 -21983
rect 20892 -22051 20904 -22017
rect 20938 -22051 20950 -22017
rect 20892 -22085 20950 -22051
rect 20892 -22119 20904 -22085
rect 20938 -22119 20950 -22085
rect 20892 -22153 20950 -22119
rect 20892 -22187 20904 -22153
rect 20938 -22187 20950 -22153
rect 20892 -22232 20950 -22187
rect 21910 -21677 21968 -21632
rect 21910 -21711 21922 -21677
rect 21956 -21711 21968 -21677
rect 21910 -21745 21968 -21711
rect 21910 -21779 21922 -21745
rect 21956 -21779 21968 -21745
rect 21910 -21813 21968 -21779
rect 21910 -21847 21922 -21813
rect 21956 -21847 21968 -21813
rect 21910 -21881 21968 -21847
rect 21910 -21915 21922 -21881
rect 21956 -21915 21968 -21881
rect 21910 -21949 21968 -21915
rect 21910 -21983 21922 -21949
rect 21956 -21983 21968 -21949
rect 21910 -22017 21968 -21983
rect 21910 -22051 21922 -22017
rect 21956 -22051 21968 -22017
rect 21910 -22085 21968 -22051
rect 21910 -22119 21922 -22085
rect 21956 -22119 21968 -22085
rect 21910 -22153 21968 -22119
rect 21910 -22187 21922 -22153
rect 21956 -22187 21968 -22153
rect 21910 -22232 21968 -22187
rect 22928 -21677 22986 -21632
rect 22928 -21711 22940 -21677
rect 22974 -21711 22986 -21677
rect 22928 -21745 22986 -21711
rect 22928 -21779 22940 -21745
rect 22974 -21779 22986 -21745
rect 22928 -21813 22986 -21779
rect 22928 -21847 22940 -21813
rect 22974 -21847 22986 -21813
rect 22928 -21881 22986 -21847
rect 22928 -21915 22940 -21881
rect 22974 -21915 22986 -21881
rect 22928 -21949 22986 -21915
rect 22928 -21983 22940 -21949
rect 22974 -21983 22986 -21949
rect 22928 -22017 22986 -21983
rect 22928 -22051 22940 -22017
rect 22974 -22051 22986 -22017
rect 22928 -22085 22986 -22051
rect 22928 -22119 22940 -22085
rect 22974 -22119 22986 -22085
rect 22928 -22153 22986 -22119
rect 22928 -22187 22940 -22153
rect 22974 -22187 22986 -22153
rect 22928 -22232 22986 -22187
rect 2568 -22909 2626 -22864
rect 2568 -22943 2580 -22909
rect 2614 -22943 2626 -22909
rect 2568 -22977 2626 -22943
rect 2568 -23011 2580 -22977
rect 2614 -23011 2626 -22977
rect 2568 -23045 2626 -23011
rect 2568 -23079 2580 -23045
rect 2614 -23079 2626 -23045
rect 2568 -23113 2626 -23079
rect 2568 -23147 2580 -23113
rect 2614 -23147 2626 -23113
rect 2568 -23181 2626 -23147
rect 2568 -23215 2580 -23181
rect 2614 -23215 2626 -23181
rect 2568 -23249 2626 -23215
rect 2568 -23283 2580 -23249
rect 2614 -23283 2626 -23249
rect 2568 -23317 2626 -23283
rect 2568 -23351 2580 -23317
rect 2614 -23351 2626 -23317
rect 2568 -23385 2626 -23351
rect 2568 -23419 2580 -23385
rect 2614 -23419 2626 -23385
rect 2568 -23464 2626 -23419
rect 3586 -22909 3644 -22864
rect 3586 -22943 3598 -22909
rect 3632 -22943 3644 -22909
rect 3586 -22977 3644 -22943
rect 3586 -23011 3598 -22977
rect 3632 -23011 3644 -22977
rect 3586 -23045 3644 -23011
rect 3586 -23079 3598 -23045
rect 3632 -23079 3644 -23045
rect 3586 -23113 3644 -23079
rect 3586 -23147 3598 -23113
rect 3632 -23147 3644 -23113
rect 3586 -23181 3644 -23147
rect 3586 -23215 3598 -23181
rect 3632 -23215 3644 -23181
rect 3586 -23249 3644 -23215
rect 3586 -23283 3598 -23249
rect 3632 -23283 3644 -23249
rect 3586 -23317 3644 -23283
rect 3586 -23351 3598 -23317
rect 3632 -23351 3644 -23317
rect 3586 -23385 3644 -23351
rect 3586 -23419 3598 -23385
rect 3632 -23419 3644 -23385
rect 3586 -23464 3644 -23419
rect 4604 -22909 4662 -22864
rect 4604 -22943 4616 -22909
rect 4650 -22943 4662 -22909
rect 4604 -22977 4662 -22943
rect 4604 -23011 4616 -22977
rect 4650 -23011 4662 -22977
rect 4604 -23045 4662 -23011
rect 4604 -23079 4616 -23045
rect 4650 -23079 4662 -23045
rect 4604 -23113 4662 -23079
rect 4604 -23147 4616 -23113
rect 4650 -23147 4662 -23113
rect 4604 -23181 4662 -23147
rect 4604 -23215 4616 -23181
rect 4650 -23215 4662 -23181
rect 4604 -23249 4662 -23215
rect 4604 -23283 4616 -23249
rect 4650 -23283 4662 -23249
rect 4604 -23317 4662 -23283
rect 4604 -23351 4616 -23317
rect 4650 -23351 4662 -23317
rect 4604 -23385 4662 -23351
rect 4604 -23419 4616 -23385
rect 4650 -23419 4662 -23385
rect 4604 -23464 4662 -23419
rect 5622 -22909 5680 -22864
rect 5622 -22943 5634 -22909
rect 5668 -22943 5680 -22909
rect 5622 -22977 5680 -22943
rect 5622 -23011 5634 -22977
rect 5668 -23011 5680 -22977
rect 5622 -23045 5680 -23011
rect 5622 -23079 5634 -23045
rect 5668 -23079 5680 -23045
rect 5622 -23113 5680 -23079
rect 5622 -23147 5634 -23113
rect 5668 -23147 5680 -23113
rect 5622 -23181 5680 -23147
rect 5622 -23215 5634 -23181
rect 5668 -23215 5680 -23181
rect 5622 -23249 5680 -23215
rect 5622 -23283 5634 -23249
rect 5668 -23283 5680 -23249
rect 5622 -23317 5680 -23283
rect 5622 -23351 5634 -23317
rect 5668 -23351 5680 -23317
rect 5622 -23385 5680 -23351
rect 5622 -23419 5634 -23385
rect 5668 -23419 5680 -23385
rect 5622 -23464 5680 -23419
rect 6640 -22909 6698 -22864
rect 6640 -22943 6652 -22909
rect 6686 -22943 6698 -22909
rect 6640 -22977 6698 -22943
rect 6640 -23011 6652 -22977
rect 6686 -23011 6698 -22977
rect 6640 -23045 6698 -23011
rect 6640 -23079 6652 -23045
rect 6686 -23079 6698 -23045
rect 6640 -23113 6698 -23079
rect 6640 -23147 6652 -23113
rect 6686 -23147 6698 -23113
rect 6640 -23181 6698 -23147
rect 6640 -23215 6652 -23181
rect 6686 -23215 6698 -23181
rect 6640 -23249 6698 -23215
rect 6640 -23283 6652 -23249
rect 6686 -23283 6698 -23249
rect 6640 -23317 6698 -23283
rect 6640 -23351 6652 -23317
rect 6686 -23351 6698 -23317
rect 6640 -23385 6698 -23351
rect 6640 -23419 6652 -23385
rect 6686 -23419 6698 -23385
rect 6640 -23464 6698 -23419
rect 7658 -22909 7716 -22864
rect 7658 -22943 7670 -22909
rect 7704 -22943 7716 -22909
rect 7658 -22977 7716 -22943
rect 7658 -23011 7670 -22977
rect 7704 -23011 7716 -22977
rect 7658 -23045 7716 -23011
rect 7658 -23079 7670 -23045
rect 7704 -23079 7716 -23045
rect 7658 -23113 7716 -23079
rect 7658 -23147 7670 -23113
rect 7704 -23147 7716 -23113
rect 7658 -23181 7716 -23147
rect 7658 -23215 7670 -23181
rect 7704 -23215 7716 -23181
rect 7658 -23249 7716 -23215
rect 7658 -23283 7670 -23249
rect 7704 -23283 7716 -23249
rect 7658 -23317 7716 -23283
rect 7658 -23351 7670 -23317
rect 7704 -23351 7716 -23317
rect 7658 -23385 7716 -23351
rect 7658 -23419 7670 -23385
rect 7704 -23419 7716 -23385
rect 7658 -23464 7716 -23419
rect 8676 -22909 8734 -22864
rect 8676 -22943 8688 -22909
rect 8722 -22943 8734 -22909
rect 8676 -22977 8734 -22943
rect 8676 -23011 8688 -22977
rect 8722 -23011 8734 -22977
rect 8676 -23045 8734 -23011
rect 8676 -23079 8688 -23045
rect 8722 -23079 8734 -23045
rect 8676 -23113 8734 -23079
rect 8676 -23147 8688 -23113
rect 8722 -23147 8734 -23113
rect 8676 -23181 8734 -23147
rect 8676 -23215 8688 -23181
rect 8722 -23215 8734 -23181
rect 8676 -23249 8734 -23215
rect 8676 -23283 8688 -23249
rect 8722 -23283 8734 -23249
rect 8676 -23317 8734 -23283
rect 8676 -23351 8688 -23317
rect 8722 -23351 8734 -23317
rect 8676 -23385 8734 -23351
rect 8676 -23419 8688 -23385
rect 8722 -23419 8734 -23385
rect 8676 -23464 8734 -23419
rect 9694 -22909 9752 -22864
rect 9694 -22943 9706 -22909
rect 9740 -22943 9752 -22909
rect 9694 -22977 9752 -22943
rect 9694 -23011 9706 -22977
rect 9740 -23011 9752 -22977
rect 9694 -23045 9752 -23011
rect 9694 -23079 9706 -23045
rect 9740 -23079 9752 -23045
rect 9694 -23113 9752 -23079
rect 9694 -23147 9706 -23113
rect 9740 -23147 9752 -23113
rect 9694 -23181 9752 -23147
rect 9694 -23215 9706 -23181
rect 9740 -23215 9752 -23181
rect 9694 -23249 9752 -23215
rect 9694 -23283 9706 -23249
rect 9740 -23283 9752 -23249
rect 9694 -23317 9752 -23283
rect 9694 -23351 9706 -23317
rect 9740 -23351 9752 -23317
rect 9694 -23385 9752 -23351
rect 9694 -23419 9706 -23385
rect 9740 -23419 9752 -23385
rect 9694 -23464 9752 -23419
rect 10712 -22909 10770 -22864
rect 10712 -22943 10724 -22909
rect 10758 -22943 10770 -22909
rect 10712 -22977 10770 -22943
rect 10712 -23011 10724 -22977
rect 10758 -23011 10770 -22977
rect 10712 -23045 10770 -23011
rect 10712 -23079 10724 -23045
rect 10758 -23079 10770 -23045
rect 10712 -23113 10770 -23079
rect 10712 -23147 10724 -23113
rect 10758 -23147 10770 -23113
rect 10712 -23181 10770 -23147
rect 10712 -23215 10724 -23181
rect 10758 -23215 10770 -23181
rect 10712 -23249 10770 -23215
rect 10712 -23283 10724 -23249
rect 10758 -23283 10770 -23249
rect 10712 -23317 10770 -23283
rect 10712 -23351 10724 -23317
rect 10758 -23351 10770 -23317
rect 10712 -23385 10770 -23351
rect 10712 -23419 10724 -23385
rect 10758 -23419 10770 -23385
rect 10712 -23464 10770 -23419
rect 11730 -22909 11788 -22864
rect 11730 -22943 11742 -22909
rect 11776 -22943 11788 -22909
rect 11730 -22977 11788 -22943
rect 11730 -23011 11742 -22977
rect 11776 -23011 11788 -22977
rect 11730 -23045 11788 -23011
rect 11730 -23079 11742 -23045
rect 11776 -23079 11788 -23045
rect 11730 -23113 11788 -23079
rect 11730 -23147 11742 -23113
rect 11776 -23147 11788 -23113
rect 11730 -23181 11788 -23147
rect 11730 -23215 11742 -23181
rect 11776 -23215 11788 -23181
rect 11730 -23249 11788 -23215
rect 11730 -23283 11742 -23249
rect 11776 -23283 11788 -23249
rect 11730 -23317 11788 -23283
rect 11730 -23351 11742 -23317
rect 11776 -23351 11788 -23317
rect 11730 -23385 11788 -23351
rect 11730 -23419 11742 -23385
rect 11776 -23419 11788 -23385
rect 11730 -23464 11788 -23419
rect 12748 -22909 12806 -22864
rect 12748 -22943 12760 -22909
rect 12794 -22943 12806 -22909
rect 12748 -22977 12806 -22943
rect 12748 -23011 12760 -22977
rect 12794 -23011 12806 -22977
rect 12748 -23045 12806 -23011
rect 12748 -23079 12760 -23045
rect 12794 -23079 12806 -23045
rect 12748 -23113 12806 -23079
rect 12748 -23147 12760 -23113
rect 12794 -23147 12806 -23113
rect 12748 -23181 12806 -23147
rect 12748 -23215 12760 -23181
rect 12794 -23215 12806 -23181
rect 12748 -23249 12806 -23215
rect 12748 -23283 12760 -23249
rect 12794 -23283 12806 -23249
rect 12748 -23317 12806 -23283
rect 12748 -23351 12760 -23317
rect 12794 -23351 12806 -23317
rect 12748 -23385 12806 -23351
rect 12748 -23419 12760 -23385
rect 12794 -23419 12806 -23385
rect 12748 -23464 12806 -23419
rect 13766 -22909 13824 -22864
rect 13766 -22943 13778 -22909
rect 13812 -22943 13824 -22909
rect 13766 -22977 13824 -22943
rect 13766 -23011 13778 -22977
rect 13812 -23011 13824 -22977
rect 13766 -23045 13824 -23011
rect 13766 -23079 13778 -23045
rect 13812 -23079 13824 -23045
rect 13766 -23113 13824 -23079
rect 13766 -23147 13778 -23113
rect 13812 -23147 13824 -23113
rect 13766 -23181 13824 -23147
rect 13766 -23215 13778 -23181
rect 13812 -23215 13824 -23181
rect 13766 -23249 13824 -23215
rect 13766 -23283 13778 -23249
rect 13812 -23283 13824 -23249
rect 13766 -23317 13824 -23283
rect 13766 -23351 13778 -23317
rect 13812 -23351 13824 -23317
rect 13766 -23385 13824 -23351
rect 13766 -23419 13778 -23385
rect 13812 -23419 13824 -23385
rect 13766 -23464 13824 -23419
rect 14784 -22909 14842 -22864
rect 14784 -22943 14796 -22909
rect 14830 -22943 14842 -22909
rect 14784 -22977 14842 -22943
rect 14784 -23011 14796 -22977
rect 14830 -23011 14842 -22977
rect 14784 -23045 14842 -23011
rect 14784 -23079 14796 -23045
rect 14830 -23079 14842 -23045
rect 14784 -23113 14842 -23079
rect 14784 -23147 14796 -23113
rect 14830 -23147 14842 -23113
rect 14784 -23181 14842 -23147
rect 14784 -23215 14796 -23181
rect 14830 -23215 14842 -23181
rect 14784 -23249 14842 -23215
rect 14784 -23283 14796 -23249
rect 14830 -23283 14842 -23249
rect 14784 -23317 14842 -23283
rect 14784 -23351 14796 -23317
rect 14830 -23351 14842 -23317
rect 14784 -23385 14842 -23351
rect 14784 -23419 14796 -23385
rect 14830 -23419 14842 -23385
rect 14784 -23464 14842 -23419
rect 15802 -22909 15860 -22864
rect 15802 -22943 15814 -22909
rect 15848 -22943 15860 -22909
rect 15802 -22977 15860 -22943
rect 15802 -23011 15814 -22977
rect 15848 -23011 15860 -22977
rect 15802 -23045 15860 -23011
rect 15802 -23079 15814 -23045
rect 15848 -23079 15860 -23045
rect 15802 -23113 15860 -23079
rect 15802 -23147 15814 -23113
rect 15848 -23147 15860 -23113
rect 15802 -23181 15860 -23147
rect 15802 -23215 15814 -23181
rect 15848 -23215 15860 -23181
rect 15802 -23249 15860 -23215
rect 15802 -23283 15814 -23249
rect 15848 -23283 15860 -23249
rect 15802 -23317 15860 -23283
rect 15802 -23351 15814 -23317
rect 15848 -23351 15860 -23317
rect 15802 -23385 15860 -23351
rect 15802 -23419 15814 -23385
rect 15848 -23419 15860 -23385
rect 15802 -23464 15860 -23419
rect 16820 -22909 16878 -22864
rect 16820 -22943 16832 -22909
rect 16866 -22943 16878 -22909
rect 16820 -22977 16878 -22943
rect 16820 -23011 16832 -22977
rect 16866 -23011 16878 -22977
rect 16820 -23045 16878 -23011
rect 16820 -23079 16832 -23045
rect 16866 -23079 16878 -23045
rect 16820 -23113 16878 -23079
rect 16820 -23147 16832 -23113
rect 16866 -23147 16878 -23113
rect 16820 -23181 16878 -23147
rect 16820 -23215 16832 -23181
rect 16866 -23215 16878 -23181
rect 16820 -23249 16878 -23215
rect 16820 -23283 16832 -23249
rect 16866 -23283 16878 -23249
rect 16820 -23317 16878 -23283
rect 16820 -23351 16832 -23317
rect 16866 -23351 16878 -23317
rect 16820 -23385 16878 -23351
rect 16820 -23419 16832 -23385
rect 16866 -23419 16878 -23385
rect 16820 -23464 16878 -23419
rect 17838 -22909 17896 -22864
rect 17838 -22943 17850 -22909
rect 17884 -22943 17896 -22909
rect 17838 -22977 17896 -22943
rect 17838 -23011 17850 -22977
rect 17884 -23011 17896 -22977
rect 17838 -23045 17896 -23011
rect 17838 -23079 17850 -23045
rect 17884 -23079 17896 -23045
rect 17838 -23113 17896 -23079
rect 17838 -23147 17850 -23113
rect 17884 -23147 17896 -23113
rect 17838 -23181 17896 -23147
rect 17838 -23215 17850 -23181
rect 17884 -23215 17896 -23181
rect 17838 -23249 17896 -23215
rect 17838 -23283 17850 -23249
rect 17884 -23283 17896 -23249
rect 17838 -23317 17896 -23283
rect 17838 -23351 17850 -23317
rect 17884 -23351 17896 -23317
rect 17838 -23385 17896 -23351
rect 17838 -23419 17850 -23385
rect 17884 -23419 17896 -23385
rect 17838 -23464 17896 -23419
rect 18856 -22909 18914 -22864
rect 18856 -22943 18868 -22909
rect 18902 -22943 18914 -22909
rect 18856 -22977 18914 -22943
rect 18856 -23011 18868 -22977
rect 18902 -23011 18914 -22977
rect 18856 -23045 18914 -23011
rect 18856 -23079 18868 -23045
rect 18902 -23079 18914 -23045
rect 18856 -23113 18914 -23079
rect 18856 -23147 18868 -23113
rect 18902 -23147 18914 -23113
rect 18856 -23181 18914 -23147
rect 18856 -23215 18868 -23181
rect 18902 -23215 18914 -23181
rect 18856 -23249 18914 -23215
rect 18856 -23283 18868 -23249
rect 18902 -23283 18914 -23249
rect 18856 -23317 18914 -23283
rect 18856 -23351 18868 -23317
rect 18902 -23351 18914 -23317
rect 18856 -23385 18914 -23351
rect 18856 -23419 18868 -23385
rect 18902 -23419 18914 -23385
rect 18856 -23464 18914 -23419
rect 19874 -22909 19932 -22864
rect 19874 -22943 19886 -22909
rect 19920 -22943 19932 -22909
rect 19874 -22977 19932 -22943
rect 19874 -23011 19886 -22977
rect 19920 -23011 19932 -22977
rect 19874 -23045 19932 -23011
rect 19874 -23079 19886 -23045
rect 19920 -23079 19932 -23045
rect 19874 -23113 19932 -23079
rect 19874 -23147 19886 -23113
rect 19920 -23147 19932 -23113
rect 19874 -23181 19932 -23147
rect 19874 -23215 19886 -23181
rect 19920 -23215 19932 -23181
rect 19874 -23249 19932 -23215
rect 19874 -23283 19886 -23249
rect 19920 -23283 19932 -23249
rect 19874 -23317 19932 -23283
rect 19874 -23351 19886 -23317
rect 19920 -23351 19932 -23317
rect 19874 -23385 19932 -23351
rect 19874 -23419 19886 -23385
rect 19920 -23419 19932 -23385
rect 19874 -23464 19932 -23419
rect 20892 -22909 20950 -22864
rect 20892 -22943 20904 -22909
rect 20938 -22943 20950 -22909
rect 20892 -22977 20950 -22943
rect 20892 -23011 20904 -22977
rect 20938 -23011 20950 -22977
rect 20892 -23045 20950 -23011
rect 20892 -23079 20904 -23045
rect 20938 -23079 20950 -23045
rect 20892 -23113 20950 -23079
rect 20892 -23147 20904 -23113
rect 20938 -23147 20950 -23113
rect 20892 -23181 20950 -23147
rect 20892 -23215 20904 -23181
rect 20938 -23215 20950 -23181
rect 20892 -23249 20950 -23215
rect 20892 -23283 20904 -23249
rect 20938 -23283 20950 -23249
rect 20892 -23317 20950 -23283
rect 20892 -23351 20904 -23317
rect 20938 -23351 20950 -23317
rect 20892 -23385 20950 -23351
rect 20892 -23419 20904 -23385
rect 20938 -23419 20950 -23385
rect 20892 -23464 20950 -23419
rect 21910 -22909 21968 -22864
rect 21910 -22943 21922 -22909
rect 21956 -22943 21968 -22909
rect 21910 -22977 21968 -22943
rect 21910 -23011 21922 -22977
rect 21956 -23011 21968 -22977
rect 21910 -23045 21968 -23011
rect 21910 -23079 21922 -23045
rect 21956 -23079 21968 -23045
rect 21910 -23113 21968 -23079
rect 21910 -23147 21922 -23113
rect 21956 -23147 21968 -23113
rect 21910 -23181 21968 -23147
rect 21910 -23215 21922 -23181
rect 21956 -23215 21968 -23181
rect 21910 -23249 21968 -23215
rect 21910 -23283 21922 -23249
rect 21956 -23283 21968 -23249
rect 21910 -23317 21968 -23283
rect 21910 -23351 21922 -23317
rect 21956 -23351 21968 -23317
rect 21910 -23385 21968 -23351
rect 21910 -23419 21922 -23385
rect 21956 -23419 21968 -23385
rect 21910 -23464 21968 -23419
rect 22928 -22909 22986 -22864
rect 22928 -22943 22940 -22909
rect 22974 -22943 22986 -22909
rect 22928 -22977 22986 -22943
rect 22928 -23011 22940 -22977
rect 22974 -23011 22986 -22977
rect 22928 -23045 22986 -23011
rect 22928 -23079 22940 -23045
rect 22974 -23079 22986 -23045
rect 22928 -23113 22986 -23079
rect 22928 -23147 22940 -23113
rect 22974 -23147 22986 -23113
rect 22928 -23181 22986 -23147
rect 22928 -23215 22940 -23181
rect 22974 -23215 22986 -23181
rect 22928 -23249 22986 -23215
rect 22928 -23283 22940 -23249
rect 22974 -23283 22986 -23249
rect 22928 -23317 22986 -23283
rect 22928 -23351 22940 -23317
rect 22974 -23351 22986 -23317
rect 22928 -23385 22986 -23351
rect 22928 -23419 22940 -23385
rect 22974 -23419 22986 -23385
rect 22928 -23464 22986 -23419
rect 2568 -24143 2626 -24098
rect 2568 -24177 2580 -24143
rect 2614 -24177 2626 -24143
rect 2568 -24211 2626 -24177
rect 2568 -24245 2580 -24211
rect 2614 -24245 2626 -24211
rect 2568 -24279 2626 -24245
rect 2568 -24313 2580 -24279
rect 2614 -24313 2626 -24279
rect 2568 -24347 2626 -24313
rect 2568 -24381 2580 -24347
rect 2614 -24381 2626 -24347
rect 2568 -24415 2626 -24381
rect 2568 -24449 2580 -24415
rect 2614 -24449 2626 -24415
rect 2568 -24483 2626 -24449
rect 2568 -24517 2580 -24483
rect 2614 -24517 2626 -24483
rect 2568 -24551 2626 -24517
rect 2568 -24585 2580 -24551
rect 2614 -24585 2626 -24551
rect 2568 -24619 2626 -24585
rect 2568 -24653 2580 -24619
rect 2614 -24653 2626 -24619
rect 2568 -24698 2626 -24653
rect 3586 -24143 3644 -24098
rect 3586 -24177 3598 -24143
rect 3632 -24177 3644 -24143
rect 3586 -24211 3644 -24177
rect 3586 -24245 3598 -24211
rect 3632 -24245 3644 -24211
rect 3586 -24279 3644 -24245
rect 3586 -24313 3598 -24279
rect 3632 -24313 3644 -24279
rect 3586 -24347 3644 -24313
rect 3586 -24381 3598 -24347
rect 3632 -24381 3644 -24347
rect 3586 -24415 3644 -24381
rect 3586 -24449 3598 -24415
rect 3632 -24449 3644 -24415
rect 3586 -24483 3644 -24449
rect 3586 -24517 3598 -24483
rect 3632 -24517 3644 -24483
rect 3586 -24551 3644 -24517
rect 3586 -24585 3598 -24551
rect 3632 -24585 3644 -24551
rect 3586 -24619 3644 -24585
rect 3586 -24653 3598 -24619
rect 3632 -24653 3644 -24619
rect 3586 -24698 3644 -24653
rect 4604 -24143 4662 -24098
rect 4604 -24177 4616 -24143
rect 4650 -24177 4662 -24143
rect 4604 -24211 4662 -24177
rect 4604 -24245 4616 -24211
rect 4650 -24245 4662 -24211
rect 4604 -24279 4662 -24245
rect 4604 -24313 4616 -24279
rect 4650 -24313 4662 -24279
rect 4604 -24347 4662 -24313
rect 4604 -24381 4616 -24347
rect 4650 -24381 4662 -24347
rect 4604 -24415 4662 -24381
rect 4604 -24449 4616 -24415
rect 4650 -24449 4662 -24415
rect 4604 -24483 4662 -24449
rect 4604 -24517 4616 -24483
rect 4650 -24517 4662 -24483
rect 4604 -24551 4662 -24517
rect 4604 -24585 4616 -24551
rect 4650 -24585 4662 -24551
rect 4604 -24619 4662 -24585
rect 4604 -24653 4616 -24619
rect 4650 -24653 4662 -24619
rect 4604 -24698 4662 -24653
rect 5622 -24143 5680 -24098
rect 5622 -24177 5634 -24143
rect 5668 -24177 5680 -24143
rect 5622 -24211 5680 -24177
rect 5622 -24245 5634 -24211
rect 5668 -24245 5680 -24211
rect 5622 -24279 5680 -24245
rect 5622 -24313 5634 -24279
rect 5668 -24313 5680 -24279
rect 5622 -24347 5680 -24313
rect 5622 -24381 5634 -24347
rect 5668 -24381 5680 -24347
rect 5622 -24415 5680 -24381
rect 5622 -24449 5634 -24415
rect 5668 -24449 5680 -24415
rect 5622 -24483 5680 -24449
rect 5622 -24517 5634 -24483
rect 5668 -24517 5680 -24483
rect 5622 -24551 5680 -24517
rect 5622 -24585 5634 -24551
rect 5668 -24585 5680 -24551
rect 5622 -24619 5680 -24585
rect 5622 -24653 5634 -24619
rect 5668 -24653 5680 -24619
rect 5622 -24698 5680 -24653
rect 6640 -24143 6698 -24098
rect 6640 -24177 6652 -24143
rect 6686 -24177 6698 -24143
rect 6640 -24211 6698 -24177
rect 6640 -24245 6652 -24211
rect 6686 -24245 6698 -24211
rect 6640 -24279 6698 -24245
rect 6640 -24313 6652 -24279
rect 6686 -24313 6698 -24279
rect 6640 -24347 6698 -24313
rect 6640 -24381 6652 -24347
rect 6686 -24381 6698 -24347
rect 6640 -24415 6698 -24381
rect 6640 -24449 6652 -24415
rect 6686 -24449 6698 -24415
rect 6640 -24483 6698 -24449
rect 6640 -24517 6652 -24483
rect 6686 -24517 6698 -24483
rect 6640 -24551 6698 -24517
rect 6640 -24585 6652 -24551
rect 6686 -24585 6698 -24551
rect 6640 -24619 6698 -24585
rect 6640 -24653 6652 -24619
rect 6686 -24653 6698 -24619
rect 6640 -24698 6698 -24653
rect 7658 -24143 7716 -24098
rect 7658 -24177 7670 -24143
rect 7704 -24177 7716 -24143
rect 7658 -24211 7716 -24177
rect 7658 -24245 7670 -24211
rect 7704 -24245 7716 -24211
rect 7658 -24279 7716 -24245
rect 7658 -24313 7670 -24279
rect 7704 -24313 7716 -24279
rect 7658 -24347 7716 -24313
rect 7658 -24381 7670 -24347
rect 7704 -24381 7716 -24347
rect 7658 -24415 7716 -24381
rect 7658 -24449 7670 -24415
rect 7704 -24449 7716 -24415
rect 7658 -24483 7716 -24449
rect 7658 -24517 7670 -24483
rect 7704 -24517 7716 -24483
rect 7658 -24551 7716 -24517
rect 7658 -24585 7670 -24551
rect 7704 -24585 7716 -24551
rect 7658 -24619 7716 -24585
rect 7658 -24653 7670 -24619
rect 7704 -24653 7716 -24619
rect 7658 -24698 7716 -24653
rect 8676 -24143 8734 -24098
rect 8676 -24177 8688 -24143
rect 8722 -24177 8734 -24143
rect 8676 -24211 8734 -24177
rect 8676 -24245 8688 -24211
rect 8722 -24245 8734 -24211
rect 8676 -24279 8734 -24245
rect 8676 -24313 8688 -24279
rect 8722 -24313 8734 -24279
rect 8676 -24347 8734 -24313
rect 8676 -24381 8688 -24347
rect 8722 -24381 8734 -24347
rect 8676 -24415 8734 -24381
rect 8676 -24449 8688 -24415
rect 8722 -24449 8734 -24415
rect 8676 -24483 8734 -24449
rect 8676 -24517 8688 -24483
rect 8722 -24517 8734 -24483
rect 8676 -24551 8734 -24517
rect 8676 -24585 8688 -24551
rect 8722 -24585 8734 -24551
rect 8676 -24619 8734 -24585
rect 8676 -24653 8688 -24619
rect 8722 -24653 8734 -24619
rect 8676 -24698 8734 -24653
rect 9694 -24143 9752 -24098
rect 9694 -24177 9706 -24143
rect 9740 -24177 9752 -24143
rect 9694 -24211 9752 -24177
rect 9694 -24245 9706 -24211
rect 9740 -24245 9752 -24211
rect 9694 -24279 9752 -24245
rect 9694 -24313 9706 -24279
rect 9740 -24313 9752 -24279
rect 9694 -24347 9752 -24313
rect 9694 -24381 9706 -24347
rect 9740 -24381 9752 -24347
rect 9694 -24415 9752 -24381
rect 9694 -24449 9706 -24415
rect 9740 -24449 9752 -24415
rect 9694 -24483 9752 -24449
rect 9694 -24517 9706 -24483
rect 9740 -24517 9752 -24483
rect 9694 -24551 9752 -24517
rect 9694 -24585 9706 -24551
rect 9740 -24585 9752 -24551
rect 9694 -24619 9752 -24585
rect 9694 -24653 9706 -24619
rect 9740 -24653 9752 -24619
rect 9694 -24698 9752 -24653
rect 10712 -24143 10770 -24098
rect 10712 -24177 10724 -24143
rect 10758 -24177 10770 -24143
rect 10712 -24211 10770 -24177
rect 10712 -24245 10724 -24211
rect 10758 -24245 10770 -24211
rect 10712 -24279 10770 -24245
rect 10712 -24313 10724 -24279
rect 10758 -24313 10770 -24279
rect 10712 -24347 10770 -24313
rect 10712 -24381 10724 -24347
rect 10758 -24381 10770 -24347
rect 10712 -24415 10770 -24381
rect 10712 -24449 10724 -24415
rect 10758 -24449 10770 -24415
rect 10712 -24483 10770 -24449
rect 10712 -24517 10724 -24483
rect 10758 -24517 10770 -24483
rect 10712 -24551 10770 -24517
rect 10712 -24585 10724 -24551
rect 10758 -24585 10770 -24551
rect 10712 -24619 10770 -24585
rect 10712 -24653 10724 -24619
rect 10758 -24653 10770 -24619
rect 10712 -24698 10770 -24653
rect 11730 -24143 11788 -24098
rect 11730 -24177 11742 -24143
rect 11776 -24177 11788 -24143
rect 11730 -24211 11788 -24177
rect 11730 -24245 11742 -24211
rect 11776 -24245 11788 -24211
rect 11730 -24279 11788 -24245
rect 11730 -24313 11742 -24279
rect 11776 -24313 11788 -24279
rect 11730 -24347 11788 -24313
rect 11730 -24381 11742 -24347
rect 11776 -24381 11788 -24347
rect 11730 -24415 11788 -24381
rect 11730 -24449 11742 -24415
rect 11776 -24449 11788 -24415
rect 11730 -24483 11788 -24449
rect 11730 -24517 11742 -24483
rect 11776 -24517 11788 -24483
rect 11730 -24551 11788 -24517
rect 11730 -24585 11742 -24551
rect 11776 -24585 11788 -24551
rect 11730 -24619 11788 -24585
rect 11730 -24653 11742 -24619
rect 11776 -24653 11788 -24619
rect 11730 -24698 11788 -24653
rect 12748 -24143 12806 -24098
rect 12748 -24177 12760 -24143
rect 12794 -24177 12806 -24143
rect 12748 -24211 12806 -24177
rect 12748 -24245 12760 -24211
rect 12794 -24245 12806 -24211
rect 12748 -24279 12806 -24245
rect 12748 -24313 12760 -24279
rect 12794 -24313 12806 -24279
rect 12748 -24347 12806 -24313
rect 12748 -24381 12760 -24347
rect 12794 -24381 12806 -24347
rect 12748 -24415 12806 -24381
rect 12748 -24449 12760 -24415
rect 12794 -24449 12806 -24415
rect 12748 -24483 12806 -24449
rect 12748 -24517 12760 -24483
rect 12794 -24517 12806 -24483
rect 12748 -24551 12806 -24517
rect 12748 -24585 12760 -24551
rect 12794 -24585 12806 -24551
rect 12748 -24619 12806 -24585
rect 12748 -24653 12760 -24619
rect 12794 -24653 12806 -24619
rect 12748 -24698 12806 -24653
rect 13766 -24143 13824 -24098
rect 13766 -24177 13778 -24143
rect 13812 -24177 13824 -24143
rect 13766 -24211 13824 -24177
rect 13766 -24245 13778 -24211
rect 13812 -24245 13824 -24211
rect 13766 -24279 13824 -24245
rect 13766 -24313 13778 -24279
rect 13812 -24313 13824 -24279
rect 13766 -24347 13824 -24313
rect 13766 -24381 13778 -24347
rect 13812 -24381 13824 -24347
rect 13766 -24415 13824 -24381
rect 13766 -24449 13778 -24415
rect 13812 -24449 13824 -24415
rect 13766 -24483 13824 -24449
rect 13766 -24517 13778 -24483
rect 13812 -24517 13824 -24483
rect 13766 -24551 13824 -24517
rect 13766 -24585 13778 -24551
rect 13812 -24585 13824 -24551
rect 13766 -24619 13824 -24585
rect 13766 -24653 13778 -24619
rect 13812 -24653 13824 -24619
rect 13766 -24698 13824 -24653
rect 14784 -24143 14842 -24098
rect 14784 -24177 14796 -24143
rect 14830 -24177 14842 -24143
rect 14784 -24211 14842 -24177
rect 14784 -24245 14796 -24211
rect 14830 -24245 14842 -24211
rect 14784 -24279 14842 -24245
rect 14784 -24313 14796 -24279
rect 14830 -24313 14842 -24279
rect 14784 -24347 14842 -24313
rect 14784 -24381 14796 -24347
rect 14830 -24381 14842 -24347
rect 14784 -24415 14842 -24381
rect 14784 -24449 14796 -24415
rect 14830 -24449 14842 -24415
rect 14784 -24483 14842 -24449
rect 14784 -24517 14796 -24483
rect 14830 -24517 14842 -24483
rect 14784 -24551 14842 -24517
rect 14784 -24585 14796 -24551
rect 14830 -24585 14842 -24551
rect 14784 -24619 14842 -24585
rect 14784 -24653 14796 -24619
rect 14830 -24653 14842 -24619
rect 14784 -24698 14842 -24653
rect 15802 -24143 15860 -24098
rect 15802 -24177 15814 -24143
rect 15848 -24177 15860 -24143
rect 15802 -24211 15860 -24177
rect 15802 -24245 15814 -24211
rect 15848 -24245 15860 -24211
rect 15802 -24279 15860 -24245
rect 15802 -24313 15814 -24279
rect 15848 -24313 15860 -24279
rect 15802 -24347 15860 -24313
rect 15802 -24381 15814 -24347
rect 15848 -24381 15860 -24347
rect 15802 -24415 15860 -24381
rect 15802 -24449 15814 -24415
rect 15848 -24449 15860 -24415
rect 15802 -24483 15860 -24449
rect 15802 -24517 15814 -24483
rect 15848 -24517 15860 -24483
rect 15802 -24551 15860 -24517
rect 15802 -24585 15814 -24551
rect 15848 -24585 15860 -24551
rect 15802 -24619 15860 -24585
rect 15802 -24653 15814 -24619
rect 15848 -24653 15860 -24619
rect 15802 -24698 15860 -24653
rect 16820 -24143 16878 -24098
rect 16820 -24177 16832 -24143
rect 16866 -24177 16878 -24143
rect 16820 -24211 16878 -24177
rect 16820 -24245 16832 -24211
rect 16866 -24245 16878 -24211
rect 16820 -24279 16878 -24245
rect 16820 -24313 16832 -24279
rect 16866 -24313 16878 -24279
rect 16820 -24347 16878 -24313
rect 16820 -24381 16832 -24347
rect 16866 -24381 16878 -24347
rect 16820 -24415 16878 -24381
rect 16820 -24449 16832 -24415
rect 16866 -24449 16878 -24415
rect 16820 -24483 16878 -24449
rect 16820 -24517 16832 -24483
rect 16866 -24517 16878 -24483
rect 16820 -24551 16878 -24517
rect 16820 -24585 16832 -24551
rect 16866 -24585 16878 -24551
rect 16820 -24619 16878 -24585
rect 16820 -24653 16832 -24619
rect 16866 -24653 16878 -24619
rect 16820 -24698 16878 -24653
rect 17838 -24143 17896 -24098
rect 17838 -24177 17850 -24143
rect 17884 -24177 17896 -24143
rect 17838 -24211 17896 -24177
rect 17838 -24245 17850 -24211
rect 17884 -24245 17896 -24211
rect 17838 -24279 17896 -24245
rect 17838 -24313 17850 -24279
rect 17884 -24313 17896 -24279
rect 17838 -24347 17896 -24313
rect 17838 -24381 17850 -24347
rect 17884 -24381 17896 -24347
rect 17838 -24415 17896 -24381
rect 17838 -24449 17850 -24415
rect 17884 -24449 17896 -24415
rect 17838 -24483 17896 -24449
rect 17838 -24517 17850 -24483
rect 17884 -24517 17896 -24483
rect 17838 -24551 17896 -24517
rect 17838 -24585 17850 -24551
rect 17884 -24585 17896 -24551
rect 17838 -24619 17896 -24585
rect 17838 -24653 17850 -24619
rect 17884 -24653 17896 -24619
rect 17838 -24698 17896 -24653
rect 18856 -24143 18914 -24098
rect 18856 -24177 18868 -24143
rect 18902 -24177 18914 -24143
rect 18856 -24211 18914 -24177
rect 18856 -24245 18868 -24211
rect 18902 -24245 18914 -24211
rect 18856 -24279 18914 -24245
rect 18856 -24313 18868 -24279
rect 18902 -24313 18914 -24279
rect 18856 -24347 18914 -24313
rect 18856 -24381 18868 -24347
rect 18902 -24381 18914 -24347
rect 18856 -24415 18914 -24381
rect 18856 -24449 18868 -24415
rect 18902 -24449 18914 -24415
rect 18856 -24483 18914 -24449
rect 18856 -24517 18868 -24483
rect 18902 -24517 18914 -24483
rect 18856 -24551 18914 -24517
rect 18856 -24585 18868 -24551
rect 18902 -24585 18914 -24551
rect 18856 -24619 18914 -24585
rect 18856 -24653 18868 -24619
rect 18902 -24653 18914 -24619
rect 18856 -24698 18914 -24653
rect 19874 -24143 19932 -24098
rect 19874 -24177 19886 -24143
rect 19920 -24177 19932 -24143
rect 19874 -24211 19932 -24177
rect 19874 -24245 19886 -24211
rect 19920 -24245 19932 -24211
rect 19874 -24279 19932 -24245
rect 19874 -24313 19886 -24279
rect 19920 -24313 19932 -24279
rect 19874 -24347 19932 -24313
rect 19874 -24381 19886 -24347
rect 19920 -24381 19932 -24347
rect 19874 -24415 19932 -24381
rect 19874 -24449 19886 -24415
rect 19920 -24449 19932 -24415
rect 19874 -24483 19932 -24449
rect 19874 -24517 19886 -24483
rect 19920 -24517 19932 -24483
rect 19874 -24551 19932 -24517
rect 19874 -24585 19886 -24551
rect 19920 -24585 19932 -24551
rect 19874 -24619 19932 -24585
rect 19874 -24653 19886 -24619
rect 19920 -24653 19932 -24619
rect 19874 -24698 19932 -24653
rect 20892 -24143 20950 -24098
rect 20892 -24177 20904 -24143
rect 20938 -24177 20950 -24143
rect 20892 -24211 20950 -24177
rect 20892 -24245 20904 -24211
rect 20938 -24245 20950 -24211
rect 20892 -24279 20950 -24245
rect 20892 -24313 20904 -24279
rect 20938 -24313 20950 -24279
rect 20892 -24347 20950 -24313
rect 20892 -24381 20904 -24347
rect 20938 -24381 20950 -24347
rect 20892 -24415 20950 -24381
rect 20892 -24449 20904 -24415
rect 20938 -24449 20950 -24415
rect 20892 -24483 20950 -24449
rect 20892 -24517 20904 -24483
rect 20938 -24517 20950 -24483
rect 20892 -24551 20950 -24517
rect 20892 -24585 20904 -24551
rect 20938 -24585 20950 -24551
rect 20892 -24619 20950 -24585
rect 20892 -24653 20904 -24619
rect 20938 -24653 20950 -24619
rect 20892 -24698 20950 -24653
rect 21910 -24143 21968 -24098
rect 21910 -24177 21922 -24143
rect 21956 -24177 21968 -24143
rect 21910 -24211 21968 -24177
rect 21910 -24245 21922 -24211
rect 21956 -24245 21968 -24211
rect 21910 -24279 21968 -24245
rect 21910 -24313 21922 -24279
rect 21956 -24313 21968 -24279
rect 21910 -24347 21968 -24313
rect 21910 -24381 21922 -24347
rect 21956 -24381 21968 -24347
rect 21910 -24415 21968 -24381
rect 21910 -24449 21922 -24415
rect 21956 -24449 21968 -24415
rect 21910 -24483 21968 -24449
rect 21910 -24517 21922 -24483
rect 21956 -24517 21968 -24483
rect 21910 -24551 21968 -24517
rect 21910 -24585 21922 -24551
rect 21956 -24585 21968 -24551
rect 21910 -24619 21968 -24585
rect 21910 -24653 21922 -24619
rect 21956 -24653 21968 -24619
rect 21910 -24698 21968 -24653
rect 22928 -24143 22986 -24098
rect 22928 -24177 22940 -24143
rect 22974 -24177 22986 -24143
rect 22928 -24211 22986 -24177
rect 22928 -24245 22940 -24211
rect 22974 -24245 22986 -24211
rect 22928 -24279 22986 -24245
rect 22928 -24313 22940 -24279
rect 22974 -24313 22986 -24279
rect 22928 -24347 22986 -24313
rect 22928 -24381 22940 -24347
rect 22974 -24381 22986 -24347
rect 22928 -24415 22986 -24381
rect 22928 -24449 22940 -24415
rect 22974 -24449 22986 -24415
rect 22928 -24483 22986 -24449
rect 22928 -24517 22940 -24483
rect 22974 -24517 22986 -24483
rect 22928 -24551 22986 -24517
rect 22928 -24585 22940 -24551
rect 22974 -24585 22986 -24551
rect 22928 -24619 22986 -24585
rect 22928 -24653 22940 -24619
rect 22974 -24653 22986 -24619
rect 22928 -24698 22986 -24653
<< ndiffc >>
rect -9184 -12591 -9150 -12557
rect -9184 -12659 -9150 -12625
rect -9184 -12727 -9150 -12693
rect -9184 -12795 -9150 -12761
rect -9184 -12863 -9150 -12829
rect -9184 -12931 -9150 -12897
rect -9184 -12999 -9150 -12965
rect -9184 -13067 -9150 -13033
rect -8166 -12591 -8132 -12557
rect -8166 -12659 -8132 -12625
rect -8166 -12727 -8132 -12693
rect -8166 -12795 -8132 -12761
rect -8166 -12863 -8132 -12829
rect -8166 -12931 -8132 -12897
rect -8166 -12999 -8132 -12965
rect -8166 -13067 -8132 -13033
rect -7148 -12591 -7114 -12557
rect -7148 -12659 -7114 -12625
rect -7148 -12727 -7114 -12693
rect -7148 -12795 -7114 -12761
rect -7148 -12863 -7114 -12829
rect -7148 -12931 -7114 -12897
rect -7148 -12999 -7114 -12965
rect -7148 -13067 -7114 -13033
rect -6130 -12591 -6096 -12557
rect -6130 -12659 -6096 -12625
rect -6130 -12727 -6096 -12693
rect -6130 -12795 -6096 -12761
rect -6130 -12863 -6096 -12829
rect -6130 -12931 -6096 -12897
rect -6130 -12999 -6096 -12965
rect -6130 -13067 -6096 -13033
rect -5112 -12591 -5078 -12557
rect -5112 -12659 -5078 -12625
rect -5112 -12727 -5078 -12693
rect -5112 -12795 -5078 -12761
rect -5112 -12863 -5078 -12829
rect -5112 -12931 -5078 -12897
rect -5112 -12999 -5078 -12965
rect -5112 -13067 -5078 -13033
rect -4094 -12591 -4060 -12557
rect -4094 -12659 -4060 -12625
rect -4094 -12727 -4060 -12693
rect -4094 -12795 -4060 -12761
rect -4094 -12863 -4060 -12829
rect -4094 -12931 -4060 -12897
rect -4094 -12999 -4060 -12965
rect -4094 -13067 -4060 -13033
rect -3076 -12591 -3042 -12557
rect -3076 -12659 -3042 -12625
rect -3076 -12727 -3042 -12693
rect -3076 -12795 -3042 -12761
rect -3076 -12863 -3042 -12829
rect -3076 -12931 -3042 -12897
rect -3076 -12999 -3042 -12965
rect -3076 -13067 -3042 -13033
rect -2058 -12591 -2024 -12557
rect -2058 -12659 -2024 -12625
rect -2058 -12727 -2024 -12693
rect -2058 -12795 -2024 -12761
rect -2058 -12863 -2024 -12829
rect -2058 -12931 -2024 -12897
rect -2058 -12999 -2024 -12965
rect -2058 -13067 -2024 -13033
rect -1040 -12591 -1006 -12557
rect -1040 -12659 -1006 -12625
rect -1040 -12727 -1006 -12693
rect -1040 -12795 -1006 -12761
rect -1040 -12863 -1006 -12829
rect -1040 -12931 -1006 -12897
rect -1040 -12999 -1006 -12965
rect -1040 -13067 -1006 -13033
rect -22 -12591 12 -12557
rect -22 -12659 12 -12625
rect -22 -12727 12 -12693
rect -22 -12795 12 -12761
rect -22 -12863 12 -12829
rect -22 -12931 12 -12897
rect -22 -12999 12 -12965
rect -22 -13067 12 -13033
rect -9184 -13409 -9150 -13375
rect -9184 -13477 -9150 -13443
rect -9184 -13545 -9150 -13511
rect -9184 -13613 -9150 -13579
rect -9184 -13681 -9150 -13647
rect -9184 -13749 -9150 -13715
rect -9184 -13817 -9150 -13783
rect -9184 -13885 -9150 -13851
rect -8166 -13409 -8132 -13375
rect -8166 -13477 -8132 -13443
rect -8166 -13545 -8132 -13511
rect -8166 -13613 -8132 -13579
rect -8166 -13681 -8132 -13647
rect -8166 -13749 -8132 -13715
rect -8166 -13817 -8132 -13783
rect -8166 -13885 -8132 -13851
rect -7148 -13409 -7114 -13375
rect -7148 -13477 -7114 -13443
rect -7148 -13545 -7114 -13511
rect -7148 -13613 -7114 -13579
rect -7148 -13681 -7114 -13647
rect -7148 -13749 -7114 -13715
rect -7148 -13817 -7114 -13783
rect -7148 -13885 -7114 -13851
rect -6130 -13409 -6096 -13375
rect -6130 -13477 -6096 -13443
rect -6130 -13545 -6096 -13511
rect -6130 -13613 -6096 -13579
rect -6130 -13681 -6096 -13647
rect -6130 -13749 -6096 -13715
rect -6130 -13817 -6096 -13783
rect -6130 -13885 -6096 -13851
rect -5112 -13409 -5078 -13375
rect -5112 -13477 -5078 -13443
rect -5112 -13545 -5078 -13511
rect -5112 -13613 -5078 -13579
rect -5112 -13681 -5078 -13647
rect -5112 -13749 -5078 -13715
rect -5112 -13817 -5078 -13783
rect -5112 -13885 -5078 -13851
rect -4094 -13409 -4060 -13375
rect -4094 -13477 -4060 -13443
rect -4094 -13545 -4060 -13511
rect -4094 -13613 -4060 -13579
rect -4094 -13681 -4060 -13647
rect -4094 -13749 -4060 -13715
rect -4094 -13817 -4060 -13783
rect -4094 -13885 -4060 -13851
rect -3076 -13409 -3042 -13375
rect -3076 -13477 -3042 -13443
rect -3076 -13545 -3042 -13511
rect -3076 -13613 -3042 -13579
rect -3076 -13681 -3042 -13647
rect -3076 -13749 -3042 -13715
rect -3076 -13817 -3042 -13783
rect -3076 -13885 -3042 -13851
rect -2058 -13409 -2024 -13375
rect -2058 -13477 -2024 -13443
rect -2058 -13545 -2024 -13511
rect -2058 -13613 -2024 -13579
rect -2058 -13681 -2024 -13647
rect -2058 -13749 -2024 -13715
rect -2058 -13817 -2024 -13783
rect -2058 -13885 -2024 -13851
rect -1040 -13409 -1006 -13375
rect -1040 -13477 -1006 -13443
rect -1040 -13545 -1006 -13511
rect -1040 -13613 -1006 -13579
rect -1040 -13681 -1006 -13647
rect -1040 -13749 -1006 -13715
rect -1040 -13817 -1006 -13783
rect -1040 -13885 -1006 -13851
rect -22 -13409 12 -13375
rect -22 -13477 12 -13443
rect -22 -13545 12 -13511
rect -22 -13613 12 -13579
rect -22 -13681 12 -13647
rect -22 -13749 12 -13715
rect -22 -13817 12 -13783
rect -22 -13885 12 -13851
rect -9184 -14227 -9150 -14193
rect -9184 -14295 -9150 -14261
rect -9184 -14363 -9150 -14329
rect -9184 -14431 -9150 -14397
rect -9184 -14499 -9150 -14465
rect -9184 -14567 -9150 -14533
rect -9184 -14635 -9150 -14601
rect -9184 -14703 -9150 -14669
rect -8166 -14227 -8132 -14193
rect -8166 -14295 -8132 -14261
rect -8166 -14363 -8132 -14329
rect -8166 -14431 -8132 -14397
rect -8166 -14499 -8132 -14465
rect -8166 -14567 -8132 -14533
rect -8166 -14635 -8132 -14601
rect -8166 -14703 -8132 -14669
rect -7148 -14227 -7114 -14193
rect -7148 -14295 -7114 -14261
rect -7148 -14363 -7114 -14329
rect -7148 -14431 -7114 -14397
rect -7148 -14499 -7114 -14465
rect -7148 -14567 -7114 -14533
rect -7148 -14635 -7114 -14601
rect -7148 -14703 -7114 -14669
rect -6130 -14227 -6096 -14193
rect -6130 -14295 -6096 -14261
rect -6130 -14363 -6096 -14329
rect -6130 -14431 -6096 -14397
rect -6130 -14499 -6096 -14465
rect -6130 -14567 -6096 -14533
rect -6130 -14635 -6096 -14601
rect -6130 -14703 -6096 -14669
rect -5112 -14227 -5078 -14193
rect -5112 -14295 -5078 -14261
rect -5112 -14363 -5078 -14329
rect -5112 -14431 -5078 -14397
rect -5112 -14499 -5078 -14465
rect -5112 -14567 -5078 -14533
rect -5112 -14635 -5078 -14601
rect -5112 -14703 -5078 -14669
rect -4094 -14227 -4060 -14193
rect -4094 -14295 -4060 -14261
rect -4094 -14363 -4060 -14329
rect -4094 -14431 -4060 -14397
rect -4094 -14499 -4060 -14465
rect -4094 -14567 -4060 -14533
rect -4094 -14635 -4060 -14601
rect -4094 -14703 -4060 -14669
rect -3076 -14227 -3042 -14193
rect -3076 -14295 -3042 -14261
rect -3076 -14363 -3042 -14329
rect -3076 -14431 -3042 -14397
rect -3076 -14499 -3042 -14465
rect -3076 -14567 -3042 -14533
rect -3076 -14635 -3042 -14601
rect -3076 -14703 -3042 -14669
rect -2058 -14227 -2024 -14193
rect -2058 -14295 -2024 -14261
rect -2058 -14363 -2024 -14329
rect -2058 -14431 -2024 -14397
rect -2058 -14499 -2024 -14465
rect -2058 -14567 -2024 -14533
rect -2058 -14635 -2024 -14601
rect -2058 -14703 -2024 -14669
rect -1040 -14227 -1006 -14193
rect -1040 -14295 -1006 -14261
rect -1040 -14363 -1006 -14329
rect -1040 -14431 -1006 -14397
rect -1040 -14499 -1006 -14465
rect -1040 -14567 -1006 -14533
rect -1040 -14635 -1006 -14601
rect -1040 -14703 -1006 -14669
rect -22 -14227 12 -14193
rect -22 -14295 12 -14261
rect -22 -14363 12 -14329
rect -22 -14431 12 -14397
rect -22 -14499 12 -14465
rect -22 -14567 12 -14533
rect -22 -14635 12 -14601
rect -22 -14703 12 -14669
rect 2582 -14311 2616 -14277
rect 2582 -14379 2616 -14345
rect 2582 -14447 2616 -14413
rect 2582 -14515 2616 -14481
rect 2582 -14583 2616 -14549
rect 2582 -14651 2616 -14617
rect 2582 -14719 2616 -14685
rect 2582 -14787 2616 -14753
rect 3600 -14311 3634 -14277
rect 3600 -14379 3634 -14345
rect 3600 -14447 3634 -14413
rect 3600 -14515 3634 -14481
rect 3600 -14583 3634 -14549
rect 3600 -14651 3634 -14617
rect 3600 -14719 3634 -14685
rect 3600 -14787 3634 -14753
rect 4618 -14311 4652 -14277
rect 4618 -14379 4652 -14345
rect 4618 -14447 4652 -14413
rect 4618 -14515 4652 -14481
rect 4618 -14583 4652 -14549
rect 4618 -14651 4652 -14617
rect 4618 -14719 4652 -14685
rect 4618 -14787 4652 -14753
rect 5636 -14311 5670 -14277
rect 5636 -14379 5670 -14345
rect 5636 -14447 5670 -14413
rect 5636 -14515 5670 -14481
rect 5636 -14583 5670 -14549
rect 5636 -14651 5670 -14617
rect 5636 -14719 5670 -14685
rect 5636 -14787 5670 -14753
rect 6654 -14311 6688 -14277
rect 6654 -14379 6688 -14345
rect 6654 -14447 6688 -14413
rect 6654 -14515 6688 -14481
rect 6654 -14583 6688 -14549
rect 6654 -14651 6688 -14617
rect 6654 -14719 6688 -14685
rect 6654 -14787 6688 -14753
rect 7672 -14311 7706 -14277
rect 7672 -14379 7706 -14345
rect 7672 -14447 7706 -14413
rect 7672 -14515 7706 -14481
rect 7672 -14583 7706 -14549
rect 7672 -14651 7706 -14617
rect 7672 -14719 7706 -14685
rect 7672 -14787 7706 -14753
rect 8690 -14311 8724 -14277
rect 8690 -14379 8724 -14345
rect 8690 -14447 8724 -14413
rect 8690 -14515 8724 -14481
rect 8690 -14583 8724 -14549
rect 8690 -14651 8724 -14617
rect 8690 -14719 8724 -14685
rect 8690 -14787 8724 -14753
rect 9708 -14311 9742 -14277
rect 9708 -14379 9742 -14345
rect 9708 -14447 9742 -14413
rect 9708 -14515 9742 -14481
rect 9708 -14583 9742 -14549
rect 9708 -14651 9742 -14617
rect 9708 -14719 9742 -14685
rect 9708 -14787 9742 -14753
rect 10726 -14311 10760 -14277
rect 10726 -14379 10760 -14345
rect 10726 -14447 10760 -14413
rect 10726 -14515 10760 -14481
rect 10726 -14583 10760 -14549
rect 10726 -14651 10760 -14617
rect 10726 -14719 10760 -14685
rect 10726 -14787 10760 -14753
rect 11744 -14311 11778 -14277
rect 11744 -14379 11778 -14345
rect 11744 -14447 11778 -14413
rect 11744 -14515 11778 -14481
rect 11744 -14583 11778 -14549
rect 11744 -14651 11778 -14617
rect 11744 -14719 11778 -14685
rect 11744 -14787 11778 -14753
rect 12762 -14311 12796 -14277
rect 12762 -14379 12796 -14345
rect 12762 -14447 12796 -14413
rect 12762 -14515 12796 -14481
rect 12762 -14583 12796 -14549
rect 12762 -14651 12796 -14617
rect 12762 -14719 12796 -14685
rect 12762 -14787 12796 -14753
rect 13780 -14311 13814 -14277
rect 13780 -14379 13814 -14345
rect 13780 -14447 13814 -14413
rect 13780 -14515 13814 -14481
rect 13780 -14583 13814 -14549
rect 13780 -14651 13814 -14617
rect 13780 -14719 13814 -14685
rect 13780 -14787 13814 -14753
rect 14798 -14311 14832 -14277
rect 14798 -14379 14832 -14345
rect 14798 -14447 14832 -14413
rect 14798 -14515 14832 -14481
rect 14798 -14583 14832 -14549
rect 14798 -14651 14832 -14617
rect 14798 -14719 14832 -14685
rect 14798 -14787 14832 -14753
rect 15816 -14311 15850 -14277
rect 15816 -14379 15850 -14345
rect 15816 -14447 15850 -14413
rect 15816 -14515 15850 -14481
rect 15816 -14583 15850 -14549
rect 15816 -14651 15850 -14617
rect 15816 -14719 15850 -14685
rect 15816 -14787 15850 -14753
rect 16834 -14311 16868 -14277
rect 16834 -14379 16868 -14345
rect 16834 -14447 16868 -14413
rect 16834 -14515 16868 -14481
rect 16834 -14583 16868 -14549
rect 16834 -14651 16868 -14617
rect 16834 -14719 16868 -14685
rect 16834 -14787 16868 -14753
rect 17852 -14311 17886 -14277
rect 17852 -14379 17886 -14345
rect 17852 -14447 17886 -14413
rect 17852 -14515 17886 -14481
rect 17852 -14583 17886 -14549
rect 17852 -14651 17886 -14617
rect 17852 -14719 17886 -14685
rect 17852 -14787 17886 -14753
rect 18870 -14311 18904 -14277
rect 18870 -14379 18904 -14345
rect 18870 -14447 18904 -14413
rect 18870 -14515 18904 -14481
rect 18870 -14583 18904 -14549
rect 18870 -14651 18904 -14617
rect 18870 -14719 18904 -14685
rect 18870 -14787 18904 -14753
rect 19888 -14311 19922 -14277
rect 19888 -14379 19922 -14345
rect 19888 -14447 19922 -14413
rect 19888 -14515 19922 -14481
rect 19888 -14583 19922 -14549
rect 19888 -14651 19922 -14617
rect 19888 -14719 19922 -14685
rect 19888 -14787 19922 -14753
rect 20906 -14311 20940 -14277
rect 20906 -14379 20940 -14345
rect 20906 -14447 20940 -14413
rect 20906 -14515 20940 -14481
rect 20906 -14583 20940 -14549
rect 20906 -14651 20940 -14617
rect 20906 -14719 20940 -14685
rect 20906 -14787 20940 -14753
rect 21924 -14311 21958 -14277
rect 21924 -14379 21958 -14345
rect 21924 -14447 21958 -14413
rect 21924 -14515 21958 -14481
rect 21924 -14583 21958 -14549
rect 21924 -14651 21958 -14617
rect 21924 -14719 21958 -14685
rect 21924 -14787 21958 -14753
rect 22942 -14311 22976 -14277
rect 22942 -14379 22976 -14345
rect 22942 -14447 22976 -14413
rect 22942 -14515 22976 -14481
rect 22942 -14583 22976 -14549
rect 22942 -14651 22976 -14617
rect 22942 -14719 22976 -14685
rect 22942 -14787 22976 -14753
rect -9184 -15045 -9150 -15011
rect -9184 -15113 -9150 -15079
rect -9184 -15181 -9150 -15147
rect -9184 -15249 -9150 -15215
rect -9184 -15317 -9150 -15283
rect -9184 -15385 -9150 -15351
rect -9184 -15453 -9150 -15419
rect -9184 -15521 -9150 -15487
rect -8166 -15045 -8132 -15011
rect -8166 -15113 -8132 -15079
rect -8166 -15181 -8132 -15147
rect -8166 -15249 -8132 -15215
rect -8166 -15317 -8132 -15283
rect -8166 -15385 -8132 -15351
rect -8166 -15453 -8132 -15419
rect -8166 -15521 -8132 -15487
rect -7148 -15045 -7114 -15011
rect -7148 -15113 -7114 -15079
rect -7148 -15181 -7114 -15147
rect -7148 -15249 -7114 -15215
rect -7148 -15317 -7114 -15283
rect -7148 -15385 -7114 -15351
rect -7148 -15453 -7114 -15419
rect -7148 -15521 -7114 -15487
rect -6130 -15045 -6096 -15011
rect -6130 -15113 -6096 -15079
rect -6130 -15181 -6096 -15147
rect -6130 -15249 -6096 -15215
rect -6130 -15317 -6096 -15283
rect -6130 -15385 -6096 -15351
rect -6130 -15453 -6096 -15419
rect -6130 -15521 -6096 -15487
rect -5112 -15045 -5078 -15011
rect -5112 -15113 -5078 -15079
rect -5112 -15181 -5078 -15147
rect -5112 -15249 -5078 -15215
rect -5112 -15317 -5078 -15283
rect -5112 -15385 -5078 -15351
rect -5112 -15453 -5078 -15419
rect -5112 -15521 -5078 -15487
rect -4094 -15045 -4060 -15011
rect -4094 -15113 -4060 -15079
rect -4094 -15181 -4060 -15147
rect -4094 -15249 -4060 -15215
rect -4094 -15317 -4060 -15283
rect -4094 -15385 -4060 -15351
rect -4094 -15453 -4060 -15419
rect -4094 -15521 -4060 -15487
rect -3076 -15045 -3042 -15011
rect -3076 -15113 -3042 -15079
rect -3076 -15181 -3042 -15147
rect -3076 -15249 -3042 -15215
rect -3076 -15317 -3042 -15283
rect -3076 -15385 -3042 -15351
rect -3076 -15453 -3042 -15419
rect -3076 -15521 -3042 -15487
rect -2058 -15045 -2024 -15011
rect -2058 -15113 -2024 -15079
rect -2058 -15181 -2024 -15147
rect -2058 -15249 -2024 -15215
rect -2058 -15317 -2024 -15283
rect -2058 -15385 -2024 -15351
rect -2058 -15453 -2024 -15419
rect -2058 -15521 -2024 -15487
rect -1040 -15045 -1006 -15011
rect -1040 -15113 -1006 -15079
rect -1040 -15181 -1006 -15147
rect -1040 -15249 -1006 -15215
rect -1040 -15317 -1006 -15283
rect -1040 -15385 -1006 -15351
rect -1040 -15453 -1006 -15419
rect -1040 -15521 -1006 -15487
rect -22 -15045 12 -15011
rect -22 -15113 12 -15079
rect -22 -15181 12 -15147
rect -22 -15249 12 -15215
rect -22 -15317 12 -15283
rect -22 -15385 12 -15351
rect -22 -15453 12 -15419
rect -22 -15521 12 -15487
rect 2582 -15543 2616 -15509
rect 2582 -15611 2616 -15577
rect 2582 -15679 2616 -15645
rect 2582 -15747 2616 -15713
rect -9184 -15863 -9150 -15829
rect -9184 -15931 -9150 -15897
rect -9184 -15999 -9150 -15965
rect -9184 -16067 -9150 -16033
rect -9184 -16135 -9150 -16101
rect -9184 -16203 -9150 -16169
rect -9184 -16271 -9150 -16237
rect -9184 -16339 -9150 -16305
rect -8166 -15863 -8132 -15829
rect -8166 -15931 -8132 -15897
rect -8166 -15999 -8132 -15965
rect -8166 -16067 -8132 -16033
rect -8166 -16135 -8132 -16101
rect -8166 -16203 -8132 -16169
rect -8166 -16271 -8132 -16237
rect -8166 -16339 -8132 -16305
rect -7148 -15863 -7114 -15829
rect -7148 -15931 -7114 -15897
rect -7148 -15999 -7114 -15965
rect -7148 -16067 -7114 -16033
rect -7148 -16135 -7114 -16101
rect -7148 -16203 -7114 -16169
rect -7148 -16271 -7114 -16237
rect -7148 -16339 -7114 -16305
rect -6130 -15863 -6096 -15829
rect -6130 -15931 -6096 -15897
rect -6130 -15999 -6096 -15965
rect -6130 -16067 -6096 -16033
rect -6130 -16135 -6096 -16101
rect -6130 -16203 -6096 -16169
rect -6130 -16271 -6096 -16237
rect -6130 -16339 -6096 -16305
rect -5112 -15863 -5078 -15829
rect -5112 -15931 -5078 -15897
rect -5112 -15999 -5078 -15965
rect -5112 -16067 -5078 -16033
rect -5112 -16135 -5078 -16101
rect -5112 -16203 -5078 -16169
rect -5112 -16271 -5078 -16237
rect -5112 -16339 -5078 -16305
rect -4094 -15863 -4060 -15829
rect -4094 -15931 -4060 -15897
rect -4094 -15999 -4060 -15965
rect -4094 -16067 -4060 -16033
rect -4094 -16135 -4060 -16101
rect -4094 -16203 -4060 -16169
rect -4094 -16271 -4060 -16237
rect -4094 -16339 -4060 -16305
rect -3076 -15863 -3042 -15829
rect -3076 -15931 -3042 -15897
rect -3076 -15999 -3042 -15965
rect -3076 -16067 -3042 -16033
rect -3076 -16135 -3042 -16101
rect -3076 -16203 -3042 -16169
rect -3076 -16271 -3042 -16237
rect -3076 -16339 -3042 -16305
rect -2058 -15863 -2024 -15829
rect -2058 -15931 -2024 -15897
rect -2058 -15999 -2024 -15965
rect -2058 -16067 -2024 -16033
rect -2058 -16135 -2024 -16101
rect -2058 -16203 -2024 -16169
rect -2058 -16271 -2024 -16237
rect -2058 -16339 -2024 -16305
rect -1040 -15863 -1006 -15829
rect -1040 -15931 -1006 -15897
rect -1040 -15999 -1006 -15965
rect -1040 -16067 -1006 -16033
rect -1040 -16135 -1006 -16101
rect -1040 -16203 -1006 -16169
rect -1040 -16271 -1006 -16237
rect -1040 -16339 -1006 -16305
rect -22 -15863 12 -15829
rect -22 -15931 12 -15897
rect -22 -15999 12 -15965
rect -22 -16067 12 -16033
rect 2582 -15815 2616 -15781
rect 2582 -15883 2616 -15849
rect 2582 -15951 2616 -15917
rect 2582 -16019 2616 -15985
rect 3600 -15543 3634 -15509
rect 3600 -15611 3634 -15577
rect 3600 -15679 3634 -15645
rect 3600 -15747 3634 -15713
rect 3600 -15815 3634 -15781
rect 3600 -15883 3634 -15849
rect 3600 -15951 3634 -15917
rect 3600 -16019 3634 -15985
rect 4618 -15543 4652 -15509
rect 4618 -15611 4652 -15577
rect 4618 -15679 4652 -15645
rect 4618 -15747 4652 -15713
rect 4618 -15815 4652 -15781
rect 4618 -15883 4652 -15849
rect 4618 -15951 4652 -15917
rect 4618 -16019 4652 -15985
rect 5636 -15543 5670 -15509
rect 5636 -15611 5670 -15577
rect 5636 -15679 5670 -15645
rect 5636 -15747 5670 -15713
rect 5636 -15815 5670 -15781
rect 5636 -15883 5670 -15849
rect 5636 -15951 5670 -15917
rect 5636 -16019 5670 -15985
rect 6654 -15543 6688 -15509
rect 6654 -15611 6688 -15577
rect 6654 -15679 6688 -15645
rect 6654 -15747 6688 -15713
rect 6654 -15815 6688 -15781
rect 6654 -15883 6688 -15849
rect 6654 -15951 6688 -15917
rect 6654 -16019 6688 -15985
rect 7672 -15543 7706 -15509
rect 7672 -15611 7706 -15577
rect 7672 -15679 7706 -15645
rect 7672 -15747 7706 -15713
rect 7672 -15815 7706 -15781
rect 7672 -15883 7706 -15849
rect 7672 -15951 7706 -15917
rect 7672 -16019 7706 -15985
rect 8690 -15543 8724 -15509
rect 8690 -15611 8724 -15577
rect 8690 -15679 8724 -15645
rect 8690 -15747 8724 -15713
rect 8690 -15815 8724 -15781
rect 8690 -15883 8724 -15849
rect 8690 -15951 8724 -15917
rect 8690 -16019 8724 -15985
rect 9708 -15543 9742 -15509
rect 9708 -15611 9742 -15577
rect 9708 -15679 9742 -15645
rect 9708 -15747 9742 -15713
rect 9708 -15815 9742 -15781
rect 9708 -15883 9742 -15849
rect 9708 -15951 9742 -15917
rect 9708 -16019 9742 -15985
rect 10726 -15543 10760 -15509
rect 10726 -15611 10760 -15577
rect 10726 -15679 10760 -15645
rect 10726 -15747 10760 -15713
rect 10726 -15815 10760 -15781
rect 10726 -15883 10760 -15849
rect 10726 -15951 10760 -15917
rect 10726 -16019 10760 -15985
rect 11744 -15543 11778 -15509
rect 11744 -15611 11778 -15577
rect 11744 -15679 11778 -15645
rect 11744 -15747 11778 -15713
rect 11744 -15815 11778 -15781
rect 11744 -15883 11778 -15849
rect 11744 -15951 11778 -15917
rect 11744 -16019 11778 -15985
rect 12762 -15543 12796 -15509
rect 12762 -15611 12796 -15577
rect 12762 -15679 12796 -15645
rect 12762 -15747 12796 -15713
rect 12762 -15815 12796 -15781
rect 12762 -15883 12796 -15849
rect 12762 -15951 12796 -15917
rect 12762 -16019 12796 -15985
rect 13780 -15543 13814 -15509
rect 13780 -15611 13814 -15577
rect 13780 -15679 13814 -15645
rect 13780 -15747 13814 -15713
rect 13780 -15815 13814 -15781
rect 13780 -15883 13814 -15849
rect 13780 -15951 13814 -15917
rect 13780 -16019 13814 -15985
rect 14798 -15543 14832 -15509
rect 14798 -15611 14832 -15577
rect 14798 -15679 14832 -15645
rect 14798 -15747 14832 -15713
rect 14798 -15815 14832 -15781
rect 14798 -15883 14832 -15849
rect 14798 -15951 14832 -15917
rect 14798 -16019 14832 -15985
rect 15816 -15543 15850 -15509
rect 15816 -15611 15850 -15577
rect 15816 -15679 15850 -15645
rect 15816 -15747 15850 -15713
rect 15816 -15815 15850 -15781
rect 15816 -15883 15850 -15849
rect 15816 -15951 15850 -15917
rect 15816 -16019 15850 -15985
rect 16834 -15543 16868 -15509
rect 16834 -15611 16868 -15577
rect 16834 -15679 16868 -15645
rect 16834 -15747 16868 -15713
rect 16834 -15815 16868 -15781
rect 16834 -15883 16868 -15849
rect 16834 -15951 16868 -15917
rect 16834 -16019 16868 -15985
rect 17852 -15543 17886 -15509
rect 17852 -15611 17886 -15577
rect 17852 -15679 17886 -15645
rect 17852 -15747 17886 -15713
rect 17852 -15815 17886 -15781
rect 17852 -15883 17886 -15849
rect 17852 -15951 17886 -15917
rect 17852 -16019 17886 -15985
rect 18870 -15543 18904 -15509
rect 18870 -15611 18904 -15577
rect 18870 -15679 18904 -15645
rect 18870 -15747 18904 -15713
rect 18870 -15815 18904 -15781
rect 18870 -15883 18904 -15849
rect 18870 -15951 18904 -15917
rect 18870 -16019 18904 -15985
rect 19888 -15543 19922 -15509
rect 19888 -15611 19922 -15577
rect 19888 -15679 19922 -15645
rect 19888 -15747 19922 -15713
rect 19888 -15815 19922 -15781
rect 19888 -15883 19922 -15849
rect 19888 -15951 19922 -15917
rect 19888 -16019 19922 -15985
rect 20906 -15543 20940 -15509
rect 20906 -15611 20940 -15577
rect 20906 -15679 20940 -15645
rect 20906 -15747 20940 -15713
rect 20906 -15815 20940 -15781
rect 20906 -15883 20940 -15849
rect 20906 -15951 20940 -15917
rect 20906 -16019 20940 -15985
rect 21924 -15543 21958 -15509
rect 21924 -15611 21958 -15577
rect 21924 -15679 21958 -15645
rect 21924 -15747 21958 -15713
rect 21924 -15815 21958 -15781
rect 21924 -15883 21958 -15849
rect 21924 -15951 21958 -15917
rect 21924 -16019 21958 -15985
rect 22942 -15543 22976 -15509
rect 22942 -15611 22976 -15577
rect 22942 -15679 22976 -15645
rect 22942 -15747 22976 -15713
rect 22942 -15815 22976 -15781
rect 22942 -15883 22976 -15849
rect 22942 -15951 22976 -15917
rect 22942 -16019 22976 -15985
rect -22 -16135 12 -16101
rect -22 -16203 12 -16169
rect -22 -16271 12 -16237
rect -22 -16339 12 -16305
rect -9184 -16681 -9150 -16647
rect -9184 -16749 -9150 -16715
rect -9184 -16817 -9150 -16783
rect -9184 -16885 -9150 -16851
rect -9184 -16953 -9150 -16919
rect -9184 -17021 -9150 -16987
rect -9184 -17089 -9150 -17055
rect -9184 -17157 -9150 -17123
rect -8166 -16681 -8132 -16647
rect -8166 -16749 -8132 -16715
rect -8166 -16817 -8132 -16783
rect -8166 -16885 -8132 -16851
rect -8166 -16953 -8132 -16919
rect -8166 -17021 -8132 -16987
rect -8166 -17089 -8132 -17055
rect -8166 -17157 -8132 -17123
rect -7148 -16681 -7114 -16647
rect -7148 -16749 -7114 -16715
rect -7148 -16817 -7114 -16783
rect -7148 -16885 -7114 -16851
rect -7148 -16953 -7114 -16919
rect -7148 -17021 -7114 -16987
rect -7148 -17089 -7114 -17055
rect -7148 -17157 -7114 -17123
rect -6130 -16681 -6096 -16647
rect -6130 -16749 -6096 -16715
rect -6130 -16817 -6096 -16783
rect -6130 -16885 -6096 -16851
rect -6130 -16953 -6096 -16919
rect -6130 -17021 -6096 -16987
rect -6130 -17089 -6096 -17055
rect -6130 -17157 -6096 -17123
rect -5112 -16681 -5078 -16647
rect -5112 -16749 -5078 -16715
rect -5112 -16817 -5078 -16783
rect -5112 -16885 -5078 -16851
rect -5112 -16953 -5078 -16919
rect -5112 -17021 -5078 -16987
rect -5112 -17089 -5078 -17055
rect -5112 -17157 -5078 -17123
rect -4094 -16681 -4060 -16647
rect -4094 -16749 -4060 -16715
rect -4094 -16817 -4060 -16783
rect -4094 -16885 -4060 -16851
rect -4094 -16953 -4060 -16919
rect -4094 -17021 -4060 -16987
rect -4094 -17089 -4060 -17055
rect -4094 -17157 -4060 -17123
rect -3076 -16681 -3042 -16647
rect -3076 -16749 -3042 -16715
rect -3076 -16817 -3042 -16783
rect -3076 -16885 -3042 -16851
rect -3076 -16953 -3042 -16919
rect -3076 -17021 -3042 -16987
rect -3076 -17089 -3042 -17055
rect -3076 -17157 -3042 -17123
rect -2058 -16681 -2024 -16647
rect -2058 -16749 -2024 -16715
rect -2058 -16817 -2024 -16783
rect -2058 -16885 -2024 -16851
rect -2058 -16953 -2024 -16919
rect -2058 -17021 -2024 -16987
rect -2058 -17089 -2024 -17055
rect -2058 -17157 -2024 -17123
rect -1040 -16681 -1006 -16647
rect -1040 -16749 -1006 -16715
rect -1040 -16817 -1006 -16783
rect -1040 -16885 -1006 -16851
rect -1040 -16953 -1006 -16919
rect -1040 -17021 -1006 -16987
rect -1040 -17089 -1006 -17055
rect -1040 -17157 -1006 -17123
rect -22 -16681 12 -16647
rect -22 -16749 12 -16715
rect -22 -16817 12 -16783
rect -22 -16885 12 -16851
rect -22 -16953 12 -16919
rect -22 -17021 12 -16987
rect -22 -17089 12 -17055
rect -22 -17157 12 -17123
rect 2580 -16777 2614 -16743
rect 2580 -16845 2614 -16811
rect 2580 -16913 2614 -16879
rect 2580 -16981 2614 -16947
rect 2580 -17049 2614 -17015
rect 2580 -17117 2614 -17083
rect 2580 -17185 2614 -17151
rect 2580 -17253 2614 -17219
rect 3598 -16777 3632 -16743
rect 3598 -16845 3632 -16811
rect 3598 -16913 3632 -16879
rect 3598 -16981 3632 -16947
rect 3598 -17049 3632 -17015
rect 3598 -17117 3632 -17083
rect 3598 -17185 3632 -17151
rect 3598 -17253 3632 -17219
rect 4616 -16777 4650 -16743
rect 4616 -16845 4650 -16811
rect 4616 -16913 4650 -16879
rect 4616 -16981 4650 -16947
rect 4616 -17049 4650 -17015
rect 4616 -17117 4650 -17083
rect 4616 -17185 4650 -17151
rect 4616 -17253 4650 -17219
rect 5634 -16777 5668 -16743
rect 5634 -16845 5668 -16811
rect 5634 -16913 5668 -16879
rect 5634 -16981 5668 -16947
rect 5634 -17049 5668 -17015
rect 5634 -17117 5668 -17083
rect 5634 -17185 5668 -17151
rect 5634 -17253 5668 -17219
rect 6652 -16777 6686 -16743
rect 6652 -16845 6686 -16811
rect 6652 -16913 6686 -16879
rect 6652 -16981 6686 -16947
rect 6652 -17049 6686 -17015
rect 6652 -17117 6686 -17083
rect 6652 -17185 6686 -17151
rect 6652 -17253 6686 -17219
rect 7670 -16777 7704 -16743
rect 7670 -16845 7704 -16811
rect 7670 -16913 7704 -16879
rect 7670 -16981 7704 -16947
rect 7670 -17049 7704 -17015
rect 7670 -17117 7704 -17083
rect 7670 -17185 7704 -17151
rect 7670 -17253 7704 -17219
rect 8688 -16777 8722 -16743
rect 8688 -16845 8722 -16811
rect 8688 -16913 8722 -16879
rect 8688 -16981 8722 -16947
rect 8688 -17049 8722 -17015
rect 8688 -17117 8722 -17083
rect 8688 -17185 8722 -17151
rect 8688 -17253 8722 -17219
rect 9706 -16777 9740 -16743
rect 9706 -16845 9740 -16811
rect 9706 -16913 9740 -16879
rect 9706 -16981 9740 -16947
rect 9706 -17049 9740 -17015
rect 9706 -17117 9740 -17083
rect 9706 -17185 9740 -17151
rect 9706 -17253 9740 -17219
rect 10724 -16777 10758 -16743
rect 10724 -16845 10758 -16811
rect 10724 -16913 10758 -16879
rect 10724 -16981 10758 -16947
rect 10724 -17049 10758 -17015
rect 10724 -17117 10758 -17083
rect 10724 -17185 10758 -17151
rect 10724 -17253 10758 -17219
rect 11742 -16777 11776 -16743
rect 11742 -16845 11776 -16811
rect 11742 -16913 11776 -16879
rect 11742 -16981 11776 -16947
rect 11742 -17049 11776 -17015
rect 11742 -17117 11776 -17083
rect 11742 -17185 11776 -17151
rect 11742 -17253 11776 -17219
rect 12760 -16777 12794 -16743
rect 12760 -16845 12794 -16811
rect 12760 -16913 12794 -16879
rect 12760 -16981 12794 -16947
rect 12760 -17049 12794 -17015
rect 12760 -17117 12794 -17083
rect 12760 -17185 12794 -17151
rect 12760 -17253 12794 -17219
rect 13778 -16777 13812 -16743
rect 13778 -16845 13812 -16811
rect 13778 -16913 13812 -16879
rect 13778 -16981 13812 -16947
rect 13778 -17049 13812 -17015
rect 13778 -17117 13812 -17083
rect 13778 -17185 13812 -17151
rect 13778 -17253 13812 -17219
rect 14796 -16777 14830 -16743
rect 14796 -16845 14830 -16811
rect 14796 -16913 14830 -16879
rect 14796 -16981 14830 -16947
rect 14796 -17049 14830 -17015
rect 14796 -17117 14830 -17083
rect 14796 -17185 14830 -17151
rect 14796 -17253 14830 -17219
rect 15814 -16777 15848 -16743
rect 15814 -16845 15848 -16811
rect 15814 -16913 15848 -16879
rect 15814 -16981 15848 -16947
rect 15814 -17049 15848 -17015
rect 15814 -17117 15848 -17083
rect 15814 -17185 15848 -17151
rect 15814 -17253 15848 -17219
rect 16832 -16777 16866 -16743
rect 16832 -16845 16866 -16811
rect 16832 -16913 16866 -16879
rect 16832 -16981 16866 -16947
rect 16832 -17049 16866 -17015
rect 16832 -17117 16866 -17083
rect 16832 -17185 16866 -17151
rect 16832 -17253 16866 -17219
rect 17850 -16777 17884 -16743
rect 17850 -16845 17884 -16811
rect 17850 -16913 17884 -16879
rect 17850 -16981 17884 -16947
rect 17850 -17049 17884 -17015
rect 17850 -17117 17884 -17083
rect 17850 -17185 17884 -17151
rect 17850 -17253 17884 -17219
rect 18868 -16777 18902 -16743
rect 18868 -16845 18902 -16811
rect 18868 -16913 18902 -16879
rect 18868 -16981 18902 -16947
rect 18868 -17049 18902 -17015
rect 18868 -17117 18902 -17083
rect 18868 -17185 18902 -17151
rect 18868 -17253 18902 -17219
rect 19886 -16777 19920 -16743
rect 19886 -16845 19920 -16811
rect 19886 -16913 19920 -16879
rect 19886 -16981 19920 -16947
rect 19886 -17049 19920 -17015
rect 19886 -17117 19920 -17083
rect 19886 -17185 19920 -17151
rect 19886 -17253 19920 -17219
rect 20904 -16777 20938 -16743
rect 20904 -16845 20938 -16811
rect 20904 -16913 20938 -16879
rect 20904 -16981 20938 -16947
rect 20904 -17049 20938 -17015
rect 20904 -17117 20938 -17083
rect 20904 -17185 20938 -17151
rect 20904 -17253 20938 -17219
rect 21922 -16777 21956 -16743
rect 21922 -16845 21956 -16811
rect 21922 -16913 21956 -16879
rect 21922 -16981 21956 -16947
rect 21922 -17049 21956 -17015
rect 21922 -17117 21956 -17083
rect 21922 -17185 21956 -17151
rect 21922 -17253 21956 -17219
rect 22940 -16777 22974 -16743
rect 22940 -16845 22974 -16811
rect 22940 -16913 22974 -16879
rect 22940 -16981 22974 -16947
rect 22940 -17049 22974 -17015
rect 22940 -17117 22974 -17083
rect 22940 -17185 22974 -17151
rect 22940 -17253 22974 -17219
rect -9184 -17499 -9150 -17465
rect -9184 -17567 -9150 -17533
rect -9184 -17635 -9150 -17601
rect -9184 -17703 -9150 -17669
rect -9184 -17771 -9150 -17737
rect -9184 -17839 -9150 -17805
rect -9184 -17907 -9150 -17873
rect -9184 -17975 -9150 -17941
rect -8166 -17499 -8132 -17465
rect -8166 -17567 -8132 -17533
rect -8166 -17635 -8132 -17601
rect -8166 -17703 -8132 -17669
rect -8166 -17771 -8132 -17737
rect -8166 -17839 -8132 -17805
rect -8166 -17907 -8132 -17873
rect -8166 -17975 -8132 -17941
rect -7148 -17499 -7114 -17465
rect -7148 -17567 -7114 -17533
rect -7148 -17635 -7114 -17601
rect -7148 -17703 -7114 -17669
rect -7148 -17771 -7114 -17737
rect -7148 -17839 -7114 -17805
rect -7148 -17907 -7114 -17873
rect -7148 -17975 -7114 -17941
rect -6130 -17499 -6096 -17465
rect -6130 -17567 -6096 -17533
rect -6130 -17635 -6096 -17601
rect -6130 -17703 -6096 -17669
rect -6130 -17771 -6096 -17737
rect -6130 -17839 -6096 -17805
rect -6130 -17907 -6096 -17873
rect -6130 -17975 -6096 -17941
rect -5112 -17499 -5078 -17465
rect -5112 -17567 -5078 -17533
rect -5112 -17635 -5078 -17601
rect -5112 -17703 -5078 -17669
rect -5112 -17771 -5078 -17737
rect -5112 -17839 -5078 -17805
rect -5112 -17907 -5078 -17873
rect -5112 -17975 -5078 -17941
rect -4094 -17499 -4060 -17465
rect -4094 -17567 -4060 -17533
rect -4094 -17635 -4060 -17601
rect -4094 -17703 -4060 -17669
rect -4094 -17771 -4060 -17737
rect -4094 -17839 -4060 -17805
rect -4094 -17907 -4060 -17873
rect -4094 -17975 -4060 -17941
rect -3076 -17499 -3042 -17465
rect -3076 -17567 -3042 -17533
rect -3076 -17635 -3042 -17601
rect -3076 -17703 -3042 -17669
rect -3076 -17771 -3042 -17737
rect -3076 -17839 -3042 -17805
rect -3076 -17907 -3042 -17873
rect -3076 -17975 -3042 -17941
rect -2058 -17499 -2024 -17465
rect -2058 -17567 -2024 -17533
rect -2058 -17635 -2024 -17601
rect -2058 -17703 -2024 -17669
rect -2058 -17771 -2024 -17737
rect -2058 -17839 -2024 -17805
rect -2058 -17907 -2024 -17873
rect -2058 -17975 -2024 -17941
rect -1040 -17499 -1006 -17465
rect -1040 -17567 -1006 -17533
rect -1040 -17635 -1006 -17601
rect -1040 -17703 -1006 -17669
rect -1040 -17771 -1006 -17737
rect -1040 -17839 -1006 -17805
rect -1040 -17907 -1006 -17873
rect -1040 -17975 -1006 -17941
rect -22 -17499 12 -17465
rect -22 -17567 12 -17533
rect -22 -17635 12 -17601
rect -22 -17703 12 -17669
rect -22 -17771 12 -17737
rect -22 -17839 12 -17805
rect -22 -17907 12 -17873
rect -22 -17975 12 -17941
rect 2580 -18011 2614 -17977
rect 2580 -18079 2614 -18045
rect 2580 -18147 2614 -18113
rect 2580 -18215 2614 -18181
rect -9184 -18317 -9150 -18283
rect -9184 -18385 -9150 -18351
rect -9184 -18453 -9150 -18419
rect -9184 -18521 -9150 -18487
rect -9184 -18589 -9150 -18555
rect -9184 -18657 -9150 -18623
rect -9184 -18725 -9150 -18691
rect -9184 -18793 -9150 -18759
rect -8166 -18317 -8132 -18283
rect -8166 -18385 -8132 -18351
rect -8166 -18453 -8132 -18419
rect -8166 -18521 -8132 -18487
rect -8166 -18589 -8132 -18555
rect -8166 -18657 -8132 -18623
rect -8166 -18725 -8132 -18691
rect -8166 -18793 -8132 -18759
rect -7148 -18317 -7114 -18283
rect -7148 -18385 -7114 -18351
rect -7148 -18453 -7114 -18419
rect -7148 -18521 -7114 -18487
rect -7148 -18589 -7114 -18555
rect -7148 -18657 -7114 -18623
rect -7148 -18725 -7114 -18691
rect -7148 -18793 -7114 -18759
rect -6130 -18317 -6096 -18283
rect -6130 -18385 -6096 -18351
rect -6130 -18453 -6096 -18419
rect -6130 -18521 -6096 -18487
rect -6130 -18589 -6096 -18555
rect -6130 -18657 -6096 -18623
rect -6130 -18725 -6096 -18691
rect -6130 -18793 -6096 -18759
rect -5112 -18317 -5078 -18283
rect -5112 -18385 -5078 -18351
rect -5112 -18453 -5078 -18419
rect -5112 -18521 -5078 -18487
rect -5112 -18589 -5078 -18555
rect -5112 -18657 -5078 -18623
rect -5112 -18725 -5078 -18691
rect -5112 -18793 -5078 -18759
rect -4094 -18317 -4060 -18283
rect -4094 -18385 -4060 -18351
rect -4094 -18453 -4060 -18419
rect -4094 -18521 -4060 -18487
rect -4094 -18589 -4060 -18555
rect -4094 -18657 -4060 -18623
rect -4094 -18725 -4060 -18691
rect -4094 -18793 -4060 -18759
rect -3076 -18317 -3042 -18283
rect -3076 -18385 -3042 -18351
rect -3076 -18453 -3042 -18419
rect -3076 -18521 -3042 -18487
rect -3076 -18589 -3042 -18555
rect -3076 -18657 -3042 -18623
rect -3076 -18725 -3042 -18691
rect -3076 -18793 -3042 -18759
rect -2058 -18317 -2024 -18283
rect -2058 -18385 -2024 -18351
rect -2058 -18453 -2024 -18419
rect -2058 -18521 -2024 -18487
rect -2058 -18589 -2024 -18555
rect -2058 -18657 -2024 -18623
rect -2058 -18725 -2024 -18691
rect -2058 -18793 -2024 -18759
rect -1040 -18317 -1006 -18283
rect -1040 -18385 -1006 -18351
rect -1040 -18453 -1006 -18419
rect -1040 -18521 -1006 -18487
rect -1040 -18589 -1006 -18555
rect -1040 -18657 -1006 -18623
rect -1040 -18725 -1006 -18691
rect -1040 -18793 -1006 -18759
rect -22 -18317 12 -18283
rect -22 -18385 12 -18351
rect -22 -18453 12 -18419
rect -22 -18521 12 -18487
rect 2580 -18283 2614 -18249
rect 2580 -18351 2614 -18317
rect 2580 -18419 2614 -18385
rect 2580 -18487 2614 -18453
rect 3598 -18011 3632 -17977
rect 3598 -18079 3632 -18045
rect 3598 -18147 3632 -18113
rect 3598 -18215 3632 -18181
rect 3598 -18283 3632 -18249
rect 3598 -18351 3632 -18317
rect 3598 -18419 3632 -18385
rect 3598 -18487 3632 -18453
rect 4616 -18011 4650 -17977
rect 4616 -18079 4650 -18045
rect 4616 -18147 4650 -18113
rect 4616 -18215 4650 -18181
rect 4616 -18283 4650 -18249
rect 4616 -18351 4650 -18317
rect 4616 -18419 4650 -18385
rect 4616 -18487 4650 -18453
rect 5634 -18011 5668 -17977
rect 5634 -18079 5668 -18045
rect 5634 -18147 5668 -18113
rect 5634 -18215 5668 -18181
rect 5634 -18283 5668 -18249
rect 5634 -18351 5668 -18317
rect 5634 -18419 5668 -18385
rect 5634 -18487 5668 -18453
rect 6652 -18011 6686 -17977
rect 6652 -18079 6686 -18045
rect 6652 -18147 6686 -18113
rect 6652 -18215 6686 -18181
rect 6652 -18283 6686 -18249
rect 6652 -18351 6686 -18317
rect 6652 -18419 6686 -18385
rect 6652 -18487 6686 -18453
rect 7670 -18011 7704 -17977
rect 7670 -18079 7704 -18045
rect 7670 -18147 7704 -18113
rect 7670 -18215 7704 -18181
rect 7670 -18283 7704 -18249
rect 7670 -18351 7704 -18317
rect 7670 -18419 7704 -18385
rect 7670 -18487 7704 -18453
rect 8688 -18011 8722 -17977
rect 8688 -18079 8722 -18045
rect 8688 -18147 8722 -18113
rect 8688 -18215 8722 -18181
rect 8688 -18283 8722 -18249
rect 8688 -18351 8722 -18317
rect 8688 -18419 8722 -18385
rect 8688 -18487 8722 -18453
rect 9706 -18011 9740 -17977
rect 9706 -18079 9740 -18045
rect 9706 -18147 9740 -18113
rect 9706 -18215 9740 -18181
rect 9706 -18283 9740 -18249
rect 9706 -18351 9740 -18317
rect 9706 -18419 9740 -18385
rect 9706 -18487 9740 -18453
rect 10724 -18011 10758 -17977
rect 10724 -18079 10758 -18045
rect 10724 -18147 10758 -18113
rect 10724 -18215 10758 -18181
rect 10724 -18283 10758 -18249
rect 10724 -18351 10758 -18317
rect 10724 -18419 10758 -18385
rect 10724 -18487 10758 -18453
rect 11742 -18011 11776 -17977
rect 11742 -18079 11776 -18045
rect 11742 -18147 11776 -18113
rect 11742 -18215 11776 -18181
rect 11742 -18283 11776 -18249
rect 11742 -18351 11776 -18317
rect 11742 -18419 11776 -18385
rect 11742 -18487 11776 -18453
rect 12760 -18011 12794 -17977
rect 12760 -18079 12794 -18045
rect 12760 -18147 12794 -18113
rect 12760 -18215 12794 -18181
rect 12760 -18283 12794 -18249
rect 12760 -18351 12794 -18317
rect 12760 -18419 12794 -18385
rect 12760 -18487 12794 -18453
rect 13778 -18011 13812 -17977
rect 13778 -18079 13812 -18045
rect 13778 -18147 13812 -18113
rect 13778 -18215 13812 -18181
rect 13778 -18283 13812 -18249
rect 13778 -18351 13812 -18317
rect 13778 -18419 13812 -18385
rect 13778 -18487 13812 -18453
rect 14796 -18011 14830 -17977
rect 14796 -18079 14830 -18045
rect 14796 -18147 14830 -18113
rect 14796 -18215 14830 -18181
rect 14796 -18283 14830 -18249
rect 14796 -18351 14830 -18317
rect 14796 -18419 14830 -18385
rect 14796 -18487 14830 -18453
rect 15814 -18011 15848 -17977
rect 15814 -18079 15848 -18045
rect 15814 -18147 15848 -18113
rect 15814 -18215 15848 -18181
rect 15814 -18283 15848 -18249
rect 15814 -18351 15848 -18317
rect 15814 -18419 15848 -18385
rect 15814 -18487 15848 -18453
rect 16832 -18011 16866 -17977
rect 16832 -18079 16866 -18045
rect 16832 -18147 16866 -18113
rect 16832 -18215 16866 -18181
rect 16832 -18283 16866 -18249
rect 16832 -18351 16866 -18317
rect 16832 -18419 16866 -18385
rect 16832 -18487 16866 -18453
rect 17850 -18011 17884 -17977
rect 17850 -18079 17884 -18045
rect 17850 -18147 17884 -18113
rect 17850 -18215 17884 -18181
rect 17850 -18283 17884 -18249
rect 17850 -18351 17884 -18317
rect 17850 -18419 17884 -18385
rect 17850 -18487 17884 -18453
rect 18868 -18011 18902 -17977
rect 18868 -18079 18902 -18045
rect 18868 -18147 18902 -18113
rect 18868 -18215 18902 -18181
rect 18868 -18283 18902 -18249
rect 18868 -18351 18902 -18317
rect 18868 -18419 18902 -18385
rect 18868 -18487 18902 -18453
rect 19886 -18011 19920 -17977
rect 19886 -18079 19920 -18045
rect 19886 -18147 19920 -18113
rect 19886 -18215 19920 -18181
rect 19886 -18283 19920 -18249
rect 19886 -18351 19920 -18317
rect 19886 -18419 19920 -18385
rect 19886 -18487 19920 -18453
rect 20904 -18011 20938 -17977
rect 20904 -18079 20938 -18045
rect 20904 -18147 20938 -18113
rect 20904 -18215 20938 -18181
rect 20904 -18283 20938 -18249
rect 20904 -18351 20938 -18317
rect 20904 -18419 20938 -18385
rect 20904 -18487 20938 -18453
rect 21922 -18011 21956 -17977
rect 21922 -18079 21956 -18045
rect 21922 -18147 21956 -18113
rect 21922 -18215 21956 -18181
rect 21922 -18283 21956 -18249
rect 21922 -18351 21956 -18317
rect 21922 -18419 21956 -18385
rect 21922 -18487 21956 -18453
rect 22940 -18011 22974 -17977
rect 22940 -18079 22974 -18045
rect 22940 -18147 22974 -18113
rect 22940 -18215 22974 -18181
rect 22940 -18283 22974 -18249
rect 22940 -18351 22974 -18317
rect 22940 -18419 22974 -18385
rect 22940 -18487 22974 -18453
rect -22 -18589 12 -18555
rect -22 -18657 12 -18623
rect -22 -18725 12 -18691
rect -22 -18793 12 -18759
rect 2580 -19243 2614 -19209
rect 2580 -19311 2614 -19277
rect 2580 -19379 2614 -19345
rect 2580 -19447 2614 -19413
rect 2580 -19515 2614 -19481
rect 2580 -19583 2614 -19549
rect 2580 -19651 2614 -19617
rect 2580 -19719 2614 -19685
rect 3598 -19243 3632 -19209
rect 3598 -19311 3632 -19277
rect 3598 -19379 3632 -19345
rect 3598 -19447 3632 -19413
rect 3598 -19515 3632 -19481
rect 3598 -19583 3632 -19549
rect 3598 -19651 3632 -19617
rect 3598 -19719 3632 -19685
rect 4616 -19243 4650 -19209
rect 4616 -19311 4650 -19277
rect 4616 -19379 4650 -19345
rect 4616 -19447 4650 -19413
rect 4616 -19515 4650 -19481
rect 4616 -19583 4650 -19549
rect 4616 -19651 4650 -19617
rect 4616 -19719 4650 -19685
rect 5634 -19243 5668 -19209
rect 5634 -19311 5668 -19277
rect 5634 -19379 5668 -19345
rect 5634 -19447 5668 -19413
rect 5634 -19515 5668 -19481
rect 5634 -19583 5668 -19549
rect 5634 -19651 5668 -19617
rect 5634 -19719 5668 -19685
rect 6652 -19243 6686 -19209
rect 6652 -19311 6686 -19277
rect 6652 -19379 6686 -19345
rect 6652 -19447 6686 -19413
rect 6652 -19515 6686 -19481
rect 6652 -19583 6686 -19549
rect 6652 -19651 6686 -19617
rect 6652 -19719 6686 -19685
rect 7670 -19243 7704 -19209
rect 7670 -19311 7704 -19277
rect 7670 -19379 7704 -19345
rect 7670 -19447 7704 -19413
rect 7670 -19515 7704 -19481
rect 7670 -19583 7704 -19549
rect 7670 -19651 7704 -19617
rect 7670 -19719 7704 -19685
rect 8688 -19243 8722 -19209
rect 8688 -19311 8722 -19277
rect 8688 -19379 8722 -19345
rect 8688 -19447 8722 -19413
rect 8688 -19515 8722 -19481
rect 8688 -19583 8722 -19549
rect 8688 -19651 8722 -19617
rect 8688 -19719 8722 -19685
rect 9706 -19243 9740 -19209
rect 9706 -19311 9740 -19277
rect 9706 -19379 9740 -19345
rect 9706 -19447 9740 -19413
rect 9706 -19515 9740 -19481
rect 9706 -19583 9740 -19549
rect 9706 -19651 9740 -19617
rect 9706 -19719 9740 -19685
rect 10724 -19243 10758 -19209
rect 10724 -19311 10758 -19277
rect 10724 -19379 10758 -19345
rect 10724 -19447 10758 -19413
rect 10724 -19515 10758 -19481
rect 10724 -19583 10758 -19549
rect 10724 -19651 10758 -19617
rect 10724 -19719 10758 -19685
rect 11742 -19243 11776 -19209
rect 11742 -19311 11776 -19277
rect 11742 -19379 11776 -19345
rect 11742 -19447 11776 -19413
rect 11742 -19515 11776 -19481
rect 11742 -19583 11776 -19549
rect 11742 -19651 11776 -19617
rect 11742 -19719 11776 -19685
rect 12760 -19243 12794 -19209
rect 12760 -19311 12794 -19277
rect 12760 -19379 12794 -19345
rect 12760 -19447 12794 -19413
rect 12760 -19515 12794 -19481
rect 12760 -19583 12794 -19549
rect 12760 -19651 12794 -19617
rect 12760 -19719 12794 -19685
rect 13778 -19243 13812 -19209
rect 13778 -19311 13812 -19277
rect 13778 -19379 13812 -19345
rect 13778 -19447 13812 -19413
rect 13778 -19515 13812 -19481
rect 13778 -19583 13812 -19549
rect 13778 -19651 13812 -19617
rect 13778 -19719 13812 -19685
rect 14796 -19243 14830 -19209
rect 14796 -19311 14830 -19277
rect 14796 -19379 14830 -19345
rect 14796 -19447 14830 -19413
rect 14796 -19515 14830 -19481
rect 14796 -19583 14830 -19549
rect 14796 -19651 14830 -19617
rect 14796 -19719 14830 -19685
rect 15814 -19243 15848 -19209
rect 15814 -19311 15848 -19277
rect 15814 -19379 15848 -19345
rect 15814 -19447 15848 -19413
rect 15814 -19515 15848 -19481
rect 15814 -19583 15848 -19549
rect 15814 -19651 15848 -19617
rect 15814 -19719 15848 -19685
rect 16832 -19243 16866 -19209
rect 16832 -19311 16866 -19277
rect 16832 -19379 16866 -19345
rect 16832 -19447 16866 -19413
rect 16832 -19515 16866 -19481
rect 16832 -19583 16866 -19549
rect 16832 -19651 16866 -19617
rect 16832 -19719 16866 -19685
rect 17850 -19243 17884 -19209
rect 17850 -19311 17884 -19277
rect 17850 -19379 17884 -19345
rect 17850 -19447 17884 -19413
rect 17850 -19515 17884 -19481
rect 17850 -19583 17884 -19549
rect 17850 -19651 17884 -19617
rect 17850 -19719 17884 -19685
rect 18868 -19243 18902 -19209
rect 18868 -19311 18902 -19277
rect 18868 -19379 18902 -19345
rect 18868 -19447 18902 -19413
rect 18868 -19515 18902 -19481
rect 18868 -19583 18902 -19549
rect 18868 -19651 18902 -19617
rect 18868 -19719 18902 -19685
rect 19886 -19243 19920 -19209
rect 19886 -19311 19920 -19277
rect 19886 -19379 19920 -19345
rect 19886 -19447 19920 -19413
rect 19886 -19515 19920 -19481
rect 19886 -19583 19920 -19549
rect 19886 -19651 19920 -19617
rect 19886 -19719 19920 -19685
rect 20904 -19243 20938 -19209
rect 20904 -19311 20938 -19277
rect 20904 -19379 20938 -19345
rect 20904 -19447 20938 -19413
rect 20904 -19515 20938 -19481
rect 20904 -19583 20938 -19549
rect 20904 -19651 20938 -19617
rect 20904 -19719 20938 -19685
rect 21922 -19243 21956 -19209
rect 21922 -19311 21956 -19277
rect 21922 -19379 21956 -19345
rect 21922 -19447 21956 -19413
rect 21922 -19515 21956 -19481
rect 21922 -19583 21956 -19549
rect 21922 -19651 21956 -19617
rect 21922 -19719 21956 -19685
rect 22940 -19243 22974 -19209
rect 22940 -19311 22974 -19277
rect 22940 -19379 22974 -19345
rect 22940 -19447 22974 -19413
rect 22940 -19515 22974 -19481
rect 22940 -19583 22974 -19549
rect 22940 -19651 22974 -19617
rect 22940 -19719 22974 -19685
rect 2580 -20477 2614 -20443
rect 2580 -20545 2614 -20511
rect 2580 -20613 2614 -20579
rect 2580 -20681 2614 -20647
rect 2580 -20749 2614 -20715
rect 2580 -20817 2614 -20783
rect 2580 -20885 2614 -20851
rect 2580 -20953 2614 -20919
rect 3598 -20477 3632 -20443
rect 3598 -20545 3632 -20511
rect 3598 -20613 3632 -20579
rect 3598 -20681 3632 -20647
rect 3598 -20749 3632 -20715
rect 3598 -20817 3632 -20783
rect 3598 -20885 3632 -20851
rect 3598 -20953 3632 -20919
rect 4616 -20477 4650 -20443
rect 4616 -20545 4650 -20511
rect 4616 -20613 4650 -20579
rect 4616 -20681 4650 -20647
rect 4616 -20749 4650 -20715
rect 4616 -20817 4650 -20783
rect 4616 -20885 4650 -20851
rect 4616 -20953 4650 -20919
rect 5634 -20477 5668 -20443
rect 5634 -20545 5668 -20511
rect 5634 -20613 5668 -20579
rect 5634 -20681 5668 -20647
rect 5634 -20749 5668 -20715
rect 5634 -20817 5668 -20783
rect 5634 -20885 5668 -20851
rect 5634 -20953 5668 -20919
rect 6652 -20477 6686 -20443
rect 6652 -20545 6686 -20511
rect 6652 -20613 6686 -20579
rect 6652 -20681 6686 -20647
rect 6652 -20749 6686 -20715
rect 6652 -20817 6686 -20783
rect 6652 -20885 6686 -20851
rect 6652 -20953 6686 -20919
rect 7670 -20477 7704 -20443
rect 7670 -20545 7704 -20511
rect 7670 -20613 7704 -20579
rect 7670 -20681 7704 -20647
rect 7670 -20749 7704 -20715
rect 7670 -20817 7704 -20783
rect 7670 -20885 7704 -20851
rect 7670 -20953 7704 -20919
rect 8688 -20477 8722 -20443
rect 8688 -20545 8722 -20511
rect 8688 -20613 8722 -20579
rect 8688 -20681 8722 -20647
rect 8688 -20749 8722 -20715
rect 8688 -20817 8722 -20783
rect 8688 -20885 8722 -20851
rect 8688 -20953 8722 -20919
rect 9706 -20477 9740 -20443
rect 9706 -20545 9740 -20511
rect 9706 -20613 9740 -20579
rect 9706 -20681 9740 -20647
rect 9706 -20749 9740 -20715
rect 9706 -20817 9740 -20783
rect 9706 -20885 9740 -20851
rect 9706 -20953 9740 -20919
rect 10724 -20477 10758 -20443
rect 10724 -20545 10758 -20511
rect 10724 -20613 10758 -20579
rect 10724 -20681 10758 -20647
rect 10724 -20749 10758 -20715
rect 10724 -20817 10758 -20783
rect 10724 -20885 10758 -20851
rect 10724 -20953 10758 -20919
rect 11742 -20477 11776 -20443
rect 11742 -20545 11776 -20511
rect 11742 -20613 11776 -20579
rect 11742 -20681 11776 -20647
rect 11742 -20749 11776 -20715
rect 11742 -20817 11776 -20783
rect 11742 -20885 11776 -20851
rect 11742 -20953 11776 -20919
rect 12760 -20477 12794 -20443
rect 12760 -20545 12794 -20511
rect 12760 -20613 12794 -20579
rect 12760 -20681 12794 -20647
rect 12760 -20749 12794 -20715
rect 12760 -20817 12794 -20783
rect 12760 -20885 12794 -20851
rect 12760 -20953 12794 -20919
rect 13778 -20477 13812 -20443
rect 13778 -20545 13812 -20511
rect 13778 -20613 13812 -20579
rect 13778 -20681 13812 -20647
rect 13778 -20749 13812 -20715
rect 13778 -20817 13812 -20783
rect 13778 -20885 13812 -20851
rect 13778 -20953 13812 -20919
rect 14796 -20477 14830 -20443
rect 14796 -20545 14830 -20511
rect 14796 -20613 14830 -20579
rect 14796 -20681 14830 -20647
rect 14796 -20749 14830 -20715
rect 14796 -20817 14830 -20783
rect 14796 -20885 14830 -20851
rect 14796 -20953 14830 -20919
rect 15814 -20477 15848 -20443
rect 15814 -20545 15848 -20511
rect 15814 -20613 15848 -20579
rect 15814 -20681 15848 -20647
rect 15814 -20749 15848 -20715
rect 15814 -20817 15848 -20783
rect 15814 -20885 15848 -20851
rect 15814 -20953 15848 -20919
rect 16832 -20477 16866 -20443
rect 16832 -20545 16866 -20511
rect 16832 -20613 16866 -20579
rect 16832 -20681 16866 -20647
rect 16832 -20749 16866 -20715
rect 16832 -20817 16866 -20783
rect 16832 -20885 16866 -20851
rect 16832 -20953 16866 -20919
rect 17850 -20477 17884 -20443
rect 17850 -20545 17884 -20511
rect 17850 -20613 17884 -20579
rect 17850 -20681 17884 -20647
rect 17850 -20749 17884 -20715
rect 17850 -20817 17884 -20783
rect 17850 -20885 17884 -20851
rect 17850 -20953 17884 -20919
rect 18868 -20477 18902 -20443
rect 18868 -20545 18902 -20511
rect 18868 -20613 18902 -20579
rect 18868 -20681 18902 -20647
rect 18868 -20749 18902 -20715
rect 18868 -20817 18902 -20783
rect 18868 -20885 18902 -20851
rect 18868 -20953 18902 -20919
rect 19886 -20477 19920 -20443
rect 19886 -20545 19920 -20511
rect 19886 -20613 19920 -20579
rect 19886 -20681 19920 -20647
rect 19886 -20749 19920 -20715
rect 19886 -20817 19920 -20783
rect 19886 -20885 19920 -20851
rect 19886 -20953 19920 -20919
rect 20904 -20477 20938 -20443
rect 20904 -20545 20938 -20511
rect 20904 -20613 20938 -20579
rect 20904 -20681 20938 -20647
rect 20904 -20749 20938 -20715
rect 20904 -20817 20938 -20783
rect 20904 -20885 20938 -20851
rect 20904 -20953 20938 -20919
rect 21922 -20477 21956 -20443
rect 21922 -20545 21956 -20511
rect 21922 -20613 21956 -20579
rect 21922 -20681 21956 -20647
rect 21922 -20749 21956 -20715
rect 21922 -20817 21956 -20783
rect 21922 -20885 21956 -20851
rect 21922 -20953 21956 -20919
rect 22940 -20477 22974 -20443
rect 22940 -20545 22974 -20511
rect 22940 -20613 22974 -20579
rect 22940 -20681 22974 -20647
rect 22940 -20749 22974 -20715
rect 22940 -20817 22974 -20783
rect 22940 -20885 22974 -20851
rect 22940 -20953 22974 -20919
rect 2580 -21711 2614 -21677
rect 2580 -21779 2614 -21745
rect 2580 -21847 2614 -21813
rect 2580 -21915 2614 -21881
rect 2580 -21983 2614 -21949
rect 2580 -22051 2614 -22017
rect 2580 -22119 2614 -22085
rect 2580 -22187 2614 -22153
rect 3598 -21711 3632 -21677
rect 3598 -21779 3632 -21745
rect 3598 -21847 3632 -21813
rect 3598 -21915 3632 -21881
rect 3598 -21983 3632 -21949
rect 3598 -22051 3632 -22017
rect 3598 -22119 3632 -22085
rect 3598 -22187 3632 -22153
rect 4616 -21711 4650 -21677
rect 4616 -21779 4650 -21745
rect 4616 -21847 4650 -21813
rect 4616 -21915 4650 -21881
rect 4616 -21983 4650 -21949
rect 4616 -22051 4650 -22017
rect 4616 -22119 4650 -22085
rect 4616 -22187 4650 -22153
rect 5634 -21711 5668 -21677
rect 5634 -21779 5668 -21745
rect 5634 -21847 5668 -21813
rect 5634 -21915 5668 -21881
rect 5634 -21983 5668 -21949
rect 5634 -22051 5668 -22017
rect 5634 -22119 5668 -22085
rect 5634 -22187 5668 -22153
rect 6652 -21711 6686 -21677
rect 6652 -21779 6686 -21745
rect 6652 -21847 6686 -21813
rect 6652 -21915 6686 -21881
rect 6652 -21983 6686 -21949
rect 6652 -22051 6686 -22017
rect 6652 -22119 6686 -22085
rect 6652 -22187 6686 -22153
rect 7670 -21711 7704 -21677
rect 7670 -21779 7704 -21745
rect 7670 -21847 7704 -21813
rect 7670 -21915 7704 -21881
rect 7670 -21983 7704 -21949
rect 7670 -22051 7704 -22017
rect 7670 -22119 7704 -22085
rect 7670 -22187 7704 -22153
rect 8688 -21711 8722 -21677
rect 8688 -21779 8722 -21745
rect 8688 -21847 8722 -21813
rect 8688 -21915 8722 -21881
rect 8688 -21983 8722 -21949
rect 8688 -22051 8722 -22017
rect 8688 -22119 8722 -22085
rect 8688 -22187 8722 -22153
rect 9706 -21711 9740 -21677
rect 9706 -21779 9740 -21745
rect 9706 -21847 9740 -21813
rect 9706 -21915 9740 -21881
rect 9706 -21983 9740 -21949
rect 9706 -22051 9740 -22017
rect 9706 -22119 9740 -22085
rect 9706 -22187 9740 -22153
rect 10724 -21711 10758 -21677
rect 10724 -21779 10758 -21745
rect 10724 -21847 10758 -21813
rect 10724 -21915 10758 -21881
rect 10724 -21983 10758 -21949
rect 10724 -22051 10758 -22017
rect 10724 -22119 10758 -22085
rect 10724 -22187 10758 -22153
rect 11742 -21711 11776 -21677
rect 11742 -21779 11776 -21745
rect 11742 -21847 11776 -21813
rect 11742 -21915 11776 -21881
rect 11742 -21983 11776 -21949
rect 11742 -22051 11776 -22017
rect 11742 -22119 11776 -22085
rect 11742 -22187 11776 -22153
rect 12760 -21711 12794 -21677
rect 12760 -21779 12794 -21745
rect 12760 -21847 12794 -21813
rect 12760 -21915 12794 -21881
rect 12760 -21983 12794 -21949
rect 12760 -22051 12794 -22017
rect 12760 -22119 12794 -22085
rect 12760 -22187 12794 -22153
rect 13778 -21711 13812 -21677
rect 13778 -21779 13812 -21745
rect 13778 -21847 13812 -21813
rect 13778 -21915 13812 -21881
rect 13778 -21983 13812 -21949
rect 13778 -22051 13812 -22017
rect 13778 -22119 13812 -22085
rect 13778 -22187 13812 -22153
rect 14796 -21711 14830 -21677
rect 14796 -21779 14830 -21745
rect 14796 -21847 14830 -21813
rect 14796 -21915 14830 -21881
rect 14796 -21983 14830 -21949
rect 14796 -22051 14830 -22017
rect 14796 -22119 14830 -22085
rect 14796 -22187 14830 -22153
rect 15814 -21711 15848 -21677
rect 15814 -21779 15848 -21745
rect 15814 -21847 15848 -21813
rect 15814 -21915 15848 -21881
rect 15814 -21983 15848 -21949
rect 15814 -22051 15848 -22017
rect 15814 -22119 15848 -22085
rect 15814 -22187 15848 -22153
rect 16832 -21711 16866 -21677
rect 16832 -21779 16866 -21745
rect 16832 -21847 16866 -21813
rect 16832 -21915 16866 -21881
rect 16832 -21983 16866 -21949
rect 16832 -22051 16866 -22017
rect 16832 -22119 16866 -22085
rect 16832 -22187 16866 -22153
rect 17850 -21711 17884 -21677
rect 17850 -21779 17884 -21745
rect 17850 -21847 17884 -21813
rect 17850 -21915 17884 -21881
rect 17850 -21983 17884 -21949
rect 17850 -22051 17884 -22017
rect 17850 -22119 17884 -22085
rect 17850 -22187 17884 -22153
rect 18868 -21711 18902 -21677
rect 18868 -21779 18902 -21745
rect 18868 -21847 18902 -21813
rect 18868 -21915 18902 -21881
rect 18868 -21983 18902 -21949
rect 18868 -22051 18902 -22017
rect 18868 -22119 18902 -22085
rect 18868 -22187 18902 -22153
rect 19886 -21711 19920 -21677
rect 19886 -21779 19920 -21745
rect 19886 -21847 19920 -21813
rect 19886 -21915 19920 -21881
rect 19886 -21983 19920 -21949
rect 19886 -22051 19920 -22017
rect 19886 -22119 19920 -22085
rect 19886 -22187 19920 -22153
rect 20904 -21711 20938 -21677
rect 20904 -21779 20938 -21745
rect 20904 -21847 20938 -21813
rect 20904 -21915 20938 -21881
rect 20904 -21983 20938 -21949
rect 20904 -22051 20938 -22017
rect 20904 -22119 20938 -22085
rect 20904 -22187 20938 -22153
rect 21922 -21711 21956 -21677
rect 21922 -21779 21956 -21745
rect 21922 -21847 21956 -21813
rect 21922 -21915 21956 -21881
rect 21922 -21983 21956 -21949
rect 21922 -22051 21956 -22017
rect 21922 -22119 21956 -22085
rect 21922 -22187 21956 -22153
rect 22940 -21711 22974 -21677
rect 22940 -21779 22974 -21745
rect 22940 -21847 22974 -21813
rect 22940 -21915 22974 -21881
rect 22940 -21983 22974 -21949
rect 22940 -22051 22974 -22017
rect 22940 -22119 22974 -22085
rect 22940 -22187 22974 -22153
rect 2580 -22943 2614 -22909
rect 2580 -23011 2614 -22977
rect 2580 -23079 2614 -23045
rect 2580 -23147 2614 -23113
rect 2580 -23215 2614 -23181
rect 2580 -23283 2614 -23249
rect 2580 -23351 2614 -23317
rect 2580 -23419 2614 -23385
rect 3598 -22943 3632 -22909
rect 3598 -23011 3632 -22977
rect 3598 -23079 3632 -23045
rect 3598 -23147 3632 -23113
rect 3598 -23215 3632 -23181
rect 3598 -23283 3632 -23249
rect 3598 -23351 3632 -23317
rect 3598 -23419 3632 -23385
rect 4616 -22943 4650 -22909
rect 4616 -23011 4650 -22977
rect 4616 -23079 4650 -23045
rect 4616 -23147 4650 -23113
rect 4616 -23215 4650 -23181
rect 4616 -23283 4650 -23249
rect 4616 -23351 4650 -23317
rect 4616 -23419 4650 -23385
rect 5634 -22943 5668 -22909
rect 5634 -23011 5668 -22977
rect 5634 -23079 5668 -23045
rect 5634 -23147 5668 -23113
rect 5634 -23215 5668 -23181
rect 5634 -23283 5668 -23249
rect 5634 -23351 5668 -23317
rect 5634 -23419 5668 -23385
rect 6652 -22943 6686 -22909
rect 6652 -23011 6686 -22977
rect 6652 -23079 6686 -23045
rect 6652 -23147 6686 -23113
rect 6652 -23215 6686 -23181
rect 6652 -23283 6686 -23249
rect 6652 -23351 6686 -23317
rect 6652 -23419 6686 -23385
rect 7670 -22943 7704 -22909
rect 7670 -23011 7704 -22977
rect 7670 -23079 7704 -23045
rect 7670 -23147 7704 -23113
rect 7670 -23215 7704 -23181
rect 7670 -23283 7704 -23249
rect 7670 -23351 7704 -23317
rect 7670 -23419 7704 -23385
rect 8688 -22943 8722 -22909
rect 8688 -23011 8722 -22977
rect 8688 -23079 8722 -23045
rect 8688 -23147 8722 -23113
rect 8688 -23215 8722 -23181
rect 8688 -23283 8722 -23249
rect 8688 -23351 8722 -23317
rect 8688 -23419 8722 -23385
rect 9706 -22943 9740 -22909
rect 9706 -23011 9740 -22977
rect 9706 -23079 9740 -23045
rect 9706 -23147 9740 -23113
rect 9706 -23215 9740 -23181
rect 9706 -23283 9740 -23249
rect 9706 -23351 9740 -23317
rect 9706 -23419 9740 -23385
rect 10724 -22943 10758 -22909
rect 10724 -23011 10758 -22977
rect 10724 -23079 10758 -23045
rect 10724 -23147 10758 -23113
rect 10724 -23215 10758 -23181
rect 10724 -23283 10758 -23249
rect 10724 -23351 10758 -23317
rect 10724 -23419 10758 -23385
rect 11742 -22943 11776 -22909
rect 11742 -23011 11776 -22977
rect 11742 -23079 11776 -23045
rect 11742 -23147 11776 -23113
rect 11742 -23215 11776 -23181
rect 11742 -23283 11776 -23249
rect 11742 -23351 11776 -23317
rect 11742 -23419 11776 -23385
rect 12760 -22943 12794 -22909
rect 12760 -23011 12794 -22977
rect 12760 -23079 12794 -23045
rect 12760 -23147 12794 -23113
rect 12760 -23215 12794 -23181
rect 12760 -23283 12794 -23249
rect 12760 -23351 12794 -23317
rect 12760 -23419 12794 -23385
rect 13778 -22943 13812 -22909
rect 13778 -23011 13812 -22977
rect 13778 -23079 13812 -23045
rect 13778 -23147 13812 -23113
rect 13778 -23215 13812 -23181
rect 13778 -23283 13812 -23249
rect 13778 -23351 13812 -23317
rect 13778 -23419 13812 -23385
rect 14796 -22943 14830 -22909
rect 14796 -23011 14830 -22977
rect 14796 -23079 14830 -23045
rect 14796 -23147 14830 -23113
rect 14796 -23215 14830 -23181
rect 14796 -23283 14830 -23249
rect 14796 -23351 14830 -23317
rect 14796 -23419 14830 -23385
rect 15814 -22943 15848 -22909
rect 15814 -23011 15848 -22977
rect 15814 -23079 15848 -23045
rect 15814 -23147 15848 -23113
rect 15814 -23215 15848 -23181
rect 15814 -23283 15848 -23249
rect 15814 -23351 15848 -23317
rect 15814 -23419 15848 -23385
rect 16832 -22943 16866 -22909
rect 16832 -23011 16866 -22977
rect 16832 -23079 16866 -23045
rect 16832 -23147 16866 -23113
rect 16832 -23215 16866 -23181
rect 16832 -23283 16866 -23249
rect 16832 -23351 16866 -23317
rect 16832 -23419 16866 -23385
rect 17850 -22943 17884 -22909
rect 17850 -23011 17884 -22977
rect 17850 -23079 17884 -23045
rect 17850 -23147 17884 -23113
rect 17850 -23215 17884 -23181
rect 17850 -23283 17884 -23249
rect 17850 -23351 17884 -23317
rect 17850 -23419 17884 -23385
rect 18868 -22943 18902 -22909
rect 18868 -23011 18902 -22977
rect 18868 -23079 18902 -23045
rect 18868 -23147 18902 -23113
rect 18868 -23215 18902 -23181
rect 18868 -23283 18902 -23249
rect 18868 -23351 18902 -23317
rect 18868 -23419 18902 -23385
rect 19886 -22943 19920 -22909
rect 19886 -23011 19920 -22977
rect 19886 -23079 19920 -23045
rect 19886 -23147 19920 -23113
rect 19886 -23215 19920 -23181
rect 19886 -23283 19920 -23249
rect 19886 -23351 19920 -23317
rect 19886 -23419 19920 -23385
rect 20904 -22943 20938 -22909
rect 20904 -23011 20938 -22977
rect 20904 -23079 20938 -23045
rect 20904 -23147 20938 -23113
rect 20904 -23215 20938 -23181
rect 20904 -23283 20938 -23249
rect 20904 -23351 20938 -23317
rect 20904 -23419 20938 -23385
rect 21922 -22943 21956 -22909
rect 21922 -23011 21956 -22977
rect 21922 -23079 21956 -23045
rect 21922 -23147 21956 -23113
rect 21922 -23215 21956 -23181
rect 21922 -23283 21956 -23249
rect 21922 -23351 21956 -23317
rect 21922 -23419 21956 -23385
rect 22940 -22943 22974 -22909
rect 22940 -23011 22974 -22977
rect 22940 -23079 22974 -23045
rect 22940 -23147 22974 -23113
rect 22940 -23215 22974 -23181
rect 22940 -23283 22974 -23249
rect 22940 -23351 22974 -23317
rect 22940 -23419 22974 -23385
rect 2580 -24177 2614 -24143
rect 2580 -24245 2614 -24211
rect 2580 -24313 2614 -24279
rect 2580 -24381 2614 -24347
rect 2580 -24449 2614 -24415
rect 2580 -24517 2614 -24483
rect 2580 -24585 2614 -24551
rect 2580 -24653 2614 -24619
rect 3598 -24177 3632 -24143
rect 3598 -24245 3632 -24211
rect 3598 -24313 3632 -24279
rect 3598 -24381 3632 -24347
rect 3598 -24449 3632 -24415
rect 3598 -24517 3632 -24483
rect 3598 -24585 3632 -24551
rect 3598 -24653 3632 -24619
rect 4616 -24177 4650 -24143
rect 4616 -24245 4650 -24211
rect 4616 -24313 4650 -24279
rect 4616 -24381 4650 -24347
rect 4616 -24449 4650 -24415
rect 4616 -24517 4650 -24483
rect 4616 -24585 4650 -24551
rect 4616 -24653 4650 -24619
rect 5634 -24177 5668 -24143
rect 5634 -24245 5668 -24211
rect 5634 -24313 5668 -24279
rect 5634 -24381 5668 -24347
rect 5634 -24449 5668 -24415
rect 5634 -24517 5668 -24483
rect 5634 -24585 5668 -24551
rect 5634 -24653 5668 -24619
rect 6652 -24177 6686 -24143
rect 6652 -24245 6686 -24211
rect 6652 -24313 6686 -24279
rect 6652 -24381 6686 -24347
rect 6652 -24449 6686 -24415
rect 6652 -24517 6686 -24483
rect 6652 -24585 6686 -24551
rect 6652 -24653 6686 -24619
rect 7670 -24177 7704 -24143
rect 7670 -24245 7704 -24211
rect 7670 -24313 7704 -24279
rect 7670 -24381 7704 -24347
rect 7670 -24449 7704 -24415
rect 7670 -24517 7704 -24483
rect 7670 -24585 7704 -24551
rect 7670 -24653 7704 -24619
rect 8688 -24177 8722 -24143
rect 8688 -24245 8722 -24211
rect 8688 -24313 8722 -24279
rect 8688 -24381 8722 -24347
rect 8688 -24449 8722 -24415
rect 8688 -24517 8722 -24483
rect 8688 -24585 8722 -24551
rect 8688 -24653 8722 -24619
rect 9706 -24177 9740 -24143
rect 9706 -24245 9740 -24211
rect 9706 -24313 9740 -24279
rect 9706 -24381 9740 -24347
rect 9706 -24449 9740 -24415
rect 9706 -24517 9740 -24483
rect 9706 -24585 9740 -24551
rect 9706 -24653 9740 -24619
rect 10724 -24177 10758 -24143
rect 10724 -24245 10758 -24211
rect 10724 -24313 10758 -24279
rect 10724 -24381 10758 -24347
rect 10724 -24449 10758 -24415
rect 10724 -24517 10758 -24483
rect 10724 -24585 10758 -24551
rect 10724 -24653 10758 -24619
rect 11742 -24177 11776 -24143
rect 11742 -24245 11776 -24211
rect 11742 -24313 11776 -24279
rect 11742 -24381 11776 -24347
rect 11742 -24449 11776 -24415
rect 11742 -24517 11776 -24483
rect 11742 -24585 11776 -24551
rect 11742 -24653 11776 -24619
rect 12760 -24177 12794 -24143
rect 12760 -24245 12794 -24211
rect 12760 -24313 12794 -24279
rect 12760 -24381 12794 -24347
rect 12760 -24449 12794 -24415
rect 12760 -24517 12794 -24483
rect 12760 -24585 12794 -24551
rect 12760 -24653 12794 -24619
rect 13778 -24177 13812 -24143
rect 13778 -24245 13812 -24211
rect 13778 -24313 13812 -24279
rect 13778 -24381 13812 -24347
rect 13778 -24449 13812 -24415
rect 13778 -24517 13812 -24483
rect 13778 -24585 13812 -24551
rect 13778 -24653 13812 -24619
rect 14796 -24177 14830 -24143
rect 14796 -24245 14830 -24211
rect 14796 -24313 14830 -24279
rect 14796 -24381 14830 -24347
rect 14796 -24449 14830 -24415
rect 14796 -24517 14830 -24483
rect 14796 -24585 14830 -24551
rect 14796 -24653 14830 -24619
rect 15814 -24177 15848 -24143
rect 15814 -24245 15848 -24211
rect 15814 -24313 15848 -24279
rect 15814 -24381 15848 -24347
rect 15814 -24449 15848 -24415
rect 15814 -24517 15848 -24483
rect 15814 -24585 15848 -24551
rect 15814 -24653 15848 -24619
rect 16832 -24177 16866 -24143
rect 16832 -24245 16866 -24211
rect 16832 -24313 16866 -24279
rect 16832 -24381 16866 -24347
rect 16832 -24449 16866 -24415
rect 16832 -24517 16866 -24483
rect 16832 -24585 16866 -24551
rect 16832 -24653 16866 -24619
rect 17850 -24177 17884 -24143
rect 17850 -24245 17884 -24211
rect 17850 -24313 17884 -24279
rect 17850 -24381 17884 -24347
rect 17850 -24449 17884 -24415
rect 17850 -24517 17884 -24483
rect 17850 -24585 17884 -24551
rect 17850 -24653 17884 -24619
rect 18868 -24177 18902 -24143
rect 18868 -24245 18902 -24211
rect 18868 -24313 18902 -24279
rect 18868 -24381 18902 -24347
rect 18868 -24449 18902 -24415
rect 18868 -24517 18902 -24483
rect 18868 -24585 18902 -24551
rect 18868 -24653 18902 -24619
rect 19886 -24177 19920 -24143
rect 19886 -24245 19920 -24211
rect 19886 -24313 19920 -24279
rect 19886 -24381 19920 -24347
rect 19886 -24449 19920 -24415
rect 19886 -24517 19920 -24483
rect 19886 -24585 19920 -24551
rect 19886 -24653 19920 -24619
rect 20904 -24177 20938 -24143
rect 20904 -24245 20938 -24211
rect 20904 -24313 20938 -24279
rect 20904 -24381 20938 -24347
rect 20904 -24449 20938 -24415
rect 20904 -24517 20938 -24483
rect 20904 -24585 20938 -24551
rect 20904 -24653 20938 -24619
rect 21922 -24177 21956 -24143
rect 21922 -24245 21956 -24211
rect 21922 -24313 21956 -24279
rect 21922 -24381 21956 -24347
rect 21922 -24449 21956 -24415
rect 21922 -24517 21956 -24483
rect 21922 -24585 21956 -24551
rect 21922 -24653 21956 -24619
rect 22940 -24177 22974 -24143
rect 22940 -24245 22974 -24211
rect 22940 -24313 22974 -24279
rect 22940 -24381 22974 -24347
rect 22940 -24449 22974 -24415
rect 22940 -24517 22974 -24483
rect 22940 -24585 22974 -24551
rect 22940 -24653 22974 -24619
<< psubdiff >>
rect -12322 -11211 24922 -11178
rect -12322 -11245 -12145 -11211
rect -12111 -11245 -12077 -11211
rect -12043 -11245 -12009 -11211
rect -11975 -11245 -11941 -11211
rect -11907 -11245 -11873 -11211
rect -11839 -11245 -11805 -11211
rect -11771 -11245 -11737 -11211
rect -11703 -11245 -11669 -11211
rect -11635 -11245 -11601 -11211
rect -11567 -11245 -11533 -11211
rect -11499 -11245 -11465 -11211
rect -11431 -11245 -11397 -11211
rect -11363 -11245 -11329 -11211
rect -11295 -11245 -11261 -11211
rect -11227 -11245 -11193 -11211
rect -11159 -11245 -11125 -11211
rect -11091 -11245 -11057 -11211
rect -11023 -11245 -10989 -11211
rect -10955 -11245 -10921 -11211
rect -10887 -11245 -10853 -11211
rect -10819 -11245 -10785 -11211
rect -10751 -11245 -10717 -11211
rect -10683 -11245 -10649 -11211
rect -10615 -11245 -10581 -11211
rect -10547 -11245 -10513 -11211
rect -10479 -11245 -10445 -11211
rect -10411 -11245 -10377 -11211
rect -10343 -11245 -10309 -11211
rect -10275 -11245 -10241 -11211
rect -10207 -11245 -10173 -11211
rect -10139 -11245 -10105 -11211
rect -10071 -11245 -10037 -11211
rect -10003 -11245 -9969 -11211
rect -9935 -11245 -9901 -11211
rect -9867 -11245 -9833 -11211
rect -9799 -11245 -9765 -11211
rect -9731 -11245 -9697 -11211
rect -9663 -11245 -9629 -11211
rect -9595 -11245 -9561 -11211
rect -9527 -11245 -9493 -11211
rect -9459 -11245 -9425 -11211
rect -9391 -11245 -9357 -11211
rect -9323 -11245 -9289 -11211
rect -9255 -11245 -9221 -11211
rect -9187 -11245 -9153 -11211
rect -9119 -11245 -9085 -11211
rect -9051 -11245 -9017 -11211
rect -8983 -11245 -8949 -11211
rect -8915 -11245 -8881 -11211
rect -8847 -11245 -8813 -11211
rect -8779 -11245 -8745 -11211
rect -8711 -11245 -8677 -11211
rect -8643 -11245 -8609 -11211
rect -8575 -11245 -8541 -11211
rect -8507 -11245 -8473 -11211
rect -8439 -11245 -8405 -11211
rect -8371 -11245 -8337 -11211
rect -8303 -11245 -8269 -11211
rect -8235 -11245 -8201 -11211
rect -8167 -11245 -8133 -11211
rect -8099 -11245 -8065 -11211
rect -8031 -11245 -7997 -11211
rect -7963 -11245 -7929 -11211
rect -7895 -11245 -7861 -11211
rect -7827 -11245 -7793 -11211
rect -7759 -11245 -7725 -11211
rect -7691 -11245 -7657 -11211
rect -7623 -11245 -7589 -11211
rect -7555 -11245 -7521 -11211
rect -7487 -11245 -7453 -11211
rect -7419 -11245 -7385 -11211
rect -7351 -11245 -7317 -11211
rect -7283 -11245 -7249 -11211
rect -7215 -11245 -7181 -11211
rect -7147 -11245 -7113 -11211
rect -7079 -11245 -7045 -11211
rect -7011 -11245 -6977 -11211
rect -6943 -11245 -6909 -11211
rect -6875 -11245 -6841 -11211
rect -6807 -11245 -6773 -11211
rect -6739 -11245 -6705 -11211
rect -6671 -11245 -6637 -11211
rect -6603 -11245 -6569 -11211
rect -6535 -11245 -6501 -11211
rect -6467 -11245 -6433 -11211
rect -6399 -11245 -6365 -11211
rect -6331 -11245 -6297 -11211
rect -6263 -11245 -6229 -11211
rect -6195 -11245 -6161 -11211
rect -6127 -11245 -6093 -11211
rect -6059 -11245 -6025 -11211
rect -5991 -11245 -5957 -11211
rect -5923 -11245 -5889 -11211
rect -5855 -11245 -5821 -11211
rect -5787 -11245 -5753 -11211
rect -5719 -11245 -5685 -11211
rect -5651 -11245 -5617 -11211
rect -5583 -11245 -5549 -11211
rect -5515 -11245 -5481 -11211
rect -5447 -11245 -5413 -11211
rect -5379 -11245 -5345 -11211
rect -5311 -11245 -5277 -11211
rect -5243 -11245 -5209 -11211
rect -5175 -11245 -5141 -11211
rect -5107 -11245 -5073 -11211
rect -5039 -11245 -5005 -11211
rect -4971 -11245 -4937 -11211
rect -4903 -11245 -4869 -11211
rect -4835 -11245 -4801 -11211
rect -4767 -11245 -4733 -11211
rect -4699 -11245 -4665 -11211
rect -4631 -11245 -4597 -11211
rect -4563 -11245 -4529 -11211
rect -4495 -11245 -4461 -11211
rect -4427 -11245 -4393 -11211
rect -4359 -11245 -4325 -11211
rect -4291 -11245 -4257 -11211
rect -4223 -11245 -4189 -11211
rect -4155 -11245 -4121 -11211
rect -4087 -11245 -4053 -11211
rect -4019 -11245 -3985 -11211
rect -3951 -11245 -3917 -11211
rect -3883 -11245 -3849 -11211
rect -3815 -11245 -3781 -11211
rect -3747 -11245 -3713 -11211
rect -3679 -11245 -3645 -11211
rect -3611 -11245 -3577 -11211
rect -3543 -11245 -3509 -11211
rect -3475 -11245 -3441 -11211
rect -3407 -11245 -3373 -11211
rect -3339 -11245 -3305 -11211
rect -3271 -11245 -3237 -11211
rect -3203 -11245 -3169 -11211
rect -3135 -11245 -3101 -11211
rect -3067 -11245 -3033 -11211
rect -2999 -11245 -2965 -11211
rect -2931 -11245 -2897 -11211
rect -2863 -11245 -2829 -11211
rect -2795 -11245 -2761 -11211
rect -2727 -11245 -2693 -11211
rect -2659 -11245 -2625 -11211
rect -2591 -11245 -2557 -11211
rect -2523 -11245 -2489 -11211
rect -2455 -11245 -2421 -11211
rect -2387 -11245 -2353 -11211
rect -2319 -11245 -2285 -11211
rect -2251 -11245 -2217 -11211
rect -2183 -11245 -2149 -11211
rect -2115 -11245 -2081 -11211
rect -2047 -11245 -2013 -11211
rect -1979 -11245 -1945 -11211
rect -1911 -11245 -1877 -11211
rect -1843 -11245 -1809 -11211
rect -1775 -11245 -1741 -11211
rect -1707 -11245 -1673 -11211
rect -1639 -11245 -1605 -11211
rect -1571 -11245 -1537 -11211
rect -1503 -11245 -1469 -11211
rect -1435 -11245 -1401 -11211
rect -1367 -11245 -1333 -11211
rect -1299 -11245 -1265 -11211
rect -1231 -11245 -1197 -11211
rect -1163 -11245 -1129 -11211
rect -1095 -11245 -1061 -11211
rect -1027 -11245 -993 -11211
rect -959 -11245 -925 -11211
rect -891 -11245 -857 -11211
rect -823 -11245 -789 -11211
rect -755 -11245 -721 -11211
rect -687 -11245 -653 -11211
rect -619 -11245 -585 -11211
rect -551 -11245 -517 -11211
rect -483 -11245 -449 -11211
rect -415 -11245 -381 -11211
rect -347 -11245 -313 -11211
rect -279 -11245 -245 -11211
rect -211 -11245 -177 -11211
rect -143 -11245 -109 -11211
rect -75 -11245 -41 -11211
rect -7 -11245 27 -11211
rect 61 -11245 95 -11211
rect 129 -11245 163 -11211
rect 197 -11245 231 -11211
rect 265 -11245 299 -11211
rect 333 -11245 367 -11211
rect 401 -11245 435 -11211
rect 469 -11245 503 -11211
rect 537 -11245 571 -11211
rect 605 -11245 639 -11211
rect 673 -11245 707 -11211
rect 741 -11245 775 -11211
rect 809 -11245 843 -11211
rect 877 -11245 911 -11211
rect 945 -11245 979 -11211
rect 1013 -11245 1047 -11211
rect 1081 -11245 1115 -11211
rect 1149 -11245 1183 -11211
rect 1217 -11245 1251 -11211
rect 1285 -11245 1319 -11211
rect 1353 -11245 1387 -11211
rect 1421 -11245 1455 -11211
rect 1489 -11245 1523 -11211
rect 1557 -11245 1591 -11211
rect 1625 -11245 1659 -11211
rect 1693 -11245 1727 -11211
rect 1761 -11245 1795 -11211
rect 1829 -11245 1863 -11211
rect 1897 -11245 1931 -11211
rect 1965 -11245 1999 -11211
rect 2033 -11245 2067 -11211
rect 2101 -11245 2135 -11211
rect 2169 -11245 2203 -11211
rect 2237 -11245 2271 -11211
rect 2305 -11245 2339 -11211
rect 2373 -11245 2407 -11211
rect 2441 -11245 2475 -11211
rect 2509 -11245 2543 -11211
rect 2577 -11245 2611 -11211
rect 2645 -11245 2679 -11211
rect 2713 -11245 2747 -11211
rect 2781 -11245 2815 -11211
rect 2849 -11245 2883 -11211
rect 2917 -11245 2951 -11211
rect 2985 -11245 3019 -11211
rect 3053 -11245 3087 -11211
rect 3121 -11245 3155 -11211
rect 3189 -11245 3223 -11211
rect 3257 -11245 3291 -11211
rect 3325 -11245 3359 -11211
rect 3393 -11245 3427 -11211
rect 3461 -11245 3495 -11211
rect 3529 -11245 3563 -11211
rect 3597 -11245 3631 -11211
rect 3665 -11245 3699 -11211
rect 3733 -11245 3767 -11211
rect 3801 -11245 3835 -11211
rect 3869 -11245 3903 -11211
rect 3937 -11245 3971 -11211
rect 4005 -11245 4039 -11211
rect 4073 -11245 4107 -11211
rect 4141 -11245 4175 -11211
rect 4209 -11245 4243 -11211
rect 4277 -11245 4311 -11211
rect 4345 -11245 4379 -11211
rect 4413 -11245 4447 -11211
rect 4481 -11245 4515 -11211
rect 4549 -11245 4583 -11211
rect 4617 -11245 4651 -11211
rect 4685 -11245 4719 -11211
rect 4753 -11245 4787 -11211
rect 4821 -11245 4855 -11211
rect 4889 -11245 4923 -11211
rect 4957 -11245 4991 -11211
rect 5025 -11245 5059 -11211
rect 5093 -11245 5127 -11211
rect 5161 -11245 5195 -11211
rect 5229 -11245 5263 -11211
rect 5297 -11245 5331 -11211
rect 5365 -11245 5399 -11211
rect 5433 -11245 5467 -11211
rect 5501 -11245 5535 -11211
rect 5569 -11245 5603 -11211
rect 5637 -11245 5671 -11211
rect 5705 -11245 5739 -11211
rect 5773 -11245 5807 -11211
rect 5841 -11245 5875 -11211
rect 5909 -11245 5943 -11211
rect 5977 -11245 6011 -11211
rect 6045 -11245 6079 -11211
rect 6113 -11245 6147 -11211
rect 6181 -11245 6215 -11211
rect 6249 -11245 6283 -11211
rect 6317 -11245 6351 -11211
rect 6385 -11245 6419 -11211
rect 6453 -11245 6487 -11211
rect 6521 -11245 6555 -11211
rect 6589 -11245 6623 -11211
rect 6657 -11245 6691 -11211
rect 6725 -11245 6759 -11211
rect 6793 -11245 6827 -11211
rect 6861 -11245 6895 -11211
rect 6929 -11245 6963 -11211
rect 6997 -11245 7031 -11211
rect 7065 -11245 7099 -11211
rect 7133 -11245 7167 -11211
rect 7201 -11245 7235 -11211
rect 7269 -11245 7303 -11211
rect 7337 -11245 7371 -11211
rect 7405 -11245 7439 -11211
rect 7473 -11245 7507 -11211
rect 7541 -11245 7575 -11211
rect 7609 -11245 7643 -11211
rect 7677 -11245 7711 -11211
rect 7745 -11245 7779 -11211
rect 7813 -11245 7847 -11211
rect 7881 -11245 7915 -11211
rect 7949 -11245 7983 -11211
rect 8017 -11245 8051 -11211
rect 8085 -11245 8119 -11211
rect 8153 -11245 8187 -11211
rect 8221 -11245 8255 -11211
rect 8289 -11245 8323 -11211
rect 8357 -11245 8391 -11211
rect 8425 -11245 8459 -11211
rect 8493 -11245 8527 -11211
rect 8561 -11245 8595 -11211
rect 8629 -11245 8663 -11211
rect 8697 -11245 8731 -11211
rect 8765 -11245 8799 -11211
rect 8833 -11245 8867 -11211
rect 8901 -11245 8935 -11211
rect 8969 -11245 9003 -11211
rect 9037 -11245 9071 -11211
rect 9105 -11245 9139 -11211
rect 9173 -11245 9207 -11211
rect 9241 -11245 9275 -11211
rect 9309 -11245 9343 -11211
rect 9377 -11245 9411 -11211
rect 9445 -11245 9479 -11211
rect 9513 -11245 9547 -11211
rect 9581 -11245 9615 -11211
rect 9649 -11245 9683 -11211
rect 9717 -11245 9751 -11211
rect 9785 -11245 9819 -11211
rect 9853 -11245 9887 -11211
rect 9921 -11245 9955 -11211
rect 9989 -11245 10023 -11211
rect 10057 -11245 10091 -11211
rect 10125 -11245 10159 -11211
rect 10193 -11245 10227 -11211
rect 10261 -11245 10295 -11211
rect 10329 -11245 10363 -11211
rect 10397 -11245 10431 -11211
rect 10465 -11245 10499 -11211
rect 10533 -11245 10567 -11211
rect 10601 -11245 10635 -11211
rect 10669 -11245 10703 -11211
rect 10737 -11245 10771 -11211
rect 10805 -11245 10839 -11211
rect 10873 -11245 10907 -11211
rect 10941 -11245 10975 -11211
rect 11009 -11245 11043 -11211
rect 11077 -11245 11111 -11211
rect 11145 -11245 11179 -11211
rect 11213 -11245 11247 -11211
rect 11281 -11245 11315 -11211
rect 11349 -11245 11383 -11211
rect 11417 -11245 11451 -11211
rect 11485 -11245 11519 -11211
rect 11553 -11245 11587 -11211
rect 11621 -11245 11655 -11211
rect 11689 -11245 11723 -11211
rect 11757 -11245 11791 -11211
rect 11825 -11245 11859 -11211
rect 11893 -11245 11927 -11211
rect 11961 -11245 11995 -11211
rect 12029 -11245 12063 -11211
rect 12097 -11245 12131 -11211
rect 12165 -11245 12199 -11211
rect 12233 -11245 12267 -11211
rect 12301 -11245 12335 -11211
rect 12369 -11245 12403 -11211
rect 12437 -11245 12471 -11211
rect 12505 -11245 12539 -11211
rect 12573 -11245 12607 -11211
rect 12641 -11245 12675 -11211
rect 12709 -11245 12743 -11211
rect 12777 -11245 12811 -11211
rect 12845 -11245 12879 -11211
rect 12913 -11245 12947 -11211
rect 12981 -11245 13015 -11211
rect 13049 -11245 13083 -11211
rect 13117 -11245 13151 -11211
rect 13185 -11245 13219 -11211
rect 13253 -11245 13287 -11211
rect 13321 -11245 13355 -11211
rect 13389 -11245 13423 -11211
rect 13457 -11245 13491 -11211
rect 13525 -11245 13559 -11211
rect 13593 -11245 13627 -11211
rect 13661 -11245 13695 -11211
rect 13729 -11245 13763 -11211
rect 13797 -11245 13831 -11211
rect 13865 -11245 13899 -11211
rect 13933 -11245 13967 -11211
rect 14001 -11245 14035 -11211
rect 14069 -11245 14103 -11211
rect 14137 -11245 14171 -11211
rect 14205 -11245 14239 -11211
rect 14273 -11245 14307 -11211
rect 14341 -11245 14375 -11211
rect 14409 -11245 14443 -11211
rect 14477 -11245 14511 -11211
rect 14545 -11245 14579 -11211
rect 14613 -11245 14647 -11211
rect 14681 -11245 14715 -11211
rect 14749 -11245 14783 -11211
rect 14817 -11245 14851 -11211
rect 14885 -11245 14919 -11211
rect 14953 -11245 14987 -11211
rect 15021 -11245 15055 -11211
rect 15089 -11245 15123 -11211
rect 15157 -11245 15191 -11211
rect 15225 -11245 15259 -11211
rect 15293 -11245 15327 -11211
rect 15361 -11245 15395 -11211
rect 15429 -11245 15463 -11211
rect 15497 -11245 15531 -11211
rect 15565 -11245 15599 -11211
rect 15633 -11245 15667 -11211
rect 15701 -11245 15735 -11211
rect 15769 -11245 15803 -11211
rect 15837 -11245 15871 -11211
rect 15905 -11245 15939 -11211
rect 15973 -11245 16007 -11211
rect 16041 -11245 16075 -11211
rect 16109 -11245 16143 -11211
rect 16177 -11245 16211 -11211
rect 16245 -11245 16279 -11211
rect 16313 -11245 16347 -11211
rect 16381 -11245 16415 -11211
rect 16449 -11245 16483 -11211
rect 16517 -11245 16551 -11211
rect 16585 -11245 16619 -11211
rect 16653 -11245 16687 -11211
rect 16721 -11245 16755 -11211
rect 16789 -11245 16823 -11211
rect 16857 -11245 16891 -11211
rect 16925 -11245 16959 -11211
rect 16993 -11245 17027 -11211
rect 17061 -11245 17095 -11211
rect 17129 -11245 17163 -11211
rect 17197 -11245 17231 -11211
rect 17265 -11245 17299 -11211
rect 17333 -11245 17367 -11211
rect 17401 -11245 17435 -11211
rect 17469 -11245 17503 -11211
rect 17537 -11245 17571 -11211
rect 17605 -11245 17639 -11211
rect 17673 -11245 17707 -11211
rect 17741 -11245 17775 -11211
rect 17809 -11245 17843 -11211
rect 17877 -11245 17911 -11211
rect 17945 -11245 17979 -11211
rect 18013 -11245 18047 -11211
rect 18081 -11245 18115 -11211
rect 18149 -11245 18183 -11211
rect 18217 -11245 18251 -11211
rect 18285 -11245 18319 -11211
rect 18353 -11245 18387 -11211
rect 18421 -11245 18455 -11211
rect 18489 -11245 18523 -11211
rect 18557 -11245 18591 -11211
rect 18625 -11245 18659 -11211
rect 18693 -11245 18727 -11211
rect 18761 -11245 18795 -11211
rect 18829 -11245 18863 -11211
rect 18897 -11245 18931 -11211
rect 18965 -11245 18999 -11211
rect 19033 -11245 19067 -11211
rect 19101 -11245 19135 -11211
rect 19169 -11245 19203 -11211
rect 19237 -11245 19271 -11211
rect 19305 -11245 19339 -11211
rect 19373 -11245 19407 -11211
rect 19441 -11245 19475 -11211
rect 19509 -11245 19543 -11211
rect 19577 -11245 19611 -11211
rect 19645 -11245 19679 -11211
rect 19713 -11245 19747 -11211
rect 19781 -11245 19815 -11211
rect 19849 -11245 19883 -11211
rect 19917 -11245 19951 -11211
rect 19985 -11245 20019 -11211
rect 20053 -11245 20087 -11211
rect 20121 -11245 20155 -11211
rect 20189 -11245 20223 -11211
rect 20257 -11245 20291 -11211
rect 20325 -11245 20359 -11211
rect 20393 -11245 20427 -11211
rect 20461 -11245 20495 -11211
rect 20529 -11245 20563 -11211
rect 20597 -11245 20631 -11211
rect 20665 -11245 20699 -11211
rect 20733 -11245 20767 -11211
rect 20801 -11245 20835 -11211
rect 20869 -11245 20903 -11211
rect 20937 -11245 20971 -11211
rect 21005 -11245 21039 -11211
rect 21073 -11245 21107 -11211
rect 21141 -11245 21175 -11211
rect 21209 -11245 21243 -11211
rect 21277 -11245 21311 -11211
rect 21345 -11245 21379 -11211
rect 21413 -11245 21447 -11211
rect 21481 -11245 21515 -11211
rect 21549 -11245 21583 -11211
rect 21617 -11245 21651 -11211
rect 21685 -11245 21719 -11211
rect 21753 -11245 21787 -11211
rect 21821 -11245 21855 -11211
rect 21889 -11245 21923 -11211
rect 21957 -11245 21991 -11211
rect 22025 -11245 22059 -11211
rect 22093 -11245 22127 -11211
rect 22161 -11245 22195 -11211
rect 22229 -11245 22263 -11211
rect 22297 -11245 22331 -11211
rect 22365 -11245 22399 -11211
rect 22433 -11245 22467 -11211
rect 22501 -11245 22535 -11211
rect 22569 -11245 22603 -11211
rect 22637 -11245 22671 -11211
rect 22705 -11245 22739 -11211
rect 22773 -11245 22807 -11211
rect 22841 -11245 22875 -11211
rect 22909 -11245 22943 -11211
rect 22977 -11245 23011 -11211
rect 23045 -11245 23079 -11211
rect 23113 -11245 23147 -11211
rect 23181 -11245 23215 -11211
rect 23249 -11245 23283 -11211
rect 23317 -11245 23351 -11211
rect 23385 -11245 23419 -11211
rect 23453 -11245 23487 -11211
rect 23521 -11245 23555 -11211
rect 23589 -11245 23623 -11211
rect 23657 -11245 23691 -11211
rect 23725 -11245 23759 -11211
rect 23793 -11245 23827 -11211
rect 23861 -11245 23895 -11211
rect 23929 -11245 23963 -11211
rect 23997 -11245 24031 -11211
rect 24065 -11245 24099 -11211
rect 24133 -11245 24167 -11211
rect 24201 -11245 24235 -11211
rect 24269 -11245 24303 -11211
rect 24337 -11245 24371 -11211
rect 24405 -11245 24439 -11211
rect 24473 -11245 24507 -11211
rect 24541 -11245 24575 -11211
rect 24609 -11245 24643 -11211
rect 24677 -11245 24711 -11211
rect 24745 -11245 24922 -11211
rect -12322 -11278 24922 -11245
rect -12322 -11363 -12222 -11278
rect -12322 -11397 -12289 -11363
rect -12255 -11397 -12222 -11363
rect -12322 -11431 -12222 -11397
rect -12322 -11465 -12289 -11431
rect -12255 -11465 -12222 -11431
rect -12322 -11499 -12222 -11465
rect -12322 -11533 -12289 -11499
rect -12255 -11533 -12222 -11499
rect -12322 -11567 -12222 -11533
rect -12322 -11601 -12289 -11567
rect -12255 -11601 -12222 -11567
rect -12322 -11635 -12222 -11601
rect -12322 -11669 -12289 -11635
rect -12255 -11669 -12222 -11635
rect -12322 -11703 -12222 -11669
rect -12322 -11737 -12289 -11703
rect -12255 -11737 -12222 -11703
rect -12322 -11771 -12222 -11737
rect -12322 -11805 -12289 -11771
rect -12255 -11805 -12222 -11771
rect -12322 -11839 -12222 -11805
rect -12322 -11873 -12289 -11839
rect -12255 -11873 -12222 -11839
rect -12322 -11907 -12222 -11873
rect -12322 -11941 -12289 -11907
rect -12255 -11941 -12222 -11907
rect -12322 -11975 -12222 -11941
rect -12322 -12009 -12289 -11975
rect -12255 -12009 -12222 -11975
rect -12322 -12043 -12222 -12009
rect -12322 -12077 -12289 -12043
rect -12255 -12077 -12222 -12043
rect -12322 -12111 -12222 -12077
rect -12322 -12145 -12289 -12111
rect -12255 -12145 -12222 -12111
rect -12322 -12179 -12222 -12145
rect -12322 -12213 -12289 -12179
rect -12255 -12213 -12222 -12179
rect -12322 -12247 -12222 -12213
rect -12322 -12281 -12289 -12247
rect -12255 -12281 -12222 -12247
rect -12322 -12315 -12222 -12281
rect -12322 -12349 -12289 -12315
rect -12255 -12349 -12222 -12315
rect -12322 -12383 -12222 -12349
rect -12322 -12417 -12289 -12383
rect -12255 -12417 -12222 -12383
rect -12322 -12451 -12222 -12417
rect 24822 -11363 24922 -11278
rect 24822 -11397 24855 -11363
rect 24889 -11397 24922 -11363
rect 24822 -11431 24922 -11397
rect 24822 -11465 24855 -11431
rect 24889 -11465 24922 -11431
rect 24822 -11499 24922 -11465
rect 24822 -11533 24855 -11499
rect 24889 -11533 24922 -11499
rect 24822 -11567 24922 -11533
rect 24822 -11601 24855 -11567
rect 24889 -11601 24922 -11567
rect 24822 -11635 24922 -11601
rect 24822 -11669 24855 -11635
rect 24889 -11669 24922 -11635
rect 24822 -11703 24922 -11669
rect 24822 -11737 24855 -11703
rect 24889 -11737 24922 -11703
rect 24822 -11771 24922 -11737
rect 24822 -11805 24855 -11771
rect 24889 -11805 24922 -11771
rect 24822 -11839 24922 -11805
rect 24822 -11873 24855 -11839
rect 24889 -11873 24922 -11839
rect 24822 -11907 24922 -11873
rect 24822 -11941 24855 -11907
rect 24889 -11941 24922 -11907
rect 24822 -11975 24922 -11941
rect 24822 -12009 24855 -11975
rect 24889 -12009 24922 -11975
rect 24822 -12043 24922 -12009
rect 24822 -12077 24855 -12043
rect 24889 -12077 24922 -12043
rect 24822 -12111 24922 -12077
rect 24822 -12145 24855 -12111
rect 24889 -12145 24922 -12111
rect 24822 -12179 24922 -12145
rect 24822 -12213 24855 -12179
rect 24889 -12213 24922 -12179
rect 24822 -12247 24922 -12213
rect 24822 -12281 24855 -12247
rect 24889 -12281 24922 -12247
rect 24822 -12315 24922 -12281
rect 24822 -12349 24855 -12315
rect 24889 -12349 24922 -12315
rect 24822 -12383 24922 -12349
rect 24822 -12417 24855 -12383
rect 24889 -12417 24922 -12383
rect -12322 -12485 -12289 -12451
rect -12255 -12485 -12222 -12451
rect -12322 -12519 -12222 -12485
rect 24822 -12451 24922 -12417
rect 24822 -12485 24855 -12451
rect 24889 -12485 24922 -12451
rect -12322 -12553 -12289 -12519
rect -12255 -12553 -12222 -12519
rect -12322 -12587 -12222 -12553
rect -12322 -12621 -12289 -12587
rect -12255 -12621 -12222 -12587
rect -12322 -12655 -12222 -12621
rect -12322 -12689 -12289 -12655
rect -12255 -12689 -12222 -12655
rect -12322 -12723 -12222 -12689
rect -12322 -12757 -12289 -12723
rect -12255 -12757 -12222 -12723
rect -12322 -12791 -12222 -12757
rect -12322 -12825 -12289 -12791
rect -12255 -12825 -12222 -12791
rect -12322 -12859 -12222 -12825
rect -12322 -12893 -12289 -12859
rect -12255 -12893 -12222 -12859
rect -12322 -12927 -12222 -12893
rect -12322 -12961 -12289 -12927
rect -12255 -12961 -12222 -12927
rect -12322 -12995 -12222 -12961
rect -12322 -13029 -12289 -12995
rect -12255 -13029 -12222 -12995
rect -12322 -13063 -12222 -13029
rect -12322 -13097 -12289 -13063
rect -12255 -13097 -12222 -13063
rect -12322 -13131 -12222 -13097
rect 24822 -12519 24922 -12485
rect 24822 -12553 24855 -12519
rect 24889 -12553 24922 -12519
rect 24822 -12587 24922 -12553
rect 24822 -12621 24855 -12587
rect 24889 -12621 24922 -12587
rect 24822 -12655 24922 -12621
rect 24822 -12689 24855 -12655
rect 24889 -12689 24922 -12655
rect 24822 -12723 24922 -12689
rect 24822 -12757 24855 -12723
rect 24889 -12757 24922 -12723
rect 24822 -12791 24922 -12757
rect 24822 -12825 24855 -12791
rect 24889 -12825 24922 -12791
rect 24822 -12859 24922 -12825
rect 24822 -12893 24855 -12859
rect 24889 -12893 24922 -12859
rect 24822 -12927 24922 -12893
rect 24822 -12961 24855 -12927
rect 24889 -12961 24922 -12927
rect 24822 -12995 24922 -12961
rect 24822 -13029 24855 -12995
rect 24889 -13029 24922 -12995
rect 24822 -13063 24922 -13029
rect 24822 -13097 24855 -13063
rect 24889 -13097 24922 -13063
rect -12322 -13165 -12289 -13131
rect -12255 -13165 -12222 -13131
rect -12322 -13199 -12222 -13165
rect -12322 -13233 -12289 -13199
rect -12255 -13233 -12222 -13199
rect 24822 -13131 24922 -13097
rect 24822 -13165 24855 -13131
rect 24889 -13165 24922 -13131
rect 24822 -13199 24922 -13165
rect -12322 -13267 -12222 -13233
rect 24822 -13233 24855 -13199
rect 24889 -13233 24922 -13199
rect -12322 -13301 -12289 -13267
rect -12255 -13301 -12222 -13267
rect -12322 -13335 -12222 -13301
rect 24822 -13267 24922 -13233
rect 24822 -13301 24855 -13267
rect 24889 -13301 24922 -13267
rect -12322 -13369 -12289 -13335
rect -12255 -13369 -12222 -13335
rect -12322 -13403 -12222 -13369
rect -12322 -13437 -12289 -13403
rect -12255 -13437 -12222 -13403
rect -12322 -13471 -12222 -13437
rect -12322 -13505 -12289 -13471
rect -12255 -13505 -12222 -13471
rect -12322 -13539 -12222 -13505
rect -12322 -13573 -12289 -13539
rect -12255 -13573 -12222 -13539
rect -12322 -13607 -12222 -13573
rect -12322 -13641 -12289 -13607
rect -12255 -13641 -12222 -13607
rect -12322 -13675 -12222 -13641
rect -12322 -13709 -12289 -13675
rect -12255 -13709 -12222 -13675
rect -12322 -13743 -12222 -13709
rect -12322 -13777 -12289 -13743
rect -12255 -13777 -12222 -13743
rect -12322 -13811 -12222 -13777
rect -12322 -13845 -12289 -13811
rect -12255 -13845 -12222 -13811
rect -12322 -13879 -12222 -13845
rect -12322 -13913 -12289 -13879
rect -12255 -13913 -12222 -13879
rect -12322 -13947 -12222 -13913
rect 24822 -13335 24922 -13301
rect 24822 -13369 24855 -13335
rect 24889 -13369 24922 -13335
rect 24822 -13403 24922 -13369
rect 24822 -13437 24855 -13403
rect 24889 -13437 24922 -13403
rect 24822 -13471 24922 -13437
rect 24822 -13505 24855 -13471
rect 24889 -13505 24922 -13471
rect 24822 -13539 24922 -13505
rect 24822 -13573 24855 -13539
rect 24889 -13573 24922 -13539
rect 24822 -13607 24922 -13573
rect 24822 -13641 24855 -13607
rect 24889 -13641 24922 -13607
rect 24822 -13675 24922 -13641
rect 24822 -13709 24855 -13675
rect 24889 -13709 24922 -13675
rect 24822 -13743 24922 -13709
rect 24822 -13777 24855 -13743
rect 24889 -13777 24922 -13743
rect 24822 -13811 24922 -13777
rect 24822 -13845 24855 -13811
rect 24889 -13845 24922 -13811
rect 24822 -13879 24922 -13845
rect 24822 -13913 24855 -13879
rect 24889 -13913 24922 -13879
rect -12322 -13981 -12289 -13947
rect -12255 -13981 -12222 -13947
rect -12322 -14015 -12222 -13981
rect -12322 -14049 -12289 -14015
rect -12255 -14049 -12222 -14015
rect 24822 -13947 24922 -13913
rect 24822 -13981 24855 -13947
rect 24889 -13981 24922 -13947
rect 24822 -14015 24922 -13981
rect -12322 -14083 -12222 -14049
rect 24822 -14049 24855 -14015
rect 24889 -14049 24922 -14015
rect -12322 -14117 -12289 -14083
rect -12255 -14117 -12222 -14083
rect -12322 -14151 -12222 -14117
rect 24822 -14083 24922 -14049
rect 24822 -14117 24855 -14083
rect 24889 -14117 24922 -14083
rect -12322 -14185 -12289 -14151
rect -12255 -14185 -12222 -14151
rect -12322 -14219 -12222 -14185
rect -12322 -14253 -12289 -14219
rect -12255 -14253 -12222 -14219
rect -12322 -14287 -12222 -14253
rect -12322 -14321 -12289 -14287
rect -12255 -14321 -12222 -14287
rect -12322 -14355 -12222 -14321
rect -12322 -14389 -12289 -14355
rect -12255 -14389 -12222 -14355
rect -12322 -14423 -12222 -14389
rect -12322 -14457 -12289 -14423
rect -12255 -14457 -12222 -14423
rect -12322 -14491 -12222 -14457
rect -12322 -14525 -12289 -14491
rect -12255 -14525 -12222 -14491
rect -12322 -14559 -12222 -14525
rect -12322 -14593 -12289 -14559
rect -12255 -14593 -12222 -14559
rect -12322 -14627 -12222 -14593
rect -12322 -14661 -12289 -14627
rect -12255 -14661 -12222 -14627
rect -12322 -14695 -12222 -14661
rect -12322 -14729 -12289 -14695
rect -12255 -14729 -12222 -14695
rect -12322 -14763 -12222 -14729
rect 24822 -14151 24922 -14117
rect 24822 -14185 24855 -14151
rect 24889 -14185 24922 -14151
rect 24822 -14219 24922 -14185
rect -12322 -14797 -12289 -14763
rect -12255 -14797 -12222 -14763
rect -12322 -14831 -12222 -14797
rect -12322 -14865 -12289 -14831
rect -12255 -14865 -12222 -14831
rect 24822 -14253 24855 -14219
rect 24889 -14253 24922 -14219
rect 24822 -14287 24922 -14253
rect 24822 -14321 24855 -14287
rect 24889 -14321 24922 -14287
rect 24822 -14355 24922 -14321
rect 24822 -14389 24855 -14355
rect 24889 -14389 24922 -14355
rect 24822 -14423 24922 -14389
rect 24822 -14457 24855 -14423
rect 24889 -14457 24922 -14423
rect 24822 -14491 24922 -14457
rect 24822 -14525 24855 -14491
rect 24889 -14525 24922 -14491
rect 24822 -14559 24922 -14525
rect 24822 -14593 24855 -14559
rect 24889 -14593 24922 -14559
rect 24822 -14627 24922 -14593
rect 24822 -14661 24855 -14627
rect 24889 -14661 24922 -14627
rect 24822 -14695 24922 -14661
rect 24822 -14729 24855 -14695
rect 24889 -14729 24922 -14695
rect 24822 -14763 24922 -14729
rect 24822 -14797 24855 -14763
rect 24889 -14797 24922 -14763
rect 24822 -14831 24922 -14797
rect -12322 -14899 -12222 -14865
rect -12322 -14933 -12289 -14899
rect -12255 -14933 -12222 -14899
rect -12322 -14967 -12222 -14933
rect 24822 -14865 24855 -14831
rect 24889 -14865 24922 -14831
rect 24822 -14899 24922 -14865
rect 24822 -14933 24855 -14899
rect 24889 -14933 24922 -14899
rect -12322 -15001 -12289 -14967
rect -12255 -15001 -12222 -14967
rect -12322 -15035 -12222 -15001
rect -12322 -15069 -12289 -15035
rect -12255 -15069 -12222 -15035
rect -12322 -15103 -12222 -15069
rect -12322 -15137 -12289 -15103
rect -12255 -15137 -12222 -15103
rect -12322 -15171 -12222 -15137
rect -12322 -15205 -12289 -15171
rect -12255 -15205 -12222 -15171
rect -12322 -15239 -12222 -15205
rect -12322 -15273 -12289 -15239
rect -12255 -15273 -12222 -15239
rect -12322 -15307 -12222 -15273
rect -12322 -15341 -12289 -15307
rect -12255 -15341 -12222 -15307
rect -12322 -15375 -12222 -15341
rect -12322 -15409 -12289 -15375
rect -12255 -15409 -12222 -15375
rect -12322 -15443 -12222 -15409
rect -12322 -15477 -12289 -15443
rect -12255 -15477 -12222 -15443
rect -12322 -15511 -12222 -15477
rect -12322 -15545 -12289 -15511
rect -12255 -15545 -12222 -15511
rect -12322 -15579 -12222 -15545
rect 24822 -14967 24922 -14933
rect 24822 -15001 24855 -14967
rect 24889 -15001 24922 -14967
rect 24822 -15035 24922 -15001
rect 24822 -15069 24855 -15035
rect 24889 -15069 24922 -15035
rect 24822 -15103 24922 -15069
rect 24822 -15137 24855 -15103
rect 24889 -15137 24922 -15103
rect 24822 -15171 24922 -15137
rect 24822 -15205 24855 -15171
rect 24889 -15205 24922 -15171
rect 24822 -15239 24922 -15205
rect 24822 -15273 24855 -15239
rect 24889 -15273 24922 -15239
rect 24822 -15307 24922 -15273
rect 24822 -15341 24855 -15307
rect 24889 -15341 24922 -15307
rect 24822 -15375 24922 -15341
rect 24822 -15409 24855 -15375
rect 24889 -15409 24922 -15375
rect 24822 -15443 24922 -15409
rect -12322 -15613 -12289 -15579
rect -12255 -15613 -12222 -15579
rect -12322 -15647 -12222 -15613
rect -12322 -15681 -12289 -15647
rect -12255 -15681 -12222 -15647
rect -12322 -15715 -12222 -15681
rect -12322 -15749 -12289 -15715
rect -12255 -15749 -12222 -15715
rect -12322 -15783 -12222 -15749
rect -12322 -15817 -12289 -15783
rect -12255 -15817 -12222 -15783
rect -12322 -15851 -12222 -15817
rect -12322 -15885 -12289 -15851
rect -12255 -15885 -12222 -15851
rect -12322 -15919 -12222 -15885
rect -12322 -15953 -12289 -15919
rect -12255 -15953 -12222 -15919
rect -12322 -15987 -12222 -15953
rect -12322 -16021 -12289 -15987
rect -12255 -16021 -12222 -15987
rect -12322 -16055 -12222 -16021
rect -12322 -16089 -12289 -16055
rect -12255 -16089 -12222 -16055
rect -12322 -16123 -12222 -16089
rect -12322 -16157 -12289 -16123
rect -12255 -16157 -12222 -16123
rect -12322 -16191 -12222 -16157
rect -12322 -16225 -12289 -16191
rect -12255 -16225 -12222 -16191
rect -12322 -16259 -12222 -16225
rect -12322 -16293 -12289 -16259
rect -12255 -16293 -12222 -16259
rect -12322 -16327 -12222 -16293
rect -12322 -16361 -12289 -16327
rect -12255 -16361 -12222 -16327
rect -12322 -16395 -12222 -16361
rect 24822 -15477 24855 -15443
rect 24889 -15477 24922 -15443
rect 24822 -15511 24922 -15477
rect 24822 -15545 24855 -15511
rect 24889 -15545 24922 -15511
rect 24822 -15579 24922 -15545
rect 24822 -15613 24855 -15579
rect 24889 -15613 24922 -15579
rect 24822 -15647 24922 -15613
rect 24822 -15681 24855 -15647
rect 24889 -15681 24922 -15647
rect 24822 -15715 24922 -15681
rect 24822 -15749 24855 -15715
rect 24889 -15749 24922 -15715
rect 24822 -15783 24922 -15749
rect 24822 -15817 24855 -15783
rect 24889 -15817 24922 -15783
rect 24822 -15851 24922 -15817
rect 24822 -15885 24855 -15851
rect 24889 -15885 24922 -15851
rect 24822 -15919 24922 -15885
rect 24822 -15953 24855 -15919
rect 24889 -15953 24922 -15919
rect 24822 -15987 24922 -15953
rect 24822 -16021 24855 -15987
rect 24889 -16021 24922 -15987
rect 24822 -16055 24922 -16021
rect 24822 -16089 24855 -16055
rect 24889 -16089 24922 -16055
rect 24822 -16123 24922 -16089
rect 24822 -16157 24855 -16123
rect 24889 -16157 24922 -16123
rect 24822 -16191 24922 -16157
rect 24822 -16225 24855 -16191
rect 24889 -16225 24922 -16191
rect 24822 -16259 24922 -16225
rect 24822 -16293 24855 -16259
rect 24889 -16293 24922 -16259
rect 24822 -16327 24922 -16293
rect 24822 -16361 24855 -16327
rect 24889 -16361 24922 -16327
rect -12322 -16429 -12289 -16395
rect -12255 -16429 -12222 -16395
rect -12322 -16463 -12222 -16429
rect -12322 -16497 -12289 -16463
rect -12255 -16497 -12222 -16463
rect 24822 -16395 24922 -16361
rect 24822 -16429 24855 -16395
rect 24889 -16429 24922 -16395
rect 24822 -16463 24922 -16429
rect -12322 -16531 -12222 -16497
rect 24822 -16497 24855 -16463
rect 24889 -16497 24922 -16463
rect -12322 -16565 -12289 -16531
rect -12255 -16565 -12222 -16531
rect -12322 -16599 -12222 -16565
rect -12322 -16633 -12289 -16599
rect -12255 -16633 -12222 -16599
rect 24822 -16531 24922 -16497
rect 24822 -16565 24855 -16531
rect 24889 -16565 24922 -16531
rect 24822 -16599 24922 -16565
rect -12322 -16667 -12222 -16633
rect -12322 -16701 -12289 -16667
rect -12255 -16701 -12222 -16667
rect -12322 -16735 -12222 -16701
rect -12322 -16769 -12289 -16735
rect -12255 -16769 -12222 -16735
rect -12322 -16803 -12222 -16769
rect -12322 -16837 -12289 -16803
rect -12255 -16837 -12222 -16803
rect -12322 -16871 -12222 -16837
rect -12322 -16905 -12289 -16871
rect -12255 -16905 -12222 -16871
rect -12322 -16939 -12222 -16905
rect -12322 -16973 -12289 -16939
rect -12255 -16973 -12222 -16939
rect -12322 -17007 -12222 -16973
rect -12322 -17041 -12289 -17007
rect -12255 -17041 -12222 -17007
rect -12322 -17075 -12222 -17041
rect -12322 -17109 -12289 -17075
rect -12255 -17109 -12222 -17075
rect -12322 -17143 -12222 -17109
rect -12322 -17177 -12289 -17143
rect -12255 -17177 -12222 -17143
rect -12322 -17211 -12222 -17177
rect 24822 -16633 24855 -16599
rect 24889 -16633 24922 -16599
rect 24822 -16667 24922 -16633
rect -12322 -17245 -12289 -17211
rect -12255 -17245 -12222 -17211
rect -12322 -17279 -12222 -17245
rect -12322 -17313 -12289 -17279
rect -12255 -17313 -12222 -17279
rect 24822 -16701 24855 -16667
rect 24889 -16701 24922 -16667
rect 24822 -16735 24922 -16701
rect 24822 -16769 24855 -16735
rect 24889 -16769 24922 -16735
rect 24822 -16803 24922 -16769
rect 24822 -16837 24855 -16803
rect 24889 -16837 24922 -16803
rect 24822 -16871 24922 -16837
rect 24822 -16905 24855 -16871
rect 24889 -16905 24922 -16871
rect 24822 -16939 24922 -16905
rect 24822 -16973 24855 -16939
rect 24889 -16973 24922 -16939
rect 24822 -17007 24922 -16973
rect 24822 -17041 24855 -17007
rect 24889 -17041 24922 -17007
rect 24822 -17075 24922 -17041
rect 24822 -17109 24855 -17075
rect 24889 -17109 24922 -17075
rect 24822 -17143 24922 -17109
rect 24822 -17177 24855 -17143
rect 24889 -17177 24922 -17143
rect 24822 -17211 24922 -17177
rect 24822 -17245 24855 -17211
rect 24889 -17245 24922 -17211
rect 24822 -17279 24922 -17245
rect -12322 -17347 -12222 -17313
rect -12322 -17381 -12289 -17347
rect -12255 -17381 -12222 -17347
rect -12322 -17415 -12222 -17381
rect -12322 -17449 -12289 -17415
rect -12255 -17449 -12222 -17415
rect 24822 -17313 24855 -17279
rect 24889 -17313 24922 -17279
rect 24822 -17347 24922 -17313
rect 24822 -17381 24855 -17347
rect 24889 -17381 24922 -17347
rect 24822 -17415 24922 -17381
rect -12322 -17483 -12222 -17449
rect -12322 -17517 -12289 -17483
rect -12255 -17517 -12222 -17483
rect -12322 -17551 -12222 -17517
rect -12322 -17585 -12289 -17551
rect -12255 -17585 -12222 -17551
rect -12322 -17619 -12222 -17585
rect -12322 -17653 -12289 -17619
rect -12255 -17653 -12222 -17619
rect -12322 -17687 -12222 -17653
rect -12322 -17721 -12289 -17687
rect -12255 -17721 -12222 -17687
rect -12322 -17755 -12222 -17721
rect -12322 -17789 -12289 -17755
rect -12255 -17789 -12222 -17755
rect -12322 -17823 -12222 -17789
rect -12322 -17857 -12289 -17823
rect -12255 -17857 -12222 -17823
rect -12322 -17891 -12222 -17857
rect -12322 -17925 -12289 -17891
rect -12255 -17925 -12222 -17891
rect -12322 -17959 -12222 -17925
rect -12322 -17993 -12289 -17959
rect -12255 -17993 -12222 -17959
rect -12322 -18027 -12222 -17993
rect 24822 -17449 24855 -17415
rect 24889 -17449 24922 -17415
rect 24822 -17483 24922 -17449
rect 24822 -17517 24855 -17483
rect 24889 -17517 24922 -17483
rect 24822 -17551 24922 -17517
rect 24822 -17585 24855 -17551
rect 24889 -17585 24922 -17551
rect 24822 -17619 24922 -17585
rect 24822 -17653 24855 -17619
rect 24889 -17653 24922 -17619
rect 24822 -17687 24922 -17653
rect 24822 -17721 24855 -17687
rect 24889 -17721 24922 -17687
rect 24822 -17755 24922 -17721
rect 24822 -17789 24855 -17755
rect 24889 -17789 24922 -17755
rect 24822 -17823 24922 -17789
rect 24822 -17857 24855 -17823
rect 24889 -17857 24922 -17823
rect 24822 -17891 24922 -17857
rect 24822 -17925 24855 -17891
rect 24889 -17925 24922 -17891
rect -12322 -18061 -12289 -18027
rect -12255 -18061 -12222 -18027
rect -12322 -18095 -12222 -18061
rect -12322 -18129 -12289 -18095
rect -12255 -18129 -12222 -18095
rect -12322 -18163 -12222 -18129
rect -12322 -18197 -12289 -18163
rect -12255 -18197 -12222 -18163
rect -12322 -18231 -12222 -18197
rect -12322 -18265 -12289 -18231
rect -12255 -18265 -12222 -18231
rect -12322 -18299 -12222 -18265
rect -12322 -18333 -12289 -18299
rect -12255 -18333 -12222 -18299
rect -12322 -18367 -12222 -18333
rect -12322 -18401 -12289 -18367
rect -12255 -18401 -12222 -18367
rect -12322 -18435 -12222 -18401
rect -12322 -18469 -12289 -18435
rect -12255 -18469 -12222 -18435
rect -12322 -18503 -12222 -18469
rect -12322 -18537 -12289 -18503
rect -12255 -18537 -12222 -18503
rect -12322 -18571 -12222 -18537
rect -12322 -18605 -12289 -18571
rect -12255 -18605 -12222 -18571
rect -12322 -18639 -12222 -18605
rect -12322 -18673 -12289 -18639
rect -12255 -18673 -12222 -18639
rect -12322 -18707 -12222 -18673
rect -12322 -18741 -12289 -18707
rect -12255 -18741 -12222 -18707
rect -12322 -18775 -12222 -18741
rect -12322 -18809 -12289 -18775
rect -12255 -18809 -12222 -18775
rect -12322 -18843 -12222 -18809
rect 24822 -17959 24922 -17925
rect 24822 -17993 24855 -17959
rect 24889 -17993 24922 -17959
rect 24822 -18027 24922 -17993
rect 24822 -18061 24855 -18027
rect 24889 -18061 24922 -18027
rect 24822 -18095 24922 -18061
rect 24822 -18129 24855 -18095
rect 24889 -18129 24922 -18095
rect 24822 -18163 24922 -18129
rect 24822 -18197 24855 -18163
rect 24889 -18197 24922 -18163
rect 24822 -18231 24922 -18197
rect 24822 -18265 24855 -18231
rect 24889 -18265 24922 -18231
rect 24822 -18299 24922 -18265
rect 24822 -18333 24855 -18299
rect 24889 -18333 24922 -18299
rect 24822 -18367 24922 -18333
rect 24822 -18401 24855 -18367
rect 24889 -18401 24922 -18367
rect 24822 -18435 24922 -18401
rect 24822 -18469 24855 -18435
rect 24889 -18469 24922 -18435
rect 24822 -18503 24922 -18469
rect 24822 -18537 24855 -18503
rect 24889 -18537 24922 -18503
rect 24822 -18571 24922 -18537
rect 24822 -18605 24855 -18571
rect 24889 -18605 24922 -18571
rect 24822 -18639 24922 -18605
rect 24822 -18673 24855 -18639
rect 24889 -18673 24922 -18639
rect 24822 -18707 24922 -18673
rect 24822 -18741 24855 -18707
rect 24889 -18741 24922 -18707
rect 24822 -18775 24922 -18741
rect 24822 -18809 24855 -18775
rect 24889 -18809 24922 -18775
rect -12322 -18877 -12289 -18843
rect -12255 -18877 -12222 -18843
rect -12322 -18911 -12222 -18877
rect -12322 -18945 -12289 -18911
rect -12255 -18945 -12222 -18911
rect 24822 -18843 24922 -18809
rect 24822 -18877 24855 -18843
rect 24889 -18877 24922 -18843
rect 24822 -18911 24922 -18877
rect -12322 -18979 -12222 -18945
rect -12322 -19013 -12289 -18979
rect -12255 -19013 -12222 -18979
rect -12322 -19047 -12222 -19013
rect -12322 -19081 -12289 -19047
rect -12255 -19081 -12222 -19047
rect 24822 -18945 24855 -18911
rect 24889 -18945 24922 -18911
rect 24822 -18979 24922 -18945
rect 24822 -19013 24855 -18979
rect 24889 -19013 24922 -18979
rect 24822 -19047 24922 -19013
rect -12322 -19115 -12222 -19081
rect -12322 -19149 -12289 -19115
rect -12255 -19149 -12222 -19115
rect -12322 -19183 -12222 -19149
rect 24822 -19081 24855 -19047
rect 24889 -19081 24922 -19047
rect 24822 -19115 24922 -19081
rect 24822 -19149 24855 -19115
rect 24889 -19149 24922 -19115
rect -12322 -19217 -12289 -19183
rect -12255 -19217 -12222 -19183
rect -12322 -19251 -12222 -19217
rect -12322 -19285 -12289 -19251
rect -12255 -19285 -12222 -19251
rect -12322 -19319 -12222 -19285
rect -12322 -19353 -12289 -19319
rect -12255 -19353 -12222 -19319
rect -12322 -19387 -12222 -19353
rect -12322 -19421 -12289 -19387
rect -12255 -19421 -12222 -19387
rect -12322 -19455 -12222 -19421
rect -12322 -19489 -12289 -19455
rect -12255 -19489 -12222 -19455
rect -12322 -19523 -12222 -19489
rect -12322 -19557 -12289 -19523
rect -12255 -19557 -12222 -19523
rect -12322 -19591 -12222 -19557
rect -12322 -19625 -12289 -19591
rect -12255 -19625 -12222 -19591
rect -12322 -19659 -12222 -19625
rect -12322 -19693 -12289 -19659
rect -12255 -19693 -12222 -19659
rect -12322 -19727 -12222 -19693
rect -12322 -19761 -12289 -19727
rect -12255 -19761 -12222 -19727
rect -12322 -19795 -12222 -19761
rect 24822 -19183 24922 -19149
rect 24822 -19217 24855 -19183
rect 24889 -19217 24922 -19183
rect 24822 -19251 24922 -19217
rect 24822 -19285 24855 -19251
rect 24889 -19285 24922 -19251
rect 24822 -19319 24922 -19285
rect 24822 -19353 24855 -19319
rect 24889 -19353 24922 -19319
rect 24822 -19387 24922 -19353
rect 24822 -19421 24855 -19387
rect 24889 -19421 24922 -19387
rect 24822 -19455 24922 -19421
rect 24822 -19489 24855 -19455
rect 24889 -19489 24922 -19455
rect 24822 -19523 24922 -19489
rect 24822 -19557 24855 -19523
rect 24889 -19557 24922 -19523
rect 24822 -19591 24922 -19557
rect 24822 -19625 24855 -19591
rect 24889 -19625 24922 -19591
rect 24822 -19659 24922 -19625
rect 24822 -19693 24855 -19659
rect 24889 -19693 24922 -19659
rect 24822 -19727 24922 -19693
rect 24822 -19761 24855 -19727
rect 24889 -19761 24922 -19727
rect -12322 -19829 -12289 -19795
rect -12255 -19829 -12222 -19795
rect -12322 -19863 -12222 -19829
rect 24822 -19795 24922 -19761
rect 24822 -19829 24855 -19795
rect 24889 -19829 24922 -19795
rect -12322 -19897 -12289 -19863
rect -12255 -19897 -12222 -19863
rect -12322 -19931 -12222 -19897
rect -12322 -19965 -12289 -19931
rect -12255 -19965 -12222 -19931
rect -12322 -19999 -12222 -19965
rect -12322 -20033 -12289 -19999
rect -12255 -20033 -12222 -19999
rect -12322 -20067 -12222 -20033
rect -12322 -20101 -12289 -20067
rect -12255 -20101 -12222 -20067
rect -12322 -20135 -12222 -20101
rect -12322 -20169 -12289 -20135
rect -12255 -20169 -12222 -20135
rect -12322 -20203 -12222 -20169
rect -12322 -20237 -12289 -20203
rect -12255 -20237 -12222 -20203
rect -12322 -20271 -12222 -20237
rect -12322 -20305 -12289 -20271
rect -12255 -20305 -12222 -20271
rect -12322 -20339 -12222 -20305
rect 24822 -19863 24922 -19829
rect 24822 -19897 24855 -19863
rect 24889 -19897 24922 -19863
rect 24822 -19931 24922 -19897
rect 24822 -19965 24855 -19931
rect 24889 -19965 24922 -19931
rect 24822 -19999 24922 -19965
rect 24822 -20033 24855 -19999
rect 24889 -20033 24922 -19999
rect 24822 -20067 24922 -20033
rect 24822 -20101 24855 -20067
rect 24889 -20101 24922 -20067
rect 24822 -20135 24922 -20101
rect 24822 -20169 24855 -20135
rect 24889 -20169 24922 -20135
rect 24822 -20203 24922 -20169
rect 24822 -20237 24855 -20203
rect 24889 -20237 24922 -20203
rect 24822 -20271 24922 -20237
rect 24822 -20305 24855 -20271
rect 24889 -20305 24922 -20271
rect -12322 -20373 -12289 -20339
rect -12255 -20373 -12222 -20339
rect -12322 -20407 -12222 -20373
rect 24822 -20339 24922 -20305
rect 24822 -20373 24855 -20339
rect 24889 -20373 24922 -20339
rect -12322 -20441 -12289 -20407
rect -12255 -20441 -12222 -20407
rect -12322 -20475 -12222 -20441
rect -12322 -20509 -12289 -20475
rect -12255 -20509 -12222 -20475
rect -12322 -20543 -12222 -20509
rect -12322 -20577 -12289 -20543
rect -12255 -20577 -12222 -20543
rect -12322 -20611 -12222 -20577
rect -12322 -20645 -12289 -20611
rect -12255 -20645 -12222 -20611
rect -12322 -20679 -12222 -20645
rect -12322 -20713 -12289 -20679
rect -12255 -20713 -12222 -20679
rect -12322 -20747 -12222 -20713
rect -12322 -20781 -12289 -20747
rect -12255 -20781 -12222 -20747
rect -12322 -20815 -12222 -20781
rect -12322 -20849 -12289 -20815
rect -12255 -20849 -12222 -20815
rect -12322 -20883 -12222 -20849
rect -12322 -20917 -12289 -20883
rect -12255 -20917 -12222 -20883
rect -12322 -20951 -12222 -20917
rect -12322 -20985 -12289 -20951
rect -12255 -20985 -12222 -20951
rect -12322 -21019 -12222 -20985
rect 24822 -20407 24922 -20373
rect 24822 -20441 24855 -20407
rect 24889 -20441 24922 -20407
rect 24822 -20475 24922 -20441
rect 24822 -20509 24855 -20475
rect 24889 -20509 24922 -20475
rect 24822 -20543 24922 -20509
rect 24822 -20577 24855 -20543
rect 24889 -20577 24922 -20543
rect 24822 -20611 24922 -20577
rect 24822 -20645 24855 -20611
rect 24889 -20645 24922 -20611
rect 24822 -20679 24922 -20645
rect 24822 -20713 24855 -20679
rect 24889 -20713 24922 -20679
rect 24822 -20747 24922 -20713
rect 24822 -20781 24855 -20747
rect 24889 -20781 24922 -20747
rect 24822 -20815 24922 -20781
rect 24822 -20849 24855 -20815
rect 24889 -20849 24922 -20815
rect 24822 -20883 24922 -20849
rect 24822 -20917 24855 -20883
rect 24889 -20917 24922 -20883
rect 24822 -20951 24922 -20917
rect 24822 -20985 24855 -20951
rect 24889 -20985 24922 -20951
rect -12322 -21053 -12289 -21019
rect -12255 -21053 -12222 -21019
rect -12322 -21087 -12222 -21053
rect 24822 -21019 24922 -20985
rect 24822 -21053 24855 -21019
rect 24889 -21053 24922 -21019
rect -12322 -21121 -12289 -21087
rect -12255 -21121 -12222 -21087
rect -12322 -21155 -12222 -21121
rect -12322 -21189 -12289 -21155
rect -12255 -21189 -12222 -21155
rect -12322 -21223 -12222 -21189
rect -12322 -21257 -12289 -21223
rect -12255 -21257 -12222 -21223
rect -12322 -21291 -12222 -21257
rect -12322 -21325 -12289 -21291
rect -12255 -21325 -12222 -21291
rect -12322 -21359 -12222 -21325
rect -12322 -21393 -12289 -21359
rect -12255 -21393 -12222 -21359
rect -12322 -21427 -12222 -21393
rect -12322 -21461 -12289 -21427
rect -12255 -21461 -12222 -21427
rect -12322 -21495 -12222 -21461
rect -12322 -21529 -12289 -21495
rect -12255 -21529 -12222 -21495
rect -12322 -21563 -12222 -21529
rect 24822 -21087 24922 -21053
rect 24822 -21121 24855 -21087
rect 24889 -21121 24922 -21087
rect 24822 -21155 24922 -21121
rect 24822 -21189 24855 -21155
rect 24889 -21189 24922 -21155
rect 24822 -21223 24922 -21189
rect 24822 -21257 24855 -21223
rect 24889 -21257 24922 -21223
rect 24822 -21291 24922 -21257
rect 24822 -21325 24855 -21291
rect 24889 -21325 24922 -21291
rect 24822 -21359 24922 -21325
rect 24822 -21393 24855 -21359
rect 24889 -21393 24922 -21359
rect 24822 -21427 24922 -21393
rect 24822 -21461 24855 -21427
rect 24889 -21461 24922 -21427
rect 24822 -21495 24922 -21461
rect 24822 -21529 24855 -21495
rect 24889 -21529 24922 -21495
rect -12322 -21597 -12289 -21563
rect -12255 -21597 -12222 -21563
rect -12322 -21631 -12222 -21597
rect -12322 -21665 -12289 -21631
rect -12255 -21665 -12222 -21631
rect 24822 -21563 24922 -21529
rect 24822 -21597 24855 -21563
rect 24889 -21597 24922 -21563
rect 24822 -21631 24922 -21597
rect -12322 -21699 -12222 -21665
rect -12322 -21733 -12289 -21699
rect -12255 -21733 -12222 -21699
rect -12322 -21767 -12222 -21733
rect -12322 -21801 -12289 -21767
rect -12255 -21801 -12222 -21767
rect -12322 -21835 -12222 -21801
rect -12322 -21869 -12289 -21835
rect -12255 -21869 -12222 -21835
rect -12322 -21903 -12222 -21869
rect -12322 -21937 -12289 -21903
rect -12255 -21937 -12222 -21903
rect -12322 -21971 -12222 -21937
rect -12322 -22005 -12289 -21971
rect -12255 -22005 -12222 -21971
rect -12322 -22039 -12222 -22005
rect -12322 -22073 -12289 -22039
rect -12255 -22073 -12222 -22039
rect -12322 -22107 -12222 -22073
rect -12322 -22141 -12289 -22107
rect -12255 -22141 -12222 -22107
rect -12322 -22175 -12222 -22141
rect -12322 -22209 -12289 -22175
rect -12255 -22209 -12222 -22175
rect -12322 -22243 -12222 -22209
rect 24822 -21665 24855 -21631
rect 24889 -21665 24922 -21631
rect 24822 -21699 24922 -21665
rect 24822 -21733 24855 -21699
rect 24889 -21733 24922 -21699
rect 24822 -21767 24922 -21733
rect 24822 -21801 24855 -21767
rect 24889 -21801 24922 -21767
rect 24822 -21835 24922 -21801
rect 24822 -21869 24855 -21835
rect 24889 -21869 24922 -21835
rect 24822 -21903 24922 -21869
rect 24822 -21937 24855 -21903
rect 24889 -21937 24922 -21903
rect 24822 -21971 24922 -21937
rect 24822 -22005 24855 -21971
rect 24889 -22005 24922 -21971
rect 24822 -22039 24922 -22005
rect 24822 -22073 24855 -22039
rect 24889 -22073 24922 -22039
rect 24822 -22107 24922 -22073
rect 24822 -22141 24855 -22107
rect 24889 -22141 24922 -22107
rect 24822 -22175 24922 -22141
rect 24822 -22209 24855 -22175
rect 24889 -22209 24922 -22175
rect -12322 -22277 -12289 -22243
rect -12255 -22277 -12222 -22243
rect -12322 -22311 -12222 -22277
rect -12322 -22345 -12289 -22311
rect -12255 -22345 -12222 -22311
rect 24822 -22243 24922 -22209
rect 24822 -22277 24855 -22243
rect 24889 -22277 24922 -22243
rect 24822 -22311 24922 -22277
rect -12322 -22379 -12222 -22345
rect -12322 -22413 -12289 -22379
rect -12255 -22413 -12222 -22379
rect -12322 -22447 -12222 -22413
rect -12322 -22481 -12289 -22447
rect -12255 -22481 -12222 -22447
rect -12322 -22515 -12222 -22481
rect -12322 -22549 -12289 -22515
rect -12255 -22549 -12222 -22515
rect -12322 -22583 -12222 -22549
rect -12322 -22617 -12289 -22583
rect -12255 -22617 -12222 -22583
rect -12322 -22651 -12222 -22617
rect -12322 -22685 -12289 -22651
rect -12255 -22685 -12222 -22651
rect -12322 -22719 -12222 -22685
rect -12322 -22753 -12289 -22719
rect -12255 -22753 -12222 -22719
rect -12322 -22787 -12222 -22753
rect 24822 -22345 24855 -22311
rect 24889 -22345 24922 -22311
rect 24822 -22379 24922 -22345
rect 24822 -22413 24855 -22379
rect 24889 -22413 24922 -22379
rect 24822 -22447 24922 -22413
rect 24822 -22481 24855 -22447
rect 24889 -22481 24922 -22447
rect 24822 -22515 24922 -22481
rect 24822 -22549 24855 -22515
rect 24889 -22549 24922 -22515
rect 24822 -22583 24922 -22549
rect 24822 -22617 24855 -22583
rect 24889 -22617 24922 -22583
rect 24822 -22651 24922 -22617
rect 24822 -22685 24855 -22651
rect 24889 -22685 24922 -22651
rect 24822 -22719 24922 -22685
rect 24822 -22753 24855 -22719
rect 24889 -22753 24922 -22719
rect -12322 -22821 -12289 -22787
rect -12255 -22821 -12222 -22787
rect -12322 -22855 -12222 -22821
rect -12322 -22889 -12289 -22855
rect -12255 -22889 -12222 -22855
rect 24822 -22787 24922 -22753
rect 24822 -22821 24855 -22787
rect 24889 -22821 24922 -22787
rect 24822 -22855 24922 -22821
rect -12322 -22923 -12222 -22889
rect -12322 -22957 -12289 -22923
rect -12255 -22957 -12222 -22923
rect -12322 -22991 -12222 -22957
rect -12322 -23025 -12289 -22991
rect -12255 -23025 -12222 -22991
rect -12322 -23059 -12222 -23025
rect -12322 -23093 -12289 -23059
rect -12255 -23093 -12222 -23059
rect -12322 -23127 -12222 -23093
rect -12322 -23161 -12289 -23127
rect -12255 -23161 -12222 -23127
rect -12322 -23195 -12222 -23161
rect -12322 -23229 -12289 -23195
rect -12255 -23229 -12222 -23195
rect -12322 -23263 -12222 -23229
rect -12322 -23297 -12289 -23263
rect -12255 -23297 -12222 -23263
rect -12322 -23331 -12222 -23297
rect -12322 -23365 -12289 -23331
rect -12255 -23365 -12222 -23331
rect -12322 -23399 -12222 -23365
rect -12322 -23433 -12289 -23399
rect -12255 -23433 -12222 -23399
rect -12322 -23467 -12222 -23433
rect 24822 -22889 24855 -22855
rect 24889 -22889 24922 -22855
rect 24822 -22923 24922 -22889
rect 24822 -22957 24855 -22923
rect 24889 -22957 24922 -22923
rect 24822 -22991 24922 -22957
rect 24822 -23025 24855 -22991
rect 24889 -23025 24922 -22991
rect 24822 -23059 24922 -23025
rect 24822 -23093 24855 -23059
rect 24889 -23093 24922 -23059
rect 24822 -23127 24922 -23093
rect 24822 -23161 24855 -23127
rect 24889 -23161 24922 -23127
rect 24822 -23195 24922 -23161
rect 24822 -23229 24855 -23195
rect 24889 -23229 24922 -23195
rect 24822 -23263 24922 -23229
rect 24822 -23297 24855 -23263
rect 24889 -23297 24922 -23263
rect 24822 -23331 24922 -23297
rect 24822 -23365 24855 -23331
rect 24889 -23365 24922 -23331
rect 24822 -23399 24922 -23365
rect 24822 -23433 24855 -23399
rect 24889 -23433 24922 -23399
rect -12322 -23501 -12289 -23467
rect -12255 -23501 -12222 -23467
rect -12322 -23535 -12222 -23501
rect -12322 -23569 -12289 -23535
rect -12255 -23569 -12222 -23535
rect 24822 -23467 24922 -23433
rect 24822 -23501 24855 -23467
rect 24889 -23501 24922 -23467
rect 24822 -23535 24922 -23501
rect -12322 -23603 -12222 -23569
rect -12322 -23637 -12289 -23603
rect -12255 -23637 -12222 -23603
rect -12322 -23671 -12222 -23637
rect -12322 -23705 -12289 -23671
rect -12255 -23705 -12222 -23671
rect -12322 -23739 -12222 -23705
rect -12322 -23773 -12289 -23739
rect -12255 -23773 -12222 -23739
rect -12322 -23807 -12222 -23773
rect -12322 -23841 -12289 -23807
rect -12255 -23841 -12222 -23807
rect -12322 -23875 -12222 -23841
rect -12322 -23909 -12289 -23875
rect -12255 -23909 -12222 -23875
rect -12322 -23943 -12222 -23909
rect -12322 -23977 -12289 -23943
rect -12255 -23977 -12222 -23943
rect -12322 -24011 -12222 -23977
rect 24822 -23569 24855 -23535
rect 24889 -23569 24922 -23535
rect 24822 -23603 24922 -23569
rect 24822 -23637 24855 -23603
rect 24889 -23637 24922 -23603
rect 24822 -23671 24922 -23637
rect 24822 -23705 24855 -23671
rect 24889 -23705 24922 -23671
rect 24822 -23739 24922 -23705
rect 24822 -23773 24855 -23739
rect 24889 -23773 24922 -23739
rect 24822 -23807 24922 -23773
rect 24822 -23841 24855 -23807
rect 24889 -23841 24922 -23807
rect 24822 -23875 24922 -23841
rect 24822 -23909 24855 -23875
rect 24889 -23909 24922 -23875
rect 24822 -23943 24922 -23909
rect 24822 -23977 24855 -23943
rect 24889 -23977 24922 -23943
rect -12322 -24045 -12289 -24011
rect -12255 -24045 -12222 -24011
rect -12322 -24079 -12222 -24045
rect -12322 -24113 -12289 -24079
rect -12255 -24113 -12222 -24079
rect 24822 -24011 24922 -23977
rect 24822 -24045 24855 -24011
rect 24889 -24045 24922 -24011
rect 24822 -24079 24922 -24045
rect -12322 -24147 -12222 -24113
rect -12322 -24181 -12289 -24147
rect -12255 -24181 -12222 -24147
rect -12322 -24215 -12222 -24181
rect -12322 -24249 -12289 -24215
rect -12255 -24249 -12222 -24215
rect -12322 -24283 -12222 -24249
rect -12322 -24317 -12289 -24283
rect -12255 -24317 -12222 -24283
rect -12322 -24351 -12222 -24317
rect -12322 -24385 -12289 -24351
rect -12255 -24385 -12222 -24351
rect -12322 -24419 -12222 -24385
rect -12322 -24453 -12289 -24419
rect -12255 -24453 -12222 -24419
rect -12322 -24487 -12222 -24453
rect -12322 -24521 -12289 -24487
rect -12255 -24521 -12222 -24487
rect -12322 -24555 -12222 -24521
rect -12322 -24589 -12289 -24555
rect -12255 -24589 -12222 -24555
rect -12322 -24623 -12222 -24589
rect -12322 -24657 -12289 -24623
rect -12255 -24657 -12222 -24623
rect -12322 -24691 -12222 -24657
rect -12322 -24725 -12289 -24691
rect -12255 -24725 -12222 -24691
rect 24822 -24113 24855 -24079
rect 24889 -24113 24922 -24079
rect 24822 -24147 24922 -24113
rect 24822 -24181 24855 -24147
rect 24889 -24181 24922 -24147
rect 24822 -24215 24922 -24181
rect 24822 -24249 24855 -24215
rect 24889 -24249 24922 -24215
rect 24822 -24283 24922 -24249
rect 24822 -24317 24855 -24283
rect 24889 -24317 24922 -24283
rect 24822 -24351 24922 -24317
rect 24822 -24385 24855 -24351
rect 24889 -24385 24922 -24351
rect 24822 -24419 24922 -24385
rect 24822 -24453 24855 -24419
rect 24889 -24453 24922 -24419
rect 24822 -24487 24922 -24453
rect 24822 -24521 24855 -24487
rect 24889 -24521 24922 -24487
rect 24822 -24555 24922 -24521
rect 24822 -24589 24855 -24555
rect 24889 -24589 24922 -24555
rect 24822 -24623 24922 -24589
rect 24822 -24657 24855 -24623
rect 24889 -24657 24922 -24623
rect 24822 -24691 24922 -24657
rect -12322 -24759 -12222 -24725
rect -12322 -24793 -12289 -24759
rect -12255 -24793 -12222 -24759
rect 24822 -24725 24855 -24691
rect 24889 -24725 24922 -24691
rect 24822 -24759 24922 -24725
rect -12322 -24827 -12222 -24793
rect -12322 -24861 -12289 -24827
rect -12255 -24861 -12222 -24827
rect -12322 -24895 -12222 -24861
rect -12322 -24929 -12289 -24895
rect -12255 -24929 -12222 -24895
rect -12322 -24963 -12222 -24929
rect -12322 -24997 -12289 -24963
rect -12255 -24997 -12222 -24963
rect -12322 -25031 -12222 -24997
rect -12322 -25065 -12289 -25031
rect -12255 -25065 -12222 -25031
rect -12322 -25099 -12222 -25065
rect -12322 -25133 -12289 -25099
rect -12255 -25133 -12222 -25099
rect -12322 -25167 -12222 -25133
rect -12322 -25201 -12289 -25167
rect -12255 -25201 -12222 -25167
rect -12322 -25235 -12222 -25201
rect -12322 -25269 -12289 -25235
rect -12255 -25269 -12222 -25235
rect -12322 -25303 -12222 -25269
rect -12322 -25337 -12289 -25303
rect -12255 -25337 -12222 -25303
rect -12322 -25371 -12222 -25337
rect -12322 -25405 -12289 -25371
rect -12255 -25405 -12222 -25371
rect -12322 -25439 -12222 -25405
rect -12322 -25473 -12289 -25439
rect -12255 -25473 -12222 -25439
rect -12322 -25507 -12222 -25473
rect -12322 -25541 -12289 -25507
rect -12255 -25541 -12222 -25507
rect -12322 -25575 -12222 -25541
rect -12322 -25609 -12289 -25575
rect -12255 -25609 -12222 -25575
rect -12322 -25643 -12222 -25609
rect -12322 -25677 -12289 -25643
rect -12255 -25677 -12222 -25643
rect -12322 -25711 -12222 -25677
rect -12322 -25745 -12289 -25711
rect -12255 -25745 -12222 -25711
rect -12322 -25779 -12222 -25745
rect -12322 -25813 -12289 -25779
rect -12255 -25813 -12222 -25779
rect -12322 -25847 -12222 -25813
rect -12322 -25881 -12289 -25847
rect -12255 -25881 -12222 -25847
rect -12322 -25915 -12222 -25881
rect -12322 -25949 -12289 -25915
rect -12255 -25949 -12222 -25915
rect -12322 -25983 -12222 -25949
rect -12322 -26017 -12289 -25983
rect -12255 -26017 -12222 -25983
rect -12322 -26051 -12222 -26017
rect -12322 -26085 -12289 -26051
rect -12255 -26085 -12222 -26051
rect -12322 -26119 -12222 -26085
rect -12322 -26153 -12289 -26119
rect -12255 -26153 -12222 -26119
rect -12322 -26187 -12222 -26153
rect -12322 -26221 -12289 -26187
rect -12255 -26221 -12222 -26187
rect -12322 -26255 -12222 -26221
rect -12322 -26289 -12289 -26255
rect -12255 -26289 -12222 -26255
rect -12322 -26323 -12222 -26289
rect -12322 -26357 -12289 -26323
rect -12255 -26357 -12222 -26323
rect -12322 -26391 -12222 -26357
rect -12322 -26425 -12289 -26391
rect -12255 -26425 -12222 -26391
rect -12322 -26459 -12222 -26425
rect -12322 -26493 -12289 -26459
rect -12255 -26493 -12222 -26459
rect -12322 -26527 -12222 -26493
rect -12322 -26561 -12289 -26527
rect -12255 -26561 -12222 -26527
rect -12322 -26595 -12222 -26561
rect -12322 -26629 -12289 -26595
rect -12255 -26629 -12222 -26595
rect -12322 -26663 -12222 -26629
rect -12322 -26697 -12289 -26663
rect -12255 -26697 -12222 -26663
rect -12322 -26731 -12222 -26697
rect -12322 -26765 -12289 -26731
rect -12255 -26765 -12222 -26731
rect -12322 -26799 -12222 -26765
rect -12322 -26833 -12289 -26799
rect -12255 -26833 -12222 -26799
rect -12322 -26867 -12222 -26833
rect -12322 -26901 -12289 -26867
rect -12255 -26901 -12222 -26867
rect -12322 -26935 -12222 -26901
rect -12322 -26969 -12289 -26935
rect -12255 -26969 -12222 -26935
rect -12322 -27003 -12222 -26969
rect -12322 -27037 -12289 -27003
rect -12255 -27037 -12222 -27003
rect -12322 -27122 -12222 -27037
rect 24822 -24793 24855 -24759
rect 24889 -24793 24922 -24759
rect 24822 -24827 24922 -24793
rect 24822 -24861 24855 -24827
rect 24889 -24861 24922 -24827
rect 24822 -24895 24922 -24861
rect 24822 -24929 24855 -24895
rect 24889 -24929 24922 -24895
rect 24822 -24963 24922 -24929
rect 24822 -24997 24855 -24963
rect 24889 -24997 24922 -24963
rect 24822 -25031 24922 -24997
rect 24822 -25065 24855 -25031
rect 24889 -25065 24922 -25031
rect 24822 -25099 24922 -25065
rect 24822 -25133 24855 -25099
rect 24889 -25133 24922 -25099
rect 24822 -25167 24922 -25133
rect 24822 -25201 24855 -25167
rect 24889 -25201 24922 -25167
rect 24822 -25235 24922 -25201
rect 24822 -25269 24855 -25235
rect 24889 -25269 24922 -25235
rect 24822 -25303 24922 -25269
rect 24822 -25337 24855 -25303
rect 24889 -25337 24922 -25303
rect 24822 -25371 24922 -25337
rect 24822 -25405 24855 -25371
rect 24889 -25405 24922 -25371
rect 24822 -25439 24922 -25405
rect 24822 -25473 24855 -25439
rect 24889 -25473 24922 -25439
rect 24822 -25507 24922 -25473
rect 24822 -25541 24855 -25507
rect 24889 -25541 24922 -25507
rect 24822 -25575 24922 -25541
rect 24822 -25609 24855 -25575
rect 24889 -25609 24922 -25575
rect 24822 -25643 24922 -25609
rect 24822 -25677 24855 -25643
rect 24889 -25677 24922 -25643
rect 24822 -25711 24922 -25677
rect 24822 -25745 24855 -25711
rect 24889 -25745 24922 -25711
rect 24822 -25779 24922 -25745
rect 24822 -25813 24855 -25779
rect 24889 -25813 24922 -25779
rect 24822 -25847 24922 -25813
rect 24822 -25881 24855 -25847
rect 24889 -25881 24922 -25847
rect 24822 -25915 24922 -25881
rect 24822 -25949 24855 -25915
rect 24889 -25949 24922 -25915
rect 24822 -25983 24922 -25949
rect 24822 -26017 24855 -25983
rect 24889 -26017 24922 -25983
rect 24822 -26051 24922 -26017
rect 24822 -26085 24855 -26051
rect 24889 -26085 24922 -26051
rect 24822 -26119 24922 -26085
rect 24822 -26153 24855 -26119
rect 24889 -26153 24922 -26119
rect 24822 -26187 24922 -26153
rect 24822 -26221 24855 -26187
rect 24889 -26221 24922 -26187
rect 24822 -26255 24922 -26221
rect 24822 -26289 24855 -26255
rect 24889 -26289 24922 -26255
rect 24822 -26323 24922 -26289
rect 24822 -26357 24855 -26323
rect 24889 -26357 24922 -26323
rect 24822 -26391 24922 -26357
rect 24822 -26425 24855 -26391
rect 24889 -26425 24922 -26391
rect 24822 -26459 24922 -26425
rect 24822 -26493 24855 -26459
rect 24889 -26493 24922 -26459
rect 24822 -26527 24922 -26493
rect 24822 -26561 24855 -26527
rect 24889 -26561 24922 -26527
rect 24822 -26595 24922 -26561
rect 24822 -26629 24855 -26595
rect 24889 -26629 24922 -26595
rect 24822 -26663 24922 -26629
rect 24822 -26697 24855 -26663
rect 24889 -26697 24922 -26663
rect 24822 -26731 24922 -26697
rect 24822 -26765 24855 -26731
rect 24889 -26765 24922 -26731
rect 24822 -26799 24922 -26765
rect 24822 -26833 24855 -26799
rect 24889 -26833 24922 -26799
rect 24822 -26867 24922 -26833
rect 24822 -26901 24855 -26867
rect 24889 -26901 24922 -26867
rect 24822 -26935 24922 -26901
rect 24822 -26969 24855 -26935
rect 24889 -26969 24922 -26935
rect 24822 -27003 24922 -26969
rect 24822 -27037 24855 -27003
rect 24889 -27037 24922 -27003
rect 24822 -27122 24922 -27037
rect -12322 -27155 24922 -27122
rect -12322 -27189 -12145 -27155
rect -12111 -27189 -12077 -27155
rect -12043 -27189 -12009 -27155
rect -11975 -27189 -11941 -27155
rect -11907 -27189 -11873 -27155
rect -11839 -27189 -11805 -27155
rect -11771 -27189 -11737 -27155
rect -11703 -27189 -11669 -27155
rect -11635 -27189 -11601 -27155
rect -11567 -27189 -11533 -27155
rect -11499 -27189 -11465 -27155
rect -11431 -27189 -11397 -27155
rect -11363 -27189 -11329 -27155
rect -11295 -27189 -11261 -27155
rect -11227 -27189 -11193 -27155
rect -11159 -27189 -11125 -27155
rect -11091 -27189 -11057 -27155
rect -11023 -27189 -10989 -27155
rect -10955 -27189 -10921 -27155
rect -10887 -27189 -10853 -27155
rect -10819 -27189 -10785 -27155
rect -10751 -27189 -10717 -27155
rect -10683 -27189 -10649 -27155
rect -10615 -27189 -10581 -27155
rect -10547 -27189 -10513 -27155
rect -10479 -27189 -10445 -27155
rect -10411 -27189 -10377 -27155
rect -10343 -27189 -10309 -27155
rect -10275 -27189 -10241 -27155
rect -10207 -27189 -10173 -27155
rect -10139 -27189 -10105 -27155
rect -10071 -27189 -10037 -27155
rect -10003 -27189 -9969 -27155
rect -9935 -27189 -9901 -27155
rect -9867 -27189 -9833 -27155
rect -9799 -27189 -9765 -27155
rect -9731 -27189 -9697 -27155
rect -9663 -27189 -9629 -27155
rect -9595 -27189 -9561 -27155
rect -9527 -27189 -9493 -27155
rect -9459 -27189 -9425 -27155
rect -9391 -27189 -9357 -27155
rect -9323 -27189 -9289 -27155
rect -9255 -27189 -9221 -27155
rect -9187 -27189 -9153 -27155
rect -9119 -27189 -9085 -27155
rect -9051 -27189 -9017 -27155
rect -8983 -27189 -8949 -27155
rect -8915 -27189 -8881 -27155
rect -8847 -27189 -8813 -27155
rect -8779 -27189 -8745 -27155
rect -8711 -27189 -8677 -27155
rect -8643 -27189 -8609 -27155
rect -8575 -27189 -8541 -27155
rect -8507 -27189 -8473 -27155
rect -8439 -27189 -8405 -27155
rect -8371 -27189 -8337 -27155
rect -8303 -27189 -8269 -27155
rect -8235 -27189 -8201 -27155
rect -8167 -27189 -8133 -27155
rect -8099 -27189 -8065 -27155
rect -8031 -27189 -7997 -27155
rect -7963 -27189 -7929 -27155
rect -7895 -27189 -7861 -27155
rect -7827 -27189 -7793 -27155
rect -7759 -27189 -7725 -27155
rect -7691 -27189 -7657 -27155
rect -7623 -27189 -7589 -27155
rect -7555 -27189 -7521 -27155
rect -7487 -27189 -7453 -27155
rect -7419 -27189 -7385 -27155
rect -7351 -27189 -7317 -27155
rect -7283 -27189 -7249 -27155
rect -7215 -27189 -7181 -27155
rect -7147 -27189 -7113 -27155
rect -7079 -27189 -7045 -27155
rect -7011 -27189 -6977 -27155
rect -6943 -27189 -6909 -27155
rect -6875 -27189 -6841 -27155
rect -6807 -27189 -6773 -27155
rect -6739 -27189 -6705 -27155
rect -6671 -27189 -6637 -27155
rect -6603 -27189 -6569 -27155
rect -6535 -27189 -6501 -27155
rect -6467 -27189 -6433 -27155
rect -6399 -27189 -6365 -27155
rect -6331 -27189 -6297 -27155
rect -6263 -27189 -6229 -27155
rect -6195 -27189 -6161 -27155
rect -6127 -27189 -6093 -27155
rect -6059 -27189 -6025 -27155
rect -5991 -27189 -5957 -27155
rect -5923 -27189 -5889 -27155
rect -5855 -27189 -5821 -27155
rect -5787 -27189 -5753 -27155
rect -5719 -27189 -5685 -27155
rect -5651 -27189 -5617 -27155
rect -5583 -27189 -5549 -27155
rect -5515 -27189 -5481 -27155
rect -5447 -27189 -5413 -27155
rect -5379 -27189 -5345 -27155
rect -5311 -27189 -5277 -27155
rect -5243 -27189 -5209 -27155
rect -5175 -27189 -5141 -27155
rect -5107 -27189 -5073 -27155
rect -5039 -27189 -5005 -27155
rect -4971 -27189 -4937 -27155
rect -4903 -27189 -4869 -27155
rect -4835 -27189 -4801 -27155
rect -4767 -27189 -4733 -27155
rect -4699 -27189 -4665 -27155
rect -4631 -27189 -4597 -27155
rect -4563 -27189 -4529 -27155
rect -4495 -27189 -4461 -27155
rect -4427 -27189 -4393 -27155
rect -4359 -27189 -4325 -27155
rect -4291 -27189 -4257 -27155
rect -4223 -27189 -4189 -27155
rect -4155 -27189 -4121 -27155
rect -4087 -27189 -4053 -27155
rect -4019 -27189 -3985 -27155
rect -3951 -27189 -3917 -27155
rect -3883 -27189 -3849 -27155
rect -3815 -27189 -3781 -27155
rect -3747 -27189 -3713 -27155
rect -3679 -27189 -3645 -27155
rect -3611 -27189 -3577 -27155
rect -3543 -27189 -3509 -27155
rect -3475 -27189 -3441 -27155
rect -3407 -27189 -3373 -27155
rect -3339 -27189 -3305 -27155
rect -3271 -27189 -3237 -27155
rect -3203 -27189 -3169 -27155
rect -3135 -27189 -3101 -27155
rect -3067 -27189 -3033 -27155
rect -2999 -27189 -2965 -27155
rect -2931 -27189 -2897 -27155
rect -2863 -27189 -2829 -27155
rect -2795 -27189 -2761 -27155
rect -2727 -27189 -2693 -27155
rect -2659 -27189 -2625 -27155
rect -2591 -27189 -2557 -27155
rect -2523 -27189 -2489 -27155
rect -2455 -27189 -2421 -27155
rect -2387 -27189 -2353 -27155
rect -2319 -27189 -2285 -27155
rect -2251 -27189 -2217 -27155
rect -2183 -27189 -2149 -27155
rect -2115 -27189 -2081 -27155
rect -2047 -27189 -2013 -27155
rect -1979 -27189 -1945 -27155
rect -1911 -27189 -1877 -27155
rect -1843 -27189 -1809 -27155
rect -1775 -27189 -1741 -27155
rect -1707 -27189 -1673 -27155
rect -1639 -27189 -1605 -27155
rect -1571 -27189 -1537 -27155
rect -1503 -27189 -1469 -27155
rect -1435 -27189 -1401 -27155
rect -1367 -27189 -1333 -27155
rect -1299 -27189 -1265 -27155
rect -1231 -27189 -1197 -27155
rect -1163 -27189 -1129 -27155
rect -1095 -27189 -1061 -27155
rect -1027 -27189 -993 -27155
rect -959 -27189 -925 -27155
rect -891 -27189 -857 -27155
rect -823 -27189 -789 -27155
rect -755 -27189 -721 -27155
rect -687 -27189 -653 -27155
rect -619 -27189 -585 -27155
rect -551 -27189 -517 -27155
rect -483 -27189 -449 -27155
rect -415 -27189 -381 -27155
rect -347 -27189 -313 -27155
rect -279 -27189 -245 -27155
rect -211 -27189 -177 -27155
rect -143 -27189 -109 -27155
rect -75 -27189 -41 -27155
rect -7 -27189 27 -27155
rect 61 -27189 95 -27155
rect 129 -27189 163 -27155
rect 197 -27189 231 -27155
rect 265 -27189 299 -27155
rect 333 -27189 367 -27155
rect 401 -27189 435 -27155
rect 469 -27189 503 -27155
rect 537 -27189 571 -27155
rect 605 -27189 639 -27155
rect 673 -27189 707 -27155
rect 741 -27189 775 -27155
rect 809 -27189 843 -27155
rect 877 -27189 911 -27155
rect 945 -27189 979 -27155
rect 1013 -27189 1047 -27155
rect 1081 -27189 1115 -27155
rect 1149 -27189 1183 -27155
rect 1217 -27189 1251 -27155
rect 1285 -27189 1319 -27155
rect 1353 -27189 1387 -27155
rect 1421 -27189 1455 -27155
rect 1489 -27189 1523 -27155
rect 1557 -27189 1591 -27155
rect 1625 -27189 1659 -27155
rect 1693 -27189 1727 -27155
rect 1761 -27189 1795 -27155
rect 1829 -27189 1863 -27155
rect 1897 -27189 1931 -27155
rect 1965 -27189 1999 -27155
rect 2033 -27189 2067 -27155
rect 2101 -27189 2135 -27155
rect 2169 -27189 2203 -27155
rect 2237 -27189 2271 -27155
rect 2305 -27189 2339 -27155
rect 2373 -27189 2407 -27155
rect 2441 -27189 2475 -27155
rect 2509 -27189 2543 -27155
rect 2577 -27189 2611 -27155
rect 2645 -27189 2679 -27155
rect 2713 -27189 2747 -27155
rect 2781 -27189 2815 -27155
rect 2849 -27189 2883 -27155
rect 2917 -27189 2951 -27155
rect 2985 -27189 3019 -27155
rect 3053 -27189 3087 -27155
rect 3121 -27189 3155 -27155
rect 3189 -27189 3223 -27155
rect 3257 -27189 3291 -27155
rect 3325 -27189 3359 -27155
rect 3393 -27189 3427 -27155
rect 3461 -27189 3495 -27155
rect 3529 -27189 3563 -27155
rect 3597 -27189 3631 -27155
rect 3665 -27189 3699 -27155
rect 3733 -27189 3767 -27155
rect 3801 -27189 3835 -27155
rect 3869 -27189 3903 -27155
rect 3937 -27189 3971 -27155
rect 4005 -27189 4039 -27155
rect 4073 -27189 4107 -27155
rect 4141 -27189 4175 -27155
rect 4209 -27189 4243 -27155
rect 4277 -27189 4311 -27155
rect 4345 -27189 4379 -27155
rect 4413 -27189 4447 -27155
rect 4481 -27189 4515 -27155
rect 4549 -27189 4583 -27155
rect 4617 -27189 4651 -27155
rect 4685 -27189 4719 -27155
rect 4753 -27189 4787 -27155
rect 4821 -27189 4855 -27155
rect 4889 -27189 4923 -27155
rect 4957 -27189 4991 -27155
rect 5025 -27189 5059 -27155
rect 5093 -27189 5127 -27155
rect 5161 -27189 5195 -27155
rect 5229 -27189 5263 -27155
rect 5297 -27189 5331 -27155
rect 5365 -27189 5399 -27155
rect 5433 -27189 5467 -27155
rect 5501 -27189 5535 -27155
rect 5569 -27189 5603 -27155
rect 5637 -27189 5671 -27155
rect 5705 -27189 5739 -27155
rect 5773 -27189 5807 -27155
rect 5841 -27189 5875 -27155
rect 5909 -27189 5943 -27155
rect 5977 -27189 6011 -27155
rect 6045 -27189 6079 -27155
rect 6113 -27189 6147 -27155
rect 6181 -27189 6215 -27155
rect 6249 -27189 6283 -27155
rect 6317 -27189 6351 -27155
rect 6385 -27189 6419 -27155
rect 6453 -27189 6487 -27155
rect 6521 -27189 6555 -27155
rect 6589 -27189 6623 -27155
rect 6657 -27189 6691 -27155
rect 6725 -27189 6759 -27155
rect 6793 -27189 6827 -27155
rect 6861 -27189 6895 -27155
rect 6929 -27189 6963 -27155
rect 6997 -27189 7031 -27155
rect 7065 -27189 7099 -27155
rect 7133 -27189 7167 -27155
rect 7201 -27189 7235 -27155
rect 7269 -27189 7303 -27155
rect 7337 -27189 7371 -27155
rect 7405 -27189 7439 -27155
rect 7473 -27189 7507 -27155
rect 7541 -27189 7575 -27155
rect 7609 -27189 7643 -27155
rect 7677 -27189 7711 -27155
rect 7745 -27189 7779 -27155
rect 7813 -27189 7847 -27155
rect 7881 -27189 7915 -27155
rect 7949 -27189 7983 -27155
rect 8017 -27189 8051 -27155
rect 8085 -27189 8119 -27155
rect 8153 -27189 8187 -27155
rect 8221 -27189 8255 -27155
rect 8289 -27189 8323 -27155
rect 8357 -27189 8391 -27155
rect 8425 -27189 8459 -27155
rect 8493 -27189 8527 -27155
rect 8561 -27189 8595 -27155
rect 8629 -27189 8663 -27155
rect 8697 -27189 8731 -27155
rect 8765 -27189 8799 -27155
rect 8833 -27189 8867 -27155
rect 8901 -27189 8935 -27155
rect 8969 -27189 9003 -27155
rect 9037 -27189 9071 -27155
rect 9105 -27189 9139 -27155
rect 9173 -27189 9207 -27155
rect 9241 -27189 9275 -27155
rect 9309 -27189 9343 -27155
rect 9377 -27189 9411 -27155
rect 9445 -27189 9479 -27155
rect 9513 -27189 9547 -27155
rect 9581 -27189 9615 -27155
rect 9649 -27189 9683 -27155
rect 9717 -27189 9751 -27155
rect 9785 -27189 9819 -27155
rect 9853 -27189 9887 -27155
rect 9921 -27189 9955 -27155
rect 9989 -27189 10023 -27155
rect 10057 -27189 10091 -27155
rect 10125 -27189 10159 -27155
rect 10193 -27189 10227 -27155
rect 10261 -27189 10295 -27155
rect 10329 -27189 10363 -27155
rect 10397 -27189 10431 -27155
rect 10465 -27189 10499 -27155
rect 10533 -27189 10567 -27155
rect 10601 -27189 10635 -27155
rect 10669 -27189 10703 -27155
rect 10737 -27189 10771 -27155
rect 10805 -27189 10839 -27155
rect 10873 -27189 10907 -27155
rect 10941 -27189 10975 -27155
rect 11009 -27189 11043 -27155
rect 11077 -27189 11111 -27155
rect 11145 -27189 11179 -27155
rect 11213 -27189 11247 -27155
rect 11281 -27189 11315 -27155
rect 11349 -27189 11383 -27155
rect 11417 -27189 11451 -27155
rect 11485 -27189 11519 -27155
rect 11553 -27189 11587 -27155
rect 11621 -27189 11655 -27155
rect 11689 -27189 11723 -27155
rect 11757 -27189 11791 -27155
rect 11825 -27189 11859 -27155
rect 11893 -27189 11927 -27155
rect 11961 -27189 11995 -27155
rect 12029 -27189 12063 -27155
rect 12097 -27189 12131 -27155
rect 12165 -27189 12199 -27155
rect 12233 -27189 12267 -27155
rect 12301 -27189 12335 -27155
rect 12369 -27189 12403 -27155
rect 12437 -27189 12471 -27155
rect 12505 -27189 12539 -27155
rect 12573 -27189 12607 -27155
rect 12641 -27189 12675 -27155
rect 12709 -27189 12743 -27155
rect 12777 -27189 12811 -27155
rect 12845 -27189 12879 -27155
rect 12913 -27189 12947 -27155
rect 12981 -27189 13015 -27155
rect 13049 -27189 13083 -27155
rect 13117 -27189 13151 -27155
rect 13185 -27189 13219 -27155
rect 13253 -27189 13287 -27155
rect 13321 -27189 13355 -27155
rect 13389 -27189 13423 -27155
rect 13457 -27189 13491 -27155
rect 13525 -27189 13559 -27155
rect 13593 -27189 13627 -27155
rect 13661 -27189 13695 -27155
rect 13729 -27189 13763 -27155
rect 13797 -27189 13831 -27155
rect 13865 -27189 13899 -27155
rect 13933 -27189 13967 -27155
rect 14001 -27189 14035 -27155
rect 14069 -27189 14103 -27155
rect 14137 -27189 14171 -27155
rect 14205 -27189 14239 -27155
rect 14273 -27189 14307 -27155
rect 14341 -27189 14375 -27155
rect 14409 -27189 14443 -27155
rect 14477 -27189 14511 -27155
rect 14545 -27189 14579 -27155
rect 14613 -27189 14647 -27155
rect 14681 -27189 14715 -27155
rect 14749 -27189 14783 -27155
rect 14817 -27189 14851 -27155
rect 14885 -27189 14919 -27155
rect 14953 -27189 14987 -27155
rect 15021 -27189 15055 -27155
rect 15089 -27189 15123 -27155
rect 15157 -27189 15191 -27155
rect 15225 -27189 15259 -27155
rect 15293 -27189 15327 -27155
rect 15361 -27189 15395 -27155
rect 15429 -27189 15463 -27155
rect 15497 -27189 15531 -27155
rect 15565 -27189 15599 -27155
rect 15633 -27189 15667 -27155
rect 15701 -27189 15735 -27155
rect 15769 -27189 15803 -27155
rect 15837 -27189 15871 -27155
rect 15905 -27189 15939 -27155
rect 15973 -27189 16007 -27155
rect 16041 -27189 16075 -27155
rect 16109 -27189 16143 -27155
rect 16177 -27189 16211 -27155
rect 16245 -27189 16279 -27155
rect 16313 -27189 16347 -27155
rect 16381 -27189 16415 -27155
rect 16449 -27189 16483 -27155
rect 16517 -27189 16551 -27155
rect 16585 -27189 16619 -27155
rect 16653 -27189 16687 -27155
rect 16721 -27189 16755 -27155
rect 16789 -27189 16823 -27155
rect 16857 -27189 16891 -27155
rect 16925 -27189 16959 -27155
rect 16993 -27189 17027 -27155
rect 17061 -27189 17095 -27155
rect 17129 -27189 17163 -27155
rect 17197 -27189 17231 -27155
rect 17265 -27189 17299 -27155
rect 17333 -27189 17367 -27155
rect 17401 -27189 17435 -27155
rect 17469 -27189 17503 -27155
rect 17537 -27189 17571 -27155
rect 17605 -27189 17639 -27155
rect 17673 -27189 17707 -27155
rect 17741 -27189 17775 -27155
rect 17809 -27189 17843 -27155
rect 17877 -27189 17911 -27155
rect 17945 -27189 17979 -27155
rect 18013 -27189 18047 -27155
rect 18081 -27189 18115 -27155
rect 18149 -27189 18183 -27155
rect 18217 -27189 18251 -27155
rect 18285 -27189 18319 -27155
rect 18353 -27189 18387 -27155
rect 18421 -27189 18455 -27155
rect 18489 -27189 18523 -27155
rect 18557 -27189 18591 -27155
rect 18625 -27189 18659 -27155
rect 18693 -27189 18727 -27155
rect 18761 -27189 18795 -27155
rect 18829 -27189 18863 -27155
rect 18897 -27189 18931 -27155
rect 18965 -27189 18999 -27155
rect 19033 -27189 19067 -27155
rect 19101 -27189 19135 -27155
rect 19169 -27189 19203 -27155
rect 19237 -27189 19271 -27155
rect 19305 -27189 19339 -27155
rect 19373 -27189 19407 -27155
rect 19441 -27189 19475 -27155
rect 19509 -27189 19543 -27155
rect 19577 -27189 19611 -27155
rect 19645 -27189 19679 -27155
rect 19713 -27189 19747 -27155
rect 19781 -27189 19815 -27155
rect 19849 -27189 19883 -27155
rect 19917 -27189 19951 -27155
rect 19985 -27189 20019 -27155
rect 20053 -27189 20087 -27155
rect 20121 -27189 20155 -27155
rect 20189 -27189 20223 -27155
rect 20257 -27189 20291 -27155
rect 20325 -27189 20359 -27155
rect 20393 -27189 20427 -27155
rect 20461 -27189 20495 -27155
rect 20529 -27189 20563 -27155
rect 20597 -27189 20631 -27155
rect 20665 -27189 20699 -27155
rect 20733 -27189 20767 -27155
rect 20801 -27189 20835 -27155
rect 20869 -27189 20903 -27155
rect 20937 -27189 20971 -27155
rect 21005 -27189 21039 -27155
rect 21073 -27189 21107 -27155
rect 21141 -27189 21175 -27155
rect 21209 -27189 21243 -27155
rect 21277 -27189 21311 -27155
rect 21345 -27189 21379 -27155
rect 21413 -27189 21447 -27155
rect 21481 -27189 21515 -27155
rect 21549 -27189 21583 -27155
rect 21617 -27189 21651 -27155
rect 21685 -27189 21719 -27155
rect 21753 -27189 21787 -27155
rect 21821 -27189 21855 -27155
rect 21889 -27189 21923 -27155
rect 21957 -27189 21991 -27155
rect 22025 -27189 22059 -27155
rect 22093 -27189 22127 -27155
rect 22161 -27189 22195 -27155
rect 22229 -27189 22263 -27155
rect 22297 -27189 22331 -27155
rect 22365 -27189 22399 -27155
rect 22433 -27189 22467 -27155
rect 22501 -27189 22535 -27155
rect 22569 -27189 22603 -27155
rect 22637 -27189 22671 -27155
rect 22705 -27189 22739 -27155
rect 22773 -27189 22807 -27155
rect 22841 -27189 22875 -27155
rect 22909 -27189 22943 -27155
rect 22977 -27189 23011 -27155
rect 23045 -27189 23079 -27155
rect 23113 -27189 23147 -27155
rect 23181 -27189 23215 -27155
rect 23249 -27189 23283 -27155
rect 23317 -27189 23351 -27155
rect 23385 -27189 23419 -27155
rect 23453 -27189 23487 -27155
rect 23521 -27189 23555 -27155
rect 23589 -27189 23623 -27155
rect 23657 -27189 23691 -27155
rect 23725 -27189 23759 -27155
rect 23793 -27189 23827 -27155
rect 23861 -27189 23895 -27155
rect 23929 -27189 23963 -27155
rect 23997 -27189 24031 -27155
rect 24065 -27189 24099 -27155
rect 24133 -27189 24167 -27155
rect 24201 -27189 24235 -27155
rect 24269 -27189 24303 -27155
rect 24337 -27189 24371 -27155
rect 24405 -27189 24439 -27155
rect 24473 -27189 24507 -27155
rect 24541 -27189 24575 -27155
rect 24609 -27189 24643 -27155
rect 24677 -27189 24711 -27155
rect 24745 -27189 24922 -27155
rect -12322 -27222 24922 -27189
<< nsubdiff >>
rect 378 4289 24822 4322
rect 378 4255 547 4289
rect 581 4255 615 4289
rect 649 4255 683 4289
rect 717 4255 751 4289
rect 785 4255 819 4289
rect 853 4255 887 4289
rect 921 4255 955 4289
rect 989 4255 1023 4289
rect 1057 4255 1091 4289
rect 1125 4255 1159 4289
rect 1193 4255 1227 4289
rect 1261 4255 1295 4289
rect 1329 4255 1363 4289
rect 1397 4255 1431 4289
rect 1465 4255 1499 4289
rect 1533 4255 1567 4289
rect 1601 4255 1635 4289
rect 1669 4255 1703 4289
rect 1737 4255 1771 4289
rect 1805 4255 1839 4289
rect 1873 4255 1907 4289
rect 1941 4255 1975 4289
rect 2009 4255 2043 4289
rect 2077 4255 2111 4289
rect 2145 4255 2179 4289
rect 2213 4255 2247 4289
rect 2281 4255 2315 4289
rect 2349 4255 2383 4289
rect 2417 4255 2451 4289
rect 2485 4255 2519 4289
rect 2553 4255 2587 4289
rect 2621 4255 2655 4289
rect 2689 4255 2723 4289
rect 2757 4255 2791 4289
rect 2825 4255 2859 4289
rect 2893 4255 2927 4289
rect 2961 4255 2995 4289
rect 3029 4255 3063 4289
rect 3097 4255 3131 4289
rect 3165 4255 3199 4289
rect 3233 4255 3267 4289
rect 3301 4255 3335 4289
rect 3369 4255 3403 4289
rect 3437 4255 3471 4289
rect 3505 4255 3539 4289
rect 3573 4255 3607 4289
rect 3641 4255 3675 4289
rect 3709 4255 3743 4289
rect 3777 4255 3811 4289
rect 3845 4255 3879 4289
rect 3913 4255 3947 4289
rect 3981 4255 4015 4289
rect 4049 4255 4083 4289
rect 4117 4255 4151 4289
rect 4185 4255 4219 4289
rect 4253 4255 4287 4289
rect 4321 4255 4355 4289
rect 4389 4255 4423 4289
rect 4457 4255 4491 4289
rect 4525 4255 4559 4289
rect 4593 4255 4627 4289
rect 4661 4255 4695 4289
rect 4729 4255 4763 4289
rect 4797 4255 4831 4289
rect 4865 4255 4899 4289
rect 4933 4255 4967 4289
rect 5001 4255 5035 4289
rect 5069 4255 5103 4289
rect 5137 4255 5171 4289
rect 5205 4255 5239 4289
rect 5273 4255 5307 4289
rect 5341 4255 5375 4289
rect 5409 4255 5443 4289
rect 5477 4255 5511 4289
rect 5545 4255 5579 4289
rect 5613 4255 5647 4289
rect 5681 4255 5715 4289
rect 5749 4255 5783 4289
rect 5817 4255 5851 4289
rect 5885 4255 5919 4289
rect 5953 4255 5987 4289
rect 6021 4255 6055 4289
rect 6089 4255 6123 4289
rect 6157 4255 6191 4289
rect 6225 4255 6259 4289
rect 6293 4255 6327 4289
rect 6361 4255 6395 4289
rect 6429 4255 6463 4289
rect 6497 4255 6531 4289
rect 6565 4255 6599 4289
rect 6633 4255 6667 4289
rect 6701 4255 6735 4289
rect 6769 4255 6803 4289
rect 6837 4255 6871 4289
rect 6905 4255 6939 4289
rect 6973 4255 7007 4289
rect 7041 4255 7075 4289
rect 7109 4255 7143 4289
rect 7177 4255 7211 4289
rect 7245 4255 7279 4289
rect 7313 4255 7347 4289
rect 7381 4255 7415 4289
rect 7449 4255 7483 4289
rect 7517 4255 7551 4289
rect 7585 4255 7619 4289
rect 7653 4255 7687 4289
rect 7721 4255 7755 4289
rect 7789 4255 7823 4289
rect 7857 4255 7891 4289
rect 7925 4255 7959 4289
rect 7993 4255 8027 4289
rect 8061 4255 8095 4289
rect 8129 4255 8163 4289
rect 8197 4255 8231 4289
rect 8265 4255 8299 4289
rect 8333 4255 8367 4289
rect 8401 4255 8435 4289
rect 8469 4255 8503 4289
rect 8537 4255 8571 4289
rect 8605 4255 8639 4289
rect 8673 4255 8707 4289
rect 8741 4255 8775 4289
rect 8809 4255 8843 4289
rect 8877 4255 8911 4289
rect 8945 4255 8979 4289
rect 9013 4255 9047 4289
rect 9081 4255 9115 4289
rect 9149 4255 9183 4289
rect 9217 4255 9251 4289
rect 9285 4255 9319 4289
rect 9353 4255 9387 4289
rect 9421 4255 9455 4289
rect 9489 4255 9523 4289
rect 9557 4255 9591 4289
rect 9625 4255 9659 4289
rect 9693 4255 9727 4289
rect 9761 4255 9795 4289
rect 9829 4255 9863 4289
rect 9897 4255 9931 4289
rect 9965 4255 9999 4289
rect 10033 4255 10067 4289
rect 10101 4255 10135 4289
rect 10169 4255 10203 4289
rect 10237 4255 10271 4289
rect 10305 4255 10339 4289
rect 10373 4255 10407 4289
rect 10441 4255 10475 4289
rect 10509 4255 10543 4289
rect 10577 4255 10611 4289
rect 10645 4255 10679 4289
rect 10713 4255 10747 4289
rect 10781 4255 10815 4289
rect 10849 4255 10883 4289
rect 10917 4255 10951 4289
rect 10985 4255 11019 4289
rect 11053 4255 11087 4289
rect 11121 4255 11155 4289
rect 11189 4255 11223 4289
rect 11257 4255 11291 4289
rect 11325 4255 11359 4289
rect 11393 4255 11427 4289
rect 11461 4255 11495 4289
rect 11529 4255 11563 4289
rect 11597 4255 11631 4289
rect 11665 4255 11699 4289
rect 11733 4255 11767 4289
rect 11801 4255 11835 4289
rect 11869 4255 11903 4289
rect 11937 4255 11971 4289
rect 12005 4255 12039 4289
rect 12073 4255 12107 4289
rect 12141 4255 12175 4289
rect 12209 4255 12243 4289
rect 12277 4255 12311 4289
rect 12345 4255 12379 4289
rect 12413 4255 12447 4289
rect 12481 4255 12515 4289
rect 12549 4255 12583 4289
rect 12617 4255 12651 4289
rect 12685 4255 12719 4289
rect 12753 4255 12787 4289
rect 12821 4255 12855 4289
rect 12889 4255 12923 4289
rect 12957 4255 12991 4289
rect 13025 4255 13059 4289
rect 13093 4255 13127 4289
rect 13161 4255 13195 4289
rect 13229 4255 13263 4289
rect 13297 4255 13331 4289
rect 13365 4255 13399 4289
rect 13433 4255 13467 4289
rect 13501 4255 13535 4289
rect 13569 4255 13603 4289
rect 13637 4255 13671 4289
rect 13705 4255 13739 4289
rect 13773 4255 13807 4289
rect 13841 4255 13875 4289
rect 13909 4255 13943 4289
rect 13977 4255 14011 4289
rect 14045 4255 14079 4289
rect 14113 4255 14147 4289
rect 14181 4255 14215 4289
rect 14249 4255 14283 4289
rect 14317 4255 14351 4289
rect 14385 4255 14419 4289
rect 14453 4255 14487 4289
rect 14521 4255 14555 4289
rect 14589 4255 14623 4289
rect 14657 4255 14691 4289
rect 14725 4255 14759 4289
rect 14793 4255 14827 4289
rect 14861 4255 14895 4289
rect 14929 4255 14963 4289
rect 14997 4255 15031 4289
rect 15065 4255 15099 4289
rect 15133 4255 15167 4289
rect 15201 4255 15235 4289
rect 15269 4255 15303 4289
rect 15337 4255 15371 4289
rect 15405 4255 15439 4289
rect 15473 4255 15507 4289
rect 15541 4255 15575 4289
rect 15609 4255 15643 4289
rect 15677 4255 15711 4289
rect 15745 4255 15779 4289
rect 15813 4255 15847 4289
rect 15881 4255 15915 4289
rect 15949 4255 15983 4289
rect 16017 4255 16051 4289
rect 16085 4255 16119 4289
rect 16153 4255 16187 4289
rect 16221 4255 16255 4289
rect 16289 4255 16323 4289
rect 16357 4255 16391 4289
rect 16425 4255 16459 4289
rect 16493 4255 16527 4289
rect 16561 4255 16595 4289
rect 16629 4255 16663 4289
rect 16697 4255 16731 4289
rect 16765 4255 16799 4289
rect 16833 4255 16867 4289
rect 16901 4255 16935 4289
rect 16969 4255 17003 4289
rect 17037 4255 17071 4289
rect 17105 4255 17139 4289
rect 17173 4255 17207 4289
rect 17241 4255 17275 4289
rect 17309 4255 17343 4289
rect 17377 4255 17411 4289
rect 17445 4255 17479 4289
rect 17513 4255 17547 4289
rect 17581 4255 17615 4289
rect 17649 4255 17683 4289
rect 17717 4255 17751 4289
rect 17785 4255 17819 4289
rect 17853 4255 17887 4289
rect 17921 4255 17955 4289
rect 17989 4255 18023 4289
rect 18057 4255 18091 4289
rect 18125 4255 18159 4289
rect 18193 4255 18227 4289
rect 18261 4255 18295 4289
rect 18329 4255 18363 4289
rect 18397 4255 18431 4289
rect 18465 4255 18499 4289
rect 18533 4255 18567 4289
rect 18601 4255 18635 4289
rect 18669 4255 18703 4289
rect 18737 4255 18771 4289
rect 18805 4255 18839 4289
rect 18873 4255 18907 4289
rect 18941 4255 18975 4289
rect 19009 4255 19043 4289
rect 19077 4255 19111 4289
rect 19145 4255 19179 4289
rect 19213 4255 19247 4289
rect 19281 4255 19315 4289
rect 19349 4255 19383 4289
rect 19417 4255 19451 4289
rect 19485 4255 19519 4289
rect 19553 4255 19587 4289
rect 19621 4255 19655 4289
rect 19689 4255 19723 4289
rect 19757 4255 19791 4289
rect 19825 4255 19859 4289
rect 19893 4255 19927 4289
rect 19961 4255 19995 4289
rect 20029 4255 20063 4289
rect 20097 4255 20131 4289
rect 20165 4255 20199 4289
rect 20233 4255 20267 4289
rect 20301 4255 20335 4289
rect 20369 4255 20403 4289
rect 20437 4255 20471 4289
rect 20505 4255 20539 4289
rect 20573 4255 20607 4289
rect 20641 4255 20675 4289
rect 20709 4255 20743 4289
rect 20777 4255 20811 4289
rect 20845 4255 20879 4289
rect 20913 4255 20947 4289
rect 20981 4255 21015 4289
rect 21049 4255 21083 4289
rect 21117 4255 21151 4289
rect 21185 4255 21219 4289
rect 21253 4255 21287 4289
rect 21321 4255 21355 4289
rect 21389 4255 21423 4289
rect 21457 4255 21491 4289
rect 21525 4255 21559 4289
rect 21593 4255 21627 4289
rect 21661 4255 21695 4289
rect 21729 4255 21763 4289
rect 21797 4255 21831 4289
rect 21865 4255 21899 4289
rect 21933 4255 21967 4289
rect 22001 4255 22035 4289
rect 22069 4255 22103 4289
rect 22137 4255 22171 4289
rect 22205 4255 22239 4289
rect 22273 4255 22307 4289
rect 22341 4255 22375 4289
rect 22409 4255 22443 4289
rect 22477 4255 22511 4289
rect 22545 4255 22579 4289
rect 22613 4255 22647 4289
rect 22681 4255 22715 4289
rect 22749 4255 22783 4289
rect 22817 4255 22851 4289
rect 22885 4255 22919 4289
rect 22953 4255 22987 4289
rect 23021 4255 23055 4289
rect 23089 4255 23123 4289
rect 23157 4255 23191 4289
rect 23225 4255 23259 4289
rect 23293 4255 23327 4289
rect 23361 4255 23395 4289
rect 23429 4255 23463 4289
rect 23497 4255 23531 4289
rect 23565 4255 23599 4289
rect 23633 4255 23667 4289
rect 23701 4255 23735 4289
rect 23769 4255 23803 4289
rect 23837 4255 23871 4289
rect 23905 4255 23939 4289
rect 23973 4255 24007 4289
rect 24041 4255 24075 4289
rect 24109 4255 24143 4289
rect 24177 4255 24211 4289
rect 24245 4255 24279 4289
rect 24313 4255 24347 4289
rect 24381 4255 24415 4289
rect 24449 4255 24483 4289
rect 24517 4255 24551 4289
rect 24585 4255 24619 4289
rect 24653 4255 24822 4289
rect 378 4222 24822 4255
rect 378 4144 478 4222
rect 378 4110 411 4144
rect 445 4110 478 4144
rect 378 4076 478 4110
rect 378 4042 411 4076
rect 445 4042 478 4076
rect 378 4008 478 4042
rect 378 3974 411 4008
rect 445 3974 478 4008
rect 378 3940 478 3974
rect 378 3906 411 3940
rect 445 3906 478 3940
rect 378 3872 478 3906
rect 378 3838 411 3872
rect 445 3838 478 3872
rect 378 3804 478 3838
rect 378 3770 411 3804
rect 445 3770 478 3804
rect 378 3736 478 3770
rect 378 3702 411 3736
rect 445 3702 478 3736
rect 378 3668 478 3702
rect 378 3634 411 3668
rect 445 3634 478 3668
rect 378 3600 478 3634
rect 378 3566 411 3600
rect 445 3566 478 3600
rect 378 3532 478 3566
rect 378 3498 411 3532
rect 445 3498 478 3532
rect 378 3464 478 3498
rect 378 3430 411 3464
rect 445 3430 478 3464
rect 378 3396 478 3430
rect 378 3362 411 3396
rect 445 3362 478 3396
rect 378 3328 478 3362
rect 378 3294 411 3328
rect 445 3294 478 3328
rect 378 3260 478 3294
rect 378 3226 411 3260
rect 445 3226 478 3260
rect 378 3192 478 3226
rect 378 3158 411 3192
rect 445 3158 478 3192
rect 378 3124 478 3158
rect 378 3090 411 3124
rect 445 3090 478 3124
rect 378 3056 478 3090
rect 378 3022 411 3056
rect 445 3022 478 3056
rect 378 2988 478 3022
rect 378 2954 411 2988
rect 445 2954 478 2988
rect 378 2920 478 2954
rect 378 2886 411 2920
rect 445 2886 478 2920
rect 378 2852 478 2886
rect 378 2818 411 2852
rect 445 2818 478 2852
rect 378 2784 478 2818
rect 378 2750 411 2784
rect 445 2750 478 2784
rect 378 2716 478 2750
rect 378 2682 411 2716
rect 445 2682 478 2716
rect 378 2648 478 2682
rect 378 2614 411 2648
rect 445 2614 478 2648
rect 378 2580 478 2614
rect 378 2546 411 2580
rect 445 2546 478 2580
rect 378 2512 478 2546
rect 378 2478 411 2512
rect 445 2478 478 2512
rect 378 2444 478 2478
rect 378 2410 411 2444
rect 445 2410 478 2444
rect 378 2376 478 2410
rect 378 2342 411 2376
rect 445 2342 478 2376
rect 378 2308 478 2342
rect 378 2274 411 2308
rect 445 2274 478 2308
rect 378 2240 478 2274
rect 378 2206 411 2240
rect 445 2206 478 2240
rect 378 2172 478 2206
rect 378 2138 411 2172
rect 445 2138 478 2172
rect 378 2104 478 2138
rect 378 2070 411 2104
rect 445 2070 478 2104
rect 378 2036 478 2070
rect 378 2002 411 2036
rect 445 2002 478 2036
rect 378 1968 478 2002
rect 378 1934 411 1968
rect 445 1934 478 1968
rect 378 1900 478 1934
rect 378 1866 411 1900
rect 445 1866 478 1900
rect 378 1832 478 1866
rect 378 1798 411 1832
rect 445 1798 478 1832
rect 378 1764 478 1798
rect 378 1730 411 1764
rect 445 1730 478 1764
rect 378 1696 478 1730
rect 378 1662 411 1696
rect 445 1662 478 1696
rect 378 1628 478 1662
rect 378 1594 411 1628
rect 445 1594 478 1628
rect 378 1560 478 1594
rect 378 1526 411 1560
rect 445 1526 478 1560
rect 378 1492 478 1526
rect 378 1458 411 1492
rect 445 1458 478 1492
rect 378 1424 478 1458
rect 378 1390 411 1424
rect 445 1390 478 1424
rect 378 1356 478 1390
rect 378 1322 411 1356
rect 445 1322 478 1356
rect 378 1288 478 1322
rect 378 1254 411 1288
rect 445 1254 478 1288
rect 378 1220 478 1254
rect 378 1186 411 1220
rect 445 1186 478 1220
rect 378 1152 478 1186
rect 378 1118 411 1152
rect 445 1118 478 1152
rect 378 1084 478 1118
rect 378 1050 411 1084
rect 445 1050 478 1084
rect 378 1016 478 1050
rect 378 982 411 1016
rect 445 982 478 1016
rect 378 948 478 982
rect 378 914 411 948
rect 445 914 478 948
rect 378 880 478 914
rect 378 846 411 880
rect 445 846 478 880
rect 378 812 478 846
rect 378 778 411 812
rect 445 778 478 812
rect 378 744 478 778
rect 378 710 411 744
rect 445 710 478 744
rect 378 676 478 710
rect 378 642 411 676
rect 445 642 478 676
rect 378 608 478 642
rect 378 574 411 608
rect 445 574 478 608
rect 378 540 478 574
rect 378 506 411 540
rect 445 506 478 540
rect 378 472 478 506
rect 378 438 411 472
rect 445 438 478 472
rect 378 404 478 438
rect 378 370 411 404
rect 445 370 478 404
rect 378 336 478 370
rect 378 302 411 336
rect 445 302 478 336
rect 378 268 478 302
rect 378 234 411 268
rect 445 234 478 268
rect 378 200 478 234
rect 378 166 411 200
rect 445 166 478 200
rect 378 132 478 166
rect 378 98 411 132
rect 445 98 478 132
rect 378 64 478 98
rect 378 30 411 64
rect 445 30 478 64
rect 378 -4 478 30
rect 378 -38 411 -4
rect 445 -38 478 -4
rect 378 -72 478 -38
rect 378 -106 411 -72
rect 445 -106 478 -72
rect 378 -140 478 -106
rect 378 -174 411 -140
rect 445 -174 478 -140
rect 378 -208 478 -174
rect 378 -242 411 -208
rect 445 -242 478 -208
rect 378 -276 478 -242
rect 378 -310 411 -276
rect 445 -310 478 -276
rect 378 -344 478 -310
rect 378 -378 411 -344
rect 445 -378 478 -344
rect 378 -412 478 -378
rect 378 -446 411 -412
rect 445 -446 478 -412
rect 378 -480 478 -446
rect 378 -514 411 -480
rect 445 -514 478 -480
rect 378 -548 478 -514
rect 378 -582 411 -548
rect 445 -582 478 -548
rect 378 -616 478 -582
rect 378 -650 411 -616
rect 445 -650 478 -616
rect 378 -684 478 -650
rect 378 -718 411 -684
rect 445 -718 478 -684
rect 378 -752 478 -718
rect 378 -786 411 -752
rect 445 -786 478 -752
rect 378 -820 478 -786
rect 378 -854 411 -820
rect 445 -854 478 -820
rect 378 -888 478 -854
rect 378 -922 411 -888
rect 445 -922 478 -888
rect 378 -956 478 -922
rect 378 -990 411 -956
rect 445 -990 478 -956
rect 378 -1024 478 -990
rect 378 -1058 411 -1024
rect 445 -1058 478 -1024
rect 378 -1092 478 -1058
rect 378 -1126 411 -1092
rect 445 -1126 478 -1092
rect 378 -1160 478 -1126
rect 378 -1194 411 -1160
rect 445 -1194 478 -1160
rect 378 -1228 478 -1194
rect 378 -1262 411 -1228
rect 445 -1262 478 -1228
rect 378 -1296 478 -1262
rect 378 -1330 411 -1296
rect 445 -1330 478 -1296
rect 378 -1364 478 -1330
rect 378 -1398 411 -1364
rect 445 -1398 478 -1364
rect 378 -1432 478 -1398
rect 378 -1466 411 -1432
rect 445 -1466 478 -1432
rect 378 -1500 478 -1466
rect 378 -1534 411 -1500
rect 445 -1534 478 -1500
rect 378 -1568 478 -1534
rect 378 -1602 411 -1568
rect 445 -1602 478 -1568
rect 378 -1636 478 -1602
rect 378 -1670 411 -1636
rect 445 -1670 478 -1636
rect 378 -1704 478 -1670
rect 378 -1738 411 -1704
rect 445 -1738 478 -1704
rect 378 -1772 478 -1738
rect 378 -1806 411 -1772
rect 445 -1806 478 -1772
rect 378 -1840 478 -1806
rect 378 -1874 411 -1840
rect 445 -1874 478 -1840
rect 378 -1908 478 -1874
rect 378 -1942 411 -1908
rect 445 -1942 478 -1908
rect 378 -1976 478 -1942
rect 378 -2010 411 -1976
rect 445 -2010 478 -1976
rect 378 -2044 478 -2010
rect 378 -2078 411 -2044
rect 445 -2078 478 -2044
rect 378 -2112 478 -2078
rect 378 -2146 411 -2112
rect 445 -2146 478 -2112
rect 378 -2180 478 -2146
rect 378 -2214 411 -2180
rect 445 -2214 478 -2180
rect 378 -2248 478 -2214
rect 378 -2282 411 -2248
rect 445 -2282 478 -2248
rect 378 -2316 478 -2282
rect 378 -2350 411 -2316
rect 445 -2350 478 -2316
rect 378 -2384 478 -2350
rect 378 -2418 411 -2384
rect 445 -2418 478 -2384
rect 378 -2452 478 -2418
rect 378 -2486 411 -2452
rect 445 -2486 478 -2452
rect 378 -2520 478 -2486
rect 378 -2554 411 -2520
rect 445 -2554 478 -2520
rect 378 -2588 478 -2554
rect 378 -2622 411 -2588
rect 445 -2622 478 -2588
rect 378 -2656 478 -2622
rect 378 -2690 411 -2656
rect 445 -2690 478 -2656
rect 378 -2724 478 -2690
rect 378 -2758 411 -2724
rect 445 -2758 478 -2724
rect 378 -2792 478 -2758
rect 378 -2826 411 -2792
rect 445 -2826 478 -2792
rect 378 -2860 478 -2826
rect 378 -2894 411 -2860
rect 445 -2894 478 -2860
rect 378 -2928 478 -2894
rect 378 -2962 411 -2928
rect 445 -2962 478 -2928
rect 378 -2996 478 -2962
rect 378 -3030 411 -2996
rect 445 -3030 478 -2996
rect 378 -3064 478 -3030
rect 378 -3098 411 -3064
rect 445 -3098 478 -3064
rect 378 -3132 478 -3098
rect 378 -3166 411 -3132
rect 445 -3166 478 -3132
rect 378 -3200 478 -3166
rect 378 -3234 411 -3200
rect 445 -3234 478 -3200
rect 378 -3268 478 -3234
rect 378 -3302 411 -3268
rect 445 -3302 478 -3268
rect 378 -3336 478 -3302
rect 378 -3370 411 -3336
rect 445 -3370 478 -3336
rect 378 -3404 478 -3370
rect 378 -3438 411 -3404
rect 445 -3438 478 -3404
rect 378 -3472 478 -3438
rect 378 -3506 411 -3472
rect 445 -3506 478 -3472
rect 378 -3540 478 -3506
rect 378 -3574 411 -3540
rect 445 -3574 478 -3540
rect 378 -3608 478 -3574
rect 378 -3642 411 -3608
rect 445 -3642 478 -3608
rect 378 -3676 478 -3642
rect 378 -3710 411 -3676
rect 445 -3710 478 -3676
rect 378 -3744 478 -3710
rect 378 -3778 411 -3744
rect 445 -3778 478 -3744
rect 378 -3812 478 -3778
rect 378 -3846 411 -3812
rect 445 -3846 478 -3812
rect 378 -3880 478 -3846
rect 378 -3914 411 -3880
rect 445 -3914 478 -3880
rect 378 -3948 478 -3914
rect 378 -3982 411 -3948
rect 445 -3982 478 -3948
rect 378 -4016 478 -3982
rect 378 -4050 411 -4016
rect 445 -4050 478 -4016
rect 378 -4084 478 -4050
rect 378 -4118 411 -4084
rect 445 -4118 478 -4084
rect 378 -4152 478 -4118
rect 378 -4186 411 -4152
rect 445 -4186 478 -4152
rect 378 -4220 478 -4186
rect 378 -4254 411 -4220
rect 445 -4254 478 -4220
rect 378 -4288 478 -4254
rect 378 -4322 411 -4288
rect 445 -4322 478 -4288
rect 378 -4356 478 -4322
rect 378 -4390 411 -4356
rect 445 -4390 478 -4356
rect 378 -4424 478 -4390
rect 378 -4458 411 -4424
rect 445 -4458 478 -4424
rect 378 -4492 478 -4458
rect 378 -4526 411 -4492
rect 445 -4526 478 -4492
rect 378 -4560 478 -4526
rect 378 -4594 411 -4560
rect 445 -4594 478 -4560
rect 378 -4628 478 -4594
rect 378 -4662 411 -4628
rect 445 -4662 478 -4628
rect 378 -4696 478 -4662
rect 378 -4730 411 -4696
rect 445 -4730 478 -4696
rect 378 -4764 478 -4730
rect 378 -4798 411 -4764
rect 445 -4798 478 -4764
rect 378 -4832 478 -4798
rect 378 -4866 411 -4832
rect 445 -4866 478 -4832
rect 378 -4900 478 -4866
rect 378 -4934 411 -4900
rect 445 -4934 478 -4900
rect 378 -4968 478 -4934
rect 378 -5002 411 -4968
rect 445 -5002 478 -4968
rect 378 -5036 478 -5002
rect 378 -5070 411 -5036
rect 445 -5070 478 -5036
rect 378 -5104 478 -5070
rect 378 -5138 411 -5104
rect 445 -5138 478 -5104
rect 378 -5172 478 -5138
rect 378 -5206 411 -5172
rect 445 -5206 478 -5172
rect 378 -5240 478 -5206
rect 378 -5274 411 -5240
rect 445 -5274 478 -5240
rect 378 -5308 478 -5274
rect 378 -5342 411 -5308
rect 445 -5342 478 -5308
rect 378 -5376 478 -5342
rect 378 -5410 411 -5376
rect 445 -5410 478 -5376
rect 378 -5444 478 -5410
rect 378 -5478 411 -5444
rect 445 -5478 478 -5444
rect 378 -5512 478 -5478
rect 378 -5546 411 -5512
rect 445 -5546 478 -5512
rect 378 -5580 478 -5546
rect 378 -5614 411 -5580
rect 445 -5614 478 -5580
rect 378 -5648 478 -5614
rect 378 -5682 411 -5648
rect 445 -5682 478 -5648
rect 378 -5716 478 -5682
rect 378 -5750 411 -5716
rect 445 -5750 478 -5716
rect 378 -5784 478 -5750
rect 378 -5818 411 -5784
rect 445 -5818 478 -5784
rect 378 -5852 478 -5818
rect 378 -5886 411 -5852
rect 445 -5886 478 -5852
rect 378 -5920 478 -5886
rect 378 -5954 411 -5920
rect 445 -5954 478 -5920
rect 378 -5988 478 -5954
rect 378 -6022 411 -5988
rect 445 -6022 478 -5988
rect 378 -6056 478 -6022
rect 378 -6090 411 -6056
rect 445 -6090 478 -6056
rect 378 -6124 478 -6090
rect 378 -6158 411 -6124
rect 445 -6158 478 -6124
rect 378 -6192 478 -6158
rect 378 -6226 411 -6192
rect 445 -6226 478 -6192
rect 378 -6260 478 -6226
rect 378 -6294 411 -6260
rect 445 -6294 478 -6260
rect 378 -6328 478 -6294
rect 378 -6362 411 -6328
rect 445 -6362 478 -6328
rect 378 -6396 478 -6362
rect 378 -6430 411 -6396
rect 445 -6430 478 -6396
rect 378 -6464 478 -6430
rect 378 -6498 411 -6464
rect 445 -6498 478 -6464
rect 378 -6532 478 -6498
rect 378 -6566 411 -6532
rect 445 -6566 478 -6532
rect 378 -6600 478 -6566
rect 378 -6634 411 -6600
rect 445 -6634 478 -6600
rect 378 -6668 478 -6634
rect 378 -6702 411 -6668
rect 445 -6702 478 -6668
rect 378 -6736 478 -6702
rect 378 -6770 411 -6736
rect 445 -6770 478 -6736
rect 378 -6804 478 -6770
rect 378 -6838 411 -6804
rect 445 -6838 478 -6804
rect 378 -6872 478 -6838
rect 378 -6906 411 -6872
rect 445 -6906 478 -6872
rect 378 -6940 478 -6906
rect 378 -6974 411 -6940
rect 445 -6974 478 -6940
rect 378 -7008 478 -6974
rect 378 -7042 411 -7008
rect 445 -7042 478 -7008
rect 378 -7076 478 -7042
rect 378 -7110 411 -7076
rect 445 -7110 478 -7076
rect 378 -7144 478 -7110
rect 378 -7178 411 -7144
rect 445 -7178 478 -7144
rect 378 -7212 478 -7178
rect 378 -7246 411 -7212
rect 445 -7246 478 -7212
rect 378 -7280 478 -7246
rect 378 -7314 411 -7280
rect 445 -7314 478 -7280
rect 378 -7348 478 -7314
rect 378 -7382 411 -7348
rect 445 -7382 478 -7348
rect 378 -7416 478 -7382
rect 378 -7450 411 -7416
rect 445 -7450 478 -7416
rect 378 -7484 478 -7450
rect 378 -7518 411 -7484
rect 445 -7518 478 -7484
rect 378 -7552 478 -7518
rect 378 -7586 411 -7552
rect 445 -7586 478 -7552
rect 378 -7620 478 -7586
rect 378 -7654 411 -7620
rect 445 -7654 478 -7620
rect 378 -7688 478 -7654
rect 378 -7722 411 -7688
rect 445 -7722 478 -7688
rect 378 -7756 478 -7722
rect 378 -7790 411 -7756
rect 445 -7790 478 -7756
rect 378 -7824 478 -7790
rect 378 -7858 411 -7824
rect 445 -7858 478 -7824
rect 378 -7892 478 -7858
rect 378 -7926 411 -7892
rect 445 -7926 478 -7892
rect 378 -7960 478 -7926
rect 378 -7994 411 -7960
rect 445 -7994 478 -7960
rect 378 -8028 478 -7994
rect 378 -8062 411 -8028
rect 445 -8062 478 -8028
rect 378 -8096 478 -8062
rect 378 -8130 411 -8096
rect 445 -8130 478 -8096
rect 378 -8164 478 -8130
rect 378 -8198 411 -8164
rect 445 -8198 478 -8164
rect 378 -8232 478 -8198
rect 378 -8266 411 -8232
rect 445 -8266 478 -8232
rect 378 -8300 478 -8266
rect 378 -8334 411 -8300
rect 445 -8334 478 -8300
rect 378 -8368 478 -8334
rect 378 -8402 411 -8368
rect 445 -8402 478 -8368
rect 378 -8436 478 -8402
rect 378 -8470 411 -8436
rect 445 -8470 478 -8436
rect 378 -8504 478 -8470
rect 378 -8538 411 -8504
rect 445 -8538 478 -8504
rect 378 -8572 478 -8538
rect 378 -8606 411 -8572
rect 445 -8606 478 -8572
rect 378 -8640 478 -8606
rect 378 -8674 411 -8640
rect 445 -8674 478 -8640
rect 378 -8708 478 -8674
rect 378 -8742 411 -8708
rect 445 -8742 478 -8708
rect 378 -8776 478 -8742
rect 378 -8810 411 -8776
rect 445 -8810 478 -8776
rect 378 -8844 478 -8810
rect 378 -8878 411 -8844
rect 445 -8878 478 -8844
rect 378 -8912 478 -8878
rect 378 -8946 411 -8912
rect 445 -8946 478 -8912
rect 378 -8980 478 -8946
rect 378 -9014 411 -8980
rect 445 -9014 478 -8980
rect 378 -9048 478 -9014
rect 378 -9082 411 -9048
rect 445 -9082 478 -9048
rect 378 -9116 478 -9082
rect 378 -9150 411 -9116
rect 445 -9150 478 -9116
rect 378 -9184 478 -9150
rect 378 -9218 411 -9184
rect 445 -9218 478 -9184
rect 378 -9252 478 -9218
rect 378 -9286 411 -9252
rect 445 -9286 478 -9252
rect 378 -9320 478 -9286
rect 378 -9354 411 -9320
rect 445 -9354 478 -9320
rect 378 -9388 478 -9354
rect 378 -9422 411 -9388
rect 445 -9422 478 -9388
rect 378 -9456 478 -9422
rect 378 -9490 411 -9456
rect 445 -9490 478 -9456
rect 378 -9524 478 -9490
rect 378 -9558 411 -9524
rect 445 -9558 478 -9524
rect 378 -9592 478 -9558
rect 378 -9626 411 -9592
rect 445 -9626 478 -9592
rect 378 -9660 478 -9626
rect 378 -9694 411 -9660
rect 445 -9694 478 -9660
rect 378 -9728 478 -9694
rect 378 -9762 411 -9728
rect 445 -9762 478 -9728
rect 378 -9796 478 -9762
rect 378 -9830 411 -9796
rect 445 -9830 478 -9796
rect 378 -9864 478 -9830
rect 378 -9898 411 -9864
rect 445 -9898 478 -9864
rect 378 -9932 478 -9898
rect 378 -9966 411 -9932
rect 445 -9966 478 -9932
rect 378 -10000 478 -9966
rect 378 -10034 411 -10000
rect 445 -10034 478 -10000
rect 378 -10068 478 -10034
rect 378 -10102 411 -10068
rect 445 -10102 478 -10068
rect 378 -10136 478 -10102
rect 378 -10170 411 -10136
rect 445 -10170 478 -10136
rect 378 -10248 478 -10170
rect 24722 4144 24822 4222
rect 24722 4110 24755 4144
rect 24789 4110 24822 4144
rect 24722 4076 24822 4110
rect 24722 4042 24755 4076
rect 24789 4042 24822 4076
rect 24722 4008 24822 4042
rect 24722 3974 24755 4008
rect 24789 3974 24822 4008
rect 24722 3940 24822 3974
rect 24722 3906 24755 3940
rect 24789 3906 24822 3940
rect 24722 3872 24822 3906
rect 24722 3838 24755 3872
rect 24789 3838 24822 3872
rect 24722 3804 24822 3838
rect 24722 3770 24755 3804
rect 24789 3770 24822 3804
rect 24722 3736 24822 3770
rect 24722 3702 24755 3736
rect 24789 3702 24822 3736
rect 24722 3668 24822 3702
rect 24722 3634 24755 3668
rect 24789 3634 24822 3668
rect 24722 3600 24822 3634
rect 24722 3566 24755 3600
rect 24789 3566 24822 3600
rect 24722 3532 24822 3566
rect 24722 3498 24755 3532
rect 24789 3498 24822 3532
rect 24722 3464 24822 3498
rect 24722 3430 24755 3464
rect 24789 3430 24822 3464
rect 24722 3396 24822 3430
rect 24722 3362 24755 3396
rect 24789 3362 24822 3396
rect 24722 3328 24822 3362
rect 24722 3294 24755 3328
rect 24789 3294 24822 3328
rect 24722 3260 24822 3294
rect 24722 3226 24755 3260
rect 24789 3226 24822 3260
rect 24722 3192 24822 3226
rect 24722 3158 24755 3192
rect 24789 3158 24822 3192
rect 24722 3124 24822 3158
rect 24722 3090 24755 3124
rect 24789 3090 24822 3124
rect 24722 3056 24822 3090
rect 24722 3022 24755 3056
rect 24789 3022 24822 3056
rect 24722 2988 24822 3022
rect 24722 2954 24755 2988
rect 24789 2954 24822 2988
rect 24722 2920 24822 2954
rect 24722 2886 24755 2920
rect 24789 2886 24822 2920
rect 24722 2852 24822 2886
rect 24722 2818 24755 2852
rect 24789 2818 24822 2852
rect 24722 2784 24822 2818
rect 24722 2750 24755 2784
rect 24789 2750 24822 2784
rect 24722 2716 24822 2750
rect 24722 2682 24755 2716
rect 24789 2682 24822 2716
rect 24722 2648 24822 2682
rect 24722 2614 24755 2648
rect 24789 2614 24822 2648
rect 24722 2580 24822 2614
rect 24722 2546 24755 2580
rect 24789 2546 24822 2580
rect 24722 2512 24822 2546
rect 24722 2478 24755 2512
rect 24789 2478 24822 2512
rect 24722 2444 24822 2478
rect 24722 2410 24755 2444
rect 24789 2410 24822 2444
rect 24722 2376 24822 2410
rect 24722 2342 24755 2376
rect 24789 2342 24822 2376
rect 24722 2308 24822 2342
rect 24722 2274 24755 2308
rect 24789 2274 24822 2308
rect 24722 2240 24822 2274
rect 24722 2206 24755 2240
rect 24789 2206 24822 2240
rect 24722 2172 24822 2206
rect 24722 2138 24755 2172
rect 24789 2138 24822 2172
rect 24722 2104 24822 2138
rect 24722 2070 24755 2104
rect 24789 2070 24822 2104
rect 24722 2036 24822 2070
rect 24722 2002 24755 2036
rect 24789 2002 24822 2036
rect 24722 1968 24822 2002
rect 24722 1934 24755 1968
rect 24789 1934 24822 1968
rect 24722 1900 24822 1934
rect 24722 1866 24755 1900
rect 24789 1866 24822 1900
rect 24722 1832 24822 1866
rect 24722 1798 24755 1832
rect 24789 1798 24822 1832
rect 24722 1764 24822 1798
rect 24722 1730 24755 1764
rect 24789 1730 24822 1764
rect 24722 1696 24822 1730
rect 24722 1662 24755 1696
rect 24789 1662 24822 1696
rect 24722 1628 24822 1662
rect 24722 1594 24755 1628
rect 24789 1594 24822 1628
rect 24722 1560 24822 1594
rect 24722 1526 24755 1560
rect 24789 1526 24822 1560
rect 24722 1492 24822 1526
rect 24722 1458 24755 1492
rect 24789 1458 24822 1492
rect 24722 1424 24822 1458
rect 24722 1390 24755 1424
rect 24789 1390 24822 1424
rect 24722 1356 24822 1390
rect 24722 1322 24755 1356
rect 24789 1322 24822 1356
rect 24722 1288 24822 1322
rect 24722 1254 24755 1288
rect 24789 1254 24822 1288
rect 24722 1220 24822 1254
rect 24722 1186 24755 1220
rect 24789 1186 24822 1220
rect 24722 1152 24822 1186
rect 24722 1118 24755 1152
rect 24789 1118 24822 1152
rect 24722 1084 24822 1118
rect 24722 1050 24755 1084
rect 24789 1050 24822 1084
rect 24722 1016 24822 1050
rect 24722 982 24755 1016
rect 24789 982 24822 1016
rect 24722 948 24822 982
rect 24722 914 24755 948
rect 24789 914 24822 948
rect 24722 880 24822 914
rect 24722 846 24755 880
rect 24789 846 24822 880
rect 24722 812 24822 846
rect 24722 778 24755 812
rect 24789 778 24822 812
rect 24722 744 24822 778
rect 24722 710 24755 744
rect 24789 710 24822 744
rect 24722 676 24822 710
rect 24722 642 24755 676
rect 24789 642 24822 676
rect 24722 608 24822 642
rect 24722 574 24755 608
rect 24789 574 24822 608
rect 24722 540 24822 574
rect 24722 506 24755 540
rect 24789 506 24822 540
rect 24722 472 24822 506
rect 24722 438 24755 472
rect 24789 438 24822 472
rect 24722 404 24822 438
rect 24722 370 24755 404
rect 24789 370 24822 404
rect 24722 336 24822 370
rect 24722 302 24755 336
rect 24789 302 24822 336
rect 24722 268 24822 302
rect 24722 234 24755 268
rect 24789 234 24822 268
rect 24722 200 24822 234
rect 24722 166 24755 200
rect 24789 166 24822 200
rect 24722 132 24822 166
rect 24722 98 24755 132
rect 24789 98 24822 132
rect 24722 64 24822 98
rect 24722 30 24755 64
rect 24789 30 24822 64
rect 24722 -4 24822 30
rect 24722 -38 24755 -4
rect 24789 -38 24822 -4
rect 24722 -72 24822 -38
rect 24722 -106 24755 -72
rect 24789 -106 24822 -72
rect 24722 -140 24822 -106
rect 24722 -174 24755 -140
rect 24789 -174 24822 -140
rect 24722 -208 24822 -174
rect 24722 -242 24755 -208
rect 24789 -242 24822 -208
rect 24722 -276 24822 -242
rect 24722 -310 24755 -276
rect 24789 -310 24822 -276
rect 24722 -344 24822 -310
rect 24722 -378 24755 -344
rect 24789 -378 24822 -344
rect 24722 -412 24822 -378
rect 24722 -446 24755 -412
rect 24789 -446 24822 -412
rect 24722 -480 24822 -446
rect 24722 -514 24755 -480
rect 24789 -514 24822 -480
rect 24722 -548 24822 -514
rect 24722 -582 24755 -548
rect 24789 -582 24822 -548
rect 24722 -616 24822 -582
rect 24722 -650 24755 -616
rect 24789 -650 24822 -616
rect 24722 -684 24822 -650
rect 24722 -718 24755 -684
rect 24789 -718 24822 -684
rect 24722 -752 24822 -718
rect 24722 -786 24755 -752
rect 24789 -786 24822 -752
rect 24722 -820 24822 -786
rect 24722 -854 24755 -820
rect 24789 -854 24822 -820
rect 24722 -888 24822 -854
rect 24722 -922 24755 -888
rect 24789 -922 24822 -888
rect 24722 -956 24822 -922
rect 24722 -990 24755 -956
rect 24789 -990 24822 -956
rect 24722 -1024 24822 -990
rect 24722 -1058 24755 -1024
rect 24789 -1058 24822 -1024
rect 24722 -1092 24822 -1058
rect 24722 -1126 24755 -1092
rect 24789 -1126 24822 -1092
rect 24722 -1160 24822 -1126
rect 24722 -1194 24755 -1160
rect 24789 -1194 24822 -1160
rect 24722 -1228 24822 -1194
rect 24722 -1262 24755 -1228
rect 24789 -1262 24822 -1228
rect 24722 -1296 24822 -1262
rect 24722 -1330 24755 -1296
rect 24789 -1330 24822 -1296
rect 24722 -1364 24822 -1330
rect 24722 -1398 24755 -1364
rect 24789 -1398 24822 -1364
rect 24722 -1432 24822 -1398
rect 24722 -1466 24755 -1432
rect 24789 -1466 24822 -1432
rect 24722 -1500 24822 -1466
rect 24722 -1534 24755 -1500
rect 24789 -1534 24822 -1500
rect 24722 -1568 24822 -1534
rect 24722 -1602 24755 -1568
rect 24789 -1602 24822 -1568
rect 24722 -1636 24822 -1602
rect 24722 -1670 24755 -1636
rect 24789 -1670 24822 -1636
rect 24722 -1704 24822 -1670
rect 24722 -1738 24755 -1704
rect 24789 -1738 24822 -1704
rect 24722 -1772 24822 -1738
rect 24722 -1806 24755 -1772
rect 24789 -1806 24822 -1772
rect 24722 -1840 24822 -1806
rect 24722 -1874 24755 -1840
rect 24789 -1874 24822 -1840
rect 24722 -1908 24822 -1874
rect 24722 -1942 24755 -1908
rect 24789 -1942 24822 -1908
rect 24722 -1976 24822 -1942
rect 24722 -2010 24755 -1976
rect 24789 -2010 24822 -1976
rect 24722 -2044 24822 -2010
rect 24722 -2078 24755 -2044
rect 24789 -2078 24822 -2044
rect 24722 -2112 24822 -2078
rect 24722 -2146 24755 -2112
rect 24789 -2146 24822 -2112
rect 24722 -2180 24822 -2146
rect 24722 -2214 24755 -2180
rect 24789 -2214 24822 -2180
rect 24722 -2248 24822 -2214
rect 24722 -2282 24755 -2248
rect 24789 -2282 24822 -2248
rect 24722 -2316 24822 -2282
rect 24722 -2350 24755 -2316
rect 24789 -2350 24822 -2316
rect 24722 -2384 24822 -2350
rect 24722 -2418 24755 -2384
rect 24789 -2418 24822 -2384
rect 24722 -2452 24822 -2418
rect 24722 -2486 24755 -2452
rect 24789 -2486 24822 -2452
rect 24722 -2520 24822 -2486
rect 24722 -2554 24755 -2520
rect 24789 -2554 24822 -2520
rect 24722 -2588 24822 -2554
rect 24722 -2622 24755 -2588
rect 24789 -2622 24822 -2588
rect 24722 -2656 24822 -2622
rect 24722 -2690 24755 -2656
rect 24789 -2690 24822 -2656
rect 24722 -2724 24822 -2690
rect 24722 -2758 24755 -2724
rect 24789 -2758 24822 -2724
rect 24722 -2792 24822 -2758
rect 24722 -2826 24755 -2792
rect 24789 -2826 24822 -2792
rect 24722 -2860 24822 -2826
rect 24722 -2894 24755 -2860
rect 24789 -2894 24822 -2860
rect 24722 -2928 24822 -2894
rect 24722 -2962 24755 -2928
rect 24789 -2962 24822 -2928
rect 24722 -2996 24822 -2962
rect 24722 -3030 24755 -2996
rect 24789 -3030 24822 -2996
rect 24722 -3064 24822 -3030
rect 24722 -3098 24755 -3064
rect 24789 -3098 24822 -3064
rect 24722 -3132 24822 -3098
rect 24722 -3166 24755 -3132
rect 24789 -3166 24822 -3132
rect 24722 -3200 24822 -3166
rect 24722 -3234 24755 -3200
rect 24789 -3234 24822 -3200
rect 24722 -3268 24822 -3234
rect 24722 -3302 24755 -3268
rect 24789 -3302 24822 -3268
rect 24722 -3336 24822 -3302
rect 24722 -3370 24755 -3336
rect 24789 -3370 24822 -3336
rect 24722 -3404 24822 -3370
rect 24722 -3438 24755 -3404
rect 24789 -3438 24822 -3404
rect 24722 -3472 24822 -3438
rect 24722 -3506 24755 -3472
rect 24789 -3506 24822 -3472
rect 24722 -3540 24822 -3506
rect 24722 -3574 24755 -3540
rect 24789 -3574 24822 -3540
rect 24722 -3608 24822 -3574
rect 24722 -3642 24755 -3608
rect 24789 -3642 24822 -3608
rect 24722 -3676 24822 -3642
rect 24722 -3710 24755 -3676
rect 24789 -3710 24822 -3676
rect 24722 -3744 24822 -3710
rect 24722 -3778 24755 -3744
rect 24789 -3778 24822 -3744
rect 24722 -3812 24822 -3778
rect 24722 -3846 24755 -3812
rect 24789 -3846 24822 -3812
rect 24722 -3880 24822 -3846
rect 24722 -3914 24755 -3880
rect 24789 -3914 24822 -3880
rect 24722 -3948 24822 -3914
rect 24722 -3982 24755 -3948
rect 24789 -3982 24822 -3948
rect 24722 -4016 24822 -3982
rect 24722 -4050 24755 -4016
rect 24789 -4050 24822 -4016
rect 24722 -4084 24822 -4050
rect 24722 -4118 24755 -4084
rect 24789 -4118 24822 -4084
rect 24722 -4152 24822 -4118
rect 24722 -4186 24755 -4152
rect 24789 -4186 24822 -4152
rect 24722 -4220 24822 -4186
rect 24722 -4254 24755 -4220
rect 24789 -4254 24822 -4220
rect 24722 -4288 24822 -4254
rect 24722 -4322 24755 -4288
rect 24789 -4322 24822 -4288
rect 24722 -4356 24822 -4322
rect 24722 -4390 24755 -4356
rect 24789 -4390 24822 -4356
rect 24722 -4424 24822 -4390
rect 24722 -4458 24755 -4424
rect 24789 -4458 24822 -4424
rect 24722 -4492 24822 -4458
rect 24722 -4526 24755 -4492
rect 24789 -4526 24822 -4492
rect 24722 -4560 24822 -4526
rect 24722 -4594 24755 -4560
rect 24789 -4594 24822 -4560
rect 24722 -4628 24822 -4594
rect 24722 -4662 24755 -4628
rect 24789 -4662 24822 -4628
rect 24722 -4696 24822 -4662
rect 24722 -4730 24755 -4696
rect 24789 -4730 24822 -4696
rect 24722 -4764 24822 -4730
rect 24722 -4798 24755 -4764
rect 24789 -4798 24822 -4764
rect 24722 -4832 24822 -4798
rect 24722 -4866 24755 -4832
rect 24789 -4866 24822 -4832
rect 24722 -4900 24822 -4866
rect 24722 -4934 24755 -4900
rect 24789 -4934 24822 -4900
rect 24722 -4968 24822 -4934
rect 24722 -5002 24755 -4968
rect 24789 -5002 24822 -4968
rect 24722 -5036 24822 -5002
rect 24722 -5070 24755 -5036
rect 24789 -5070 24822 -5036
rect 24722 -5104 24822 -5070
rect 24722 -5138 24755 -5104
rect 24789 -5138 24822 -5104
rect 24722 -5172 24822 -5138
rect 24722 -5206 24755 -5172
rect 24789 -5206 24822 -5172
rect 24722 -5240 24822 -5206
rect 24722 -5274 24755 -5240
rect 24789 -5274 24822 -5240
rect 24722 -5308 24822 -5274
rect 24722 -5342 24755 -5308
rect 24789 -5342 24822 -5308
rect 24722 -5376 24822 -5342
rect 24722 -5410 24755 -5376
rect 24789 -5410 24822 -5376
rect 24722 -5444 24822 -5410
rect 24722 -5478 24755 -5444
rect 24789 -5478 24822 -5444
rect 24722 -5512 24822 -5478
rect 24722 -5546 24755 -5512
rect 24789 -5546 24822 -5512
rect 24722 -5580 24822 -5546
rect 24722 -5614 24755 -5580
rect 24789 -5614 24822 -5580
rect 24722 -5648 24822 -5614
rect 24722 -5682 24755 -5648
rect 24789 -5682 24822 -5648
rect 24722 -5716 24822 -5682
rect 24722 -5750 24755 -5716
rect 24789 -5750 24822 -5716
rect 24722 -5784 24822 -5750
rect 24722 -5818 24755 -5784
rect 24789 -5818 24822 -5784
rect 24722 -5852 24822 -5818
rect 24722 -5886 24755 -5852
rect 24789 -5886 24822 -5852
rect 24722 -5920 24822 -5886
rect 24722 -5954 24755 -5920
rect 24789 -5954 24822 -5920
rect 24722 -5988 24822 -5954
rect 24722 -6022 24755 -5988
rect 24789 -6022 24822 -5988
rect 24722 -6056 24822 -6022
rect 24722 -6090 24755 -6056
rect 24789 -6090 24822 -6056
rect 24722 -6124 24822 -6090
rect 24722 -6158 24755 -6124
rect 24789 -6158 24822 -6124
rect 24722 -6192 24822 -6158
rect 24722 -6226 24755 -6192
rect 24789 -6226 24822 -6192
rect 24722 -6260 24822 -6226
rect 24722 -6294 24755 -6260
rect 24789 -6294 24822 -6260
rect 24722 -6328 24822 -6294
rect 24722 -6362 24755 -6328
rect 24789 -6362 24822 -6328
rect 24722 -6396 24822 -6362
rect 24722 -6430 24755 -6396
rect 24789 -6430 24822 -6396
rect 24722 -6464 24822 -6430
rect 24722 -6498 24755 -6464
rect 24789 -6498 24822 -6464
rect 24722 -6532 24822 -6498
rect 24722 -6566 24755 -6532
rect 24789 -6566 24822 -6532
rect 24722 -6600 24822 -6566
rect 24722 -6634 24755 -6600
rect 24789 -6634 24822 -6600
rect 24722 -6668 24822 -6634
rect 24722 -6702 24755 -6668
rect 24789 -6702 24822 -6668
rect 24722 -6736 24822 -6702
rect 24722 -6770 24755 -6736
rect 24789 -6770 24822 -6736
rect 24722 -6804 24822 -6770
rect 24722 -6838 24755 -6804
rect 24789 -6838 24822 -6804
rect 24722 -6872 24822 -6838
rect 24722 -6906 24755 -6872
rect 24789 -6906 24822 -6872
rect 24722 -6940 24822 -6906
rect 24722 -6974 24755 -6940
rect 24789 -6974 24822 -6940
rect 24722 -7008 24822 -6974
rect 24722 -7042 24755 -7008
rect 24789 -7042 24822 -7008
rect 24722 -7076 24822 -7042
rect 24722 -7110 24755 -7076
rect 24789 -7110 24822 -7076
rect 24722 -7144 24822 -7110
rect 24722 -7178 24755 -7144
rect 24789 -7178 24822 -7144
rect 24722 -7212 24822 -7178
rect 24722 -7246 24755 -7212
rect 24789 -7246 24822 -7212
rect 24722 -7280 24822 -7246
rect 24722 -7314 24755 -7280
rect 24789 -7314 24822 -7280
rect 24722 -7348 24822 -7314
rect 24722 -7382 24755 -7348
rect 24789 -7382 24822 -7348
rect 24722 -7416 24822 -7382
rect 24722 -7450 24755 -7416
rect 24789 -7450 24822 -7416
rect 24722 -7484 24822 -7450
rect 24722 -7518 24755 -7484
rect 24789 -7518 24822 -7484
rect 24722 -7552 24822 -7518
rect 24722 -7586 24755 -7552
rect 24789 -7586 24822 -7552
rect 24722 -7620 24822 -7586
rect 24722 -7654 24755 -7620
rect 24789 -7654 24822 -7620
rect 24722 -7688 24822 -7654
rect 24722 -7722 24755 -7688
rect 24789 -7722 24822 -7688
rect 24722 -7756 24822 -7722
rect 24722 -7790 24755 -7756
rect 24789 -7790 24822 -7756
rect 24722 -7824 24822 -7790
rect 24722 -7858 24755 -7824
rect 24789 -7858 24822 -7824
rect 24722 -7892 24822 -7858
rect 24722 -7926 24755 -7892
rect 24789 -7926 24822 -7892
rect 24722 -7960 24822 -7926
rect 24722 -7994 24755 -7960
rect 24789 -7994 24822 -7960
rect 24722 -8028 24822 -7994
rect 24722 -8062 24755 -8028
rect 24789 -8062 24822 -8028
rect 24722 -8096 24822 -8062
rect 24722 -8130 24755 -8096
rect 24789 -8130 24822 -8096
rect 24722 -8164 24822 -8130
rect 24722 -8198 24755 -8164
rect 24789 -8198 24822 -8164
rect 24722 -8232 24822 -8198
rect 24722 -8266 24755 -8232
rect 24789 -8266 24822 -8232
rect 24722 -8300 24822 -8266
rect 24722 -8334 24755 -8300
rect 24789 -8334 24822 -8300
rect 24722 -8368 24822 -8334
rect 24722 -8402 24755 -8368
rect 24789 -8402 24822 -8368
rect 24722 -8436 24822 -8402
rect 24722 -8470 24755 -8436
rect 24789 -8470 24822 -8436
rect 24722 -8504 24822 -8470
rect 24722 -8538 24755 -8504
rect 24789 -8538 24822 -8504
rect 24722 -8572 24822 -8538
rect 24722 -8606 24755 -8572
rect 24789 -8606 24822 -8572
rect 24722 -8640 24822 -8606
rect 24722 -8674 24755 -8640
rect 24789 -8674 24822 -8640
rect 24722 -8708 24822 -8674
rect 24722 -8742 24755 -8708
rect 24789 -8742 24822 -8708
rect 24722 -8776 24822 -8742
rect 24722 -8810 24755 -8776
rect 24789 -8810 24822 -8776
rect 24722 -8844 24822 -8810
rect 24722 -8878 24755 -8844
rect 24789 -8878 24822 -8844
rect 24722 -8912 24822 -8878
rect 24722 -8946 24755 -8912
rect 24789 -8946 24822 -8912
rect 24722 -8980 24822 -8946
rect 24722 -9014 24755 -8980
rect 24789 -9014 24822 -8980
rect 24722 -9048 24822 -9014
rect 24722 -9082 24755 -9048
rect 24789 -9082 24822 -9048
rect 24722 -9116 24822 -9082
rect 24722 -9150 24755 -9116
rect 24789 -9150 24822 -9116
rect 24722 -9184 24822 -9150
rect 24722 -9218 24755 -9184
rect 24789 -9218 24822 -9184
rect 24722 -9252 24822 -9218
rect 24722 -9286 24755 -9252
rect 24789 -9286 24822 -9252
rect 24722 -9320 24822 -9286
rect 24722 -9354 24755 -9320
rect 24789 -9354 24822 -9320
rect 24722 -9388 24822 -9354
rect 24722 -9422 24755 -9388
rect 24789 -9422 24822 -9388
rect 24722 -9456 24822 -9422
rect 24722 -9490 24755 -9456
rect 24789 -9490 24822 -9456
rect 24722 -9524 24822 -9490
rect 24722 -9558 24755 -9524
rect 24789 -9558 24822 -9524
rect 24722 -9592 24822 -9558
rect 24722 -9626 24755 -9592
rect 24789 -9626 24822 -9592
rect 24722 -9660 24822 -9626
rect 24722 -9694 24755 -9660
rect 24789 -9694 24822 -9660
rect 24722 -9728 24822 -9694
rect 24722 -9762 24755 -9728
rect 24789 -9762 24822 -9728
rect 24722 -9796 24822 -9762
rect 24722 -9830 24755 -9796
rect 24789 -9830 24822 -9796
rect 24722 -9864 24822 -9830
rect 24722 -9898 24755 -9864
rect 24789 -9898 24822 -9864
rect 24722 -9932 24822 -9898
rect 24722 -9966 24755 -9932
rect 24789 -9966 24822 -9932
rect 24722 -10000 24822 -9966
rect 24722 -10034 24755 -10000
rect 24789 -10034 24822 -10000
rect 24722 -10068 24822 -10034
rect 24722 -10102 24755 -10068
rect 24789 -10102 24822 -10068
rect 24722 -10136 24822 -10102
rect 24722 -10170 24755 -10136
rect 24789 -10170 24822 -10136
rect 24722 -10248 24822 -10170
rect 378 -10281 24822 -10248
rect 378 -10315 547 -10281
rect 581 -10315 615 -10281
rect 649 -10315 683 -10281
rect 717 -10315 751 -10281
rect 785 -10315 819 -10281
rect 853 -10315 887 -10281
rect 921 -10315 955 -10281
rect 989 -10315 1023 -10281
rect 1057 -10315 1091 -10281
rect 1125 -10315 1159 -10281
rect 1193 -10315 1227 -10281
rect 1261 -10315 1295 -10281
rect 1329 -10315 1363 -10281
rect 1397 -10315 1431 -10281
rect 1465 -10315 1499 -10281
rect 1533 -10315 1567 -10281
rect 1601 -10315 1635 -10281
rect 1669 -10315 1703 -10281
rect 1737 -10315 1771 -10281
rect 1805 -10315 1839 -10281
rect 1873 -10315 1907 -10281
rect 1941 -10315 1975 -10281
rect 2009 -10315 2043 -10281
rect 2077 -10315 2111 -10281
rect 2145 -10315 2179 -10281
rect 2213 -10315 2247 -10281
rect 2281 -10315 2315 -10281
rect 2349 -10315 2383 -10281
rect 2417 -10315 2451 -10281
rect 2485 -10315 2519 -10281
rect 2553 -10315 2587 -10281
rect 2621 -10315 2655 -10281
rect 2689 -10315 2723 -10281
rect 2757 -10315 2791 -10281
rect 2825 -10315 2859 -10281
rect 2893 -10315 2927 -10281
rect 2961 -10315 2995 -10281
rect 3029 -10315 3063 -10281
rect 3097 -10315 3131 -10281
rect 3165 -10315 3199 -10281
rect 3233 -10315 3267 -10281
rect 3301 -10315 3335 -10281
rect 3369 -10315 3403 -10281
rect 3437 -10315 3471 -10281
rect 3505 -10315 3539 -10281
rect 3573 -10315 3607 -10281
rect 3641 -10315 3675 -10281
rect 3709 -10315 3743 -10281
rect 3777 -10315 3811 -10281
rect 3845 -10315 3879 -10281
rect 3913 -10315 3947 -10281
rect 3981 -10315 4015 -10281
rect 4049 -10315 4083 -10281
rect 4117 -10315 4151 -10281
rect 4185 -10315 4219 -10281
rect 4253 -10315 4287 -10281
rect 4321 -10315 4355 -10281
rect 4389 -10315 4423 -10281
rect 4457 -10315 4491 -10281
rect 4525 -10315 4559 -10281
rect 4593 -10315 4627 -10281
rect 4661 -10315 4695 -10281
rect 4729 -10315 4763 -10281
rect 4797 -10315 4831 -10281
rect 4865 -10315 4899 -10281
rect 4933 -10315 4967 -10281
rect 5001 -10315 5035 -10281
rect 5069 -10315 5103 -10281
rect 5137 -10315 5171 -10281
rect 5205 -10315 5239 -10281
rect 5273 -10315 5307 -10281
rect 5341 -10315 5375 -10281
rect 5409 -10315 5443 -10281
rect 5477 -10315 5511 -10281
rect 5545 -10315 5579 -10281
rect 5613 -10315 5647 -10281
rect 5681 -10315 5715 -10281
rect 5749 -10315 5783 -10281
rect 5817 -10315 5851 -10281
rect 5885 -10315 5919 -10281
rect 5953 -10315 5987 -10281
rect 6021 -10315 6055 -10281
rect 6089 -10315 6123 -10281
rect 6157 -10315 6191 -10281
rect 6225 -10315 6259 -10281
rect 6293 -10315 6327 -10281
rect 6361 -10315 6395 -10281
rect 6429 -10315 6463 -10281
rect 6497 -10315 6531 -10281
rect 6565 -10315 6599 -10281
rect 6633 -10315 6667 -10281
rect 6701 -10315 6735 -10281
rect 6769 -10315 6803 -10281
rect 6837 -10315 6871 -10281
rect 6905 -10315 6939 -10281
rect 6973 -10315 7007 -10281
rect 7041 -10315 7075 -10281
rect 7109 -10315 7143 -10281
rect 7177 -10315 7211 -10281
rect 7245 -10315 7279 -10281
rect 7313 -10315 7347 -10281
rect 7381 -10315 7415 -10281
rect 7449 -10315 7483 -10281
rect 7517 -10315 7551 -10281
rect 7585 -10315 7619 -10281
rect 7653 -10315 7687 -10281
rect 7721 -10315 7755 -10281
rect 7789 -10315 7823 -10281
rect 7857 -10315 7891 -10281
rect 7925 -10315 7959 -10281
rect 7993 -10315 8027 -10281
rect 8061 -10315 8095 -10281
rect 8129 -10315 8163 -10281
rect 8197 -10315 8231 -10281
rect 8265 -10315 8299 -10281
rect 8333 -10315 8367 -10281
rect 8401 -10315 8435 -10281
rect 8469 -10315 8503 -10281
rect 8537 -10315 8571 -10281
rect 8605 -10315 8639 -10281
rect 8673 -10315 8707 -10281
rect 8741 -10315 8775 -10281
rect 8809 -10315 8843 -10281
rect 8877 -10315 8911 -10281
rect 8945 -10315 8979 -10281
rect 9013 -10315 9047 -10281
rect 9081 -10315 9115 -10281
rect 9149 -10315 9183 -10281
rect 9217 -10315 9251 -10281
rect 9285 -10315 9319 -10281
rect 9353 -10315 9387 -10281
rect 9421 -10315 9455 -10281
rect 9489 -10315 9523 -10281
rect 9557 -10315 9591 -10281
rect 9625 -10315 9659 -10281
rect 9693 -10315 9727 -10281
rect 9761 -10315 9795 -10281
rect 9829 -10315 9863 -10281
rect 9897 -10315 9931 -10281
rect 9965 -10315 9999 -10281
rect 10033 -10315 10067 -10281
rect 10101 -10315 10135 -10281
rect 10169 -10315 10203 -10281
rect 10237 -10315 10271 -10281
rect 10305 -10315 10339 -10281
rect 10373 -10315 10407 -10281
rect 10441 -10315 10475 -10281
rect 10509 -10315 10543 -10281
rect 10577 -10315 10611 -10281
rect 10645 -10315 10679 -10281
rect 10713 -10315 10747 -10281
rect 10781 -10315 10815 -10281
rect 10849 -10315 10883 -10281
rect 10917 -10315 10951 -10281
rect 10985 -10315 11019 -10281
rect 11053 -10315 11087 -10281
rect 11121 -10315 11155 -10281
rect 11189 -10315 11223 -10281
rect 11257 -10315 11291 -10281
rect 11325 -10315 11359 -10281
rect 11393 -10315 11427 -10281
rect 11461 -10315 11495 -10281
rect 11529 -10315 11563 -10281
rect 11597 -10315 11631 -10281
rect 11665 -10315 11699 -10281
rect 11733 -10315 11767 -10281
rect 11801 -10315 11835 -10281
rect 11869 -10315 11903 -10281
rect 11937 -10315 11971 -10281
rect 12005 -10315 12039 -10281
rect 12073 -10315 12107 -10281
rect 12141 -10315 12175 -10281
rect 12209 -10315 12243 -10281
rect 12277 -10315 12311 -10281
rect 12345 -10315 12379 -10281
rect 12413 -10315 12447 -10281
rect 12481 -10315 12515 -10281
rect 12549 -10315 12583 -10281
rect 12617 -10315 12651 -10281
rect 12685 -10315 12719 -10281
rect 12753 -10315 12787 -10281
rect 12821 -10315 12855 -10281
rect 12889 -10315 12923 -10281
rect 12957 -10315 12991 -10281
rect 13025 -10315 13059 -10281
rect 13093 -10315 13127 -10281
rect 13161 -10315 13195 -10281
rect 13229 -10315 13263 -10281
rect 13297 -10315 13331 -10281
rect 13365 -10315 13399 -10281
rect 13433 -10315 13467 -10281
rect 13501 -10315 13535 -10281
rect 13569 -10315 13603 -10281
rect 13637 -10315 13671 -10281
rect 13705 -10315 13739 -10281
rect 13773 -10315 13807 -10281
rect 13841 -10315 13875 -10281
rect 13909 -10315 13943 -10281
rect 13977 -10315 14011 -10281
rect 14045 -10315 14079 -10281
rect 14113 -10315 14147 -10281
rect 14181 -10315 14215 -10281
rect 14249 -10315 14283 -10281
rect 14317 -10315 14351 -10281
rect 14385 -10315 14419 -10281
rect 14453 -10315 14487 -10281
rect 14521 -10315 14555 -10281
rect 14589 -10315 14623 -10281
rect 14657 -10315 14691 -10281
rect 14725 -10315 14759 -10281
rect 14793 -10315 14827 -10281
rect 14861 -10315 14895 -10281
rect 14929 -10315 14963 -10281
rect 14997 -10315 15031 -10281
rect 15065 -10315 15099 -10281
rect 15133 -10315 15167 -10281
rect 15201 -10315 15235 -10281
rect 15269 -10315 15303 -10281
rect 15337 -10315 15371 -10281
rect 15405 -10315 15439 -10281
rect 15473 -10315 15507 -10281
rect 15541 -10315 15575 -10281
rect 15609 -10315 15643 -10281
rect 15677 -10315 15711 -10281
rect 15745 -10315 15779 -10281
rect 15813 -10315 15847 -10281
rect 15881 -10315 15915 -10281
rect 15949 -10315 15983 -10281
rect 16017 -10315 16051 -10281
rect 16085 -10315 16119 -10281
rect 16153 -10315 16187 -10281
rect 16221 -10315 16255 -10281
rect 16289 -10315 16323 -10281
rect 16357 -10315 16391 -10281
rect 16425 -10315 16459 -10281
rect 16493 -10315 16527 -10281
rect 16561 -10315 16595 -10281
rect 16629 -10315 16663 -10281
rect 16697 -10315 16731 -10281
rect 16765 -10315 16799 -10281
rect 16833 -10315 16867 -10281
rect 16901 -10315 16935 -10281
rect 16969 -10315 17003 -10281
rect 17037 -10315 17071 -10281
rect 17105 -10315 17139 -10281
rect 17173 -10315 17207 -10281
rect 17241 -10315 17275 -10281
rect 17309 -10315 17343 -10281
rect 17377 -10315 17411 -10281
rect 17445 -10315 17479 -10281
rect 17513 -10315 17547 -10281
rect 17581 -10315 17615 -10281
rect 17649 -10315 17683 -10281
rect 17717 -10315 17751 -10281
rect 17785 -10315 17819 -10281
rect 17853 -10315 17887 -10281
rect 17921 -10315 17955 -10281
rect 17989 -10315 18023 -10281
rect 18057 -10315 18091 -10281
rect 18125 -10315 18159 -10281
rect 18193 -10315 18227 -10281
rect 18261 -10315 18295 -10281
rect 18329 -10315 18363 -10281
rect 18397 -10315 18431 -10281
rect 18465 -10315 18499 -10281
rect 18533 -10315 18567 -10281
rect 18601 -10315 18635 -10281
rect 18669 -10315 18703 -10281
rect 18737 -10315 18771 -10281
rect 18805 -10315 18839 -10281
rect 18873 -10315 18907 -10281
rect 18941 -10315 18975 -10281
rect 19009 -10315 19043 -10281
rect 19077 -10315 19111 -10281
rect 19145 -10315 19179 -10281
rect 19213 -10315 19247 -10281
rect 19281 -10315 19315 -10281
rect 19349 -10315 19383 -10281
rect 19417 -10315 19451 -10281
rect 19485 -10315 19519 -10281
rect 19553 -10315 19587 -10281
rect 19621 -10315 19655 -10281
rect 19689 -10315 19723 -10281
rect 19757 -10315 19791 -10281
rect 19825 -10315 19859 -10281
rect 19893 -10315 19927 -10281
rect 19961 -10315 19995 -10281
rect 20029 -10315 20063 -10281
rect 20097 -10315 20131 -10281
rect 20165 -10315 20199 -10281
rect 20233 -10315 20267 -10281
rect 20301 -10315 20335 -10281
rect 20369 -10315 20403 -10281
rect 20437 -10315 20471 -10281
rect 20505 -10315 20539 -10281
rect 20573 -10315 20607 -10281
rect 20641 -10315 20675 -10281
rect 20709 -10315 20743 -10281
rect 20777 -10315 20811 -10281
rect 20845 -10315 20879 -10281
rect 20913 -10315 20947 -10281
rect 20981 -10315 21015 -10281
rect 21049 -10315 21083 -10281
rect 21117 -10315 21151 -10281
rect 21185 -10315 21219 -10281
rect 21253 -10315 21287 -10281
rect 21321 -10315 21355 -10281
rect 21389 -10315 21423 -10281
rect 21457 -10315 21491 -10281
rect 21525 -10315 21559 -10281
rect 21593 -10315 21627 -10281
rect 21661 -10315 21695 -10281
rect 21729 -10315 21763 -10281
rect 21797 -10315 21831 -10281
rect 21865 -10315 21899 -10281
rect 21933 -10315 21967 -10281
rect 22001 -10315 22035 -10281
rect 22069 -10315 22103 -10281
rect 22137 -10315 22171 -10281
rect 22205 -10315 22239 -10281
rect 22273 -10315 22307 -10281
rect 22341 -10315 22375 -10281
rect 22409 -10315 22443 -10281
rect 22477 -10315 22511 -10281
rect 22545 -10315 22579 -10281
rect 22613 -10315 22647 -10281
rect 22681 -10315 22715 -10281
rect 22749 -10315 22783 -10281
rect 22817 -10315 22851 -10281
rect 22885 -10315 22919 -10281
rect 22953 -10315 22987 -10281
rect 23021 -10315 23055 -10281
rect 23089 -10315 23123 -10281
rect 23157 -10315 23191 -10281
rect 23225 -10315 23259 -10281
rect 23293 -10315 23327 -10281
rect 23361 -10315 23395 -10281
rect 23429 -10315 23463 -10281
rect 23497 -10315 23531 -10281
rect 23565 -10315 23599 -10281
rect 23633 -10315 23667 -10281
rect 23701 -10315 23735 -10281
rect 23769 -10315 23803 -10281
rect 23837 -10315 23871 -10281
rect 23905 -10315 23939 -10281
rect 23973 -10315 24007 -10281
rect 24041 -10315 24075 -10281
rect 24109 -10315 24143 -10281
rect 24177 -10315 24211 -10281
rect 24245 -10315 24279 -10281
rect 24313 -10315 24347 -10281
rect 24381 -10315 24415 -10281
rect 24449 -10315 24483 -10281
rect 24517 -10315 24551 -10281
rect 24585 -10315 24619 -10281
rect 24653 -10315 24822 -10281
rect 378 -10348 24822 -10315
<< psubdiffcont >>
rect -12145 -11245 -12111 -11211
rect -12077 -11245 -12043 -11211
rect -12009 -11245 -11975 -11211
rect -11941 -11245 -11907 -11211
rect -11873 -11245 -11839 -11211
rect -11805 -11245 -11771 -11211
rect -11737 -11245 -11703 -11211
rect -11669 -11245 -11635 -11211
rect -11601 -11245 -11567 -11211
rect -11533 -11245 -11499 -11211
rect -11465 -11245 -11431 -11211
rect -11397 -11245 -11363 -11211
rect -11329 -11245 -11295 -11211
rect -11261 -11245 -11227 -11211
rect -11193 -11245 -11159 -11211
rect -11125 -11245 -11091 -11211
rect -11057 -11245 -11023 -11211
rect -10989 -11245 -10955 -11211
rect -10921 -11245 -10887 -11211
rect -10853 -11245 -10819 -11211
rect -10785 -11245 -10751 -11211
rect -10717 -11245 -10683 -11211
rect -10649 -11245 -10615 -11211
rect -10581 -11245 -10547 -11211
rect -10513 -11245 -10479 -11211
rect -10445 -11245 -10411 -11211
rect -10377 -11245 -10343 -11211
rect -10309 -11245 -10275 -11211
rect -10241 -11245 -10207 -11211
rect -10173 -11245 -10139 -11211
rect -10105 -11245 -10071 -11211
rect -10037 -11245 -10003 -11211
rect -9969 -11245 -9935 -11211
rect -9901 -11245 -9867 -11211
rect -9833 -11245 -9799 -11211
rect -9765 -11245 -9731 -11211
rect -9697 -11245 -9663 -11211
rect -9629 -11245 -9595 -11211
rect -9561 -11245 -9527 -11211
rect -9493 -11245 -9459 -11211
rect -9425 -11245 -9391 -11211
rect -9357 -11245 -9323 -11211
rect -9289 -11245 -9255 -11211
rect -9221 -11245 -9187 -11211
rect -9153 -11245 -9119 -11211
rect -9085 -11245 -9051 -11211
rect -9017 -11245 -8983 -11211
rect -8949 -11245 -8915 -11211
rect -8881 -11245 -8847 -11211
rect -8813 -11245 -8779 -11211
rect -8745 -11245 -8711 -11211
rect -8677 -11245 -8643 -11211
rect -8609 -11245 -8575 -11211
rect -8541 -11245 -8507 -11211
rect -8473 -11245 -8439 -11211
rect -8405 -11245 -8371 -11211
rect -8337 -11245 -8303 -11211
rect -8269 -11245 -8235 -11211
rect -8201 -11245 -8167 -11211
rect -8133 -11245 -8099 -11211
rect -8065 -11245 -8031 -11211
rect -7997 -11245 -7963 -11211
rect -7929 -11245 -7895 -11211
rect -7861 -11245 -7827 -11211
rect -7793 -11245 -7759 -11211
rect -7725 -11245 -7691 -11211
rect -7657 -11245 -7623 -11211
rect -7589 -11245 -7555 -11211
rect -7521 -11245 -7487 -11211
rect -7453 -11245 -7419 -11211
rect -7385 -11245 -7351 -11211
rect -7317 -11245 -7283 -11211
rect -7249 -11245 -7215 -11211
rect -7181 -11245 -7147 -11211
rect -7113 -11245 -7079 -11211
rect -7045 -11245 -7011 -11211
rect -6977 -11245 -6943 -11211
rect -6909 -11245 -6875 -11211
rect -6841 -11245 -6807 -11211
rect -6773 -11245 -6739 -11211
rect -6705 -11245 -6671 -11211
rect -6637 -11245 -6603 -11211
rect -6569 -11245 -6535 -11211
rect -6501 -11245 -6467 -11211
rect -6433 -11245 -6399 -11211
rect -6365 -11245 -6331 -11211
rect -6297 -11245 -6263 -11211
rect -6229 -11245 -6195 -11211
rect -6161 -11245 -6127 -11211
rect -6093 -11245 -6059 -11211
rect -6025 -11245 -5991 -11211
rect -5957 -11245 -5923 -11211
rect -5889 -11245 -5855 -11211
rect -5821 -11245 -5787 -11211
rect -5753 -11245 -5719 -11211
rect -5685 -11245 -5651 -11211
rect -5617 -11245 -5583 -11211
rect -5549 -11245 -5515 -11211
rect -5481 -11245 -5447 -11211
rect -5413 -11245 -5379 -11211
rect -5345 -11245 -5311 -11211
rect -5277 -11245 -5243 -11211
rect -5209 -11245 -5175 -11211
rect -5141 -11245 -5107 -11211
rect -5073 -11245 -5039 -11211
rect -5005 -11245 -4971 -11211
rect -4937 -11245 -4903 -11211
rect -4869 -11245 -4835 -11211
rect -4801 -11245 -4767 -11211
rect -4733 -11245 -4699 -11211
rect -4665 -11245 -4631 -11211
rect -4597 -11245 -4563 -11211
rect -4529 -11245 -4495 -11211
rect -4461 -11245 -4427 -11211
rect -4393 -11245 -4359 -11211
rect -4325 -11245 -4291 -11211
rect -4257 -11245 -4223 -11211
rect -4189 -11245 -4155 -11211
rect -4121 -11245 -4087 -11211
rect -4053 -11245 -4019 -11211
rect -3985 -11245 -3951 -11211
rect -3917 -11245 -3883 -11211
rect -3849 -11245 -3815 -11211
rect -3781 -11245 -3747 -11211
rect -3713 -11245 -3679 -11211
rect -3645 -11245 -3611 -11211
rect -3577 -11245 -3543 -11211
rect -3509 -11245 -3475 -11211
rect -3441 -11245 -3407 -11211
rect -3373 -11245 -3339 -11211
rect -3305 -11245 -3271 -11211
rect -3237 -11245 -3203 -11211
rect -3169 -11245 -3135 -11211
rect -3101 -11245 -3067 -11211
rect -3033 -11245 -2999 -11211
rect -2965 -11245 -2931 -11211
rect -2897 -11245 -2863 -11211
rect -2829 -11245 -2795 -11211
rect -2761 -11245 -2727 -11211
rect -2693 -11245 -2659 -11211
rect -2625 -11245 -2591 -11211
rect -2557 -11245 -2523 -11211
rect -2489 -11245 -2455 -11211
rect -2421 -11245 -2387 -11211
rect -2353 -11245 -2319 -11211
rect -2285 -11245 -2251 -11211
rect -2217 -11245 -2183 -11211
rect -2149 -11245 -2115 -11211
rect -2081 -11245 -2047 -11211
rect -2013 -11245 -1979 -11211
rect -1945 -11245 -1911 -11211
rect -1877 -11245 -1843 -11211
rect -1809 -11245 -1775 -11211
rect -1741 -11245 -1707 -11211
rect -1673 -11245 -1639 -11211
rect -1605 -11245 -1571 -11211
rect -1537 -11245 -1503 -11211
rect -1469 -11245 -1435 -11211
rect -1401 -11245 -1367 -11211
rect -1333 -11245 -1299 -11211
rect -1265 -11245 -1231 -11211
rect -1197 -11245 -1163 -11211
rect -1129 -11245 -1095 -11211
rect -1061 -11245 -1027 -11211
rect -993 -11245 -959 -11211
rect -925 -11245 -891 -11211
rect -857 -11245 -823 -11211
rect -789 -11245 -755 -11211
rect -721 -11245 -687 -11211
rect -653 -11245 -619 -11211
rect -585 -11245 -551 -11211
rect -517 -11245 -483 -11211
rect -449 -11245 -415 -11211
rect -381 -11245 -347 -11211
rect -313 -11245 -279 -11211
rect -245 -11245 -211 -11211
rect -177 -11245 -143 -11211
rect -109 -11245 -75 -11211
rect -41 -11245 -7 -11211
rect 27 -11245 61 -11211
rect 95 -11245 129 -11211
rect 163 -11245 197 -11211
rect 231 -11245 265 -11211
rect 299 -11245 333 -11211
rect 367 -11245 401 -11211
rect 435 -11245 469 -11211
rect 503 -11245 537 -11211
rect 571 -11245 605 -11211
rect 639 -11245 673 -11211
rect 707 -11245 741 -11211
rect 775 -11245 809 -11211
rect 843 -11245 877 -11211
rect 911 -11245 945 -11211
rect 979 -11245 1013 -11211
rect 1047 -11245 1081 -11211
rect 1115 -11245 1149 -11211
rect 1183 -11245 1217 -11211
rect 1251 -11245 1285 -11211
rect 1319 -11245 1353 -11211
rect 1387 -11245 1421 -11211
rect 1455 -11245 1489 -11211
rect 1523 -11245 1557 -11211
rect 1591 -11245 1625 -11211
rect 1659 -11245 1693 -11211
rect 1727 -11245 1761 -11211
rect 1795 -11245 1829 -11211
rect 1863 -11245 1897 -11211
rect 1931 -11245 1965 -11211
rect 1999 -11245 2033 -11211
rect 2067 -11245 2101 -11211
rect 2135 -11245 2169 -11211
rect 2203 -11245 2237 -11211
rect 2271 -11245 2305 -11211
rect 2339 -11245 2373 -11211
rect 2407 -11245 2441 -11211
rect 2475 -11245 2509 -11211
rect 2543 -11245 2577 -11211
rect 2611 -11245 2645 -11211
rect 2679 -11245 2713 -11211
rect 2747 -11245 2781 -11211
rect 2815 -11245 2849 -11211
rect 2883 -11245 2917 -11211
rect 2951 -11245 2985 -11211
rect 3019 -11245 3053 -11211
rect 3087 -11245 3121 -11211
rect 3155 -11245 3189 -11211
rect 3223 -11245 3257 -11211
rect 3291 -11245 3325 -11211
rect 3359 -11245 3393 -11211
rect 3427 -11245 3461 -11211
rect 3495 -11245 3529 -11211
rect 3563 -11245 3597 -11211
rect 3631 -11245 3665 -11211
rect 3699 -11245 3733 -11211
rect 3767 -11245 3801 -11211
rect 3835 -11245 3869 -11211
rect 3903 -11245 3937 -11211
rect 3971 -11245 4005 -11211
rect 4039 -11245 4073 -11211
rect 4107 -11245 4141 -11211
rect 4175 -11245 4209 -11211
rect 4243 -11245 4277 -11211
rect 4311 -11245 4345 -11211
rect 4379 -11245 4413 -11211
rect 4447 -11245 4481 -11211
rect 4515 -11245 4549 -11211
rect 4583 -11245 4617 -11211
rect 4651 -11245 4685 -11211
rect 4719 -11245 4753 -11211
rect 4787 -11245 4821 -11211
rect 4855 -11245 4889 -11211
rect 4923 -11245 4957 -11211
rect 4991 -11245 5025 -11211
rect 5059 -11245 5093 -11211
rect 5127 -11245 5161 -11211
rect 5195 -11245 5229 -11211
rect 5263 -11245 5297 -11211
rect 5331 -11245 5365 -11211
rect 5399 -11245 5433 -11211
rect 5467 -11245 5501 -11211
rect 5535 -11245 5569 -11211
rect 5603 -11245 5637 -11211
rect 5671 -11245 5705 -11211
rect 5739 -11245 5773 -11211
rect 5807 -11245 5841 -11211
rect 5875 -11245 5909 -11211
rect 5943 -11245 5977 -11211
rect 6011 -11245 6045 -11211
rect 6079 -11245 6113 -11211
rect 6147 -11245 6181 -11211
rect 6215 -11245 6249 -11211
rect 6283 -11245 6317 -11211
rect 6351 -11245 6385 -11211
rect 6419 -11245 6453 -11211
rect 6487 -11245 6521 -11211
rect 6555 -11245 6589 -11211
rect 6623 -11245 6657 -11211
rect 6691 -11245 6725 -11211
rect 6759 -11245 6793 -11211
rect 6827 -11245 6861 -11211
rect 6895 -11245 6929 -11211
rect 6963 -11245 6997 -11211
rect 7031 -11245 7065 -11211
rect 7099 -11245 7133 -11211
rect 7167 -11245 7201 -11211
rect 7235 -11245 7269 -11211
rect 7303 -11245 7337 -11211
rect 7371 -11245 7405 -11211
rect 7439 -11245 7473 -11211
rect 7507 -11245 7541 -11211
rect 7575 -11245 7609 -11211
rect 7643 -11245 7677 -11211
rect 7711 -11245 7745 -11211
rect 7779 -11245 7813 -11211
rect 7847 -11245 7881 -11211
rect 7915 -11245 7949 -11211
rect 7983 -11245 8017 -11211
rect 8051 -11245 8085 -11211
rect 8119 -11245 8153 -11211
rect 8187 -11245 8221 -11211
rect 8255 -11245 8289 -11211
rect 8323 -11245 8357 -11211
rect 8391 -11245 8425 -11211
rect 8459 -11245 8493 -11211
rect 8527 -11245 8561 -11211
rect 8595 -11245 8629 -11211
rect 8663 -11245 8697 -11211
rect 8731 -11245 8765 -11211
rect 8799 -11245 8833 -11211
rect 8867 -11245 8901 -11211
rect 8935 -11245 8969 -11211
rect 9003 -11245 9037 -11211
rect 9071 -11245 9105 -11211
rect 9139 -11245 9173 -11211
rect 9207 -11245 9241 -11211
rect 9275 -11245 9309 -11211
rect 9343 -11245 9377 -11211
rect 9411 -11245 9445 -11211
rect 9479 -11245 9513 -11211
rect 9547 -11245 9581 -11211
rect 9615 -11245 9649 -11211
rect 9683 -11245 9717 -11211
rect 9751 -11245 9785 -11211
rect 9819 -11245 9853 -11211
rect 9887 -11245 9921 -11211
rect 9955 -11245 9989 -11211
rect 10023 -11245 10057 -11211
rect 10091 -11245 10125 -11211
rect 10159 -11245 10193 -11211
rect 10227 -11245 10261 -11211
rect 10295 -11245 10329 -11211
rect 10363 -11245 10397 -11211
rect 10431 -11245 10465 -11211
rect 10499 -11245 10533 -11211
rect 10567 -11245 10601 -11211
rect 10635 -11245 10669 -11211
rect 10703 -11245 10737 -11211
rect 10771 -11245 10805 -11211
rect 10839 -11245 10873 -11211
rect 10907 -11245 10941 -11211
rect 10975 -11245 11009 -11211
rect 11043 -11245 11077 -11211
rect 11111 -11245 11145 -11211
rect 11179 -11245 11213 -11211
rect 11247 -11245 11281 -11211
rect 11315 -11245 11349 -11211
rect 11383 -11245 11417 -11211
rect 11451 -11245 11485 -11211
rect 11519 -11245 11553 -11211
rect 11587 -11245 11621 -11211
rect 11655 -11245 11689 -11211
rect 11723 -11245 11757 -11211
rect 11791 -11245 11825 -11211
rect 11859 -11245 11893 -11211
rect 11927 -11245 11961 -11211
rect 11995 -11245 12029 -11211
rect 12063 -11245 12097 -11211
rect 12131 -11245 12165 -11211
rect 12199 -11245 12233 -11211
rect 12267 -11245 12301 -11211
rect 12335 -11245 12369 -11211
rect 12403 -11245 12437 -11211
rect 12471 -11245 12505 -11211
rect 12539 -11245 12573 -11211
rect 12607 -11245 12641 -11211
rect 12675 -11245 12709 -11211
rect 12743 -11245 12777 -11211
rect 12811 -11245 12845 -11211
rect 12879 -11245 12913 -11211
rect 12947 -11245 12981 -11211
rect 13015 -11245 13049 -11211
rect 13083 -11245 13117 -11211
rect 13151 -11245 13185 -11211
rect 13219 -11245 13253 -11211
rect 13287 -11245 13321 -11211
rect 13355 -11245 13389 -11211
rect 13423 -11245 13457 -11211
rect 13491 -11245 13525 -11211
rect 13559 -11245 13593 -11211
rect 13627 -11245 13661 -11211
rect 13695 -11245 13729 -11211
rect 13763 -11245 13797 -11211
rect 13831 -11245 13865 -11211
rect 13899 -11245 13933 -11211
rect 13967 -11245 14001 -11211
rect 14035 -11245 14069 -11211
rect 14103 -11245 14137 -11211
rect 14171 -11245 14205 -11211
rect 14239 -11245 14273 -11211
rect 14307 -11245 14341 -11211
rect 14375 -11245 14409 -11211
rect 14443 -11245 14477 -11211
rect 14511 -11245 14545 -11211
rect 14579 -11245 14613 -11211
rect 14647 -11245 14681 -11211
rect 14715 -11245 14749 -11211
rect 14783 -11245 14817 -11211
rect 14851 -11245 14885 -11211
rect 14919 -11245 14953 -11211
rect 14987 -11245 15021 -11211
rect 15055 -11245 15089 -11211
rect 15123 -11245 15157 -11211
rect 15191 -11245 15225 -11211
rect 15259 -11245 15293 -11211
rect 15327 -11245 15361 -11211
rect 15395 -11245 15429 -11211
rect 15463 -11245 15497 -11211
rect 15531 -11245 15565 -11211
rect 15599 -11245 15633 -11211
rect 15667 -11245 15701 -11211
rect 15735 -11245 15769 -11211
rect 15803 -11245 15837 -11211
rect 15871 -11245 15905 -11211
rect 15939 -11245 15973 -11211
rect 16007 -11245 16041 -11211
rect 16075 -11245 16109 -11211
rect 16143 -11245 16177 -11211
rect 16211 -11245 16245 -11211
rect 16279 -11245 16313 -11211
rect 16347 -11245 16381 -11211
rect 16415 -11245 16449 -11211
rect 16483 -11245 16517 -11211
rect 16551 -11245 16585 -11211
rect 16619 -11245 16653 -11211
rect 16687 -11245 16721 -11211
rect 16755 -11245 16789 -11211
rect 16823 -11245 16857 -11211
rect 16891 -11245 16925 -11211
rect 16959 -11245 16993 -11211
rect 17027 -11245 17061 -11211
rect 17095 -11245 17129 -11211
rect 17163 -11245 17197 -11211
rect 17231 -11245 17265 -11211
rect 17299 -11245 17333 -11211
rect 17367 -11245 17401 -11211
rect 17435 -11245 17469 -11211
rect 17503 -11245 17537 -11211
rect 17571 -11245 17605 -11211
rect 17639 -11245 17673 -11211
rect 17707 -11245 17741 -11211
rect 17775 -11245 17809 -11211
rect 17843 -11245 17877 -11211
rect 17911 -11245 17945 -11211
rect 17979 -11245 18013 -11211
rect 18047 -11245 18081 -11211
rect 18115 -11245 18149 -11211
rect 18183 -11245 18217 -11211
rect 18251 -11245 18285 -11211
rect 18319 -11245 18353 -11211
rect 18387 -11245 18421 -11211
rect 18455 -11245 18489 -11211
rect 18523 -11245 18557 -11211
rect 18591 -11245 18625 -11211
rect 18659 -11245 18693 -11211
rect 18727 -11245 18761 -11211
rect 18795 -11245 18829 -11211
rect 18863 -11245 18897 -11211
rect 18931 -11245 18965 -11211
rect 18999 -11245 19033 -11211
rect 19067 -11245 19101 -11211
rect 19135 -11245 19169 -11211
rect 19203 -11245 19237 -11211
rect 19271 -11245 19305 -11211
rect 19339 -11245 19373 -11211
rect 19407 -11245 19441 -11211
rect 19475 -11245 19509 -11211
rect 19543 -11245 19577 -11211
rect 19611 -11245 19645 -11211
rect 19679 -11245 19713 -11211
rect 19747 -11245 19781 -11211
rect 19815 -11245 19849 -11211
rect 19883 -11245 19917 -11211
rect 19951 -11245 19985 -11211
rect 20019 -11245 20053 -11211
rect 20087 -11245 20121 -11211
rect 20155 -11245 20189 -11211
rect 20223 -11245 20257 -11211
rect 20291 -11245 20325 -11211
rect 20359 -11245 20393 -11211
rect 20427 -11245 20461 -11211
rect 20495 -11245 20529 -11211
rect 20563 -11245 20597 -11211
rect 20631 -11245 20665 -11211
rect 20699 -11245 20733 -11211
rect 20767 -11245 20801 -11211
rect 20835 -11245 20869 -11211
rect 20903 -11245 20937 -11211
rect 20971 -11245 21005 -11211
rect 21039 -11245 21073 -11211
rect 21107 -11245 21141 -11211
rect 21175 -11245 21209 -11211
rect 21243 -11245 21277 -11211
rect 21311 -11245 21345 -11211
rect 21379 -11245 21413 -11211
rect 21447 -11245 21481 -11211
rect 21515 -11245 21549 -11211
rect 21583 -11245 21617 -11211
rect 21651 -11245 21685 -11211
rect 21719 -11245 21753 -11211
rect 21787 -11245 21821 -11211
rect 21855 -11245 21889 -11211
rect 21923 -11245 21957 -11211
rect 21991 -11245 22025 -11211
rect 22059 -11245 22093 -11211
rect 22127 -11245 22161 -11211
rect 22195 -11245 22229 -11211
rect 22263 -11245 22297 -11211
rect 22331 -11245 22365 -11211
rect 22399 -11245 22433 -11211
rect 22467 -11245 22501 -11211
rect 22535 -11245 22569 -11211
rect 22603 -11245 22637 -11211
rect 22671 -11245 22705 -11211
rect 22739 -11245 22773 -11211
rect 22807 -11245 22841 -11211
rect 22875 -11245 22909 -11211
rect 22943 -11245 22977 -11211
rect 23011 -11245 23045 -11211
rect 23079 -11245 23113 -11211
rect 23147 -11245 23181 -11211
rect 23215 -11245 23249 -11211
rect 23283 -11245 23317 -11211
rect 23351 -11245 23385 -11211
rect 23419 -11245 23453 -11211
rect 23487 -11245 23521 -11211
rect 23555 -11245 23589 -11211
rect 23623 -11245 23657 -11211
rect 23691 -11245 23725 -11211
rect 23759 -11245 23793 -11211
rect 23827 -11245 23861 -11211
rect 23895 -11245 23929 -11211
rect 23963 -11245 23997 -11211
rect 24031 -11245 24065 -11211
rect 24099 -11245 24133 -11211
rect 24167 -11245 24201 -11211
rect 24235 -11245 24269 -11211
rect 24303 -11245 24337 -11211
rect 24371 -11245 24405 -11211
rect 24439 -11245 24473 -11211
rect 24507 -11245 24541 -11211
rect 24575 -11245 24609 -11211
rect 24643 -11245 24677 -11211
rect 24711 -11245 24745 -11211
rect -12289 -11397 -12255 -11363
rect -12289 -11465 -12255 -11431
rect -12289 -11533 -12255 -11499
rect -12289 -11601 -12255 -11567
rect -12289 -11669 -12255 -11635
rect -12289 -11737 -12255 -11703
rect -12289 -11805 -12255 -11771
rect -12289 -11873 -12255 -11839
rect -12289 -11941 -12255 -11907
rect -12289 -12009 -12255 -11975
rect -12289 -12077 -12255 -12043
rect -12289 -12145 -12255 -12111
rect -12289 -12213 -12255 -12179
rect -12289 -12281 -12255 -12247
rect -12289 -12349 -12255 -12315
rect -12289 -12417 -12255 -12383
rect 24855 -11397 24889 -11363
rect 24855 -11465 24889 -11431
rect 24855 -11533 24889 -11499
rect 24855 -11601 24889 -11567
rect 24855 -11669 24889 -11635
rect 24855 -11737 24889 -11703
rect 24855 -11805 24889 -11771
rect 24855 -11873 24889 -11839
rect 24855 -11941 24889 -11907
rect 24855 -12009 24889 -11975
rect 24855 -12077 24889 -12043
rect 24855 -12145 24889 -12111
rect 24855 -12213 24889 -12179
rect 24855 -12281 24889 -12247
rect 24855 -12349 24889 -12315
rect 24855 -12417 24889 -12383
rect -12289 -12485 -12255 -12451
rect 24855 -12485 24889 -12451
rect -12289 -12553 -12255 -12519
rect -12289 -12621 -12255 -12587
rect -12289 -12689 -12255 -12655
rect -12289 -12757 -12255 -12723
rect -12289 -12825 -12255 -12791
rect -12289 -12893 -12255 -12859
rect -12289 -12961 -12255 -12927
rect -12289 -13029 -12255 -12995
rect -12289 -13097 -12255 -13063
rect 24855 -12553 24889 -12519
rect 24855 -12621 24889 -12587
rect 24855 -12689 24889 -12655
rect 24855 -12757 24889 -12723
rect 24855 -12825 24889 -12791
rect 24855 -12893 24889 -12859
rect 24855 -12961 24889 -12927
rect 24855 -13029 24889 -12995
rect 24855 -13097 24889 -13063
rect -12289 -13165 -12255 -13131
rect -12289 -13233 -12255 -13199
rect 24855 -13165 24889 -13131
rect 24855 -13233 24889 -13199
rect -12289 -13301 -12255 -13267
rect 24855 -13301 24889 -13267
rect -12289 -13369 -12255 -13335
rect -12289 -13437 -12255 -13403
rect -12289 -13505 -12255 -13471
rect -12289 -13573 -12255 -13539
rect -12289 -13641 -12255 -13607
rect -12289 -13709 -12255 -13675
rect -12289 -13777 -12255 -13743
rect -12289 -13845 -12255 -13811
rect -12289 -13913 -12255 -13879
rect 24855 -13369 24889 -13335
rect 24855 -13437 24889 -13403
rect 24855 -13505 24889 -13471
rect 24855 -13573 24889 -13539
rect 24855 -13641 24889 -13607
rect 24855 -13709 24889 -13675
rect 24855 -13777 24889 -13743
rect 24855 -13845 24889 -13811
rect 24855 -13913 24889 -13879
rect -12289 -13981 -12255 -13947
rect -12289 -14049 -12255 -14015
rect 24855 -13981 24889 -13947
rect 24855 -14049 24889 -14015
rect -12289 -14117 -12255 -14083
rect 24855 -14117 24889 -14083
rect -12289 -14185 -12255 -14151
rect -12289 -14253 -12255 -14219
rect -12289 -14321 -12255 -14287
rect -12289 -14389 -12255 -14355
rect -12289 -14457 -12255 -14423
rect -12289 -14525 -12255 -14491
rect -12289 -14593 -12255 -14559
rect -12289 -14661 -12255 -14627
rect -12289 -14729 -12255 -14695
rect 24855 -14185 24889 -14151
rect -12289 -14797 -12255 -14763
rect -12289 -14865 -12255 -14831
rect 24855 -14253 24889 -14219
rect 24855 -14321 24889 -14287
rect 24855 -14389 24889 -14355
rect 24855 -14457 24889 -14423
rect 24855 -14525 24889 -14491
rect 24855 -14593 24889 -14559
rect 24855 -14661 24889 -14627
rect 24855 -14729 24889 -14695
rect 24855 -14797 24889 -14763
rect -12289 -14933 -12255 -14899
rect 24855 -14865 24889 -14831
rect 24855 -14933 24889 -14899
rect -12289 -15001 -12255 -14967
rect -12289 -15069 -12255 -15035
rect -12289 -15137 -12255 -15103
rect -12289 -15205 -12255 -15171
rect -12289 -15273 -12255 -15239
rect -12289 -15341 -12255 -15307
rect -12289 -15409 -12255 -15375
rect -12289 -15477 -12255 -15443
rect -12289 -15545 -12255 -15511
rect 24855 -15001 24889 -14967
rect 24855 -15069 24889 -15035
rect 24855 -15137 24889 -15103
rect 24855 -15205 24889 -15171
rect 24855 -15273 24889 -15239
rect 24855 -15341 24889 -15307
rect 24855 -15409 24889 -15375
rect -12289 -15613 -12255 -15579
rect -12289 -15681 -12255 -15647
rect -12289 -15749 -12255 -15715
rect -12289 -15817 -12255 -15783
rect -12289 -15885 -12255 -15851
rect -12289 -15953 -12255 -15919
rect -12289 -16021 -12255 -15987
rect -12289 -16089 -12255 -16055
rect -12289 -16157 -12255 -16123
rect -12289 -16225 -12255 -16191
rect -12289 -16293 -12255 -16259
rect -12289 -16361 -12255 -16327
rect 24855 -15477 24889 -15443
rect 24855 -15545 24889 -15511
rect 24855 -15613 24889 -15579
rect 24855 -15681 24889 -15647
rect 24855 -15749 24889 -15715
rect 24855 -15817 24889 -15783
rect 24855 -15885 24889 -15851
rect 24855 -15953 24889 -15919
rect 24855 -16021 24889 -15987
rect 24855 -16089 24889 -16055
rect 24855 -16157 24889 -16123
rect 24855 -16225 24889 -16191
rect 24855 -16293 24889 -16259
rect 24855 -16361 24889 -16327
rect -12289 -16429 -12255 -16395
rect -12289 -16497 -12255 -16463
rect 24855 -16429 24889 -16395
rect 24855 -16497 24889 -16463
rect -12289 -16565 -12255 -16531
rect -12289 -16633 -12255 -16599
rect 24855 -16565 24889 -16531
rect -12289 -16701 -12255 -16667
rect -12289 -16769 -12255 -16735
rect -12289 -16837 -12255 -16803
rect -12289 -16905 -12255 -16871
rect -12289 -16973 -12255 -16939
rect -12289 -17041 -12255 -17007
rect -12289 -17109 -12255 -17075
rect -12289 -17177 -12255 -17143
rect 24855 -16633 24889 -16599
rect -12289 -17245 -12255 -17211
rect -12289 -17313 -12255 -17279
rect 24855 -16701 24889 -16667
rect 24855 -16769 24889 -16735
rect 24855 -16837 24889 -16803
rect 24855 -16905 24889 -16871
rect 24855 -16973 24889 -16939
rect 24855 -17041 24889 -17007
rect 24855 -17109 24889 -17075
rect 24855 -17177 24889 -17143
rect 24855 -17245 24889 -17211
rect -12289 -17381 -12255 -17347
rect -12289 -17449 -12255 -17415
rect 24855 -17313 24889 -17279
rect 24855 -17381 24889 -17347
rect -12289 -17517 -12255 -17483
rect -12289 -17585 -12255 -17551
rect -12289 -17653 -12255 -17619
rect -12289 -17721 -12255 -17687
rect -12289 -17789 -12255 -17755
rect -12289 -17857 -12255 -17823
rect -12289 -17925 -12255 -17891
rect -12289 -17993 -12255 -17959
rect 24855 -17449 24889 -17415
rect 24855 -17517 24889 -17483
rect 24855 -17585 24889 -17551
rect 24855 -17653 24889 -17619
rect 24855 -17721 24889 -17687
rect 24855 -17789 24889 -17755
rect 24855 -17857 24889 -17823
rect 24855 -17925 24889 -17891
rect -12289 -18061 -12255 -18027
rect -12289 -18129 -12255 -18095
rect -12289 -18197 -12255 -18163
rect -12289 -18265 -12255 -18231
rect -12289 -18333 -12255 -18299
rect -12289 -18401 -12255 -18367
rect -12289 -18469 -12255 -18435
rect -12289 -18537 -12255 -18503
rect -12289 -18605 -12255 -18571
rect -12289 -18673 -12255 -18639
rect -12289 -18741 -12255 -18707
rect -12289 -18809 -12255 -18775
rect 24855 -17993 24889 -17959
rect 24855 -18061 24889 -18027
rect 24855 -18129 24889 -18095
rect 24855 -18197 24889 -18163
rect 24855 -18265 24889 -18231
rect 24855 -18333 24889 -18299
rect 24855 -18401 24889 -18367
rect 24855 -18469 24889 -18435
rect 24855 -18537 24889 -18503
rect 24855 -18605 24889 -18571
rect 24855 -18673 24889 -18639
rect 24855 -18741 24889 -18707
rect 24855 -18809 24889 -18775
rect -12289 -18877 -12255 -18843
rect -12289 -18945 -12255 -18911
rect 24855 -18877 24889 -18843
rect -12289 -19013 -12255 -18979
rect -12289 -19081 -12255 -19047
rect 24855 -18945 24889 -18911
rect 24855 -19013 24889 -18979
rect -12289 -19149 -12255 -19115
rect 24855 -19081 24889 -19047
rect 24855 -19149 24889 -19115
rect -12289 -19217 -12255 -19183
rect -12289 -19285 -12255 -19251
rect -12289 -19353 -12255 -19319
rect -12289 -19421 -12255 -19387
rect -12289 -19489 -12255 -19455
rect -12289 -19557 -12255 -19523
rect -12289 -19625 -12255 -19591
rect -12289 -19693 -12255 -19659
rect -12289 -19761 -12255 -19727
rect 24855 -19217 24889 -19183
rect 24855 -19285 24889 -19251
rect 24855 -19353 24889 -19319
rect 24855 -19421 24889 -19387
rect 24855 -19489 24889 -19455
rect 24855 -19557 24889 -19523
rect 24855 -19625 24889 -19591
rect 24855 -19693 24889 -19659
rect 24855 -19761 24889 -19727
rect -12289 -19829 -12255 -19795
rect 24855 -19829 24889 -19795
rect -12289 -19897 -12255 -19863
rect -12289 -19965 -12255 -19931
rect -12289 -20033 -12255 -19999
rect -12289 -20101 -12255 -20067
rect -12289 -20169 -12255 -20135
rect -12289 -20237 -12255 -20203
rect -12289 -20305 -12255 -20271
rect 24855 -19897 24889 -19863
rect 24855 -19965 24889 -19931
rect 24855 -20033 24889 -19999
rect 24855 -20101 24889 -20067
rect 24855 -20169 24889 -20135
rect 24855 -20237 24889 -20203
rect 24855 -20305 24889 -20271
rect -12289 -20373 -12255 -20339
rect 24855 -20373 24889 -20339
rect -12289 -20441 -12255 -20407
rect -12289 -20509 -12255 -20475
rect -12289 -20577 -12255 -20543
rect -12289 -20645 -12255 -20611
rect -12289 -20713 -12255 -20679
rect -12289 -20781 -12255 -20747
rect -12289 -20849 -12255 -20815
rect -12289 -20917 -12255 -20883
rect -12289 -20985 -12255 -20951
rect 24855 -20441 24889 -20407
rect 24855 -20509 24889 -20475
rect 24855 -20577 24889 -20543
rect 24855 -20645 24889 -20611
rect 24855 -20713 24889 -20679
rect 24855 -20781 24889 -20747
rect 24855 -20849 24889 -20815
rect 24855 -20917 24889 -20883
rect 24855 -20985 24889 -20951
rect -12289 -21053 -12255 -21019
rect 24855 -21053 24889 -21019
rect -12289 -21121 -12255 -21087
rect -12289 -21189 -12255 -21155
rect -12289 -21257 -12255 -21223
rect -12289 -21325 -12255 -21291
rect -12289 -21393 -12255 -21359
rect -12289 -21461 -12255 -21427
rect -12289 -21529 -12255 -21495
rect 24855 -21121 24889 -21087
rect 24855 -21189 24889 -21155
rect 24855 -21257 24889 -21223
rect 24855 -21325 24889 -21291
rect 24855 -21393 24889 -21359
rect 24855 -21461 24889 -21427
rect 24855 -21529 24889 -21495
rect -12289 -21597 -12255 -21563
rect -12289 -21665 -12255 -21631
rect 24855 -21597 24889 -21563
rect -12289 -21733 -12255 -21699
rect -12289 -21801 -12255 -21767
rect -12289 -21869 -12255 -21835
rect -12289 -21937 -12255 -21903
rect -12289 -22005 -12255 -21971
rect -12289 -22073 -12255 -22039
rect -12289 -22141 -12255 -22107
rect -12289 -22209 -12255 -22175
rect 24855 -21665 24889 -21631
rect 24855 -21733 24889 -21699
rect 24855 -21801 24889 -21767
rect 24855 -21869 24889 -21835
rect 24855 -21937 24889 -21903
rect 24855 -22005 24889 -21971
rect 24855 -22073 24889 -22039
rect 24855 -22141 24889 -22107
rect 24855 -22209 24889 -22175
rect -12289 -22277 -12255 -22243
rect -12289 -22345 -12255 -22311
rect 24855 -22277 24889 -22243
rect -12289 -22413 -12255 -22379
rect -12289 -22481 -12255 -22447
rect -12289 -22549 -12255 -22515
rect -12289 -22617 -12255 -22583
rect -12289 -22685 -12255 -22651
rect -12289 -22753 -12255 -22719
rect 24855 -22345 24889 -22311
rect 24855 -22413 24889 -22379
rect 24855 -22481 24889 -22447
rect 24855 -22549 24889 -22515
rect 24855 -22617 24889 -22583
rect 24855 -22685 24889 -22651
rect 24855 -22753 24889 -22719
rect -12289 -22821 -12255 -22787
rect -12289 -22889 -12255 -22855
rect 24855 -22821 24889 -22787
rect -12289 -22957 -12255 -22923
rect -12289 -23025 -12255 -22991
rect -12289 -23093 -12255 -23059
rect -12289 -23161 -12255 -23127
rect -12289 -23229 -12255 -23195
rect -12289 -23297 -12255 -23263
rect -12289 -23365 -12255 -23331
rect -12289 -23433 -12255 -23399
rect 24855 -22889 24889 -22855
rect 24855 -22957 24889 -22923
rect 24855 -23025 24889 -22991
rect 24855 -23093 24889 -23059
rect 24855 -23161 24889 -23127
rect 24855 -23229 24889 -23195
rect 24855 -23297 24889 -23263
rect 24855 -23365 24889 -23331
rect 24855 -23433 24889 -23399
rect -12289 -23501 -12255 -23467
rect -12289 -23569 -12255 -23535
rect 24855 -23501 24889 -23467
rect -12289 -23637 -12255 -23603
rect -12289 -23705 -12255 -23671
rect -12289 -23773 -12255 -23739
rect -12289 -23841 -12255 -23807
rect -12289 -23909 -12255 -23875
rect -12289 -23977 -12255 -23943
rect 24855 -23569 24889 -23535
rect 24855 -23637 24889 -23603
rect 24855 -23705 24889 -23671
rect 24855 -23773 24889 -23739
rect 24855 -23841 24889 -23807
rect 24855 -23909 24889 -23875
rect 24855 -23977 24889 -23943
rect -12289 -24045 -12255 -24011
rect -12289 -24113 -12255 -24079
rect 24855 -24045 24889 -24011
rect -12289 -24181 -12255 -24147
rect -12289 -24249 -12255 -24215
rect -12289 -24317 -12255 -24283
rect -12289 -24385 -12255 -24351
rect -12289 -24453 -12255 -24419
rect -12289 -24521 -12255 -24487
rect -12289 -24589 -12255 -24555
rect -12289 -24657 -12255 -24623
rect -12289 -24725 -12255 -24691
rect 24855 -24113 24889 -24079
rect 24855 -24181 24889 -24147
rect 24855 -24249 24889 -24215
rect 24855 -24317 24889 -24283
rect 24855 -24385 24889 -24351
rect 24855 -24453 24889 -24419
rect 24855 -24521 24889 -24487
rect 24855 -24589 24889 -24555
rect 24855 -24657 24889 -24623
rect -12289 -24793 -12255 -24759
rect 24855 -24725 24889 -24691
rect -12289 -24861 -12255 -24827
rect -12289 -24929 -12255 -24895
rect -12289 -24997 -12255 -24963
rect -12289 -25065 -12255 -25031
rect -12289 -25133 -12255 -25099
rect -12289 -25201 -12255 -25167
rect -12289 -25269 -12255 -25235
rect -12289 -25337 -12255 -25303
rect -12289 -25405 -12255 -25371
rect -12289 -25473 -12255 -25439
rect -12289 -25541 -12255 -25507
rect -12289 -25609 -12255 -25575
rect -12289 -25677 -12255 -25643
rect -12289 -25745 -12255 -25711
rect -12289 -25813 -12255 -25779
rect -12289 -25881 -12255 -25847
rect -12289 -25949 -12255 -25915
rect -12289 -26017 -12255 -25983
rect -12289 -26085 -12255 -26051
rect -12289 -26153 -12255 -26119
rect -12289 -26221 -12255 -26187
rect -12289 -26289 -12255 -26255
rect -12289 -26357 -12255 -26323
rect -12289 -26425 -12255 -26391
rect -12289 -26493 -12255 -26459
rect -12289 -26561 -12255 -26527
rect -12289 -26629 -12255 -26595
rect -12289 -26697 -12255 -26663
rect -12289 -26765 -12255 -26731
rect -12289 -26833 -12255 -26799
rect -12289 -26901 -12255 -26867
rect -12289 -26969 -12255 -26935
rect -12289 -27037 -12255 -27003
rect 24855 -24793 24889 -24759
rect 24855 -24861 24889 -24827
rect 24855 -24929 24889 -24895
rect 24855 -24997 24889 -24963
rect 24855 -25065 24889 -25031
rect 24855 -25133 24889 -25099
rect 24855 -25201 24889 -25167
rect 24855 -25269 24889 -25235
rect 24855 -25337 24889 -25303
rect 24855 -25405 24889 -25371
rect 24855 -25473 24889 -25439
rect 24855 -25541 24889 -25507
rect 24855 -25609 24889 -25575
rect 24855 -25677 24889 -25643
rect 24855 -25745 24889 -25711
rect 24855 -25813 24889 -25779
rect 24855 -25881 24889 -25847
rect 24855 -25949 24889 -25915
rect 24855 -26017 24889 -25983
rect 24855 -26085 24889 -26051
rect 24855 -26153 24889 -26119
rect 24855 -26221 24889 -26187
rect 24855 -26289 24889 -26255
rect 24855 -26357 24889 -26323
rect 24855 -26425 24889 -26391
rect 24855 -26493 24889 -26459
rect 24855 -26561 24889 -26527
rect 24855 -26629 24889 -26595
rect 24855 -26697 24889 -26663
rect 24855 -26765 24889 -26731
rect 24855 -26833 24889 -26799
rect 24855 -26901 24889 -26867
rect 24855 -26969 24889 -26935
rect 24855 -27037 24889 -27003
rect -12145 -27189 -12111 -27155
rect -12077 -27189 -12043 -27155
rect -12009 -27189 -11975 -27155
rect -11941 -27189 -11907 -27155
rect -11873 -27189 -11839 -27155
rect -11805 -27189 -11771 -27155
rect -11737 -27189 -11703 -27155
rect -11669 -27189 -11635 -27155
rect -11601 -27189 -11567 -27155
rect -11533 -27189 -11499 -27155
rect -11465 -27189 -11431 -27155
rect -11397 -27189 -11363 -27155
rect -11329 -27189 -11295 -27155
rect -11261 -27189 -11227 -27155
rect -11193 -27189 -11159 -27155
rect -11125 -27189 -11091 -27155
rect -11057 -27189 -11023 -27155
rect -10989 -27189 -10955 -27155
rect -10921 -27189 -10887 -27155
rect -10853 -27189 -10819 -27155
rect -10785 -27189 -10751 -27155
rect -10717 -27189 -10683 -27155
rect -10649 -27189 -10615 -27155
rect -10581 -27189 -10547 -27155
rect -10513 -27189 -10479 -27155
rect -10445 -27189 -10411 -27155
rect -10377 -27189 -10343 -27155
rect -10309 -27189 -10275 -27155
rect -10241 -27189 -10207 -27155
rect -10173 -27189 -10139 -27155
rect -10105 -27189 -10071 -27155
rect -10037 -27189 -10003 -27155
rect -9969 -27189 -9935 -27155
rect -9901 -27189 -9867 -27155
rect -9833 -27189 -9799 -27155
rect -9765 -27189 -9731 -27155
rect -9697 -27189 -9663 -27155
rect -9629 -27189 -9595 -27155
rect -9561 -27189 -9527 -27155
rect -9493 -27189 -9459 -27155
rect -9425 -27189 -9391 -27155
rect -9357 -27189 -9323 -27155
rect -9289 -27189 -9255 -27155
rect -9221 -27189 -9187 -27155
rect -9153 -27189 -9119 -27155
rect -9085 -27189 -9051 -27155
rect -9017 -27189 -8983 -27155
rect -8949 -27189 -8915 -27155
rect -8881 -27189 -8847 -27155
rect -8813 -27189 -8779 -27155
rect -8745 -27189 -8711 -27155
rect -8677 -27189 -8643 -27155
rect -8609 -27189 -8575 -27155
rect -8541 -27189 -8507 -27155
rect -8473 -27189 -8439 -27155
rect -8405 -27189 -8371 -27155
rect -8337 -27189 -8303 -27155
rect -8269 -27189 -8235 -27155
rect -8201 -27189 -8167 -27155
rect -8133 -27189 -8099 -27155
rect -8065 -27189 -8031 -27155
rect -7997 -27189 -7963 -27155
rect -7929 -27189 -7895 -27155
rect -7861 -27189 -7827 -27155
rect -7793 -27189 -7759 -27155
rect -7725 -27189 -7691 -27155
rect -7657 -27189 -7623 -27155
rect -7589 -27189 -7555 -27155
rect -7521 -27189 -7487 -27155
rect -7453 -27189 -7419 -27155
rect -7385 -27189 -7351 -27155
rect -7317 -27189 -7283 -27155
rect -7249 -27189 -7215 -27155
rect -7181 -27189 -7147 -27155
rect -7113 -27189 -7079 -27155
rect -7045 -27189 -7011 -27155
rect -6977 -27189 -6943 -27155
rect -6909 -27189 -6875 -27155
rect -6841 -27189 -6807 -27155
rect -6773 -27189 -6739 -27155
rect -6705 -27189 -6671 -27155
rect -6637 -27189 -6603 -27155
rect -6569 -27189 -6535 -27155
rect -6501 -27189 -6467 -27155
rect -6433 -27189 -6399 -27155
rect -6365 -27189 -6331 -27155
rect -6297 -27189 -6263 -27155
rect -6229 -27189 -6195 -27155
rect -6161 -27189 -6127 -27155
rect -6093 -27189 -6059 -27155
rect -6025 -27189 -5991 -27155
rect -5957 -27189 -5923 -27155
rect -5889 -27189 -5855 -27155
rect -5821 -27189 -5787 -27155
rect -5753 -27189 -5719 -27155
rect -5685 -27189 -5651 -27155
rect -5617 -27189 -5583 -27155
rect -5549 -27189 -5515 -27155
rect -5481 -27189 -5447 -27155
rect -5413 -27189 -5379 -27155
rect -5345 -27189 -5311 -27155
rect -5277 -27189 -5243 -27155
rect -5209 -27189 -5175 -27155
rect -5141 -27189 -5107 -27155
rect -5073 -27189 -5039 -27155
rect -5005 -27189 -4971 -27155
rect -4937 -27189 -4903 -27155
rect -4869 -27189 -4835 -27155
rect -4801 -27189 -4767 -27155
rect -4733 -27189 -4699 -27155
rect -4665 -27189 -4631 -27155
rect -4597 -27189 -4563 -27155
rect -4529 -27189 -4495 -27155
rect -4461 -27189 -4427 -27155
rect -4393 -27189 -4359 -27155
rect -4325 -27189 -4291 -27155
rect -4257 -27189 -4223 -27155
rect -4189 -27189 -4155 -27155
rect -4121 -27189 -4087 -27155
rect -4053 -27189 -4019 -27155
rect -3985 -27189 -3951 -27155
rect -3917 -27189 -3883 -27155
rect -3849 -27189 -3815 -27155
rect -3781 -27189 -3747 -27155
rect -3713 -27189 -3679 -27155
rect -3645 -27189 -3611 -27155
rect -3577 -27189 -3543 -27155
rect -3509 -27189 -3475 -27155
rect -3441 -27189 -3407 -27155
rect -3373 -27189 -3339 -27155
rect -3305 -27189 -3271 -27155
rect -3237 -27189 -3203 -27155
rect -3169 -27189 -3135 -27155
rect -3101 -27189 -3067 -27155
rect -3033 -27189 -2999 -27155
rect -2965 -27189 -2931 -27155
rect -2897 -27189 -2863 -27155
rect -2829 -27189 -2795 -27155
rect -2761 -27189 -2727 -27155
rect -2693 -27189 -2659 -27155
rect -2625 -27189 -2591 -27155
rect -2557 -27189 -2523 -27155
rect -2489 -27189 -2455 -27155
rect -2421 -27189 -2387 -27155
rect -2353 -27189 -2319 -27155
rect -2285 -27189 -2251 -27155
rect -2217 -27189 -2183 -27155
rect -2149 -27189 -2115 -27155
rect -2081 -27189 -2047 -27155
rect -2013 -27189 -1979 -27155
rect -1945 -27189 -1911 -27155
rect -1877 -27189 -1843 -27155
rect -1809 -27189 -1775 -27155
rect -1741 -27189 -1707 -27155
rect -1673 -27189 -1639 -27155
rect -1605 -27189 -1571 -27155
rect -1537 -27189 -1503 -27155
rect -1469 -27189 -1435 -27155
rect -1401 -27189 -1367 -27155
rect -1333 -27189 -1299 -27155
rect -1265 -27189 -1231 -27155
rect -1197 -27189 -1163 -27155
rect -1129 -27189 -1095 -27155
rect -1061 -27189 -1027 -27155
rect -993 -27189 -959 -27155
rect -925 -27189 -891 -27155
rect -857 -27189 -823 -27155
rect -789 -27189 -755 -27155
rect -721 -27189 -687 -27155
rect -653 -27189 -619 -27155
rect -585 -27189 -551 -27155
rect -517 -27189 -483 -27155
rect -449 -27189 -415 -27155
rect -381 -27189 -347 -27155
rect -313 -27189 -279 -27155
rect -245 -27189 -211 -27155
rect -177 -27189 -143 -27155
rect -109 -27189 -75 -27155
rect -41 -27189 -7 -27155
rect 27 -27189 61 -27155
rect 95 -27189 129 -27155
rect 163 -27189 197 -27155
rect 231 -27189 265 -27155
rect 299 -27189 333 -27155
rect 367 -27189 401 -27155
rect 435 -27189 469 -27155
rect 503 -27189 537 -27155
rect 571 -27189 605 -27155
rect 639 -27189 673 -27155
rect 707 -27189 741 -27155
rect 775 -27189 809 -27155
rect 843 -27189 877 -27155
rect 911 -27189 945 -27155
rect 979 -27189 1013 -27155
rect 1047 -27189 1081 -27155
rect 1115 -27189 1149 -27155
rect 1183 -27189 1217 -27155
rect 1251 -27189 1285 -27155
rect 1319 -27189 1353 -27155
rect 1387 -27189 1421 -27155
rect 1455 -27189 1489 -27155
rect 1523 -27189 1557 -27155
rect 1591 -27189 1625 -27155
rect 1659 -27189 1693 -27155
rect 1727 -27189 1761 -27155
rect 1795 -27189 1829 -27155
rect 1863 -27189 1897 -27155
rect 1931 -27189 1965 -27155
rect 1999 -27189 2033 -27155
rect 2067 -27189 2101 -27155
rect 2135 -27189 2169 -27155
rect 2203 -27189 2237 -27155
rect 2271 -27189 2305 -27155
rect 2339 -27189 2373 -27155
rect 2407 -27189 2441 -27155
rect 2475 -27189 2509 -27155
rect 2543 -27189 2577 -27155
rect 2611 -27189 2645 -27155
rect 2679 -27189 2713 -27155
rect 2747 -27189 2781 -27155
rect 2815 -27189 2849 -27155
rect 2883 -27189 2917 -27155
rect 2951 -27189 2985 -27155
rect 3019 -27189 3053 -27155
rect 3087 -27189 3121 -27155
rect 3155 -27189 3189 -27155
rect 3223 -27189 3257 -27155
rect 3291 -27189 3325 -27155
rect 3359 -27189 3393 -27155
rect 3427 -27189 3461 -27155
rect 3495 -27189 3529 -27155
rect 3563 -27189 3597 -27155
rect 3631 -27189 3665 -27155
rect 3699 -27189 3733 -27155
rect 3767 -27189 3801 -27155
rect 3835 -27189 3869 -27155
rect 3903 -27189 3937 -27155
rect 3971 -27189 4005 -27155
rect 4039 -27189 4073 -27155
rect 4107 -27189 4141 -27155
rect 4175 -27189 4209 -27155
rect 4243 -27189 4277 -27155
rect 4311 -27189 4345 -27155
rect 4379 -27189 4413 -27155
rect 4447 -27189 4481 -27155
rect 4515 -27189 4549 -27155
rect 4583 -27189 4617 -27155
rect 4651 -27189 4685 -27155
rect 4719 -27189 4753 -27155
rect 4787 -27189 4821 -27155
rect 4855 -27189 4889 -27155
rect 4923 -27189 4957 -27155
rect 4991 -27189 5025 -27155
rect 5059 -27189 5093 -27155
rect 5127 -27189 5161 -27155
rect 5195 -27189 5229 -27155
rect 5263 -27189 5297 -27155
rect 5331 -27189 5365 -27155
rect 5399 -27189 5433 -27155
rect 5467 -27189 5501 -27155
rect 5535 -27189 5569 -27155
rect 5603 -27189 5637 -27155
rect 5671 -27189 5705 -27155
rect 5739 -27189 5773 -27155
rect 5807 -27189 5841 -27155
rect 5875 -27189 5909 -27155
rect 5943 -27189 5977 -27155
rect 6011 -27189 6045 -27155
rect 6079 -27189 6113 -27155
rect 6147 -27189 6181 -27155
rect 6215 -27189 6249 -27155
rect 6283 -27189 6317 -27155
rect 6351 -27189 6385 -27155
rect 6419 -27189 6453 -27155
rect 6487 -27189 6521 -27155
rect 6555 -27189 6589 -27155
rect 6623 -27189 6657 -27155
rect 6691 -27189 6725 -27155
rect 6759 -27189 6793 -27155
rect 6827 -27189 6861 -27155
rect 6895 -27189 6929 -27155
rect 6963 -27189 6997 -27155
rect 7031 -27189 7065 -27155
rect 7099 -27189 7133 -27155
rect 7167 -27189 7201 -27155
rect 7235 -27189 7269 -27155
rect 7303 -27189 7337 -27155
rect 7371 -27189 7405 -27155
rect 7439 -27189 7473 -27155
rect 7507 -27189 7541 -27155
rect 7575 -27189 7609 -27155
rect 7643 -27189 7677 -27155
rect 7711 -27189 7745 -27155
rect 7779 -27189 7813 -27155
rect 7847 -27189 7881 -27155
rect 7915 -27189 7949 -27155
rect 7983 -27189 8017 -27155
rect 8051 -27189 8085 -27155
rect 8119 -27189 8153 -27155
rect 8187 -27189 8221 -27155
rect 8255 -27189 8289 -27155
rect 8323 -27189 8357 -27155
rect 8391 -27189 8425 -27155
rect 8459 -27189 8493 -27155
rect 8527 -27189 8561 -27155
rect 8595 -27189 8629 -27155
rect 8663 -27189 8697 -27155
rect 8731 -27189 8765 -27155
rect 8799 -27189 8833 -27155
rect 8867 -27189 8901 -27155
rect 8935 -27189 8969 -27155
rect 9003 -27189 9037 -27155
rect 9071 -27189 9105 -27155
rect 9139 -27189 9173 -27155
rect 9207 -27189 9241 -27155
rect 9275 -27189 9309 -27155
rect 9343 -27189 9377 -27155
rect 9411 -27189 9445 -27155
rect 9479 -27189 9513 -27155
rect 9547 -27189 9581 -27155
rect 9615 -27189 9649 -27155
rect 9683 -27189 9717 -27155
rect 9751 -27189 9785 -27155
rect 9819 -27189 9853 -27155
rect 9887 -27189 9921 -27155
rect 9955 -27189 9989 -27155
rect 10023 -27189 10057 -27155
rect 10091 -27189 10125 -27155
rect 10159 -27189 10193 -27155
rect 10227 -27189 10261 -27155
rect 10295 -27189 10329 -27155
rect 10363 -27189 10397 -27155
rect 10431 -27189 10465 -27155
rect 10499 -27189 10533 -27155
rect 10567 -27189 10601 -27155
rect 10635 -27189 10669 -27155
rect 10703 -27189 10737 -27155
rect 10771 -27189 10805 -27155
rect 10839 -27189 10873 -27155
rect 10907 -27189 10941 -27155
rect 10975 -27189 11009 -27155
rect 11043 -27189 11077 -27155
rect 11111 -27189 11145 -27155
rect 11179 -27189 11213 -27155
rect 11247 -27189 11281 -27155
rect 11315 -27189 11349 -27155
rect 11383 -27189 11417 -27155
rect 11451 -27189 11485 -27155
rect 11519 -27189 11553 -27155
rect 11587 -27189 11621 -27155
rect 11655 -27189 11689 -27155
rect 11723 -27189 11757 -27155
rect 11791 -27189 11825 -27155
rect 11859 -27189 11893 -27155
rect 11927 -27189 11961 -27155
rect 11995 -27189 12029 -27155
rect 12063 -27189 12097 -27155
rect 12131 -27189 12165 -27155
rect 12199 -27189 12233 -27155
rect 12267 -27189 12301 -27155
rect 12335 -27189 12369 -27155
rect 12403 -27189 12437 -27155
rect 12471 -27189 12505 -27155
rect 12539 -27189 12573 -27155
rect 12607 -27189 12641 -27155
rect 12675 -27189 12709 -27155
rect 12743 -27189 12777 -27155
rect 12811 -27189 12845 -27155
rect 12879 -27189 12913 -27155
rect 12947 -27189 12981 -27155
rect 13015 -27189 13049 -27155
rect 13083 -27189 13117 -27155
rect 13151 -27189 13185 -27155
rect 13219 -27189 13253 -27155
rect 13287 -27189 13321 -27155
rect 13355 -27189 13389 -27155
rect 13423 -27189 13457 -27155
rect 13491 -27189 13525 -27155
rect 13559 -27189 13593 -27155
rect 13627 -27189 13661 -27155
rect 13695 -27189 13729 -27155
rect 13763 -27189 13797 -27155
rect 13831 -27189 13865 -27155
rect 13899 -27189 13933 -27155
rect 13967 -27189 14001 -27155
rect 14035 -27189 14069 -27155
rect 14103 -27189 14137 -27155
rect 14171 -27189 14205 -27155
rect 14239 -27189 14273 -27155
rect 14307 -27189 14341 -27155
rect 14375 -27189 14409 -27155
rect 14443 -27189 14477 -27155
rect 14511 -27189 14545 -27155
rect 14579 -27189 14613 -27155
rect 14647 -27189 14681 -27155
rect 14715 -27189 14749 -27155
rect 14783 -27189 14817 -27155
rect 14851 -27189 14885 -27155
rect 14919 -27189 14953 -27155
rect 14987 -27189 15021 -27155
rect 15055 -27189 15089 -27155
rect 15123 -27189 15157 -27155
rect 15191 -27189 15225 -27155
rect 15259 -27189 15293 -27155
rect 15327 -27189 15361 -27155
rect 15395 -27189 15429 -27155
rect 15463 -27189 15497 -27155
rect 15531 -27189 15565 -27155
rect 15599 -27189 15633 -27155
rect 15667 -27189 15701 -27155
rect 15735 -27189 15769 -27155
rect 15803 -27189 15837 -27155
rect 15871 -27189 15905 -27155
rect 15939 -27189 15973 -27155
rect 16007 -27189 16041 -27155
rect 16075 -27189 16109 -27155
rect 16143 -27189 16177 -27155
rect 16211 -27189 16245 -27155
rect 16279 -27189 16313 -27155
rect 16347 -27189 16381 -27155
rect 16415 -27189 16449 -27155
rect 16483 -27189 16517 -27155
rect 16551 -27189 16585 -27155
rect 16619 -27189 16653 -27155
rect 16687 -27189 16721 -27155
rect 16755 -27189 16789 -27155
rect 16823 -27189 16857 -27155
rect 16891 -27189 16925 -27155
rect 16959 -27189 16993 -27155
rect 17027 -27189 17061 -27155
rect 17095 -27189 17129 -27155
rect 17163 -27189 17197 -27155
rect 17231 -27189 17265 -27155
rect 17299 -27189 17333 -27155
rect 17367 -27189 17401 -27155
rect 17435 -27189 17469 -27155
rect 17503 -27189 17537 -27155
rect 17571 -27189 17605 -27155
rect 17639 -27189 17673 -27155
rect 17707 -27189 17741 -27155
rect 17775 -27189 17809 -27155
rect 17843 -27189 17877 -27155
rect 17911 -27189 17945 -27155
rect 17979 -27189 18013 -27155
rect 18047 -27189 18081 -27155
rect 18115 -27189 18149 -27155
rect 18183 -27189 18217 -27155
rect 18251 -27189 18285 -27155
rect 18319 -27189 18353 -27155
rect 18387 -27189 18421 -27155
rect 18455 -27189 18489 -27155
rect 18523 -27189 18557 -27155
rect 18591 -27189 18625 -27155
rect 18659 -27189 18693 -27155
rect 18727 -27189 18761 -27155
rect 18795 -27189 18829 -27155
rect 18863 -27189 18897 -27155
rect 18931 -27189 18965 -27155
rect 18999 -27189 19033 -27155
rect 19067 -27189 19101 -27155
rect 19135 -27189 19169 -27155
rect 19203 -27189 19237 -27155
rect 19271 -27189 19305 -27155
rect 19339 -27189 19373 -27155
rect 19407 -27189 19441 -27155
rect 19475 -27189 19509 -27155
rect 19543 -27189 19577 -27155
rect 19611 -27189 19645 -27155
rect 19679 -27189 19713 -27155
rect 19747 -27189 19781 -27155
rect 19815 -27189 19849 -27155
rect 19883 -27189 19917 -27155
rect 19951 -27189 19985 -27155
rect 20019 -27189 20053 -27155
rect 20087 -27189 20121 -27155
rect 20155 -27189 20189 -27155
rect 20223 -27189 20257 -27155
rect 20291 -27189 20325 -27155
rect 20359 -27189 20393 -27155
rect 20427 -27189 20461 -27155
rect 20495 -27189 20529 -27155
rect 20563 -27189 20597 -27155
rect 20631 -27189 20665 -27155
rect 20699 -27189 20733 -27155
rect 20767 -27189 20801 -27155
rect 20835 -27189 20869 -27155
rect 20903 -27189 20937 -27155
rect 20971 -27189 21005 -27155
rect 21039 -27189 21073 -27155
rect 21107 -27189 21141 -27155
rect 21175 -27189 21209 -27155
rect 21243 -27189 21277 -27155
rect 21311 -27189 21345 -27155
rect 21379 -27189 21413 -27155
rect 21447 -27189 21481 -27155
rect 21515 -27189 21549 -27155
rect 21583 -27189 21617 -27155
rect 21651 -27189 21685 -27155
rect 21719 -27189 21753 -27155
rect 21787 -27189 21821 -27155
rect 21855 -27189 21889 -27155
rect 21923 -27189 21957 -27155
rect 21991 -27189 22025 -27155
rect 22059 -27189 22093 -27155
rect 22127 -27189 22161 -27155
rect 22195 -27189 22229 -27155
rect 22263 -27189 22297 -27155
rect 22331 -27189 22365 -27155
rect 22399 -27189 22433 -27155
rect 22467 -27189 22501 -27155
rect 22535 -27189 22569 -27155
rect 22603 -27189 22637 -27155
rect 22671 -27189 22705 -27155
rect 22739 -27189 22773 -27155
rect 22807 -27189 22841 -27155
rect 22875 -27189 22909 -27155
rect 22943 -27189 22977 -27155
rect 23011 -27189 23045 -27155
rect 23079 -27189 23113 -27155
rect 23147 -27189 23181 -27155
rect 23215 -27189 23249 -27155
rect 23283 -27189 23317 -27155
rect 23351 -27189 23385 -27155
rect 23419 -27189 23453 -27155
rect 23487 -27189 23521 -27155
rect 23555 -27189 23589 -27155
rect 23623 -27189 23657 -27155
rect 23691 -27189 23725 -27155
rect 23759 -27189 23793 -27155
rect 23827 -27189 23861 -27155
rect 23895 -27189 23929 -27155
rect 23963 -27189 23997 -27155
rect 24031 -27189 24065 -27155
rect 24099 -27189 24133 -27155
rect 24167 -27189 24201 -27155
rect 24235 -27189 24269 -27155
rect 24303 -27189 24337 -27155
rect 24371 -27189 24405 -27155
rect 24439 -27189 24473 -27155
rect 24507 -27189 24541 -27155
rect 24575 -27189 24609 -27155
rect 24643 -27189 24677 -27155
rect 24711 -27189 24745 -27155
<< nsubdiffcont >>
rect 547 4255 581 4289
rect 615 4255 649 4289
rect 683 4255 717 4289
rect 751 4255 785 4289
rect 819 4255 853 4289
rect 887 4255 921 4289
rect 955 4255 989 4289
rect 1023 4255 1057 4289
rect 1091 4255 1125 4289
rect 1159 4255 1193 4289
rect 1227 4255 1261 4289
rect 1295 4255 1329 4289
rect 1363 4255 1397 4289
rect 1431 4255 1465 4289
rect 1499 4255 1533 4289
rect 1567 4255 1601 4289
rect 1635 4255 1669 4289
rect 1703 4255 1737 4289
rect 1771 4255 1805 4289
rect 1839 4255 1873 4289
rect 1907 4255 1941 4289
rect 1975 4255 2009 4289
rect 2043 4255 2077 4289
rect 2111 4255 2145 4289
rect 2179 4255 2213 4289
rect 2247 4255 2281 4289
rect 2315 4255 2349 4289
rect 2383 4255 2417 4289
rect 2451 4255 2485 4289
rect 2519 4255 2553 4289
rect 2587 4255 2621 4289
rect 2655 4255 2689 4289
rect 2723 4255 2757 4289
rect 2791 4255 2825 4289
rect 2859 4255 2893 4289
rect 2927 4255 2961 4289
rect 2995 4255 3029 4289
rect 3063 4255 3097 4289
rect 3131 4255 3165 4289
rect 3199 4255 3233 4289
rect 3267 4255 3301 4289
rect 3335 4255 3369 4289
rect 3403 4255 3437 4289
rect 3471 4255 3505 4289
rect 3539 4255 3573 4289
rect 3607 4255 3641 4289
rect 3675 4255 3709 4289
rect 3743 4255 3777 4289
rect 3811 4255 3845 4289
rect 3879 4255 3913 4289
rect 3947 4255 3981 4289
rect 4015 4255 4049 4289
rect 4083 4255 4117 4289
rect 4151 4255 4185 4289
rect 4219 4255 4253 4289
rect 4287 4255 4321 4289
rect 4355 4255 4389 4289
rect 4423 4255 4457 4289
rect 4491 4255 4525 4289
rect 4559 4255 4593 4289
rect 4627 4255 4661 4289
rect 4695 4255 4729 4289
rect 4763 4255 4797 4289
rect 4831 4255 4865 4289
rect 4899 4255 4933 4289
rect 4967 4255 5001 4289
rect 5035 4255 5069 4289
rect 5103 4255 5137 4289
rect 5171 4255 5205 4289
rect 5239 4255 5273 4289
rect 5307 4255 5341 4289
rect 5375 4255 5409 4289
rect 5443 4255 5477 4289
rect 5511 4255 5545 4289
rect 5579 4255 5613 4289
rect 5647 4255 5681 4289
rect 5715 4255 5749 4289
rect 5783 4255 5817 4289
rect 5851 4255 5885 4289
rect 5919 4255 5953 4289
rect 5987 4255 6021 4289
rect 6055 4255 6089 4289
rect 6123 4255 6157 4289
rect 6191 4255 6225 4289
rect 6259 4255 6293 4289
rect 6327 4255 6361 4289
rect 6395 4255 6429 4289
rect 6463 4255 6497 4289
rect 6531 4255 6565 4289
rect 6599 4255 6633 4289
rect 6667 4255 6701 4289
rect 6735 4255 6769 4289
rect 6803 4255 6837 4289
rect 6871 4255 6905 4289
rect 6939 4255 6973 4289
rect 7007 4255 7041 4289
rect 7075 4255 7109 4289
rect 7143 4255 7177 4289
rect 7211 4255 7245 4289
rect 7279 4255 7313 4289
rect 7347 4255 7381 4289
rect 7415 4255 7449 4289
rect 7483 4255 7517 4289
rect 7551 4255 7585 4289
rect 7619 4255 7653 4289
rect 7687 4255 7721 4289
rect 7755 4255 7789 4289
rect 7823 4255 7857 4289
rect 7891 4255 7925 4289
rect 7959 4255 7993 4289
rect 8027 4255 8061 4289
rect 8095 4255 8129 4289
rect 8163 4255 8197 4289
rect 8231 4255 8265 4289
rect 8299 4255 8333 4289
rect 8367 4255 8401 4289
rect 8435 4255 8469 4289
rect 8503 4255 8537 4289
rect 8571 4255 8605 4289
rect 8639 4255 8673 4289
rect 8707 4255 8741 4289
rect 8775 4255 8809 4289
rect 8843 4255 8877 4289
rect 8911 4255 8945 4289
rect 8979 4255 9013 4289
rect 9047 4255 9081 4289
rect 9115 4255 9149 4289
rect 9183 4255 9217 4289
rect 9251 4255 9285 4289
rect 9319 4255 9353 4289
rect 9387 4255 9421 4289
rect 9455 4255 9489 4289
rect 9523 4255 9557 4289
rect 9591 4255 9625 4289
rect 9659 4255 9693 4289
rect 9727 4255 9761 4289
rect 9795 4255 9829 4289
rect 9863 4255 9897 4289
rect 9931 4255 9965 4289
rect 9999 4255 10033 4289
rect 10067 4255 10101 4289
rect 10135 4255 10169 4289
rect 10203 4255 10237 4289
rect 10271 4255 10305 4289
rect 10339 4255 10373 4289
rect 10407 4255 10441 4289
rect 10475 4255 10509 4289
rect 10543 4255 10577 4289
rect 10611 4255 10645 4289
rect 10679 4255 10713 4289
rect 10747 4255 10781 4289
rect 10815 4255 10849 4289
rect 10883 4255 10917 4289
rect 10951 4255 10985 4289
rect 11019 4255 11053 4289
rect 11087 4255 11121 4289
rect 11155 4255 11189 4289
rect 11223 4255 11257 4289
rect 11291 4255 11325 4289
rect 11359 4255 11393 4289
rect 11427 4255 11461 4289
rect 11495 4255 11529 4289
rect 11563 4255 11597 4289
rect 11631 4255 11665 4289
rect 11699 4255 11733 4289
rect 11767 4255 11801 4289
rect 11835 4255 11869 4289
rect 11903 4255 11937 4289
rect 11971 4255 12005 4289
rect 12039 4255 12073 4289
rect 12107 4255 12141 4289
rect 12175 4255 12209 4289
rect 12243 4255 12277 4289
rect 12311 4255 12345 4289
rect 12379 4255 12413 4289
rect 12447 4255 12481 4289
rect 12515 4255 12549 4289
rect 12583 4255 12617 4289
rect 12651 4255 12685 4289
rect 12719 4255 12753 4289
rect 12787 4255 12821 4289
rect 12855 4255 12889 4289
rect 12923 4255 12957 4289
rect 12991 4255 13025 4289
rect 13059 4255 13093 4289
rect 13127 4255 13161 4289
rect 13195 4255 13229 4289
rect 13263 4255 13297 4289
rect 13331 4255 13365 4289
rect 13399 4255 13433 4289
rect 13467 4255 13501 4289
rect 13535 4255 13569 4289
rect 13603 4255 13637 4289
rect 13671 4255 13705 4289
rect 13739 4255 13773 4289
rect 13807 4255 13841 4289
rect 13875 4255 13909 4289
rect 13943 4255 13977 4289
rect 14011 4255 14045 4289
rect 14079 4255 14113 4289
rect 14147 4255 14181 4289
rect 14215 4255 14249 4289
rect 14283 4255 14317 4289
rect 14351 4255 14385 4289
rect 14419 4255 14453 4289
rect 14487 4255 14521 4289
rect 14555 4255 14589 4289
rect 14623 4255 14657 4289
rect 14691 4255 14725 4289
rect 14759 4255 14793 4289
rect 14827 4255 14861 4289
rect 14895 4255 14929 4289
rect 14963 4255 14997 4289
rect 15031 4255 15065 4289
rect 15099 4255 15133 4289
rect 15167 4255 15201 4289
rect 15235 4255 15269 4289
rect 15303 4255 15337 4289
rect 15371 4255 15405 4289
rect 15439 4255 15473 4289
rect 15507 4255 15541 4289
rect 15575 4255 15609 4289
rect 15643 4255 15677 4289
rect 15711 4255 15745 4289
rect 15779 4255 15813 4289
rect 15847 4255 15881 4289
rect 15915 4255 15949 4289
rect 15983 4255 16017 4289
rect 16051 4255 16085 4289
rect 16119 4255 16153 4289
rect 16187 4255 16221 4289
rect 16255 4255 16289 4289
rect 16323 4255 16357 4289
rect 16391 4255 16425 4289
rect 16459 4255 16493 4289
rect 16527 4255 16561 4289
rect 16595 4255 16629 4289
rect 16663 4255 16697 4289
rect 16731 4255 16765 4289
rect 16799 4255 16833 4289
rect 16867 4255 16901 4289
rect 16935 4255 16969 4289
rect 17003 4255 17037 4289
rect 17071 4255 17105 4289
rect 17139 4255 17173 4289
rect 17207 4255 17241 4289
rect 17275 4255 17309 4289
rect 17343 4255 17377 4289
rect 17411 4255 17445 4289
rect 17479 4255 17513 4289
rect 17547 4255 17581 4289
rect 17615 4255 17649 4289
rect 17683 4255 17717 4289
rect 17751 4255 17785 4289
rect 17819 4255 17853 4289
rect 17887 4255 17921 4289
rect 17955 4255 17989 4289
rect 18023 4255 18057 4289
rect 18091 4255 18125 4289
rect 18159 4255 18193 4289
rect 18227 4255 18261 4289
rect 18295 4255 18329 4289
rect 18363 4255 18397 4289
rect 18431 4255 18465 4289
rect 18499 4255 18533 4289
rect 18567 4255 18601 4289
rect 18635 4255 18669 4289
rect 18703 4255 18737 4289
rect 18771 4255 18805 4289
rect 18839 4255 18873 4289
rect 18907 4255 18941 4289
rect 18975 4255 19009 4289
rect 19043 4255 19077 4289
rect 19111 4255 19145 4289
rect 19179 4255 19213 4289
rect 19247 4255 19281 4289
rect 19315 4255 19349 4289
rect 19383 4255 19417 4289
rect 19451 4255 19485 4289
rect 19519 4255 19553 4289
rect 19587 4255 19621 4289
rect 19655 4255 19689 4289
rect 19723 4255 19757 4289
rect 19791 4255 19825 4289
rect 19859 4255 19893 4289
rect 19927 4255 19961 4289
rect 19995 4255 20029 4289
rect 20063 4255 20097 4289
rect 20131 4255 20165 4289
rect 20199 4255 20233 4289
rect 20267 4255 20301 4289
rect 20335 4255 20369 4289
rect 20403 4255 20437 4289
rect 20471 4255 20505 4289
rect 20539 4255 20573 4289
rect 20607 4255 20641 4289
rect 20675 4255 20709 4289
rect 20743 4255 20777 4289
rect 20811 4255 20845 4289
rect 20879 4255 20913 4289
rect 20947 4255 20981 4289
rect 21015 4255 21049 4289
rect 21083 4255 21117 4289
rect 21151 4255 21185 4289
rect 21219 4255 21253 4289
rect 21287 4255 21321 4289
rect 21355 4255 21389 4289
rect 21423 4255 21457 4289
rect 21491 4255 21525 4289
rect 21559 4255 21593 4289
rect 21627 4255 21661 4289
rect 21695 4255 21729 4289
rect 21763 4255 21797 4289
rect 21831 4255 21865 4289
rect 21899 4255 21933 4289
rect 21967 4255 22001 4289
rect 22035 4255 22069 4289
rect 22103 4255 22137 4289
rect 22171 4255 22205 4289
rect 22239 4255 22273 4289
rect 22307 4255 22341 4289
rect 22375 4255 22409 4289
rect 22443 4255 22477 4289
rect 22511 4255 22545 4289
rect 22579 4255 22613 4289
rect 22647 4255 22681 4289
rect 22715 4255 22749 4289
rect 22783 4255 22817 4289
rect 22851 4255 22885 4289
rect 22919 4255 22953 4289
rect 22987 4255 23021 4289
rect 23055 4255 23089 4289
rect 23123 4255 23157 4289
rect 23191 4255 23225 4289
rect 23259 4255 23293 4289
rect 23327 4255 23361 4289
rect 23395 4255 23429 4289
rect 23463 4255 23497 4289
rect 23531 4255 23565 4289
rect 23599 4255 23633 4289
rect 23667 4255 23701 4289
rect 23735 4255 23769 4289
rect 23803 4255 23837 4289
rect 23871 4255 23905 4289
rect 23939 4255 23973 4289
rect 24007 4255 24041 4289
rect 24075 4255 24109 4289
rect 24143 4255 24177 4289
rect 24211 4255 24245 4289
rect 24279 4255 24313 4289
rect 24347 4255 24381 4289
rect 24415 4255 24449 4289
rect 24483 4255 24517 4289
rect 24551 4255 24585 4289
rect 24619 4255 24653 4289
rect 411 4110 445 4144
rect 411 4042 445 4076
rect 411 3974 445 4008
rect 411 3906 445 3940
rect 411 3838 445 3872
rect 411 3770 445 3804
rect 411 3702 445 3736
rect 411 3634 445 3668
rect 411 3566 445 3600
rect 411 3498 445 3532
rect 411 3430 445 3464
rect 411 3362 445 3396
rect 411 3294 445 3328
rect 411 3226 445 3260
rect 411 3158 445 3192
rect 411 3090 445 3124
rect 411 3022 445 3056
rect 411 2954 445 2988
rect 411 2886 445 2920
rect 411 2818 445 2852
rect 411 2750 445 2784
rect 411 2682 445 2716
rect 411 2614 445 2648
rect 411 2546 445 2580
rect 411 2478 445 2512
rect 411 2410 445 2444
rect 411 2342 445 2376
rect 411 2274 445 2308
rect 411 2206 445 2240
rect 411 2138 445 2172
rect 411 2070 445 2104
rect 411 2002 445 2036
rect 411 1934 445 1968
rect 411 1866 445 1900
rect 411 1798 445 1832
rect 411 1730 445 1764
rect 411 1662 445 1696
rect 411 1594 445 1628
rect 411 1526 445 1560
rect 411 1458 445 1492
rect 411 1390 445 1424
rect 411 1322 445 1356
rect 411 1254 445 1288
rect 411 1186 445 1220
rect 411 1118 445 1152
rect 411 1050 445 1084
rect 411 982 445 1016
rect 411 914 445 948
rect 411 846 445 880
rect 411 778 445 812
rect 411 710 445 744
rect 411 642 445 676
rect 411 574 445 608
rect 411 506 445 540
rect 411 438 445 472
rect 411 370 445 404
rect 411 302 445 336
rect 411 234 445 268
rect 411 166 445 200
rect 411 98 445 132
rect 411 30 445 64
rect 411 -38 445 -4
rect 411 -106 445 -72
rect 411 -174 445 -140
rect 411 -242 445 -208
rect 411 -310 445 -276
rect 411 -378 445 -344
rect 411 -446 445 -412
rect 411 -514 445 -480
rect 411 -582 445 -548
rect 411 -650 445 -616
rect 411 -718 445 -684
rect 411 -786 445 -752
rect 411 -854 445 -820
rect 411 -922 445 -888
rect 411 -990 445 -956
rect 411 -1058 445 -1024
rect 411 -1126 445 -1092
rect 411 -1194 445 -1160
rect 411 -1262 445 -1228
rect 411 -1330 445 -1296
rect 411 -1398 445 -1364
rect 411 -1466 445 -1432
rect 411 -1534 445 -1500
rect 411 -1602 445 -1568
rect 411 -1670 445 -1636
rect 411 -1738 445 -1704
rect 411 -1806 445 -1772
rect 411 -1874 445 -1840
rect 411 -1942 445 -1908
rect 411 -2010 445 -1976
rect 411 -2078 445 -2044
rect 411 -2146 445 -2112
rect 411 -2214 445 -2180
rect 411 -2282 445 -2248
rect 411 -2350 445 -2316
rect 411 -2418 445 -2384
rect 411 -2486 445 -2452
rect 411 -2554 445 -2520
rect 411 -2622 445 -2588
rect 411 -2690 445 -2656
rect 411 -2758 445 -2724
rect 411 -2826 445 -2792
rect 411 -2894 445 -2860
rect 411 -2962 445 -2928
rect 411 -3030 445 -2996
rect 411 -3098 445 -3064
rect 411 -3166 445 -3132
rect 411 -3234 445 -3200
rect 411 -3302 445 -3268
rect 411 -3370 445 -3336
rect 411 -3438 445 -3404
rect 411 -3506 445 -3472
rect 411 -3574 445 -3540
rect 411 -3642 445 -3608
rect 411 -3710 445 -3676
rect 411 -3778 445 -3744
rect 411 -3846 445 -3812
rect 411 -3914 445 -3880
rect 411 -3982 445 -3948
rect 411 -4050 445 -4016
rect 411 -4118 445 -4084
rect 411 -4186 445 -4152
rect 411 -4254 445 -4220
rect 411 -4322 445 -4288
rect 411 -4390 445 -4356
rect 411 -4458 445 -4424
rect 411 -4526 445 -4492
rect 411 -4594 445 -4560
rect 411 -4662 445 -4628
rect 411 -4730 445 -4696
rect 411 -4798 445 -4764
rect 411 -4866 445 -4832
rect 411 -4934 445 -4900
rect 411 -5002 445 -4968
rect 411 -5070 445 -5036
rect 411 -5138 445 -5104
rect 411 -5206 445 -5172
rect 411 -5274 445 -5240
rect 411 -5342 445 -5308
rect 411 -5410 445 -5376
rect 411 -5478 445 -5444
rect 411 -5546 445 -5512
rect 411 -5614 445 -5580
rect 411 -5682 445 -5648
rect 411 -5750 445 -5716
rect 411 -5818 445 -5784
rect 411 -5886 445 -5852
rect 411 -5954 445 -5920
rect 411 -6022 445 -5988
rect 411 -6090 445 -6056
rect 411 -6158 445 -6124
rect 411 -6226 445 -6192
rect 411 -6294 445 -6260
rect 411 -6362 445 -6328
rect 411 -6430 445 -6396
rect 411 -6498 445 -6464
rect 411 -6566 445 -6532
rect 411 -6634 445 -6600
rect 411 -6702 445 -6668
rect 411 -6770 445 -6736
rect 411 -6838 445 -6804
rect 411 -6906 445 -6872
rect 411 -6974 445 -6940
rect 411 -7042 445 -7008
rect 411 -7110 445 -7076
rect 411 -7178 445 -7144
rect 411 -7246 445 -7212
rect 411 -7314 445 -7280
rect 411 -7382 445 -7348
rect 411 -7450 445 -7416
rect 411 -7518 445 -7484
rect 411 -7586 445 -7552
rect 411 -7654 445 -7620
rect 411 -7722 445 -7688
rect 411 -7790 445 -7756
rect 411 -7858 445 -7824
rect 411 -7926 445 -7892
rect 411 -7994 445 -7960
rect 411 -8062 445 -8028
rect 411 -8130 445 -8096
rect 411 -8198 445 -8164
rect 411 -8266 445 -8232
rect 411 -8334 445 -8300
rect 411 -8402 445 -8368
rect 411 -8470 445 -8436
rect 411 -8538 445 -8504
rect 411 -8606 445 -8572
rect 411 -8674 445 -8640
rect 411 -8742 445 -8708
rect 411 -8810 445 -8776
rect 411 -8878 445 -8844
rect 411 -8946 445 -8912
rect 411 -9014 445 -8980
rect 411 -9082 445 -9048
rect 411 -9150 445 -9116
rect 411 -9218 445 -9184
rect 411 -9286 445 -9252
rect 411 -9354 445 -9320
rect 411 -9422 445 -9388
rect 411 -9490 445 -9456
rect 411 -9558 445 -9524
rect 411 -9626 445 -9592
rect 411 -9694 445 -9660
rect 411 -9762 445 -9728
rect 411 -9830 445 -9796
rect 411 -9898 445 -9864
rect 411 -9966 445 -9932
rect 411 -10034 445 -10000
rect 411 -10102 445 -10068
rect 411 -10170 445 -10136
rect 24755 4110 24789 4144
rect 24755 4042 24789 4076
rect 24755 3974 24789 4008
rect 24755 3906 24789 3940
rect 24755 3838 24789 3872
rect 24755 3770 24789 3804
rect 24755 3702 24789 3736
rect 24755 3634 24789 3668
rect 24755 3566 24789 3600
rect 24755 3498 24789 3532
rect 24755 3430 24789 3464
rect 24755 3362 24789 3396
rect 24755 3294 24789 3328
rect 24755 3226 24789 3260
rect 24755 3158 24789 3192
rect 24755 3090 24789 3124
rect 24755 3022 24789 3056
rect 24755 2954 24789 2988
rect 24755 2886 24789 2920
rect 24755 2818 24789 2852
rect 24755 2750 24789 2784
rect 24755 2682 24789 2716
rect 24755 2614 24789 2648
rect 24755 2546 24789 2580
rect 24755 2478 24789 2512
rect 24755 2410 24789 2444
rect 24755 2342 24789 2376
rect 24755 2274 24789 2308
rect 24755 2206 24789 2240
rect 24755 2138 24789 2172
rect 24755 2070 24789 2104
rect 24755 2002 24789 2036
rect 24755 1934 24789 1968
rect 24755 1866 24789 1900
rect 24755 1798 24789 1832
rect 24755 1730 24789 1764
rect 24755 1662 24789 1696
rect 24755 1594 24789 1628
rect 24755 1526 24789 1560
rect 24755 1458 24789 1492
rect 24755 1390 24789 1424
rect 24755 1322 24789 1356
rect 24755 1254 24789 1288
rect 24755 1186 24789 1220
rect 24755 1118 24789 1152
rect 24755 1050 24789 1084
rect 24755 982 24789 1016
rect 24755 914 24789 948
rect 24755 846 24789 880
rect 24755 778 24789 812
rect 24755 710 24789 744
rect 24755 642 24789 676
rect 24755 574 24789 608
rect 24755 506 24789 540
rect 24755 438 24789 472
rect 24755 370 24789 404
rect 24755 302 24789 336
rect 24755 234 24789 268
rect 24755 166 24789 200
rect 24755 98 24789 132
rect 24755 30 24789 64
rect 24755 -38 24789 -4
rect 24755 -106 24789 -72
rect 24755 -174 24789 -140
rect 24755 -242 24789 -208
rect 24755 -310 24789 -276
rect 24755 -378 24789 -344
rect 24755 -446 24789 -412
rect 24755 -514 24789 -480
rect 24755 -582 24789 -548
rect 24755 -650 24789 -616
rect 24755 -718 24789 -684
rect 24755 -786 24789 -752
rect 24755 -854 24789 -820
rect 24755 -922 24789 -888
rect 24755 -990 24789 -956
rect 24755 -1058 24789 -1024
rect 24755 -1126 24789 -1092
rect 24755 -1194 24789 -1160
rect 24755 -1262 24789 -1228
rect 24755 -1330 24789 -1296
rect 24755 -1398 24789 -1364
rect 24755 -1466 24789 -1432
rect 24755 -1534 24789 -1500
rect 24755 -1602 24789 -1568
rect 24755 -1670 24789 -1636
rect 24755 -1738 24789 -1704
rect 24755 -1806 24789 -1772
rect 24755 -1874 24789 -1840
rect 24755 -1942 24789 -1908
rect 24755 -2010 24789 -1976
rect 24755 -2078 24789 -2044
rect 24755 -2146 24789 -2112
rect 24755 -2214 24789 -2180
rect 24755 -2282 24789 -2248
rect 24755 -2350 24789 -2316
rect 24755 -2418 24789 -2384
rect 24755 -2486 24789 -2452
rect 24755 -2554 24789 -2520
rect 24755 -2622 24789 -2588
rect 24755 -2690 24789 -2656
rect 24755 -2758 24789 -2724
rect 24755 -2826 24789 -2792
rect 24755 -2894 24789 -2860
rect 24755 -2962 24789 -2928
rect 24755 -3030 24789 -2996
rect 24755 -3098 24789 -3064
rect 24755 -3166 24789 -3132
rect 24755 -3234 24789 -3200
rect 24755 -3302 24789 -3268
rect 24755 -3370 24789 -3336
rect 24755 -3438 24789 -3404
rect 24755 -3506 24789 -3472
rect 24755 -3574 24789 -3540
rect 24755 -3642 24789 -3608
rect 24755 -3710 24789 -3676
rect 24755 -3778 24789 -3744
rect 24755 -3846 24789 -3812
rect 24755 -3914 24789 -3880
rect 24755 -3982 24789 -3948
rect 24755 -4050 24789 -4016
rect 24755 -4118 24789 -4084
rect 24755 -4186 24789 -4152
rect 24755 -4254 24789 -4220
rect 24755 -4322 24789 -4288
rect 24755 -4390 24789 -4356
rect 24755 -4458 24789 -4424
rect 24755 -4526 24789 -4492
rect 24755 -4594 24789 -4560
rect 24755 -4662 24789 -4628
rect 24755 -4730 24789 -4696
rect 24755 -4798 24789 -4764
rect 24755 -4866 24789 -4832
rect 24755 -4934 24789 -4900
rect 24755 -5002 24789 -4968
rect 24755 -5070 24789 -5036
rect 24755 -5138 24789 -5104
rect 24755 -5206 24789 -5172
rect 24755 -5274 24789 -5240
rect 24755 -5342 24789 -5308
rect 24755 -5410 24789 -5376
rect 24755 -5478 24789 -5444
rect 24755 -5546 24789 -5512
rect 24755 -5614 24789 -5580
rect 24755 -5682 24789 -5648
rect 24755 -5750 24789 -5716
rect 24755 -5818 24789 -5784
rect 24755 -5886 24789 -5852
rect 24755 -5954 24789 -5920
rect 24755 -6022 24789 -5988
rect 24755 -6090 24789 -6056
rect 24755 -6158 24789 -6124
rect 24755 -6226 24789 -6192
rect 24755 -6294 24789 -6260
rect 24755 -6362 24789 -6328
rect 24755 -6430 24789 -6396
rect 24755 -6498 24789 -6464
rect 24755 -6566 24789 -6532
rect 24755 -6634 24789 -6600
rect 24755 -6702 24789 -6668
rect 24755 -6770 24789 -6736
rect 24755 -6838 24789 -6804
rect 24755 -6906 24789 -6872
rect 24755 -6974 24789 -6940
rect 24755 -7042 24789 -7008
rect 24755 -7110 24789 -7076
rect 24755 -7178 24789 -7144
rect 24755 -7246 24789 -7212
rect 24755 -7314 24789 -7280
rect 24755 -7382 24789 -7348
rect 24755 -7450 24789 -7416
rect 24755 -7518 24789 -7484
rect 24755 -7586 24789 -7552
rect 24755 -7654 24789 -7620
rect 24755 -7722 24789 -7688
rect 24755 -7790 24789 -7756
rect 24755 -7858 24789 -7824
rect 24755 -7926 24789 -7892
rect 24755 -7994 24789 -7960
rect 24755 -8062 24789 -8028
rect 24755 -8130 24789 -8096
rect 24755 -8198 24789 -8164
rect 24755 -8266 24789 -8232
rect 24755 -8334 24789 -8300
rect 24755 -8402 24789 -8368
rect 24755 -8470 24789 -8436
rect 24755 -8538 24789 -8504
rect 24755 -8606 24789 -8572
rect 24755 -8674 24789 -8640
rect 24755 -8742 24789 -8708
rect 24755 -8810 24789 -8776
rect 24755 -8878 24789 -8844
rect 24755 -8946 24789 -8912
rect 24755 -9014 24789 -8980
rect 24755 -9082 24789 -9048
rect 24755 -9150 24789 -9116
rect 24755 -9218 24789 -9184
rect 24755 -9286 24789 -9252
rect 24755 -9354 24789 -9320
rect 24755 -9422 24789 -9388
rect 24755 -9490 24789 -9456
rect 24755 -9558 24789 -9524
rect 24755 -9626 24789 -9592
rect 24755 -9694 24789 -9660
rect 24755 -9762 24789 -9728
rect 24755 -9830 24789 -9796
rect 24755 -9898 24789 -9864
rect 24755 -9966 24789 -9932
rect 24755 -10034 24789 -10000
rect 24755 -10102 24789 -10068
rect 24755 -10170 24789 -10136
rect 547 -10315 581 -10281
rect 615 -10315 649 -10281
rect 683 -10315 717 -10281
rect 751 -10315 785 -10281
rect 819 -10315 853 -10281
rect 887 -10315 921 -10281
rect 955 -10315 989 -10281
rect 1023 -10315 1057 -10281
rect 1091 -10315 1125 -10281
rect 1159 -10315 1193 -10281
rect 1227 -10315 1261 -10281
rect 1295 -10315 1329 -10281
rect 1363 -10315 1397 -10281
rect 1431 -10315 1465 -10281
rect 1499 -10315 1533 -10281
rect 1567 -10315 1601 -10281
rect 1635 -10315 1669 -10281
rect 1703 -10315 1737 -10281
rect 1771 -10315 1805 -10281
rect 1839 -10315 1873 -10281
rect 1907 -10315 1941 -10281
rect 1975 -10315 2009 -10281
rect 2043 -10315 2077 -10281
rect 2111 -10315 2145 -10281
rect 2179 -10315 2213 -10281
rect 2247 -10315 2281 -10281
rect 2315 -10315 2349 -10281
rect 2383 -10315 2417 -10281
rect 2451 -10315 2485 -10281
rect 2519 -10315 2553 -10281
rect 2587 -10315 2621 -10281
rect 2655 -10315 2689 -10281
rect 2723 -10315 2757 -10281
rect 2791 -10315 2825 -10281
rect 2859 -10315 2893 -10281
rect 2927 -10315 2961 -10281
rect 2995 -10315 3029 -10281
rect 3063 -10315 3097 -10281
rect 3131 -10315 3165 -10281
rect 3199 -10315 3233 -10281
rect 3267 -10315 3301 -10281
rect 3335 -10315 3369 -10281
rect 3403 -10315 3437 -10281
rect 3471 -10315 3505 -10281
rect 3539 -10315 3573 -10281
rect 3607 -10315 3641 -10281
rect 3675 -10315 3709 -10281
rect 3743 -10315 3777 -10281
rect 3811 -10315 3845 -10281
rect 3879 -10315 3913 -10281
rect 3947 -10315 3981 -10281
rect 4015 -10315 4049 -10281
rect 4083 -10315 4117 -10281
rect 4151 -10315 4185 -10281
rect 4219 -10315 4253 -10281
rect 4287 -10315 4321 -10281
rect 4355 -10315 4389 -10281
rect 4423 -10315 4457 -10281
rect 4491 -10315 4525 -10281
rect 4559 -10315 4593 -10281
rect 4627 -10315 4661 -10281
rect 4695 -10315 4729 -10281
rect 4763 -10315 4797 -10281
rect 4831 -10315 4865 -10281
rect 4899 -10315 4933 -10281
rect 4967 -10315 5001 -10281
rect 5035 -10315 5069 -10281
rect 5103 -10315 5137 -10281
rect 5171 -10315 5205 -10281
rect 5239 -10315 5273 -10281
rect 5307 -10315 5341 -10281
rect 5375 -10315 5409 -10281
rect 5443 -10315 5477 -10281
rect 5511 -10315 5545 -10281
rect 5579 -10315 5613 -10281
rect 5647 -10315 5681 -10281
rect 5715 -10315 5749 -10281
rect 5783 -10315 5817 -10281
rect 5851 -10315 5885 -10281
rect 5919 -10315 5953 -10281
rect 5987 -10315 6021 -10281
rect 6055 -10315 6089 -10281
rect 6123 -10315 6157 -10281
rect 6191 -10315 6225 -10281
rect 6259 -10315 6293 -10281
rect 6327 -10315 6361 -10281
rect 6395 -10315 6429 -10281
rect 6463 -10315 6497 -10281
rect 6531 -10315 6565 -10281
rect 6599 -10315 6633 -10281
rect 6667 -10315 6701 -10281
rect 6735 -10315 6769 -10281
rect 6803 -10315 6837 -10281
rect 6871 -10315 6905 -10281
rect 6939 -10315 6973 -10281
rect 7007 -10315 7041 -10281
rect 7075 -10315 7109 -10281
rect 7143 -10315 7177 -10281
rect 7211 -10315 7245 -10281
rect 7279 -10315 7313 -10281
rect 7347 -10315 7381 -10281
rect 7415 -10315 7449 -10281
rect 7483 -10315 7517 -10281
rect 7551 -10315 7585 -10281
rect 7619 -10315 7653 -10281
rect 7687 -10315 7721 -10281
rect 7755 -10315 7789 -10281
rect 7823 -10315 7857 -10281
rect 7891 -10315 7925 -10281
rect 7959 -10315 7993 -10281
rect 8027 -10315 8061 -10281
rect 8095 -10315 8129 -10281
rect 8163 -10315 8197 -10281
rect 8231 -10315 8265 -10281
rect 8299 -10315 8333 -10281
rect 8367 -10315 8401 -10281
rect 8435 -10315 8469 -10281
rect 8503 -10315 8537 -10281
rect 8571 -10315 8605 -10281
rect 8639 -10315 8673 -10281
rect 8707 -10315 8741 -10281
rect 8775 -10315 8809 -10281
rect 8843 -10315 8877 -10281
rect 8911 -10315 8945 -10281
rect 8979 -10315 9013 -10281
rect 9047 -10315 9081 -10281
rect 9115 -10315 9149 -10281
rect 9183 -10315 9217 -10281
rect 9251 -10315 9285 -10281
rect 9319 -10315 9353 -10281
rect 9387 -10315 9421 -10281
rect 9455 -10315 9489 -10281
rect 9523 -10315 9557 -10281
rect 9591 -10315 9625 -10281
rect 9659 -10315 9693 -10281
rect 9727 -10315 9761 -10281
rect 9795 -10315 9829 -10281
rect 9863 -10315 9897 -10281
rect 9931 -10315 9965 -10281
rect 9999 -10315 10033 -10281
rect 10067 -10315 10101 -10281
rect 10135 -10315 10169 -10281
rect 10203 -10315 10237 -10281
rect 10271 -10315 10305 -10281
rect 10339 -10315 10373 -10281
rect 10407 -10315 10441 -10281
rect 10475 -10315 10509 -10281
rect 10543 -10315 10577 -10281
rect 10611 -10315 10645 -10281
rect 10679 -10315 10713 -10281
rect 10747 -10315 10781 -10281
rect 10815 -10315 10849 -10281
rect 10883 -10315 10917 -10281
rect 10951 -10315 10985 -10281
rect 11019 -10315 11053 -10281
rect 11087 -10315 11121 -10281
rect 11155 -10315 11189 -10281
rect 11223 -10315 11257 -10281
rect 11291 -10315 11325 -10281
rect 11359 -10315 11393 -10281
rect 11427 -10315 11461 -10281
rect 11495 -10315 11529 -10281
rect 11563 -10315 11597 -10281
rect 11631 -10315 11665 -10281
rect 11699 -10315 11733 -10281
rect 11767 -10315 11801 -10281
rect 11835 -10315 11869 -10281
rect 11903 -10315 11937 -10281
rect 11971 -10315 12005 -10281
rect 12039 -10315 12073 -10281
rect 12107 -10315 12141 -10281
rect 12175 -10315 12209 -10281
rect 12243 -10315 12277 -10281
rect 12311 -10315 12345 -10281
rect 12379 -10315 12413 -10281
rect 12447 -10315 12481 -10281
rect 12515 -10315 12549 -10281
rect 12583 -10315 12617 -10281
rect 12651 -10315 12685 -10281
rect 12719 -10315 12753 -10281
rect 12787 -10315 12821 -10281
rect 12855 -10315 12889 -10281
rect 12923 -10315 12957 -10281
rect 12991 -10315 13025 -10281
rect 13059 -10315 13093 -10281
rect 13127 -10315 13161 -10281
rect 13195 -10315 13229 -10281
rect 13263 -10315 13297 -10281
rect 13331 -10315 13365 -10281
rect 13399 -10315 13433 -10281
rect 13467 -10315 13501 -10281
rect 13535 -10315 13569 -10281
rect 13603 -10315 13637 -10281
rect 13671 -10315 13705 -10281
rect 13739 -10315 13773 -10281
rect 13807 -10315 13841 -10281
rect 13875 -10315 13909 -10281
rect 13943 -10315 13977 -10281
rect 14011 -10315 14045 -10281
rect 14079 -10315 14113 -10281
rect 14147 -10315 14181 -10281
rect 14215 -10315 14249 -10281
rect 14283 -10315 14317 -10281
rect 14351 -10315 14385 -10281
rect 14419 -10315 14453 -10281
rect 14487 -10315 14521 -10281
rect 14555 -10315 14589 -10281
rect 14623 -10315 14657 -10281
rect 14691 -10315 14725 -10281
rect 14759 -10315 14793 -10281
rect 14827 -10315 14861 -10281
rect 14895 -10315 14929 -10281
rect 14963 -10315 14997 -10281
rect 15031 -10315 15065 -10281
rect 15099 -10315 15133 -10281
rect 15167 -10315 15201 -10281
rect 15235 -10315 15269 -10281
rect 15303 -10315 15337 -10281
rect 15371 -10315 15405 -10281
rect 15439 -10315 15473 -10281
rect 15507 -10315 15541 -10281
rect 15575 -10315 15609 -10281
rect 15643 -10315 15677 -10281
rect 15711 -10315 15745 -10281
rect 15779 -10315 15813 -10281
rect 15847 -10315 15881 -10281
rect 15915 -10315 15949 -10281
rect 15983 -10315 16017 -10281
rect 16051 -10315 16085 -10281
rect 16119 -10315 16153 -10281
rect 16187 -10315 16221 -10281
rect 16255 -10315 16289 -10281
rect 16323 -10315 16357 -10281
rect 16391 -10315 16425 -10281
rect 16459 -10315 16493 -10281
rect 16527 -10315 16561 -10281
rect 16595 -10315 16629 -10281
rect 16663 -10315 16697 -10281
rect 16731 -10315 16765 -10281
rect 16799 -10315 16833 -10281
rect 16867 -10315 16901 -10281
rect 16935 -10315 16969 -10281
rect 17003 -10315 17037 -10281
rect 17071 -10315 17105 -10281
rect 17139 -10315 17173 -10281
rect 17207 -10315 17241 -10281
rect 17275 -10315 17309 -10281
rect 17343 -10315 17377 -10281
rect 17411 -10315 17445 -10281
rect 17479 -10315 17513 -10281
rect 17547 -10315 17581 -10281
rect 17615 -10315 17649 -10281
rect 17683 -10315 17717 -10281
rect 17751 -10315 17785 -10281
rect 17819 -10315 17853 -10281
rect 17887 -10315 17921 -10281
rect 17955 -10315 17989 -10281
rect 18023 -10315 18057 -10281
rect 18091 -10315 18125 -10281
rect 18159 -10315 18193 -10281
rect 18227 -10315 18261 -10281
rect 18295 -10315 18329 -10281
rect 18363 -10315 18397 -10281
rect 18431 -10315 18465 -10281
rect 18499 -10315 18533 -10281
rect 18567 -10315 18601 -10281
rect 18635 -10315 18669 -10281
rect 18703 -10315 18737 -10281
rect 18771 -10315 18805 -10281
rect 18839 -10315 18873 -10281
rect 18907 -10315 18941 -10281
rect 18975 -10315 19009 -10281
rect 19043 -10315 19077 -10281
rect 19111 -10315 19145 -10281
rect 19179 -10315 19213 -10281
rect 19247 -10315 19281 -10281
rect 19315 -10315 19349 -10281
rect 19383 -10315 19417 -10281
rect 19451 -10315 19485 -10281
rect 19519 -10315 19553 -10281
rect 19587 -10315 19621 -10281
rect 19655 -10315 19689 -10281
rect 19723 -10315 19757 -10281
rect 19791 -10315 19825 -10281
rect 19859 -10315 19893 -10281
rect 19927 -10315 19961 -10281
rect 19995 -10315 20029 -10281
rect 20063 -10315 20097 -10281
rect 20131 -10315 20165 -10281
rect 20199 -10315 20233 -10281
rect 20267 -10315 20301 -10281
rect 20335 -10315 20369 -10281
rect 20403 -10315 20437 -10281
rect 20471 -10315 20505 -10281
rect 20539 -10315 20573 -10281
rect 20607 -10315 20641 -10281
rect 20675 -10315 20709 -10281
rect 20743 -10315 20777 -10281
rect 20811 -10315 20845 -10281
rect 20879 -10315 20913 -10281
rect 20947 -10315 20981 -10281
rect 21015 -10315 21049 -10281
rect 21083 -10315 21117 -10281
rect 21151 -10315 21185 -10281
rect 21219 -10315 21253 -10281
rect 21287 -10315 21321 -10281
rect 21355 -10315 21389 -10281
rect 21423 -10315 21457 -10281
rect 21491 -10315 21525 -10281
rect 21559 -10315 21593 -10281
rect 21627 -10315 21661 -10281
rect 21695 -10315 21729 -10281
rect 21763 -10315 21797 -10281
rect 21831 -10315 21865 -10281
rect 21899 -10315 21933 -10281
rect 21967 -10315 22001 -10281
rect 22035 -10315 22069 -10281
rect 22103 -10315 22137 -10281
rect 22171 -10315 22205 -10281
rect 22239 -10315 22273 -10281
rect 22307 -10315 22341 -10281
rect 22375 -10315 22409 -10281
rect 22443 -10315 22477 -10281
rect 22511 -10315 22545 -10281
rect 22579 -10315 22613 -10281
rect 22647 -10315 22681 -10281
rect 22715 -10315 22749 -10281
rect 22783 -10315 22817 -10281
rect 22851 -10315 22885 -10281
rect 22919 -10315 22953 -10281
rect 22987 -10315 23021 -10281
rect 23055 -10315 23089 -10281
rect 23123 -10315 23157 -10281
rect 23191 -10315 23225 -10281
rect 23259 -10315 23293 -10281
rect 23327 -10315 23361 -10281
rect 23395 -10315 23429 -10281
rect 23463 -10315 23497 -10281
rect 23531 -10315 23565 -10281
rect 23599 -10315 23633 -10281
rect 23667 -10315 23701 -10281
rect 23735 -10315 23769 -10281
rect 23803 -10315 23837 -10281
rect 23871 -10315 23905 -10281
rect 23939 -10315 23973 -10281
rect 24007 -10315 24041 -10281
rect 24075 -10315 24109 -10281
rect 24143 -10315 24177 -10281
rect 24211 -10315 24245 -10281
rect 24279 -10315 24313 -10281
rect 24347 -10315 24381 -10281
rect 24415 -10315 24449 -10281
rect 24483 -10315 24517 -10281
rect 24551 -10315 24585 -10281
rect 24619 -10315 24653 -10281
<< poly >>
rect -8952 -12440 -8364 -12424
rect -8952 -12457 -8913 -12440
rect -9138 -12474 -8913 -12457
rect -8879 -12474 -8845 -12440
rect -8811 -12474 -8777 -12440
rect -8743 -12474 -8709 -12440
rect -8675 -12474 -8641 -12440
rect -8607 -12474 -8573 -12440
rect -8539 -12474 -8505 -12440
rect -8471 -12474 -8437 -12440
rect -8403 -12457 -8364 -12440
rect -7934 -12440 -7346 -12424
rect -7934 -12457 -7895 -12440
rect -8403 -12474 -8178 -12457
rect -9138 -12512 -8178 -12474
rect -8120 -12474 -7895 -12457
rect -7861 -12474 -7827 -12440
rect -7793 -12474 -7759 -12440
rect -7725 -12474 -7691 -12440
rect -7657 -12474 -7623 -12440
rect -7589 -12474 -7555 -12440
rect -7521 -12474 -7487 -12440
rect -7453 -12474 -7419 -12440
rect -7385 -12457 -7346 -12440
rect -6916 -12440 -6328 -12424
rect -6916 -12457 -6877 -12440
rect -7385 -12474 -7160 -12457
rect -8120 -12512 -7160 -12474
rect -7102 -12474 -6877 -12457
rect -6843 -12474 -6809 -12440
rect -6775 -12474 -6741 -12440
rect -6707 -12474 -6673 -12440
rect -6639 -12474 -6605 -12440
rect -6571 -12474 -6537 -12440
rect -6503 -12474 -6469 -12440
rect -6435 -12474 -6401 -12440
rect -6367 -12457 -6328 -12440
rect -5898 -12440 -5310 -12424
rect -5898 -12457 -5859 -12440
rect -6367 -12474 -6142 -12457
rect -7102 -12512 -6142 -12474
rect -6084 -12474 -5859 -12457
rect -5825 -12474 -5791 -12440
rect -5757 -12474 -5723 -12440
rect -5689 -12474 -5655 -12440
rect -5621 -12474 -5587 -12440
rect -5553 -12474 -5519 -12440
rect -5485 -12474 -5451 -12440
rect -5417 -12474 -5383 -12440
rect -5349 -12457 -5310 -12440
rect -4880 -12440 -4292 -12424
rect -4880 -12457 -4841 -12440
rect -5349 -12474 -5124 -12457
rect -6084 -12512 -5124 -12474
rect -5066 -12474 -4841 -12457
rect -4807 -12474 -4773 -12440
rect -4739 -12474 -4705 -12440
rect -4671 -12474 -4637 -12440
rect -4603 -12474 -4569 -12440
rect -4535 -12474 -4501 -12440
rect -4467 -12474 -4433 -12440
rect -4399 -12474 -4365 -12440
rect -4331 -12457 -4292 -12440
rect -3862 -12440 -3274 -12424
rect -3862 -12457 -3823 -12440
rect -4331 -12474 -4106 -12457
rect -5066 -12512 -4106 -12474
rect -4048 -12474 -3823 -12457
rect -3789 -12474 -3755 -12440
rect -3721 -12474 -3687 -12440
rect -3653 -12474 -3619 -12440
rect -3585 -12474 -3551 -12440
rect -3517 -12474 -3483 -12440
rect -3449 -12474 -3415 -12440
rect -3381 -12474 -3347 -12440
rect -3313 -12457 -3274 -12440
rect -2844 -12440 -2256 -12424
rect -2844 -12457 -2805 -12440
rect -3313 -12474 -3088 -12457
rect -4048 -12512 -3088 -12474
rect -3030 -12474 -2805 -12457
rect -2771 -12474 -2737 -12440
rect -2703 -12474 -2669 -12440
rect -2635 -12474 -2601 -12440
rect -2567 -12474 -2533 -12440
rect -2499 -12474 -2465 -12440
rect -2431 -12474 -2397 -12440
rect -2363 -12474 -2329 -12440
rect -2295 -12457 -2256 -12440
rect -1826 -12440 -1238 -12424
rect -1826 -12457 -1787 -12440
rect -2295 -12474 -2070 -12457
rect -3030 -12512 -2070 -12474
rect -2012 -12474 -1787 -12457
rect -1753 -12474 -1719 -12440
rect -1685 -12474 -1651 -12440
rect -1617 -12474 -1583 -12440
rect -1549 -12474 -1515 -12440
rect -1481 -12474 -1447 -12440
rect -1413 -12474 -1379 -12440
rect -1345 -12474 -1311 -12440
rect -1277 -12457 -1238 -12440
rect -808 -12440 -220 -12424
rect -808 -12457 -769 -12440
rect -1277 -12474 -1052 -12457
rect -2012 -12512 -1052 -12474
rect -994 -12474 -769 -12457
rect -735 -12474 -701 -12440
rect -667 -12474 -633 -12440
rect -599 -12474 -565 -12440
rect -531 -12474 -497 -12440
rect -463 -12474 -429 -12440
rect -395 -12474 -361 -12440
rect -327 -12474 -293 -12440
rect -259 -12457 -220 -12440
rect -259 -12474 -34 -12457
rect -994 -12512 -34 -12474
rect -9138 -13150 -8178 -13112
rect -9138 -13167 -8913 -13150
rect -8952 -13184 -8913 -13167
rect -8879 -13184 -8845 -13150
rect -8811 -13184 -8777 -13150
rect -8743 -13184 -8709 -13150
rect -8675 -13184 -8641 -13150
rect -8607 -13184 -8573 -13150
rect -8539 -13184 -8505 -13150
rect -8471 -13184 -8437 -13150
rect -8403 -13167 -8178 -13150
rect -8120 -13150 -7160 -13112
rect -8120 -13167 -7895 -13150
rect -8403 -13184 -8364 -13167
rect -8952 -13200 -8364 -13184
rect -7934 -13184 -7895 -13167
rect -7861 -13184 -7827 -13150
rect -7793 -13184 -7759 -13150
rect -7725 -13184 -7691 -13150
rect -7657 -13184 -7623 -13150
rect -7589 -13184 -7555 -13150
rect -7521 -13184 -7487 -13150
rect -7453 -13184 -7419 -13150
rect -7385 -13167 -7160 -13150
rect -7102 -13150 -6142 -13112
rect -7102 -13167 -6877 -13150
rect -7385 -13184 -7346 -13167
rect -7934 -13200 -7346 -13184
rect -6916 -13184 -6877 -13167
rect -6843 -13184 -6809 -13150
rect -6775 -13184 -6741 -13150
rect -6707 -13184 -6673 -13150
rect -6639 -13184 -6605 -13150
rect -6571 -13184 -6537 -13150
rect -6503 -13184 -6469 -13150
rect -6435 -13184 -6401 -13150
rect -6367 -13167 -6142 -13150
rect -6084 -13150 -5124 -13112
rect -6084 -13167 -5859 -13150
rect -6367 -13184 -6328 -13167
rect -6916 -13200 -6328 -13184
rect -5898 -13184 -5859 -13167
rect -5825 -13184 -5791 -13150
rect -5757 -13184 -5723 -13150
rect -5689 -13184 -5655 -13150
rect -5621 -13184 -5587 -13150
rect -5553 -13184 -5519 -13150
rect -5485 -13184 -5451 -13150
rect -5417 -13184 -5383 -13150
rect -5349 -13167 -5124 -13150
rect -5066 -13150 -4106 -13112
rect -5066 -13167 -4841 -13150
rect -5349 -13184 -5310 -13167
rect -5898 -13200 -5310 -13184
rect -4880 -13184 -4841 -13167
rect -4807 -13184 -4773 -13150
rect -4739 -13184 -4705 -13150
rect -4671 -13184 -4637 -13150
rect -4603 -13184 -4569 -13150
rect -4535 -13184 -4501 -13150
rect -4467 -13184 -4433 -13150
rect -4399 -13184 -4365 -13150
rect -4331 -13167 -4106 -13150
rect -4048 -13150 -3088 -13112
rect -4048 -13167 -3823 -13150
rect -4331 -13184 -4292 -13167
rect -4880 -13200 -4292 -13184
rect -3862 -13184 -3823 -13167
rect -3789 -13184 -3755 -13150
rect -3721 -13184 -3687 -13150
rect -3653 -13184 -3619 -13150
rect -3585 -13184 -3551 -13150
rect -3517 -13184 -3483 -13150
rect -3449 -13184 -3415 -13150
rect -3381 -13184 -3347 -13150
rect -3313 -13167 -3088 -13150
rect -3030 -13150 -2070 -13112
rect -3030 -13167 -2805 -13150
rect -3313 -13184 -3274 -13167
rect -3862 -13200 -3274 -13184
rect -2844 -13184 -2805 -13167
rect -2771 -13184 -2737 -13150
rect -2703 -13184 -2669 -13150
rect -2635 -13184 -2601 -13150
rect -2567 -13184 -2533 -13150
rect -2499 -13184 -2465 -13150
rect -2431 -13184 -2397 -13150
rect -2363 -13184 -2329 -13150
rect -2295 -13167 -2070 -13150
rect -2012 -13150 -1052 -13112
rect -2012 -13167 -1787 -13150
rect -2295 -13184 -2256 -13167
rect -2844 -13200 -2256 -13184
rect -1826 -13184 -1787 -13167
rect -1753 -13184 -1719 -13150
rect -1685 -13184 -1651 -13150
rect -1617 -13184 -1583 -13150
rect -1549 -13184 -1515 -13150
rect -1481 -13184 -1447 -13150
rect -1413 -13184 -1379 -13150
rect -1345 -13184 -1311 -13150
rect -1277 -13167 -1052 -13150
rect -994 -13150 -34 -13112
rect -994 -13167 -769 -13150
rect -1277 -13184 -1238 -13167
rect -1826 -13200 -1238 -13184
rect -808 -13184 -769 -13167
rect -735 -13184 -701 -13150
rect -667 -13184 -633 -13150
rect -599 -13184 -565 -13150
rect -531 -13184 -497 -13150
rect -463 -13184 -429 -13150
rect -395 -13184 -361 -13150
rect -327 -13184 -293 -13150
rect -259 -13167 -34 -13150
rect -259 -13184 -220 -13167
rect -808 -13200 -220 -13184
rect -8952 -13258 -8364 -13242
rect -8952 -13275 -8913 -13258
rect -9138 -13292 -8913 -13275
rect -8879 -13292 -8845 -13258
rect -8811 -13292 -8777 -13258
rect -8743 -13292 -8709 -13258
rect -8675 -13292 -8641 -13258
rect -8607 -13292 -8573 -13258
rect -8539 -13292 -8505 -13258
rect -8471 -13292 -8437 -13258
rect -8403 -13275 -8364 -13258
rect -7934 -13258 -7346 -13242
rect -7934 -13275 -7895 -13258
rect -8403 -13292 -8178 -13275
rect -9138 -13330 -8178 -13292
rect -8120 -13292 -7895 -13275
rect -7861 -13292 -7827 -13258
rect -7793 -13292 -7759 -13258
rect -7725 -13292 -7691 -13258
rect -7657 -13292 -7623 -13258
rect -7589 -13292 -7555 -13258
rect -7521 -13292 -7487 -13258
rect -7453 -13292 -7419 -13258
rect -7385 -13275 -7346 -13258
rect -6916 -13258 -6328 -13242
rect -6916 -13275 -6877 -13258
rect -7385 -13292 -7160 -13275
rect -8120 -13330 -7160 -13292
rect -7102 -13292 -6877 -13275
rect -6843 -13292 -6809 -13258
rect -6775 -13292 -6741 -13258
rect -6707 -13292 -6673 -13258
rect -6639 -13292 -6605 -13258
rect -6571 -13292 -6537 -13258
rect -6503 -13292 -6469 -13258
rect -6435 -13292 -6401 -13258
rect -6367 -13275 -6328 -13258
rect -5898 -13258 -5310 -13242
rect -5898 -13275 -5859 -13258
rect -6367 -13292 -6142 -13275
rect -7102 -13330 -6142 -13292
rect -6084 -13292 -5859 -13275
rect -5825 -13292 -5791 -13258
rect -5757 -13292 -5723 -13258
rect -5689 -13292 -5655 -13258
rect -5621 -13292 -5587 -13258
rect -5553 -13292 -5519 -13258
rect -5485 -13292 -5451 -13258
rect -5417 -13292 -5383 -13258
rect -5349 -13275 -5310 -13258
rect -4880 -13258 -4292 -13242
rect -4880 -13275 -4841 -13258
rect -5349 -13292 -5124 -13275
rect -6084 -13330 -5124 -13292
rect -5066 -13292 -4841 -13275
rect -4807 -13292 -4773 -13258
rect -4739 -13292 -4705 -13258
rect -4671 -13292 -4637 -13258
rect -4603 -13292 -4569 -13258
rect -4535 -13292 -4501 -13258
rect -4467 -13292 -4433 -13258
rect -4399 -13292 -4365 -13258
rect -4331 -13275 -4292 -13258
rect -3862 -13258 -3274 -13242
rect -3862 -13275 -3823 -13258
rect -4331 -13292 -4106 -13275
rect -5066 -13330 -4106 -13292
rect -4048 -13292 -3823 -13275
rect -3789 -13292 -3755 -13258
rect -3721 -13292 -3687 -13258
rect -3653 -13292 -3619 -13258
rect -3585 -13292 -3551 -13258
rect -3517 -13292 -3483 -13258
rect -3449 -13292 -3415 -13258
rect -3381 -13292 -3347 -13258
rect -3313 -13275 -3274 -13258
rect -2844 -13258 -2256 -13242
rect -2844 -13275 -2805 -13258
rect -3313 -13292 -3088 -13275
rect -4048 -13330 -3088 -13292
rect -3030 -13292 -2805 -13275
rect -2771 -13292 -2737 -13258
rect -2703 -13292 -2669 -13258
rect -2635 -13292 -2601 -13258
rect -2567 -13292 -2533 -13258
rect -2499 -13292 -2465 -13258
rect -2431 -13292 -2397 -13258
rect -2363 -13292 -2329 -13258
rect -2295 -13275 -2256 -13258
rect -1826 -13258 -1238 -13242
rect -1826 -13275 -1787 -13258
rect -2295 -13292 -2070 -13275
rect -3030 -13330 -2070 -13292
rect -2012 -13292 -1787 -13275
rect -1753 -13292 -1719 -13258
rect -1685 -13292 -1651 -13258
rect -1617 -13292 -1583 -13258
rect -1549 -13292 -1515 -13258
rect -1481 -13292 -1447 -13258
rect -1413 -13292 -1379 -13258
rect -1345 -13292 -1311 -13258
rect -1277 -13275 -1238 -13258
rect -808 -13258 -220 -13242
rect -808 -13275 -769 -13258
rect -1277 -13292 -1052 -13275
rect -2012 -13330 -1052 -13292
rect -994 -13292 -769 -13275
rect -735 -13292 -701 -13258
rect -667 -13292 -633 -13258
rect -599 -13292 -565 -13258
rect -531 -13292 -497 -13258
rect -463 -13292 -429 -13258
rect -395 -13292 -361 -13258
rect -327 -13292 -293 -13258
rect -259 -13275 -220 -13258
rect -259 -13292 -34 -13275
rect -994 -13330 -34 -13292
rect -9138 -13968 -8178 -13930
rect -9138 -13985 -8913 -13968
rect -8952 -14002 -8913 -13985
rect -8879 -14002 -8845 -13968
rect -8811 -14002 -8777 -13968
rect -8743 -14002 -8709 -13968
rect -8675 -14002 -8641 -13968
rect -8607 -14002 -8573 -13968
rect -8539 -14002 -8505 -13968
rect -8471 -14002 -8437 -13968
rect -8403 -13985 -8178 -13968
rect -8120 -13968 -7160 -13930
rect -8120 -13985 -7895 -13968
rect -8403 -14002 -8364 -13985
rect -8952 -14018 -8364 -14002
rect -7934 -14002 -7895 -13985
rect -7861 -14002 -7827 -13968
rect -7793 -14002 -7759 -13968
rect -7725 -14002 -7691 -13968
rect -7657 -14002 -7623 -13968
rect -7589 -14002 -7555 -13968
rect -7521 -14002 -7487 -13968
rect -7453 -14002 -7419 -13968
rect -7385 -13985 -7160 -13968
rect -7102 -13968 -6142 -13930
rect -7102 -13985 -6877 -13968
rect -7385 -14002 -7346 -13985
rect -7934 -14018 -7346 -14002
rect -6916 -14002 -6877 -13985
rect -6843 -14002 -6809 -13968
rect -6775 -14002 -6741 -13968
rect -6707 -14002 -6673 -13968
rect -6639 -14002 -6605 -13968
rect -6571 -14002 -6537 -13968
rect -6503 -14002 -6469 -13968
rect -6435 -14002 -6401 -13968
rect -6367 -13985 -6142 -13968
rect -6084 -13968 -5124 -13930
rect -6084 -13985 -5859 -13968
rect -6367 -14002 -6328 -13985
rect -6916 -14018 -6328 -14002
rect -5898 -14002 -5859 -13985
rect -5825 -14002 -5791 -13968
rect -5757 -14002 -5723 -13968
rect -5689 -14002 -5655 -13968
rect -5621 -14002 -5587 -13968
rect -5553 -14002 -5519 -13968
rect -5485 -14002 -5451 -13968
rect -5417 -14002 -5383 -13968
rect -5349 -13985 -5124 -13968
rect -5066 -13968 -4106 -13930
rect -5066 -13985 -4841 -13968
rect -5349 -14002 -5310 -13985
rect -5898 -14018 -5310 -14002
rect -4880 -14002 -4841 -13985
rect -4807 -14002 -4773 -13968
rect -4739 -14002 -4705 -13968
rect -4671 -14002 -4637 -13968
rect -4603 -14002 -4569 -13968
rect -4535 -14002 -4501 -13968
rect -4467 -14002 -4433 -13968
rect -4399 -14002 -4365 -13968
rect -4331 -13985 -4106 -13968
rect -4048 -13968 -3088 -13930
rect -4048 -13985 -3823 -13968
rect -4331 -14002 -4292 -13985
rect -4880 -14018 -4292 -14002
rect -3862 -14002 -3823 -13985
rect -3789 -14002 -3755 -13968
rect -3721 -14002 -3687 -13968
rect -3653 -14002 -3619 -13968
rect -3585 -14002 -3551 -13968
rect -3517 -14002 -3483 -13968
rect -3449 -14002 -3415 -13968
rect -3381 -14002 -3347 -13968
rect -3313 -13985 -3088 -13968
rect -3030 -13968 -2070 -13930
rect -3030 -13985 -2805 -13968
rect -3313 -14002 -3274 -13985
rect -3862 -14018 -3274 -14002
rect -2844 -14002 -2805 -13985
rect -2771 -14002 -2737 -13968
rect -2703 -14002 -2669 -13968
rect -2635 -14002 -2601 -13968
rect -2567 -14002 -2533 -13968
rect -2499 -14002 -2465 -13968
rect -2431 -14002 -2397 -13968
rect -2363 -14002 -2329 -13968
rect -2295 -13985 -2070 -13968
rect -2012 -13968 -1052 -13930
rect -2012 -13985 -1787 -13968
rect -2295 -14002 -2256 -13985
rect -2844 -14018 -2256 -14002
rect -1826 -14002 -1787 -13985
rect -1753 -14002 -1719 -13968
rect -1685 -14002 -1651 -13968
rect -1617 -14002 -1583 -13968
rect -1549 -14002 -1515 -13968
rect -1481 -14002 -1447 -13968
rect -1413 -14002 -1379 -13968
rect -1345 -14002 -1311 -13968
rect -1277 -13985 -1052 -13968
rect -994 -13968 -34 -13930
rect -994 -13985 -769 -13968
rect -1277 -14002 -1238 -13985
rect -1826 -14018 -1238 -14002
rect -808 -14002 -769 -13985
rect -735 -14002 -701 -13968
rect -667 -14002 -633 -13968
rect -599 -14002 -565 -13968
rect -531 -14002 -497 -13968
rect -463 -14002 -429 -13968
rect -395 -14002 -361 -13968
rect -327 -14002 -293 -13968
rect -259 -13985 -34 -13968
rect -259 -14002 -220 -13985
rect -808 -14018 -220 -14002
rect -8952 -14076 -8364 -14060
rect -8952 -14093 -8913 -14076
rect -9138 -14110 -8913 -14093
rect -8879 -14110 -8845 -14076
rect -8811 -14110 -8777 -14076
rect -8743 -14110 -8709 -14076
rect -8675 -14110 -8641 -14076
rect -8607 -14110 -8573 -14076
rect -8539 -14110 -8505 -14076
rect -8471 -14110 -8437 -14076
rect -8403 -14093 -8364 -14076
rect -7934 -14076 -7346 -14060
rect -7934 -14093 -7895 -14076
rect -8403 -14110 -8178 -14093
rect -9138 -14148 -8178 -14110
rect -8120 -14110 -7895 -14093
rect -7861 -14110 -7827 -14076
rect -7793 -14110 -7759 -14076
rect -7725 -14110 -7691 -14076
rect -7657 -14110 -7623 -14076
rect -7589 -14110 -7555 -14076
rect -7521 -14110 -7487 -14076
rect -7453 -14110 -7419 -14076
rect -7385 -14093 -7346 -14076
rect -6916 -14076 -6328 -14060
rect -6916 -14093 -6877 -14076
rect -7385 -14110 -7160 -14093
rect -8120 -14148 -7160 -14110
rect -7102 -14110 -6877 -14093
rect -6843 -14110 -6809 -14076
rect -6775 -14110 -6741 -14076
rect -6707 -14110 -6673 -14076
rect -6639 -14110 -6605 -14076
rect -6571 -14110 -6537 -14076
rect -6503 -14110 -6469 -14076
rect -6435 -14110 -6401 -14076
rect -6367 -14093 -6328 -14076
rect -5898 -14076 -5310 -14060
rect -5898 -14093 -5859 -14076
rect -6367 -14110 -6142 -14093
rect -7102 -14148 -6142 -14110
rect -6084 -14110 -5859 -14093
rect -5825 -14110 -5791 -14076
rect -5757 -14110 -5723 -14076
rect -5689 -14110 -5655 -14076
rect -5621 -14110 -5587 -14076
rect -5553 -14110 -5519 -14076
rect -5485 -14110 -5451 -14076
rect -5417 -14110 -5383 -14076
rect -5349 -14093 -5310 -14076
rect -4880 -14076 -4292 -14060
rect -4880 -14093 -4841 -14076
rect -5349 -14110 -5124 -14093
rect -6084 -14148 -5124 -14110
rect -5066 -14110 -4841 -14093
rect -4807 -14110 -4773 -14076
rect -4739 -14110 -4705 -14076
rect -4671 -14110 -4637 -14076
rect -4603 -14110 -4569 -14076
rect -4535 -14110 -4501 -14076
rect -4467 -14110 -4433 -14076
rect -4399 -14110 -4365 -14076
rect -4331 -14093 -4292 -14076
rect -3862 -14076 -3274 -14060
rect -3862 -14093 -3823 -14076
rect -4331 -14110 -4106 -14093
rect -5066 -14148 -4106 -14110
rect -4048 -14110 -3823 -14093
rect -3789 -14110 -3755 -14076
rect -3721 -14110 -3687 -14076
rect -3653 -14110 -3619 -14076
rect -3585 -14110 -3551 -14076
rect -3517 -14110 -3483 -14076
rect -3449 -14110 -3415 -14076
rect -3381 -14110 -3347 -14076
rect -3313 -14093 -3274 -14076
rect -2844 -14076 -2256 -14060
rect -2844 -14093 -2805 -14076
rect -3313 -14110 -3088 -14093
rect -4048 -14148 -3088 -14110
rect -3030 -14110 -2805 -14093
rect -2771 -14110 -2737 -14076
rect -2703 -14110 -2669 -14076
rect -2635 -14110 -2601 -14076
rect -2567 -14110 -2533 -14076
rect -2499 -14110 -2465 -14076
rect -2431 -14110 -2397 -14076
rect -2363 -14110 -2329 -14076
rect -2295 -14093 -2256 -14076
rect -1826 -14076 -1238 -14060
rect -1826 -14093 -1787 -14076
rect -2295 -14110 -2070 -14093
rect -3030 -14148 -2070 -14110
rect -2012 -14110 -1787 -14093
rect -1753 -14110 -1719 -14076
rect -1685 -14110 -1651 -14076
rect -1617 -14110 -1583 -14076
rect -1549 -14110 -1515 -14076
rect -1481 -14110 -1447 -14076
rect -1413 -14110 -1379 -14076
rect -1345 -14110 -1311 -14076
rect -1277 -14093 -1238 -14076
rect -808 -14076 -220 -14060
rect -808 -14093 -769 -14076
rect -1277 -14110 -1052 -14093
rect -2012 -14148 -1052 -14110
rect -994 -14110 -769 -14093
rect -735 -14110 -701 -14076
rect -667 -14110 -633 -14076
rect -599 -14110 -565 -14076
rect -531 -14110 -497 -14076
rect -463 -14110 -429 -14076
rect -395 -14110 -361 -14076
rect -327 -14110 -293 -14076
rect -259 -14093 -220 -14076
rect -259 -14110 -34 -14093
rect -994 -14148 -34 -14110
rect 2814 -14160 3402 -14144
rect 2814 -14177 2853 -14160
rect 2628 -14194 2853 -14177
rect 2887 -14194 2921 -14160
rect 2955 -14194 2989 -14160
rect 3023 -14194 3057 -14160
rect 3091 -14194 3125 -14160
rect 3159 -14194 3193 -14160
rect 3227 -14194 3261 -14160
rect 3295 -14194 3329 -14160
rect 3363 -14177 3402 -14160
rect 3832 -14160 4420 -14144
rect 3832 -14177 3871 -14160
rect 3363 -14194 3588 -14177
rect 2628 -14232 3588 -14194
rect 3646 -14194 3871 -14177
rect 3905 -14194 3939 -14160
rect 3973 -14194 4007 -14160
rect 4041 -14194 4075 -14160
rect 4109 -14194 4143 -14160
rect 4177 -14194 4211 -14160
rect 4245 -14194 4279 -14160
rect 4313 -14194 4347 -14160
rect 4381 -14177 4420 -14160
rect 4850 -14160 5438 -14144
rect 4850 -14177 4889 -14160
rect 4381 -14194 4606 -14177
rect 3646 -14232 4606 -14194
rect 4664 -14194 4889 -14177
rect 4923 -14194 4957 -14160
rect 4991 -14194 5025 -14160
rect 5059 -14194 5093 -14160
rect 5127 -14194 5161 -14160
rect 5195 -14194 5229 -14160
rect 5263 -14194 5297 -14160
rect 5331 -14194 5365 -14160
rect 5399 -14177 5438 -14160
rect 5868 -14160 6456 -14144
rect 5868 -14177 5907 -14160
rect 5399 -14194 5624 -14177
rect 4664 -14232 5624 -14194
rect 5682 -14194 5907 -14177
rect 5941 -14194 5975 -14160
rect 6009 -14194 6043 -14160
rect 6077 -14194 6111 -14160
rect 6145 -14194 6179 -14160
rect 6213 -14194 6247 -14160
rect 6281 -14194 6315 -14160
rect 6349 -14194 6383 -14160
rect 6417 -14177 6456 -14160
rect 6886 -14160 7474 -14144
rect 6886 -14177 6925 -14160
rect 6417 -14194 6642 -14177
rect 5682 -14232 6642 -14194
rect 6700 -14194 6925 -14177
rect 6959 -14194 6993 -14160
rect 7027 -14194 7061 -14160
rect 7095 -14194 7129 -14160
rect 7163 -14194 7197 -14160
rect 7231 -14194 7265 -14160
rect 7299 -14194 7333 -14160
rect 7367 -14194 7401 -14160
rect 7435 -14177 7474 -14160
rect 7904 -14160 8492 -14144
rect 7904 -14177 7943 -14160
rect 7435 -14194 7660 -14177
rect 6700 -14232 7660 -14194
rect 7718 -14194 7943 -14177
rect 7977 -14194 8011 -14160
rect 8045 -14194 8079 -14160
rect 8113 -14194 8147 -14160
rect 8181 -14194 8215 -14160
rect 8249 -14194 8283 -14160
rect 8317 -14194 8351 -14160
rect 8385 -14194 8419 -14160
rect 8453 -14177 8492 -14160
rect 8922 -14160 9510 -14144
rect 8922 -14177 8961 -14160
rect 8453 -14194 8678 -14177
rect 7718 -14232 8678 -14194
rect 8736 -14194 8961 -14177
rect 8995 -14194 9029 -14160
rect 9063 -14194 9097 -14160
rect 9131 -14194 9165 -14160
rect 9199 -14194 9233 -14160
rect 9267 -14194 9301 -14160
rect 9335 -14194 9369 -14160
rect 9403 -14194 9437 -14160
rect 9471 -14177 9510 -14160
rect 9940 -14160 10528 -14144
rect 9940 -14177 9979 -14160
rect 9471 -14194 9696 -14177
rect 8736 -14232 9696 -14194
rect 9754 -14194 9979 -14177
rect 10013 -14194 10047 -14160
rect 10081 -14194 10115 -14160
rect 10149 -14194 10183 -14160
rect 10217 -14194 10251 -14160
rect 10285 -14194 10319 -14160
rect 10353 -14194 10387 -14160
rect 10421 -14194 10455 -14160
rect 10489 -14177 10528 -14160
rect 10958 -14160 11546 -14144
rect 10958 -14177 10997 -14160
rect 10489 -14194 10714 -14177
rect 9754 -14232 10714 -14194
rect 10772 -14194 10997 -14177
rect 11031 -14194 11065 -14160
rect 11099 -14194 11133 -14160
rect 11167 -14194 11201 -14160
rect 11235 -14194 11269 -14160
rect 11303 -14194 11337 -14160
rect 11371 -14194 11405 -14160
rect 11439 -14194 11473 -14160
rect 11507 -14177 11546 -14160
rect 11976 -14160 12564 -14144
rect 11976 -14177 12015 -14160
rect 11507 -14194 11732 -14177
rect 10772 -14232 11732 -14194
rect 11790 -14194 12015 -14177
rect 12049 -14194 12083 -14160
rect 12117 -14194 12151 -14160
rect 12185 -14194 12219 -14160
rect 12253 -14194 12287 -14160
rect 12321 -14194 12355 -14160
rect 12389 -14194 12423 -14160
rect 12457 -14194 12491 -14160
rect 12525 -14177 12564 -14160
rect 12994 -14160 13582 -14144
rect 12994 -14177 13033 -14160
rect 12525 -14194 12750 -14177
rect 11790 -14232 12750 -14194
rect 12808 -14194 13033 -14177
rect 13067 -14194 13101 -14160
rect 13135 -14194 13169 -14160
rect 13203 -14194 13237 -14160
rect 13271 -14194 13305 -14160
rect 13339 -14194 13373 -14160
rect 13407 -14194 13441 -14160
rect 13475 -14194 13509 -14160
rect 13543 -14177 13582 -14160
rect 14012 -14160 14600 -14144
rect 14012 -14177 14051 -14160
rect 13543 -14194 13768 -14177
rect 12808 -14232 13768 -14194
rect 13826 -14194 14051 -14177
rect 14085 -14194 14119 -14160
rect 14153 -14194 14187 -14160
rect 14221 -14194 14255 -14160
rect 14289 -14194 14323 -14160
rect 14357 -14194 14391 -14160
rect 14425 -14194 14459 -14160
rect 14493 -14194 14527 -14160
rect 14561 -14177 14600 -14160
rect 15030 -14160 15618 -14144
rect 15030 -14177 15069 -14160
rect 14561 -14194 14786 -14177
rect 13826 -14232 14786 -14194
rect 14844 -14194 15069 -14177
rect 15103 -14194 15137 -14160
rect 15171 -14194 15205 -14160
rect 15239 -14194 15273 -14160
rect 15307 -14194 15341 -14160
rect 15375 -14194 15409 -14160
rect 15443 -14194 15477 -14160
rect 15511 -14194 15545 -14160
rect 15579 -14177 15618 -14160
rect 16048 -14160 16636 -14144
rect 16048 -14177 16087 -14160
rect 15579 -14194 15804 -14177
rect 14844 -14232 15804 -14194
rect 15862 -14194 16087 -14177
rect 16121 -14194 16155 -14160
rect 16189 -14194 16223 -14160
rect 16257 -14194 16291 -14160
rect 16325 -14194 16359 -14160
rect 16393 -14194 16427 -14160
rect 16461 -14194 16495 -14160
rect 16529 -14194 16563 -14160
rect 16597 -14177 16636 -14160
rect 17066 -14160 17654 -14144
rect 17066 -14177 17105 -14160
rect 16597 -14194 16822 -14177
rect 15862 -14232 16822 -14194
rect 16880 -14194 17105 -14177
rect 17139 -14194 17173 -14160
rect 17207 -14194 17241 -14160
rect 17275 -14194 17309 -14160
rect 17343 -14194 17377 -14160
rect 17411 -14194 17445 -14160
rect 17479 -14194 17513 -14160
rect 17547 -14194 17581 -14160
rect 17615 -14177 17654 -14160
rect 18084 -14160 18672 -14144
rect 18084 -14177 18123 -14160
rect 17615 -14194 17840 -14177
rect 16880 -14232 17840 -14194
rect 17898 -14194 18123 -14177
rect 18157 -14194 18191 -14160
rect 18225 -14194 18259 -14160
rect 18293 -14194 18327 -14160
rect 18361 -14194 18395 -14160
rect 18429 -14194 18463 -14160
rect 18497 -14194 18531 -14160
rect 18565 -14194 18599 -14160
rect 18633 -14177 18672 -14160
rect 19102 -14160 19690 -14144
rect 19102 -14177 19141 -14160
rect 18633 -14194 18858 -14177
rect 17898 -14232 18858 -14194
rect 18916 -14194 19141 -14177
rect 19175 -14194 19209 -14160
rect 19243 -14194 19277 -14160
rect 19311 -14194 19345 -14160
rect 19379 -14194 19413 -14160
rect 19447 -14194 19481 -14160
rect 19515 -14194 19549 -14160
rect 19583 -14194 19617 -14160
rect 19651 -14177 19690 -14160
rect 20120 -14160 20708 -14144
rect 20120 -14177 20159 -14160
rect 19651 -14194 19876 -14177
rect 18916 -14232 19876 -14194
rect 19934 -14194 20159 -14177
rect 20193 -14194 20227 -14160
rect 20261 -14194 20295 -14160
rect 20329 -14194 20363 -14160
rect 20397 -14194 20431 -14160
rect 20465 -14194 20499 -14160
rect 20533 -14194 20567 -14160
rect 20601 -14194 20635 -14160
rect 20669 -14177 20708 -14160
rect 21138 -14160 21726 -14144
rect 21138 -14177 21177 -14160
rect 20669 -14194 20894 -14177
rect 19934 -14232 20894 -14194
rect 20952 -14194 21177 -14177
rect 21211 -14194 21245 -14160
rect 21279 -14194 21313 -14160
rect 21347 -14194 21381 -14160
rect 21415 -14194 21449 -14160
rect 21483 -14194 21517 -14160
rect 21551 -14194 21585 -14160
rect 21619 -14194 21653 -14160
rect 21687 -14177 21726 -14160
rect 22156 -14160 22744 -14144
rect 22156 -14177 22195 -14160
rect 21687 -14194 21912 -14177
rect 20952 -14232 21912 -14194
rect 21970 -14194 22195 -14177
rect 22229 -14194 22263 -14160
rect 22297 -14194 22331 -14160
rect 22365 -14194 22399 -14160
rect 22433 -14194 22467 -14160
rect 22501 -14194 22535 -14160
rect 22569 -14194 22603 -14160
rect 22637 -14194 22671 -14160
rect 22705 -14177 22744 -14160
rect 22705 -14194 22930 -14177
rect 21970 -14232 22930 -14194
rect -9138 -14786 -8178 -14748
rect -9138 -14803 -8913 -14786
rect -8952 -14820 -8913 -14803
rect -8879 -14820 -8845 -14786
rect -8811 -14820 -8777 -14786
rect -8743 -14820 -8709 -14786
rect -8675 -14820 -8641 -14786
rect -8607 -14820 -8573 -14786
rect -8539 -14820 -8505 -14786
rect -8471 -14820 -8437 -14786
rect -8403 -14803 -8178 -14786
rect -8120 -14786 -7160 -14748
rect -8120 -14803 -7895 -14786
rect -8403 -14820 -8364 -14803
rect -8952 -14836 -8364 -14820
rect -7934 -14820 -7895 -14803
rect -7861 -14820 -7827 -14786
rect -7793 -14820 -7759 -14786
rect -7725 -14820 -7691 -14786
rect -7657 -14820 -7623 -14786
rect -7589 -14820 -7555 -14786
rect -7521 -14820 -7487 -14786
rect -7453 -14820 -7419 -14786
rect -7385 -14803 -7160 -14786
rect -7102 -14786 -6142 -14748
rect -7102 -14803 -6877 -14786
rect -7385 -14820 -7346 -14803
rect -7934 -14836 -7346 -14820
rect -6916 -14820 -6877 -14803
rect -6843 -14820 -6809 -14786
rect -6775 -14820 -6741 -14786
rect -6707 -14820 -6673 -14786
rect -6639 -14820 -6605 -14786
rect -6571 -14820 -6537 -14786
rect -6503 -14820 -6469 -14786
rect -6435 -14820 -6401 -14786
rect -6367 -14803 -6142 -14786
rect -6084 -14786 -5124 -14748
rect -6084 -14803 -5859 -14786
rect -6367 -14820 -6328 -14803
rect -6916 -14836 -6328 -14820
rect -5898 -14820 -5859 -14803
rect -5825 -14820 -5791 -14786
rect -5757 -14820 -5723 -14786
rect -5689 -14820 -5655 -14786
rect -5621 -14820 -5587 -14786
rect -5553 -14820 -5519 -14786
rect -5485 -14820 -5451 -14786
rect -5417 -14820 -5383 -14786
rect -5349 -14803 -5124 -14786
rect -5066 -14786 -4106 -14748
rect -5066 -14803 -4841 -14786
rect -5349 -14820 -5310 -14803
rect -5898 -14836 -5310 -14820
rect -4880 -14820 -4841 -14803
rect -4807 -14820 -4773 -14786
rect -4739 -14820 -4705 -14786
rect -4671 -14820 -4637 -14786
rect -4603 -14820 -4569 -14786
rect -4535 -14820 -4501 -14786
rect -4467 -14820 -4433 -14786
rect -4399 -14820 -4365 -14786
rect -4331 -14803 -4106 -14786
rect -4048 -14786 -3088 -14748
rect -4048 -14803 -3823 -14786
rect -4331 -14820 -4292 -14803
rect -4880 -14836 -4292 -14820
rect -3862 -14820 -3823 -14803
rect -3789 -14820 -3755 -14786
rect -3721 -14820 -3687 -14786
rect -3653 -14820 -3619 -14786
rect -3585 -14820 -3551 -14786
rect -3517 -14820 -3483 -14786
rect -3449 -14820 -3415 -14786
rect -3381 -14820 -3347 -14786
rect -3313 -14803 -3088 -14786
rect -3030 -14786 -2070 -14748
rect -3030 -14803 -2805 -14786
rect -3313 -14820 -3274 -14803
rect -3862 -14836 -3274 -14820
rect -2844 -14820 -2805 -14803
rect -2771 -14820 -2737 -14786
rect -2703 -14820 -2669 -14786
rect -2635 -14820 -2601 -14786
rect -2567 -14820 -2533 -14786
rect -2499 -14820 -2465 -14786
rect -2431 -14820 -2397 -14786
rect -2363 -14820 -2329 -14786
rect -2295 -14803 -2070 -14786
rect -2012 -14786 -1052 -14748
rect -2012 -14803 -1787 -14786
rect -2295 -14820 -2256 -14803
rect -2844 -14836 -2256 -14820
rect -1826 -14820 -1787 -14803
rect -1753 -14820 -1719 -14786
rect -1685 -14820 -1651 -14786
rect -1617 -14820 -1583 -14786
rect -1549 -14820 -1515 -14786
rect -1481 -14820 -1447 -14786
rect -1413 -14820 -1379 -14786
rect -1345 -14820 -1311 -14786
rect -1277 -14803 -1052 -14786
rect -994 -14786 -34 -14748
rect -994 -14803 -769 -14786
rect -1277 -14820 -1238 -14803
rect -1826 -14836 -1238 -14820
rect -808 -14820 -769 -14803
rect -735 -14820 -701 -14786
rect -667 -14820 -633 -14786
rect -599 -14820 -565 -14786
rect -531 -14820 -497 -14786
rect -463 -14820 -429 -14786
rect -395 -14820 -361 -14786
rect -327 -14820 -293 -14786
rect -259 -14803 -34 -14786
rect -259 -14820 -220 -14803
rect -808 -14836 -220 -14820
rect 2628 -14870 3588 -14832
rect -8952 -14894 -8364 -14878
rect -8952 -14911 -8913 -14894
rect -9138 -14928 -8913 -14911
rect -8879 -14928 -8845 -14894
rect -8811 -14928 -8777 -14894
rect -8743 -14928 -8709 -14894
rect -8675 -14928 -8641 -14894
rect -8607 -14928 -8573 -14894
rect -8539 -14928 -8505 -14894
rect -8471 -14928 -8437 -14894
rect -8403 -14911 -8364 -14894
rect -7934 -14894 -7346 -14878
rect -7934 -14911 -7895 -14894
rect -8403 -14928 -8178 -14911
rect -9138 -14966 -8178 -14928
rect -8120 -14928 -7895 -14911
rect -7861 -14928 -7827 -14894
rect -7793 -14928 -7759 -14894
rect -7725 -14928 -7691 -14894
rect -7657 -14928 -7623 -14894
rect -7589 -14928 -7555 -14894
rect -7521 -14928 -7487 -14894
rect -7453 -14928 -7419 -14894
rect -7385 -14911 -7346 -14894
rect -6916 -14894 -6328 -14878
rect -6916 -14911 -6877 -14894
rect -7385 -14928 -7160 -14911
rect -8120 -14966 -7160 -14928
rect -7102 -14928 -6877 -14911
rect -6843 -14928 -6809 -14894
rect -6775 -14928 -6741 -14894
rect -6707 -14928 -6673 -14894
rect -6639 -14928 -6605 -14894
rect -6571 -14928 -6537 -14894
rect -6503 -14928 -6469 -14894
rect -6435 -14928 -6401 -14894
rect -6367 -14911 -6328 -14894
rect -5898 -14894 -5310 -14878
rect -5898 -14911 -5859 -14894
rect -6367 -14928 -6142 -14911
rect -7102 -14966 -6142 -14928
rect -6084 -14928 -5859 -14911
rect -5825 -14928 -5791 -14894
rect -5757 -14928 -5723 -14894
rect -5689 -14928 -5655 -14894
rect -5621 -14928 -5587 -14894
rect -5553 -14928 -5519 -14894
rect -5485 -14928 -5451 -14894
rect -5417 -14928 -5383 -14894
rect -5349 -14911 -5310 -14894
rect -4880 -14894 -4292 -14878
rect -4880 -14911 -4841 -14894
rect -5349 -14928 -5124 -14911
rect -6084 -14966 -5124 -14928
rect -5066 -14928 -4841 -14911
rect -4807 -14928 -4773 -14894
rect -4739 -14928 -4705 -14894
rect -4671 -14928 -4637 -14894
rect -4603 -14928 -4569 -14894
rect -4535 -14928 -4501 -14894
rect -4467 -14928 -4433 -14894
rect -4399 -14928 -4365 -14894
rect -4331 -14911 -4292 -14894
rect -3862 -14894 -3274 -14878
rect -3862 -14911 -3823 -14894
rect -4331 -14928 -4106 -14911
rect -5066 -14966 -4106 -14928
rect -4048 -14928 -3823 -14911
rect -3789 -14928 -3755 -14894
rect -3721 -14928 -3687 -14894
rect -3653 -14928 -3619 -14894
rect -3585 -14928 -3551 -14894
rect -3517 -14928 -3483 -14894
rect -3449 -14928 -3415 -14894
rect -3381 -14928 -3347 -14894
rect -3313 -14911 -3274 -14894
rect -2844 -14894 -2256 -14878
rect -2844 -14911 -2805 -14894
rect -3313 -14928 -3088 -14911
rect -4048 -14966 -3088 -14928
rect -3030 -14928 -2805 -14911
rect -2771 -14928 -2737 -14894
rect -2703 -14928 -2669 -14894
rect -2635 -14928 -2601 -14894
rect -2567 -14928 -2533 -14894
rect -2499 -14928 -2465 -14894
rect -2431 -14928 -2397 -14894
rect -2363 -14928 -2329 -14894
rect -2295 -14911 -2256 -14894
rect -1826 -14894 -1238 -14878
rect -1826 -14911 -1787 -14894
rect -2295 -14928 -2070 -14911
rect -3030 -14966 -2070 -14928
rect -2012 -14928 -1787 -14911
rect -1753 -14928 -1719 -14894
rect -1685 -14928 -1651 -14894
rect -1617 -14928 -1583 -14894
rect -1549 -14928 -1515 -14894
rect -1481 -14928 -1447 -14894
rect -1413 -14928 -1379 -14894
rect -1345 -14928 -1311 -14894
rect -1277 -14911 -1238 -14894
rect -808 -14894 -220 -14878
rect 2628 -14887 2853 -14870
rect -808 -14911 -769 -14894
rect -1277 -14928 -1052 -14911
rect -2012 -14966 -1052 -14928
rect -994 -14928 -769 -14911
rect -735 -14928 -701 -14894
rect -667 -14928 -633 -14894
rect -599 -14928 -565 -14894
rect -531 -14928 -497 -14894
rect -463 -14928 -429 -14894
rect -395 -14928 -361 -14894
rect -327 -14928 -293 -14894
rect -259 -14911 -220 -14894
rect 2814 -14904 2853 -14887
rect 2887 -14904 2921 -14870
rect 2955 -14904 2989 -14870
rect 3023 -14904 3057 -14870
rect 3091 -14904 3125 -14870
rect 3159 -14904 3193 -14870
rect 3227 -14904 3261 -14870
rect 3295 -14904 3329 -14870
rect 3363 -14887 3588 -14870
rect 3646 -14870 4606 -14832
rect 3646 -14887 3871 -14870
rect 3363 -14904 3402 -14887
rect -259 -14928 -34 -14911
rect 2814 -14920 3402 -14904
rect 3832 -14904 3871 -14887
rect 3905 -14904 3939 -14870
rect 3973 -14904 4007 -14870
rect 4041 -14904 4075 -14870
rect 4109 -14904 4143 -14870
rect 4177 -14904 4211 -14870
rect 4245 -14904 4279 -14870
rect 4313 -14904 4347 -14870
rect 4381 -14887 4606 -14870
rect 4664 -14870 5624 -14832
rect 4664 -14887 4889 -14870
rect 4381 -14904 4420 -14887
rect 3832 -14920 4420 -14904
rect 4850 -14904 4889 -14887
rect 4923 -14904 4957 -14870
rect 4991 -14904 5025 -14870
rect 5059 -14904 5093 -14870
rect 5127 -14904 5161 -14870
rect 5195 -14904 5229 -14870
rect 5263 -14904 5297 -14870
rect 5331 -14904 5365 -14870
rect 5399 -14887 5624 -14870
rect 5682 -14870 6642 -14832
rect 5682 -14887 5907 -14870
rect 5399 -14904 5438 -14887
rect 4850 -14920 5438 -14904
rect 5868 -14904 5907 -14887
rect 5941 -14904 5975 -14870
rect 6009 -14904 6043 -14870
rect 6077 -14904 6111 -14870
rect 6145 -14904 6179 -14870
rect 6213 -14904 6247 -14870
rect 6281 -14904 6315 -14870
rect 6349 -14904 6383 -14870
rect 6417 -14887 6642 -14870
rect 6700 -14870 7660 -14832
rect 6700 -14887 6925 -14870
rect 6417 -14904 6456 -14887
rect 5868 -14920 6456 -14904
rect 6886 -14904 6925 -14887
rect 6959 -14904 6993 -14870
rect 7027 -14904 7061 -14870
rect 7095 -14904 7129 -14870
rect 7163 -14904 7197 -14870
rect 7231 -14904 7265 -14870
rect 7299 -14904 7333 -14870
rect 7367 -14904 7401 -14870
rect 7435 -14887 7660 -14870
rect 7718 -14870 8678 -14832
rect 7718 -14887 7943 -14870
rect 7435 -14904 7474 -14887
rect 6886 -14920 7474 -14904
rect 7904 -14904 7943 -14887
rect 7977 -14904 8011 -14870
rect 8045 -14904 8079 -14870
rect 8113 -14904 8147 -14870
rect 8181 -14904 8215 -14870
rect 8249 -14904 8283 -14870
rect 8317 -14904 8351 -14870
rect 8385 -14904 8419 -14870
rect 8453 -14887 8678 -14870
rect 8736 -14870 9696 -14832
rect 8736 -14887 8961 -14870
rect 8453 -14904 8492 -14887
rect 7904 -14920 8492 -14904
rect 8922 -14904 8961 -14887
rect 8995 -14904 9029 -14870
rect 9063 -14904 9097 -14870
rect 9131 -14904 9165 -14870
rect 9199 -14904 9233 -14870
rect 9267 -14904 9301 -14870
rect 9335 -14904 9369 -14870
rect 9403 -14904 9437 -14870
rect 9471 -14887 9696 -14870
rect 9754 -14870 10714 -14832
rect 9754 -14887 9979 -14870
rect 9471 -14904 9510 -14887
rect 8922 -14920 9510 -14904
rect 9940 -14904 9979 -14887
rect 10013 -14904 10047 -14870
rect 10081 -14904 10115 -14870
rect 10149 -14904 10183 -14870
rect 10217 -14904 10251 -14870
rect 10285 -14904 10319 -14870
rect 10353 -14904 10387 -14870
rect 10421 -14904 10455 -14870
rect 10489 -14887 10714 -14870
rect 10772 -14870 11732 -14832
rect 10772 -14887 10997 -14870
rect 10489 -14904 10528 -14887
rect 9940 -14920 10528 -14904
rect 10958 -14904 10997 -14887
rect 11031 -14904 11065 -14870
rect 11099 -14904 11133 -14870
rect 11167 -14904 11201 -14870
rect 11235 -14904 11269 -14870
rect 11303 -14904 11337 -14870
rect 11371 -14904 11405 -14870
rect 11439 -14904 11473 -14870
rect 11507 -14887 11732 -14870
rect 11790 -14870 12750 -14832
rect 11790 -14887 12015 -14870
rect 11507 -14904 11546 -14887
rect 10958 -14920 11546 -14904
rect 11976 -14904 12015 -14887
rect 12049 -14904 12083 -14870
rect 12117 -14904 12151 -14870
rect 12185 -14904 12219 -14870
rect 12253 -14904 12287 -14870
rect 12321 -14904 12355 -14870
rect 12389 -14904 12423 -14870
rect 12457 -14904 12491 -14870
rect 12525 -14887 12750 -14870
rect 12808 -14870 13768 -14832
rect 12808 -14887 13033 -14870
rect 12525 -14904 12564 -14887
rect 11976 -14920 12564 -14904
rect 12994 -14904 13033 -14887
rect 13067 -14904 13101 -14870
rect 13135 -14904 13169 -14870
rect 13203 -14904 13237 -14870
rect 13271 -14904 13305 -14870
rect 13339 -14904 13373 -14870
rect 13407 -14904 13441 -14870
rect 13475 -14904 13509 -14870
rect 13543 -14887 13768 -14870
rect 13826 -14870 14786 -14832
rect 13826 -14887 14051 -14870
rect 13543 -14904 13582 -14887
rect 12994 -14920 13582 -14904
rect 14012 -14904 14051 -14887
rect 14085 -14904 14119 -14870
rect 14153 -14904 14187 -14870
rect 14221 -14904 14255 -14870
rect 14289 -14904 14323 -14870
rect 14357 -14904 14391 -14870
rect 14425 -14904 14459 -14870
rect 14493 -14904 14527 -14870
rect 14561 -14887 14786 -14870
rect 14844 -14870 15804 -14832
rect 14844 -14887 15069 -14870
rect 14561 -14904 14600 -14887
rect 14012 -14920 14600 -14904
rect 15030 -14904 15069 -14887
rect 15103 -14904 15137 -14870
rect 15171 -14904 15205 -14870
rect 15239 -14904 15273 -14870
rect 15307 -14904 15341 -14870
rect 15375 -14904 15409 -14870
rect 15443 -14904 15477 -14870
rect 15511 -14904 15545 -14870
rect 15579 -14887 15804 -14870
rect 15862 -14870 16822 -14832
rect 15862 -14887 16087 -14870
rect 15579 -14904 15618 -14887
rect 15030 -14920 15618 -14904
rect 16048 -14904 16087 -14887
rect 16121 -14904 16155 -14870
rect 16189 -14904 16223 -14870
rect 16257 -14904 16291 -14870
rect 16325 -14904 16359 -14870
rect 16393 -14904 16427 -14870
rect 16461 -14904 16495 -14870
rect 16529 -14904 16563 -14870
rect 16597 -14887 16822 -14870
rect 16880 -14870 17840 -14832
rect 16880 -14887 17105 -14870
rect 16597 -14904 16636 -14887
rect 16048 -14920 16636 -14904
rect 17066 -14904 17105 -14887
rect 17139 -14904 17173 -14870
rect 17207 -14904 17241 -14870
rect 17275 -14904 17309 -14870
rect 17343 -14904 17377 -14870
rect 17411 -14904 17445 -14870
rect 17479 -14904 17513 -14870
rect 17547 -14904 17581 -14870
rect 17615 -14887 17840 -14870
rect 17898 -14870 18858 -14832
rect 17898 -14887 18123 -14870
rect 17615 -14904 17654 -14887
rect 17066 -14920 17654 -14904
rect 18084 -14904 18123 -14887
rect 18157 -14904 18191 -14870
rect 18225 -14904 18259 -14870
rect 18293 -14904 18327 -14870
rect 18361 -14904 18395 -14870
rect 18429 -14904 18463 -14870
rect 18497 -14904 18531 -14870
rect 18565 -14904 18599 -14870
rect 18633 -14887 18858 -14870
rect 18916 -14870 19876 -14832
rect 18916 -14887 19141 -14870
rect 18633 -14904 18672 -14887
rect 18084 -14920 18672 -14904
rect 19102 -14904 19141 -14887
rect 19175 -14904 19209 -14870
rect 19243 -14904 19277 -14870
rect 19311 -14904 19345 -14870
rect 19379 -14904 19413 -14870
rect 19447 -14904 19481 -14870
rect 19515 -14904 19549 -14870
rect 19583 -14904 19617 -14870
rect 19651 -14887 19876 -14870
rect 19934 -14870 20894 -14832
rect 19934 -14887 20159 -14870
rect 19651 -14904 19690 -14887
rect 19102 -14920 19690 -14904
rect 20120 -14904 20159 -14887
rect 20193 -14904 20227 -14870
rect 20261 -14904 20295 -14870
rect 20329 -14904 20363 -14870
rect 20397 -14904 20431 -14870
rect 20465 -14904 20499 -14870
rect 20533 -14904 20567 -14870
rect 20601 -14904 20635 -14870
rect 20669 -14887 20894 -14870
rect 20952 -14870 21912 -14832
rect 20952 -14887 21177 -14870
rect 20669 -14904 20708 -14887
rect 20120 -14920 20708 -14904
rect 21138 -14904 21177 -14887
rect 21211 -14904 21245 -14870
rect 21279 -14904 21313 -14870
rect 21347 -14904 21381 -14870
rect 21415 -14904 21449 -14870
rect 21483 -14904 21517 -14870
rect 21551 -14904 21585 -14870
rect 21619 -14904 21653 -14870
rect 21687 -14887 21912 -14870
rect 21970 -14870 22930 -14832
rect 21970 -14887 22195 -14870
rect 21687 -14904 21726 -14887
rect 21138 -14920 21726 -14904
rect 22156 -14904 22195 -14887
rect 22229 -14904 22263 -14870
rect 22297 -14904 22331 -14870
rect 22365 -14904 22399 -14870
rect 22433 -14904 22467 -14870
rect 22501 -14904 22535 -14870
rect 22569 -14904 22603 -14870
rect 22637 -14904 22671 -14870
rect 22705 -14887 22930 -14870
rect 22705 -14904 22744 -14887
rect 22156 -14920 22744 -14904
rect -994 -14966 -34 -14928
rect 2814 -15392 3402 -15376
rect 2814 -15409 2853 -15392
rect 2628 -15426 2853 -15409
rect 2887 -15426 2921 -15392
rect 2955 -15426 2989 -15392
rect 3023 -15426 3057 -15392
rect 3091 -15426 3125 -15392
rect 3159 -15426 3193 -15392
rect 3227 -15426 3261 -15392
rect 3295 -15426 3329 -15392
rect 3363 -15409 3402 -15392
rect 3832 -15392 4420 -15376
rect 3832 -15409 3871 -15392
rect 3363 -15426 3588 -15409
rect 2628 -15464 3588 -15426
rect 3646 -15426 3871 -15409
rect 3905 -15426 3939 -15392
rect 3973 -15426 4007 -15392
rect 4041 -15426 4075 -15392
rect 4109 -15426 4143 -15392
rect 4177 -15426 4211 -15392
rect 4245 -15426 4279 -15392
rect 4313 -15426 4347 -15392
rect 4381 -15409 4420 -15392
rect 4850 -15392 5438 -15376
rect 4850 -15409 4889 -15392
rect 4381 -15426 4606 -15409
rect 3646 -15464 4606 -15426
rect 4664 -15426 4889 -15409
rect 4923 -15426 4957 -15392
rect 4991 -15426 5025 -15392
rect 5059 -15426 5093 -15392
rect 5127 -15426 5161 -15392
rect 5195 -15426 5229 -15392
rect 5263 -15426 5297 -15392
rect 5331 -15426 5365 -15392
rect 5399 -15409 5438 -15392
rect 5868 -15392 6456 -15376
rect 5868 -15409 5907 -15392
rect 5399 -15426 5624 -15409
rect 4664 -15464 5624 -15426
rect 5682 -15426 5907 -15409
rect 5941 -15426 5975 -15392
rect 6009 -15426 6043 -15392
rect 6077 -15426 6111 -15392
rect 6145 -15426 6179 -15392
rect 6213 -15426 6247 -15392
rect 6281 -15426 6315 -15392
rect 6349 -15426 6383 -15392
rect 6417 -15409 6456 -15392
rect 6886 -15392 7474 -15376
rect 6886 -15409 6925 -15392
rect 6417 -15426 6642 -15409
rect 5682 -15464 6642 -15426
rect 6700 -15426 6925 -15409
rect 6959 -15426 6993 -15392
rect 7027 -15426 7061 -15392
rect 7095 -15426 7129 -15392
rect 7163 -15426 7197 -15392
rect 7231 -15426 7265 -15392
rect 7299 -15426 7333 -15392
rect 7367 -15426 7401 -15392
rect 7435 -15409 7474 -15392
rect 7904 -15392 8492 -15376
rect 7904 -15409 7943 -15392
rect 7435 -15426 7660 -15409
rect 6700 -15464 7660 -15426
rect 7718 -15426 7943 -15409
rect 7977 -15426 8011 -15392
rect 8045 -15426 8079 -15392
rect 8113 -15426 8147 -15392
rect 8181 -15426 8215 -15392
rect 8249 -15426 8283 -15392
rect 8317 -15426 8351 -15392
rect 8385 -15426 8419 -15392
rect 8453 -15409 8492 -15392
rect 8922 -15392 9510 -15376
rect 8922 -15409 8961 -15392
rect 8453 -15426 8678 -15409
rect 7718 -15464 8678 -15426
rect 8736 -15426 8961 -15409
rect 8995 -15426 9029 -15392
rect 9063 -15426 9097 -15392
rect 9131 -15426 9165 -15392
rect 9199 -15426 9233 -15392
rect 9267 -15426 9301 -15392
rect 9335 -15426 9369 -15392
rect 9403 -15426 9437 -15392
rect 9471 -15409 9510 -15392
rect 9940 -15392 10528 -15376
rect 9940 -15409 9979 -15392
rect 9471 -15426 9696 -15409
rect 8736 -15464 9696 -15426
rect 9754 -15426 9979 -15409
rect 10013 -15426 10047 -15392
rect 10081 -15426 10115 -15392
rect 10149 -15426 10183 -15392
rect 10217 -15426 10251 -15392
rect 10285 -15426 10319 -15392
rect 10353 -15426 10387 -15392
rect 10421 -15426 10455 -15392
rect 10489 -15409 10528 -15392
rect 10958 -15392 11546 -15376
rect 10958 -15409 10997 -15392
rect 10489 -15426 10714 -15409
rect 9754 -15464 10714 -15426
rect 10772 -15426 10997 -15409
rect 11031 -15426 11065 -15392
rect 11099 -15426 11133 -15392
rect 11167 -15426 11201 -15392
rect 11235 -15426 11269 -15392
rect 11303 -15426 11337 -15392
rect 11371 -15426 11405 -15392
rect 11439 -15426 11473 -15392
rect 11507 -15409 11546 -15392
rect 11976 -15392 12564 -15376
rect 11976 -15409 12015 -15392
rect 11507 -15426 11732 -15409
rect 10772 -15464 11732 -15426
rect 11790 -15426 12015 -15409
rect 12049 -15426 12083 -15392
rect 12117 -15426 12151 -15392
rect 12185 -15426 12219 -15392
rect 12253 -15426 12287 -15392
rect 12321 -15426 12355 -15392
rect 12389 -15426 12423 -15392
rect 12457 -15426 12491 -15392
rect 12525 -15409 12564 -15392
rect 12994 -15392 13582 -15376
rect 12994 -15409 13033 -15392
rect 12525 -15426 12750 -15409
rect 11790 -15464 12750 -15426
rect 12808 -15426 13033 -15409
rect 13067 -15426 13101 -15392
rect 13135 -15426 13169 -15392
rect 13203 -15426 13237 -15392
rect 13271 -15426 13305 -15392
rect 13339 -15426 13373 -15392
rect 13407 -15426 13441 -15392
rect 13475 -15426 13509 -15392
rect 13543 -15409 13582 -15392
rect 14012 -15392 14600 -15376
rect 14012 -15409 14051 -15392
rect 13543 -15426 13768 -15409
rect 12808 -15464 13768 -15426
rect 13826 -15426 14051 -15409
rect 14085 -15426 14119 -15392
rect 14153 -15426 14187 -15392
rect 14221 -15426 14255 -15392
rect 14289 -15426 14323 -15392
rect 14357 -15426 14391 -15392
rect 14425 -15426 14459 -15392
rect 14493 -15426 14527 -15392
rect 14561 -15409 14600 -15392
rect 15030 -15392 15618 -15376
rect 15030 -15409 15069 -15392
rect 14561 -15426 14786 -15409
rect 13826 -15464 14786 -15426
rect 14844 -15426 15069 -15409
rect 15103 -15426 15137 -15392
rect 15171 -15426 15205 -15392
rect 15239 -15426 15273 -15392
rect 15307 -15426 15341 -15392
rect 15375 -15426 15409 -15392
rect 15443 -15426 15477 -15392
rect 15511 -15426 15545 -15392
rect 15579 -15409 15618 -15392
rect 16048 -15392 16636 -15376
rect 16048 -15409 16087 -15392
rect 15579 -15426 15804 -15409
rect 14844 -15464 15804 -15426
rect 15862 -15426 16087 -15409
rect 16121 -15426 16155 -15392
rect 16189 -15426 16223 -15392
rect 16257 -15426 16291 -15392
rect 16325 -15426 16359 -15392
rect 16393 -15426 16427 -15392
rect 16461 -15426 16495 -15392
rect 16529 -15426 16563 -15392
rect 16597 -15409 16636 -15392
rect 17066 -15392 17654 -15376
rect 17066 -15409 17105 -15392
rect 16597 -15426 16822 -15409
rect 15862 -15464 16822 -15426
rect 16880 -15426 17105 -15409
rect 17139 -15426 17173 -15392
rect 17207 -15426 17241 -15392
rect 17275 -15426 17309 -15392
rect 17343 -15426 17377 -15392
rect 17411 -15426 17445 -15392
rect 17479 -15426 17513 -15392
rect 17547 -15426 17581 -15392
rect 17615 -15409 17654 -15392
rect 18084 -15392 18672 -15376
rect 18084 -15409 18123 -15392
rect 17615 -15426 17840 -15409
rect 16880 -15464 17840 -15426
rect 17898 -15426 18123 -15409
rect 18157 -15426 18191 -15392
rect 18225 -15426 18259 -15392
rect 18293 -15426 18327 -15392
rect 18361 -15426 18395 -15392
rect 18429 -15426 18463 -15392
rect 18497 -15426 18531 -15392
rect 18565 -15426 18599 -15392
rect 18633 -15409 18672 -15392
rect 19102 -15392 19690 -15376
rect 19102 -15409 19141 -15392
rect 18633 -15426 18858 -15409
rect 17898 -15464 18858 -15426
rect 18916 -15426 19141 -15409
rect 19175 -15426 19209 -15392
rect 19243 -15426 19277 -15392
rect 19311 -15426 19345 -15392
rect 19379 -15426 19413 -15392
rect 19447 -15426 19481 -15392
rect 19515 -15426 19549 -15392
rect 19583 -15426 19617 -15392
rect 19651 -15409 19690 -15392
rect 20120 -15392 20708 -15376
rect 20120 -15409 20159 -15392
rect 19651 -15426 19876 -15409
rect 18916 -15464 19876 -15426
rect 19934 -15426 20159 -15409
rect 20193 -15426 20227 -15392
rect 20261 -15426 20295 -15392
rect 20329 -15426 20363 -15392
rect 20397 -15426 20431 -15392
rect 20465 -15426 20499 -15392
rect 20533 -15426 20567 -15392
rect 20601 -15426 20635 -15392
rect 20669 -15409 20708 -15392
rect 21138 -15392 21726 -15376
rect 21138 -15409 21177 -15392
rect 20669 -15426 20894 -15409
rect 19934 -15464 20894 -15426
rect 20952 -15426 21177 -15409
rect 21211 -15426 21245 -15392
rect 21279 -15426 21313 -15392
rect 21347 -15426 21381 -15392
rect 21415 -15426 21449 -15392
rect 21483 -15426 21517 -15392
rect 21551 -15426 21585 -15392
rect 21619 -15426 21653 -15392
rect 21687 -15409 21726 -15392
rect 22156 -15392 22744 -15376
rect 22156 -15409 22195 -15392
rect 21687 -15426 21912 -15409
rect 20952 -15464 21912 -15426
rect 21970 -15426 22195 -15409
rect 22229 -15426 22263 -15392
rect 22297 -15426 22331 -15392
rect 22365 -15426 22399 -15392
rect 22433 -15426 22467 -15392
rect 22501 -15426 22535 -15392
rect 22569 -15426 22603 -15392
rect 22637 -15426 22671 -15392
rect 22705 -15409 22744 -15392
rect 22705 -15426 22930 -15409
rect 21970 -15464 22930 -15426
rect -9138 -15604 -8178 -15566
rect -9138 -15621 -8913 -15604
rect -8952 -15638 -8913 -15621
rect -8879 -15638 -8845 -15604
rect -8811 -15638 -8777 -15604
rect -8743 -15638 -8709 -15604
rect -8675 -15638 -8641 -15604
rect -8607 -15638 -8573 -15604
rect -8539 -15638 -8505 -15604
rect -8471 -15638 -8437 -15604
rect -8403 -15621 -8178 -15604
rect -8120 -15604 -7160 -15566
rect -8120 -15621 -7895 -15604
rect -8403 -15638 -8364 -15621
rect -8952 -15654 -8364 -15638
rect -7934 -15638 -7895 -15621
rect -7861 -15638 -7827 -15604
rect -7793 -15638 -7759 -15604
rect -7725 -15638 -7691 -15604
rect -7657 -15638 -7623 -15604
rect -7589 -15638 -7555 -15604
rect -7521 -15638 -7487 -15604
rect -7453 -15638 -7419 -15604
rect -7385 -15621 -7160 -15604
rect -7102 -15604 -6142 -15566
rect -7102 -15621 -6877 -15604
rect -7385 -15638 -7346 -15621
rect -7934 -15654 -7346 -15638
rect -6916 -15638 -6877 -15621
rect -6843 -15638 -6809 -15604
rect -6775 -15638 -6741 -15604
rect -6707 -15638 -6673 -15604
rect -6639 -15638 -6605 -15604
rect -6571 -15638 -6537 -15604
rect -6503 -15638 -6469 -15604
rect -6435 -15638 -6401 -15604
rect -6367 -15621 -6142 -15604
rect -6084 -15604 -5124 -15566
rect -6084 -15621 -5859 -15604
rect -6367 -15638 -6328 -15621
rect -6916 -15654 -6328 -15638
rect -5898 -15638 -5859 -15621
rect -5825 -15638 -5791 -15604
rect -5757 -15638 -5723 -15604
rect -5689 -15638 -5655 -15604
rect -5621 -15638 -5587 -15604
rect -5553 -15638 -5519 -15604
rect -5485 -15638 -5451 -15604
rect -5417 -15638 -5383 -15604
rect -5349 -15621 -5124 -15604
rect -5066 -15604 -4106 -15566
rect -5066 -15621 -4841 -15604
rect -5349 -15638 -5310 -15621
rect -5898 -15654 -5310 -15638
rect -4880 -15638 -4841 -15621
rect -4807 -15638 -4773 -15604
rect -4739 -15638 -4705 -15604
rect -4671 -15638 -4637 -15604
rect -4603 -15638 -4569 -15604
rect -4535 -15638 -4501 -15604
rect -4467 -15638 -4433 -15604
rect -4399 -15638 -4365 -15604
rect -4331 -15621 -4106 -15604
rect -4048 -15604 -3088 -15566
rect -4048 -15621 -3823 -15604
rect -4331 -15638 -4292 -15621
rect -4880 -15654 -4292 -15638
rect -3862 -15638 -3823 -15621
rect -3789 -15638 -3755 -15604
rect -3721 -15638 -3687 -15604
rect -3653 -15638 -3619 -15604
rect -3585 -15638 -3551 -15604
rect -3517 -15638 -3483 -15604
rect -3449 -15638 -3415 -15604
rect -3381 -15638 -3347 -15604
rect -3313 -15621 -3088 -15604
rect -3030 -15604 -2070 -15566
rect -3030 -15621 -2805 -15604
rect -3313 -15638 -3274 -15621
rect -3862 -15654 -3274 -15638
rect -2844 -15638 -2805 -15621
rect -2771 -15638 -2737 -15604
rect -2703 -15638 -2669 -15604
rect -2635 -15638 -2601 -15604
rect -2567 -15638 -2533 -15604
rect -2499 -15638 -2465 -15604
rect -2431 -15638 -2397 -15604
rect -2363 -15638 -2329 -15604
rect -2295 -15621 -2070 -15604
rect -2012 -15604 -1052 -15566
rect -2012 -15621 -1787 -15604
rect -2295 -15638 -2256 -15621
rect -2844 -15654 -2256 -15638
rect -1826 -15638 -1787 -15621
rect -1753 -15638 -1719 -15604
rect -1685 -15638 -1651 -15604
rect -1617 -15638 -1583 -15604
rect -1549 -15638 -1515 -15604
rect -1481 -15638 -1447 -15604
rect -1413 -15638 -1379 -15604
rect -1345 -15638 -1311 -15604
rect -1277 -15621 -1052 -15604
rect -994 -15604 -34 -15566
rect -994 -15621 -769 -15604
rect -1277 -15638 -1238 -15621
rect -1826 -15654 -1238 -15638
rect -808 -15638 -769 -15621
rect -735 -15638 -701 -15604
rect -667 -15638 -633 -15604
rect -599 -15638 -565 -15604
rect -531 -15638 -497 -15604
rect -463 -15638 -429 -15604
rect -395 -15638 -361 -15604
rect -327 -15638 -293 -15604
rect -259 -15621 -34 -15604
rect -259 -15638 -220 -15621
rect -808 -15654 -220 -15638
rect -8952 -15712 -8364 -15696
rect -8952 -15729 -8913 -15712
rect -9138 -15746 -8913 -15729
rect -8879 -15746 -8845 -15712
rect -8811 -15746 -8777 -15712
rect -8743 -15746 -8709 -15712
rect -8675 -15746 -8641 -15712
rect -8607 -15746 -8573 -15712
rect -8539 -15746 -8505 -15712
rect -8471 -15746 -8437 -15712
rect -8403 -15729 -8364 -15712
rect -7934 -15712 -7346 -15696
rect -7934 -15729 -7895 -15712
rect -8403 -15746 -8178 -15729
rect -9138 -15784 -8178 -15746
rect -8120 -15746 -7895 -15729
rect -7861 -15746 -7827 -15712
rect -7793 -15746 -7759 -15712
rect -7725 -15746 -7691 -15712
rect -7657 -15746 -7623 -15712
rect -7589 -15746 -7555 -15712
rect -7521 -15746 -7487 -15712
rect -7453 -15746 -7419 -15712
rect -7385 -15729 -7346 -15712
rect -6916 -15712 -6328 -15696
rect -6916 -15729 -6877 -15712
rect -7385 -15746 -7160 -15729
rect -8120 -15784 -7160 -15746
rect -7102 -15746 -6877 -15729
rect -6843 -15746 -6809 -15712
rect -6775 -15746 -6741 -15712
rect -6707 -15746 -6673 -15712
rect -6639 -15746 -6605 -15712
rect -6571 -15746 -6537 -15712
rect -6503 -15746 -6469 -15712
rect -6435 -15746 -6401 -15712
rect -6367 -15729 -6328 -15712
rect -5898 -15712 -5310 -15696
rect -5898 -15729 -5859 -15712
rect -6367 -15746 -6142 -15729
rect -7102 -15784 -6142 -15746
rect -6084 -15746 -5859 -15729
rect -5825 -15746 -5791 -15712
rect -5757 -15746 -5723 -15712
rect -5689 -15746 -5655 -15712
rect -5621 -15746 -5587 -15712
rect -5553 -15746 -5519 -15712
rect -5485 -15746 -5451 -15712
rect -5417 -15746 -5383 -15712
rect -5349 -15729 -5310 -15712
rect -4880 -15712 -4292 -15696
rect -4880 -15729 -4841 -15712
rect -5349 -15746 -5124 -15729
rect -6084 -15784 -5124 -15746
rect -5066 -15746 -4841 -15729
rect -4807 -15746 -4773 -15712
rect -4739 -15746 -4705 -15712
rect -4671 -15746 -4637 -15712
rect -4603 -15746 -4569 -15712
rect -4535 -15746 -4501 -15712
rect -4467 -15746 -4433 -15712
rect -4399 -15746 -4365 -15712
rect -4331 -15729 -4292 -15712
rect -3862 -15712 -3274 -15696
rect -3862 -15729 -3823 -15712
rect -4331 -15746 -4106 -15729
rect -5066 -15784 -4106 -15746
rect -4048 -15746 -3823 -15729
rect -3789 -15746 -3755 -15712
rect -3721 -15746 -3687 -15712
rect -3653 -15746 -3619 -15712
rect -3585 -15746 -3551 -15712
rect -3517 -15746 -3483 -15712
rect -3449 -15746 -3415 -15712
rect -3381 -15746 -3347 -15712
rect -3313 -15729 -3274 -15712
rect -2844 -15712 -2256 -15696
rect -2844 -15729 -2805 -15712
rect -3313 -15746 -3088 -15729
rect -4048 -15784 -3088 -15746
rect -3030 -15746 -2805 -15729
rect -2771 -15746 -2737 -15712
rect -2703 -15746 -2669 -15712
rect -2635 -15746 -2601 -15712
rect -2567 -15746 -2533 -15712
rect -2499 -15746 -2465 -15712
rect -2431 -15746 -2397 -15712
rect -2363 -15746 -2329 -15712
rect -2295 -15729 -2256 -15712
rect -1826 -15712 -1238 -15696
rect -1826 -15729 -1787 -15712
rect -2295 -15746 -2070 -15729
rect -3030 -15784 -2070 -15746
rect -2012 -15746 -1787 -15729
rect -1753 -15746 -1719 -15712
rect -1685 -15746 -1651 -15712
rect -1617 -15746 -1583 -15712
rect -1549 -15746 -1515 -15712
rect -1481 -15746 -1447 -15712
rect -1413 -15746 -1379 -15712
rect -1345 -15746 -1311 -15712
rect -1277 -15729 -1238 -15712
rect -808 -15712 -220 -15696
rect -808 -15729 -769 -15712
rect -1277 -15746 -1052 -15729
rect -2012 -15784 -1052 -15746
rect -994 -15746 -769 -15729
rect -735 -15746 -701 -15712
rect -667 -15746 -633 -15712
rect -599 -15746 -565 -15712
rect -531 -15746 -497 -15712
rect -463 -15746 -429 -15712
rect -395 -15746 -361 -15712
rect -327 -15746 -293 -15712
rect -259 -15729 -220 -15712
rect -259 -15746 -34 -15729
rect -994 -15784 -34 -15746
rect 2628 -16102 3588 -16064
rect 2628 -16119 2853 -16102
rect 2814 -16136 2853 -16119
rect 2887 -16136 2921 -16102
rect 2955 -16136 2989 -16102
rect 3023 -16136 3057 -16102
rect 3091 -16136 3125 -16102
rect 3159 -16136 3193 -16102
rect 3227 -16136 3261 -16102
rect 3295 -16136 3329 -16102
rect 3363 -16119 3588 -16102
rect 3646 -16102 4606 -16064
rect 3646 -16119 3871 -16102
rect 3363 -16136 3402 -16119
rect 2814 -16152 3402 -16136
rect 3832 -16136 3871 -16119
rect 3905 -16136 3939 -16102
rect 3973 -16136 4007 -16102
rect 4041 -16136 4075 -16102
rect 4109 -16136 4143 -16102
rect 4177 -16136 4211 -16102
rect 4245 -16136 4279 -16102
rect 4313 -16136 4347 -16102
rect 4381 -16119 4606 -16102
rect 4664 -16102 5624 -16064
rect 4664 -16119 4889 -16102
rect 4381 -16136 4420 -16119
rect 3832 -16152 4420 -16136
rect 4850 -16136 4889 -16119
rect 4923 -16136 4957 -16102
rect 4991 -16136 5025 -16102
rect 5059 -16136 5093 -16102
rect 5127 -16136 5161 -16102
rect 5195 -16136 5229 -16102
rect 5263 -16136 5297 -16102
rect 5331 -16136 5365 -16102
rect 5399 -16119 5624 -16102
rect 5682 -16102 6642 -16064
rect 5682 -16119 5907 -16102
rect 5399 -16136 5438 -16119
rect 4850 -16152 5438 -16136
rect 5868 -16136 5907 -16119
rect 5941 -16136 5975 -16102
rect 6009 -16136 6043 -16102
rect 6077 -16136 6111 -16102
rect 6145 -16136 6179 -16102
rect 6213 -16136 6247 -16102
rect 6281 -16136 6315 -16102
rect 6349 -16136 6383 -16102
rect 6417 -16119 6642 -16102
rect 6700 -16102 7660 -16064
rect 6700 -16119 6925 -16102
rect 6417 -16136 6456 -16119
rect 5868 -16152 6456 -16136
rect 6886 -16136 6925 -16119
rect 6959 -16136 6993 -16102
rect 7027 -16136 7061 -16102
rect 7095 -16136 7129 -16102
rect 7163 -16136 7197 -16102
rect 7231 -16136 7265 -16102
rect 7299 -16136 7333 -16102
rect 7367 -16136 7401 -16102
rect 7435 -16119 7660 -16102
rect 7718 -16102 8678 -16064
rect 7718 -16119 7943 -16102
rect 7435 -16136 7474 -16119
rect 6886 -16152 7474 -16136
rect 7904 -16136 7943 -16119
rect 7977 -16136 8011 -16102
rect 8045 -16136 8079 -16102
rect 8113 -16136 8147 -16102
rect 8181 -16136 8215 -16102
rect 8249 -16136 8283 -16102
rect 8317 -16136 8351 -16102
rect 8385 -16136 8419 -16102
rect 8453 -16119 8678 -16102
rect 8736 -16102 9696 -16064
rect 8736 -16119 8961 -16102
rect 8453 -16136 8492 -16119
rect 7904 -16152 8492 -16136
rect 8922 -16136 8961 -16119
rect 8995 -16136 9029 -16102
rect 9063 -16136 9097 -16102
rect 9131 -16136 9165 -16102
rect 9199 -16136 9233 -16102
rect 9267 -16136 9301 -16102
rect 9335 -16136 9369 -16102
rect 9403 -16136 9437 -16102
rect 9471 -16119 9696 -16102
rect 9754 -16102 10714 -16064
rect 9754 -16119 9979 -16102
rect 9471 -16136 9510 -16119
rect 8922 -16152 9510 -16136
rect 9940 -16136 9979 -16119
rect 10013 -16136 10047 -16102
rect 10081 -16136 10115 -16102
rect 10149 -16136 10183 -16102
rect 10217 -16136 10251 -16102
rect 10285 -16136 10319 -16102
rect 10353 -16136 10387 -16102
rect 10421 -16136 10455 -16102
rect 10489 -16119 10714 -16102
rect 10772 -16102 11732 -16064
rect 10772 -16119 10997 -16102
rect 10489 -16136 10528 -16119
rect 9940 -16152 10528 -16136
rect 10958 -16136 10997 -16119
rect 11031 -16136 11065 -16102
rect 11099 -16136 11133 -16102
rect 11167 -16136 11201 -16102
rect 11235 -16136 11269 -16102
rect 11303 -16136 11337 -16102
rect 11371 -16136 11405 -16102
rect 11439 -16136 11473 -16102
rect 11507 -16119 11732 -16102
rect 11790 -16102 12750 -16064
rect 11790 -16119 12015 -16102
rect 11507 -16136 11546 -16119
rect 10958 -16152 11546 -16136
rect 11976 -16136 12015 -16119
rect 12049 -16136 12083 -16102
rect 12117 -16136 12151 -16102
rect 12185 -16136 12219 -16102
rect 12253 -16136 12287 -16102
rect 12321 -16136 12355 -16102
rect 12389 -16136 12423 -16102
rect 12457 -16136 12491 -16102
rect 12525 -16119 12750 -16102
rect 12808 -16102 13768 -16064
rect 12808 -16119 13033 -16102
rect 12525 -16136 12564 -16119
rect 11976 -16152 12564 -16136
rect 12994 -16136 13033 -16119
rect 13067 -16136 13101 -16102
rect 13135 -16136 13169 -16102
rect 13203 -16136 13237 -16102
rect 13271 -16136 13305 -16102
rect 13339 -16136 13373 -16102
rect 13407 -16136 13441 -16102
rect 13475 -16136 13509 -16102
rect 13543 -16119 13768 -16102
rect 13826 -16102 14786 -16064
rect 13826 -16119 14051 -16102
rect 13543 -16136 13582 -16119
rect 12994 -16152 13582 -16136
rect 14012 -16136 14051 -16119
rect 14085 -16136 14119 -16102
rect 14153 -16136 14187 -16102
rect 14221 -16136 14255 -16102
rect 14289 -16136 14323 -16102
rect 14357 -16136 14391 -16102
rect 14425 -16136 14459 -16102
rect 14493 -16136 14527 -16102
rect 14561 -16119 14786 -16102
rect 14844 -16102 15804 -16064
rect 14844 -16119 15069 -16102
rect 14561 -16136 14600 -16119
rect 14012 -16152 14600 -16136
rect 15030 -16136 15069 -16119
rect 15103 -16136 15137 -16102
rect 15171 -16136 15205 -16102
rect 15239 -16136 15273 -16102
rect 15307 -16136 15341 -16102
rect 15375 -16136 15409 -16102
rect 15443 -16136 15477 -16102
rect 15511 -16136 15545 -16102
rect 15579 -16119 15804 -16102
rect 15862 -16102 16822 -16064
rect 15862 -16119 16087 -16102
rect 15579 -16136 15618 -16119
rect 15030 -16152 15618 -16136
rect 16048 -16136 16087 -16119
rect 16121 -16136 16155 -16102
rect 16189 -16136 16223 -16102
rect 16257 -16136 16291 -16102
rect 16325 -16136 16359 -16102
rect 16393 -16136 16427 -16102
rect 16461 -16136 16495 -16102
rect 16529 -16136 16563 -16102
rect 16597 -16119 16822 -16102
rect 16880 -16102 17840 -16064
rect 16880 -16119 17105 -16102
rect 16597 -16136 16636 -16119
rect 16048 -16152 16636 -16136
rect 17066 -16136 17105 -16119
rect 17139 -16136 17173 -16102
rect 17207 -16136 17241 -16102
rect 17275 -16136 17309 -16102
rect 17343 -16136 17377 -16102
rect 17411 -16136 17445 -16102
rect 17479 -16136 17513 -16102
rect 17547 -16136 17581 -16102
rect 17615 -16119 17840 -16102
rect 17898 -16102 18858 -16064
rect 17898 -16119 18123 -16102
rect 17615 -16136 17654 -16119
rect 17066 -16152 17654 -16136
rect 18084 -16136 18123 -16119
rect 18157 -16136 18191 -16102
rect 18225 -16136 18259 -16102
rect 18293 -16136 18327 -16102
rect 18361 -16136 18395 -16102
rect 18429 -16136 18463 -16102
rect 18497 -16136 18531 -16102
rect 18565 -16136 18599 -16102
rect 18633 -16119 18858 -16102
rect 18916 -16102 19876 -16064
rect 18916 -16119 19141 -16102
rect 18633 -16136 18672 -16119
rect 18084 -16152 18672 -16136
rect 19102 -16136 19141 -16119
rect 19175 -16136 19209 -16102
rect 19243 -16136 19277 -16102
rect 19311 -16136 19345 -16102
rect 19379 -16136 19413 -16102
rect 19447 -16136 19481 -16102
rect 19515 -16136 19549 -16102
rect 19583 -16136 19617 -16102
rect 19651 -16119 19876 -16102
rect 19934 -16102 20894 -16064
rect 19934 -16119 20159 -16102
rect 19651 -16136 19690 -16119
rect 19102 -16152 19690 -16136
rect 20120 -16136 20159 -16119
rect 20193 -16136 20227 -16102
rect 20261 -16136 20295 -16102
rect 20329 -16136 20363 -16102
rect 20397 -16136 20431 -16102
rect 20465 -16136 20499 -16102
rect 20533 -16136 20567 -16102
rect 20601 -16136 20635 -16102
rect 20669 -16119 20894 -16102
rect 20952 -16102 21912 -16064
rect 20952 -16119 21177 -16102
rect 20669 -16136 20708 -16119
rect 20120 -16152 20708 -16136
rect 21138 -16136 21177 -16119
rect 21211 -16136 21245 -16102
rect 21279 -16136 21313 -16102
rect 21347 -16136 21381 -16102
rect 21415 -16136 21449 -16102
rect 21483 -16136 21517 -16102
rect 21551 -16136 21585 -16102
rect 21619 -16136 21653 -16102
rect 21687 -16119 21912 -16102
rect 21970 -16102 22930 -16064
rect 21970 -16119 22195 -16102
rect 21687 -16136 21726 -16119
rect 21138 -16152 21726 -16136
rect 22156 -16136 22195 -16119
rect 22229 -16136 22263 -16102
rect 22297 -16136 22331 -16102
rect 22365 -16136 22399 -16102
rect 22433 -16136 22467 -16102
rect 22501 -16136 22535 -16102
rect 22569 -16136 22603 -16102
rect 22637 -16136 22671 -16102
rect 22705 -16119 22930 -16102
rect 22705 -16136 22744 -16119
rect 22156 -16152 22744 -16136
rect -9138 -16422 -8178 -16384
rect -9138 -16439 -8913 -16422
rect -8952 -16456 -8913 -16439
rect -8879 -16456 -8845 -16422
rect -8811 -16456 -8777 -16422
rect -8743 -16456 -8709 -16422
rect -8675 -16456 -8641 -16422
rect -8607 -16456 -8573 -16422
rect -8539 -16456 -8505 -16422
rect -8471 -16456 -8437 -16422
rect -8403 -16439 -8178 -16422
rect -8120 -16422 -7160 -16384
rect -8120 -16439 -7895 -16422
rect -8403 -16456 -8364 -16439
rect -8952 -16472 -8364 -16456
rect -7934 -16456 -7895 -16439
rect -7861 -16456 -7827 -16422
rect -7793 -16456 -7759 -16422
rect -7725 -16456 -7691 -16422
rect -7657 -16456 -7623 -16422
rect -7589 -16456 -7555 -16422
rect -7521 -16456 -7487 -16422
rect -7453 -16456 -7419 -16422
rect -7385 -16439 -7160 -16422
rect -7102 -16422 -6142 -16384
rect -7102 -16439 -6877 -16422
rect -7385 -16456 -7346 -16439
rect -7934 -16472 -7346 -16456
rect -6916 -16456 -6877 -16439
rect -6843 -16456 -6809 -16422
rect -6775 -16456 -6741 -16422
rect -6707 -16456 -6673 -16422
rect -6639 -16456 -6605 -16422
rect -6571 -16456 -6537 -16422
rect -6503 -16456 -6469 -16422
rect -6435 -16456 -6401 -16422
rect -6367 -16439 -6142 -16422
rect -6084 -16422 -5124 -16384
rect -6084 -16439 -5859 -16422
rect -6367 -16456 -6328 -16439
rect -6916 -16472 -6328 -16456
rect -5898 -16456 -5859 -16439
rect -5825 -16456 -5791 -16422
rect -5757 -16456 -5723 -16422
rect -5689 -16456 -5655 -16422
rect -5621 -16456 -5587 -16422
rect -5553 -16456 -5519 -16422
rect -5485 -16456 -5451 -16422
rect -5417 -16456 -5383 -16422
rect -5349 -16439 -5124 -16422
rect -5066 -16422 -4106 -16384
rect -5066 -16439 -4841 -16422
rect -5349 -16456 -5310 -16439
rect -5898 -16472 -5310 -16456
rect -4880 -16456 -4841 -16439
rect -4807 -16456 -4773 -16422
rect -4739 -16456 -4705 -16422
rect -4671 -16456 -4637 -16422
rect -4603 -16456 -4569 -16422
rect -4535 -16456 -4501 -16422
rect -4467 -16456 -4433 -16422
rect -4399 -16456 -4365 -16422
rect -4331 -16439 -4106 -16422
rect -4048 -16422 -3088 -16384
rect -4048 -16439 -3823 -16422
rect -4331 -16456 -4292 -16439
rect -4880 -16472 -4292 -16456
rect -3862 -16456 -3823 -16439
rect -3789 -16456 -3755 -16422
rect -3721 -16456 -3687 -16422
rect -3653 -16456 -3619 -16422
rect -3585 -16456 -3551 -16422
rect -3517 -16456 -3483 -16422
rect -3449 -16456 -3415 -16422
rect -3381 -16456 -3347 -16422
rect -3313 -16439 -3088 -16422
rect -3030 -16422 -2070 -16384
rect -3030 -16439 -2805 -16422
rect -3313 -16456 -3274 -16439
rect -3862 -16472 -3274 -16456
rect -2844 -16456 -2805 -16439
rect -2771 -16456 -2737 -16422
rect -2703 -16456 -2669 -16422
rect -2635 -16456 -2601 -16422
rect -2567 -16456 -2533 -16422
rect -2499 -16456 -2465 -16422
rect -2431 -16456 -2397 -16422
rect -2363 -16456 -2329 -16422
rect -2295 -16439 -2070 -16422
rect -2012 -16422 -1052 -16384
rect -2012 -16439 -1787 -16422
rect -2295 -16456 -2256 -16439
rect -2844 -16472 -2256 -16456
rect -1826 -16456 -1787 -16439
rect -1753 -16456 -1719 -16422
rect -1685 -16456 -1651 -16422
rect -1617 -16456 -1583 -16422
rect -1549 -16456 -1515 -16422
rect -1481 -16456 -1447 -16422
rect -1413 -16456 -1379 -16422
rect -1345 -16456 -1311 -16422
rect -1277 -16439 -1052 -16422
rect -994 -16422 -34 -16384
rect -994 -16439 -769 -16422
rect -1277 -16456 -1238 -16439
rect -1826 -16472 -1238 -16456
rect -808 -16456 -769 -16439
rect -735 -16456 -701 -16422
rect -667 -16456 -633 -16422
rect -599 -16456 -565 -16422
rect -531 -16456 -497 -16422
rect -463 -16456 -429 -16422
rect -395 -16456 -361 -16422
rect -327 -16456 -293 -16422
rect -259 -16439 -34 -16422
rect -259 -16456 -220 -16439
rect -808 -16472 -220 -16456
rect -8952 -16530 -8364 -16514
rect -8952 -16547 -8913 -16530
rect -9138 -16564 -8913 -16547
rect -8879 -16564 -8845 -16530
rect -8811 -16564 -8777 -16530
rect -8743 -16564 -8709 -16530
rect -8675 -16564 -8641 -16530
rect -8607 -16564 -8573 -16530
rect -8539 -16564 -8505 -16530
rect -8471 -16564 -8437 -16530
rect -8403 -16547 -8364 -16530
rect -7934 -16530 -7346 -16514
rect -7934 -16547 -7895 -16530
rect -8403 -16564 -8178 -16547
rect -9138 -16602 -8178 -16564
rect -8120 -16564 -7895 -16547
rect -7861 -16564 -7827 -16530
rect -7793 -16564 -7759 -16530
rect -7725 -16564 -7691 -16530
rect -7657 -16564 -7623 -16530
rect -7589 -16564 -7555 -16530
rect -7521 -16564 -7487 -16530
rect -7453 -16564 -7419 -16530
rect -7385 -16547 -7346 -16530
rect -6916 -16530 -6328 -16514
rect -6916 -16547 -6877 -16530
rect -7385 -16564 -7160 -16547
rect -8120 -16602 -7160 -16564
rect -7102 -16564 -6877 -16547
rect -6843 -16564 -6809 -16530
rect -6775 -16564 -6741 -16530
rect -6707 -16564 -6673 -16530
rect -6639 -16564 -6605 -16530
rect -6571 -16564 -6537 -16530
rect -6503 -16564 -6469 -16530
rect -6435 -16564 -6401 -16530
rect -6367 -16547 -6328 -16530
rect -5898 -16530 -5310 -16514
rect -5898 -16547 -5859 -16530
rect -6367 -16564 -6142 -16547
rect -7102 -16602 -6142 -16564
rect -6084 -16564 -5859 -16547
rect -5825 -16564 -5791 -16530
rect -5757 -16564 -5723 -16530
rect -5689 -16564 -5655 -16530
rect -5621 -16564 -5587 -16530
rect -5553 -16564 -5519 -16530
rect -5485 -16564 -5451 -16530
rect -5417 -16564 -5383 -16530
rect -5349 -16547 -5310 -16530
rect -4880 -16530 -4292 -16514
rect -4880 -16547 -4841 -16530
rect -5349 -16564 -5124 -16547
rect -6084 -16602 -5124 -16564
rect -5066 -16564 -4841 -16547
rect -4807 -16564 -4773 -16530
rect -4739 -16564 -4705 -16530
rect -4671 -16564 -4637 -16530
rect -4603 -16564 -4569 -16530
rect -4535 -16564 -4501 -16530
rect -4467 -16564 -4433 -16530
rect -4399 -16564 -4365 -16530
rect -4331 -16547 -4292 -16530
rect -3862 -16530 -3274 -16514
rect -3862 -16547 -3823 -16530
rect -4331 -16564 -4106 -16547
rect -5066 -16602 -4106 -16564
rect -4048 -16564 -3823 -16547
rect -3789 -16564 -3755 -16530
rect -3721 -16564 -3687 -16530
rect -3653 -16564 -3619 -16530
rect -3585 -16564 -3551 -16530
rect -3517 -16564 -3483 -16530
rect -3449 -16564 -3415 -16530
rect -3381 -16564 -3347 -16530
rect -3313 -16547 -3274 -16530
rect -2844 -16530 -2256 -16514
rect -2844 -16547 -2805 -16530
rect -3313 -16564 -3088 -16547
rect -4048 -16602 -3088 -16564
rect -3030 -16564 -2805 -16547
rect -2771 -16564 -2737 -16530
rect -2703 -16564 -2669 -16530
rect -2635 -16564 -2601 -16530
rect -2567 -16564 -2533 -16530
rect -2499 -16564 -2465 -16530
rect -2431 -16564 -2397 -16530
rect -2363 -16564 -2329 -16530
rect -2295 -16547 -2256 -16530
rect -1826 -16530 -1238 -16514
rect -1826 -16547 -1787 -16530
rect -2295 -16564 -2070 -16547
rect -3030 -16602 -2070 -16564
rect -2012 -16564 -1787 -16547
rect -1753 -16564 -1719 -16530
rect -1685 -16564 -1651 -16530
rect -1617 -16564 -1583 -16530
rect -1549 -16564 -1515 -16530
rect -1481 -16564 -1447 -16530
rect -1413 -16564 -1379 -16530
rect -1345 -16564 -1311 -16530
rect -1277 -16547 -1238 -16530
rect -808 -16530 -220 -16514
rect -808 -16547 -769 -16530
rect -1277 -16564 -1052 -16547
rect -2012 -16602 -1052 -16564
rect -994 -16564 -769 -16547
rect -735 -16564 -701 -16530
rect -667 -16564 -633 -16530
rect -599 -16564 -565 -16530
rect -531 -16564 -497 -16530
rect -463 -16564 -429 -16530
rect -395 -16564 -361 -16530
rect -327 -16564 -293 -16530
rect -259 -16547 -220 -16530
rect -259 -16564 -34 -16547
rect -994 -16602 -34 -16564
rect 2812 -16626 3400 -16610
rect 2812 -16643 2851 -16626
rect 2626 -16660 2851 -16643
rect 2885 -16660 2919 -16626
rect 2953 -16660 2987 -16626
rect 3021 -16660 3055 -16626
rect 3089 -16660 3123 -16626
rect 3157 -16660 3191 -16626
rect 3225 -16660 3259 -16626
rect 3293 -16660 3327 -16626
rect 3361 -16643 3400 -16626
rect 3830 -16626 4418 -16610
rect 3830 -16643 3869 -16626
rect 3361 -16660 3586 -16643
rect 2626 -16698 3586 -16660
rect 3644 -16660 3869 -16643
rect 3903 -16660 3937 -16626
rect 3971 -16660 4005 -16626
rect 4039 -16660 4073 -16626
rect 4107 -16660 4141 -16626
rect 4175 -16660 4209 -16626
rect 4243 -16660 4277 -16626
rect 4311 -16660 4345 -16626
rect 4379 -16643 4418 -16626
rect 4848 -16626 5436 -16610
rect 4848 -16643 4887 -16626
rect 4379 -16660 4604 -16643
rect 3644 -16698 4604 -16660
rect 4662 -16660 4887 -16643
rect 4921 -16660 4955 -16626
rect 4989 -16660 5023 -16626
rect 5057 -16660 5091 -16626
rect 5125 -16660 5159 -16626
rect 5193 -16660 5227 -16626
rect 5261 -16660 5295 -16626
rect 5329 -16660 5363 -16626
rect 5397 -16643 5436 -16626
rect 5866 -16626 6454 -16610
rect 5866 -16643 5905 -16626
rect 5397 -16660 5622 -16643
rect 4662 -16698 5622 -16660
rect 5680 -16660 5905 -16643
rect 5939 -16660 5973 -16626
rect 6007 -16660 6041 -16626
rect 6075 -16660 6109 -16626
rect 6143 -16660 6177 -16626
rect 6211 -16660 6245 -16626
rect 6279 -16660 6313 -16626
rect 6347 -16660 6381 -16626
rect 6415 -16643 6454 -16626
rect 6884 -16626 7472 -16610
rect 6884 -16643 6923 -16626
rect 6415 -16660 6640 -16643
rect 5680 -16698 6640 -16660
rect 6698 -16660 6923 -16643
rect 6957 -16660 6991 -16626
rect 7025 -16660 7059 -16626
rect 7093 -16660 7127 -16626
rect 7161 -16660 7195 -16626
rect 7229 -16660 7263 -16626
rect 7297 -16660 7331 -16626
rect 7365 -16660 7399 -16626
rect 7433 -16643 7472 -16626
rect 7902 -16626 8490 -16610
rect 7902 -16643 7941 -16626
rect 7433 -16660 7658 -16643
rect 6698 -16698 7658 -16660
rect 7716 -16660 7941 -16643
rect 7975 -16660 8009 -16626
rect 8043 -16660 8077 -16626
rect 8111 -16660 8145 -16626
rect 8179 -16660 8213 -16626
rect 8247 -16660 8281 -16626
rect 8315 -16660 8349 -16626
rect 8383 -16660 8417 -16626
rect 8451 -16643 8490 -16626
rect 8920 -16626 9508 -16610
rect 8920 -16643 8959 -16626
rect 8451 -16660 8676 -16643
rect 7716 -16698 8676 -16660
rect 8734 -16660 8959 -16643
rect 8993 -16660 9027 -16626
rect 9061 -16660 9095 -16626
rect 9129 -16660 9163 -16626
rect 9197 -16660 9231 -16626
rect 9265 -16660 9299 -16626
rect 9333 -16660 9367 -16626
rect 9401 -16660 9435 -16626
rect 9469 -16643 9508 -16626
rect 9938 -16626 10526 -16610
rect 9938 -16643 9977 -16626
rect 9469 -16660 9694 -16643
rect 8734 -16698 9694 -16660
rect 9752 -16660 9977 -16643
rect 10011 -16660 10045 -16626
rect 10079 -16660 10113 -16626
rect 10147 -16660 10181 -16626
rect 10215 -16660 10249 -16626
rect 10283 -16660 10317 -16626
rect 10351 -16660 10385 -16626
rect 10419 -16660 10453 -16626
rect 10487 -16643 10526 -16626
rect 10956 -16626 11544 -16610
rect 10956 -16643 10995 -16626
rect 10487 -16660 10712 -16643
rect 9752 -16698 10712 -16660
rect 10770 -16660 10995 -16643
rect 11029 -16660 11063 -16626
rect 11097 -16660 11131 -16626
rect 11165 -16660 11199 -16626
rect 11233 -16660 11267 -16626
rect 11301 -16660 11335 -16626
rect 11369 -16660 11403 -16626
rect 11437 -16660 11471 -16626
rect 11505 -16643 11544 -16626
rect 11974 -16626 12562 -16610
rect 11974 -16643 12013 -16626
rect 11505 -16660 11730 -16643
rect 10770 -16698 11730 -16660
rect 11788 -16660 12013 -16643
rect 12047 -16660 12081 -16626
rect 12115 -16660 12149 -16626
rect 12183 -16660 12217 -16626
rect 12251 -16660 12285 -16626
rect 12319 -16660 12353 -16626
rect 12387 -16660 12421 -16626
rect 12455 -16660 12489 -16626
rect 12523 -16643 12562 -16626
rect 12992 -16626 13580 -16610
rect 12992 -16643 13031 -16626
rect 12523 -16660 12748 -16643
rect 11788 -16698 12748 -16660
rect 12806 -16660 13031 -16643
rect 13065 -16660 13099 -16626
rect 13133 -16660 13167 -16626
rect 13201 -16660 13235 -16626
rect 13269 -16660 13303 -16626
rect 13337 -16660 13371 -16626
rect 13405 -16660 13439 -16626
rect 13473 -16660 13507 -16626
rect 13541 -16643 13580 -16626
rect 14010 -16626 14598 -16610
rect 14010 -16643 14049 -16626
rect 13541 -16660 13766 -16643
rect 12806 -16698 13766 -16660
rect 13824 -16660 14049 -16643
rect 14083 -16660 14117 -16626
rect 14151 -16660 14185 -16626
rect 14219 -16660 14253 -16626
rect 14287 -16660 14321 -16626
rect 14355 -16660 14389 -16626
rect 14423 -16660 14457 -16626
rect 14491 -16660 14525 -16626
rect 14559 -16643 14598 -16626
rect 15028 -16626 15616 -16610
rect 15028 -16643 15067 -16626
rect 14559 -16660 14784 -16643
rect 13824 -16698 14784 -16660
rect 14842 -16660 15067 -16643
rect 15101 -16660 15135 -16626
rect 15169 -16660 15203 -16626
rect 15237 -16660 15271 -16626
rect 15305 -16660 15339 -16626
rect 15373 -16660 15407 -16626
rect 15441 -16660 15475 -16626
rect 15509 -16660 15543 -16626
rect 15577 -16643 15616 -16626
rect 16046 -16626 16634 -16610
rect 16046 -16643 16085 -16626
rect 15577 -16660 15802 -16643
rect 14842 -16698 15802 -16660
rect 15860 -16660 16085 -16643
rect 16119 -16660 16153 -16626
rect 16187 -16660 16221 -16626
rect 16255 -16660 16289 -16626
rect 16323 -16660 16357 -16626
rect 16391 -16660 16425 -16626
rect 16459 -16660 16493 -16626
rect 16527 -16660 16561 -16626
rect 16595 -16643 16634 -16626
rect 17064 -16626 17652 -16610
rect 17064 -16643 17103 -16626
rect 16595 -16660 16820 -16643
rect 15860 -16698 16820 -16660
rect 16878 -16660 17103 -16643
rect 17137 -16660 17171 -16626
rect 17205 -16660 17239 -16626
rect 17273 -16660 17307 -16626
rect 17341 -16660 17375 -16626
rect 17409 -16660 17443 -16626
rect 17477 -16660 17511 -16626
rect 17545 -16660 17579 -16626
rect 17613 -16643 17652 -16626
rect 18082 -16626 18670 -16610
rect 18082 -16643 18121 -16626
rect 17613 -16660 17838 -16643
rect 16878 -16698 17838 -16660
rect 17896 -16660 18121 -16643
rect 18155 -16660 18189 -16626
rect 18223 -16660 18257 -16626
rect 18291 -16660 18325 -16626
rect 18359 -16660 18393 -16626
rect 18427 -16660 18461 -16626
rect 18495 -16660 18529 -16626
rect 18563 -16660 18597 -16626
rect 18631 -16643 18670 -16626
rect 19100 -16626 19688 -16610
rect 19100 -16643 19139 -16626
rect 18631 -16660 18856 -16643
rect 17896 -16698 18856 -16660
rect 18914 -16660 19139 -16643
rect 19173 -16660 19207 -16626
rect 19241 -16660 19275 -16626
rect 19309 -16660 19343 -16626
rect 19377 -16660 19411 -16626
rect 19445 -16660 19479 -16626
rect 19513 -16660 19547 -16626
rect 19581 -16660 19615 -16626
rect 19649 -16643 19688 -16626
rect 20118 -16626 20706 -16610
rect 20118 -16643 20157 -16626
rect 19649 -16660 19874 -16643
rect 18914 -16698 19874 -16660
rect 19932 -16660 20157 -16643
rect 20191 -16660 20225 -16626
rect 20259 -16660 20293 -16626
rect 20327 -16660 20361 -16626
rect 20395 -16660 20429 -16626
rect 20463 -16660 20497 -16626
rect 20531 -16660 20565 -16626
rect 20599 -16660 20633 -16626
rect 20667 -16643 20706 -16626
rect 21136 -16626 21724 -16610
rect 21136 -16643 21175 -16626
rect 20667 -16660 20892 -16643
rect 19932 -16698 20892 -16660
rect 20950 -16660 21175 -16643
rect 21209 -16660 21243 -16626
rect 21277 -16660 21311 -16626
rect 21345 -16660 21379 -16626
rect 21413 -16660 21447 -16626
rect 21481 -16660 21515 -16626
rect 21549 -16660 21583 -16626
rect 21617 -16660 21651 -16626
rect 21685 -16643 21724 -16626
rect 22154 -16626 22742 -16610
rect 22154 -16643 22193 -16626
rect 21685 -16660 21910 -16643
rect 20950 -16698 21910 -16660
rect 21968 -16660 22193 -16643
rect 22227 -16660 22261 -16626
rect 22295 -16660 22329 -16626
rect 22363 -16660 22397 -16626
rect 22431 -16660 22465 -16626
rect 22499 -16660 22533 -16626
rect 22567 -16660 22601 -16626
rect 22635 -16660 22669 -16626
rect 22703 -16643 22742 -16626
rect 22703 -16660 22928 -16643
rect 21968 -16698 22928 -16660
rect -9138 -17240 -8178 -17202
rect -9138 -17257 -8913 -17240
rect -8952 -17274 -8913 -17257
rect -8879 -17274 -8845 -17240
rect -8811 -17274 -8777 -17240
rect -8743 -17274 -8709 -17240
rect -8675 -17274 -8641 -17240
rect -8607 -17274 -8573 -17240
rect -8539 -17274 -8505 -17240
rect -8471 -17274 -8437 -17240
rect -8403 -17257 -8178 -17240
rect -8120 -17240 -7160 -17202
rect -8120 -17257 -7895 -17240
rect -8403 -17274 -8364 -17257
rect -8952 -17290 -8364 -17274
rect -7934 -17274 -7895 -17257
rect -7861 -17274 -7827 -17240
rect -7793 -17274 -7759 -17240
rect -7725 -17274 -7691 -17240
rect -7657 -17274 -7623 -17240
rect -7589 -17274 -7555 -17240
rect -7521 -17274 -7487 -17240
rect -7453 -17274 -7419 -17240
rect -7385 -17257 -7160 -17240
rect -7102 -17240 -6142 -17202
rect -7102 -17257 -6877 -17240
rect -7385 -17274 -7346 -17257
rect -7934 -17290 -7346 -17274
rect -6916 -17274 -6877 -17257
rect -6843 -17274 -6809 -17240
rect -6775 -17274 -6741 -17240
rect -6707 -17274 -6673 -17240
rect -6639 -17274 -6605 -17240
rect -6571 -17274 -6537 -17240
rect -6503 -17274 -6469 -17240
rect -6435 -17274 -6401 -17240
rect -6367 -17257 -6142 -17240
rect -6084 -17240 -5124 -17202
rect -6084 -17257 -5859 -17240
rect -6367 -17274 -6328 -17257
rect -6916 -17290 -6328 -17274
rect -5898 -17274 -5859 -17257
rect -5825 -17274 -5791 -17240
rect -5757 -17274 -5723 -17240
rect -5689 -17274 -5655 -17240
rect -5621 -17274 -5587 -17240
rect -5553 -17274 -5519 -17240
rect -5485 -17274 -5451 -17240
rect -5417 -17274 -5383 -17240
rect -5349 -17257 -5124 -17240
rect -5066 -17240 -4106 -17202
rect -5066 -17257 -4841 -17240
rect -5349 -17274 -5310 -17257
rect -5898 -17290 -5310 -17274
rect -4880 -17274 -4841 -17257
rect -4807 -17274 -4773 -17240
rect -4739 -17274 -4705 -17240
rect -4671 -17274 -4637 -17240
rect -4603 -17274 -4569 -17240
rect -4535 -17274 -4501 -17240
rect -4467 -17274 -4433 -17240
rect -4399 -17274 -4365 -17240
rect -4331 -17257 -4106 -17240
rect -4048 -17240 -3088 -17202
rect -4048 -17257 -3823 -17240
rect -4331 -17274 -4292 -17257
rect -4880 -17290 -4292 -17274
rect -3862 -17274 -3823 -17257
rect -3789 -17274 -3755 -17240
rect -3721 -17274 -3687 -17240
rect -3653 -17274 -3619 -17240
rect -3585 -17274 -3551 -17240
rect -3517 -17274 -3483 -17240
rect -3449 -17274 -3415 -17240
rect -3381 -17274 -3347 -17240
rect -3313 -17257 -3088 -17240
rect -3030 -17240 -2070 -17202
rect -3030 -17257 -2805 -17240
rect -3313 -17274 -3274 -17257
rect -3862 -17290 -3274 -17274
rect -2844 -17274 -2805 -17257
rect -2771 -17274 -2737 -17240
rect -2703 -17274 -2669 -17240
rect -2635 -17274 -2601 -17240
rect -2567 -17274 -2533 -17240
rect -2499 -17274 -2465 -17240
rect -2431 -17274 -2397 -17240
rect -2363 -17274 -2329 -17240
rect -2295 -17257 -2070 -17240
rect -2012 -17240 -1052 -17202
rect -2012 -17257 -1787 -17240
rect -2295 -17274 -2256 -17257
rect -2844 -17290 -2256 -17274
rect -1826 -17274 -1787 -17257
rect -1753 -17274 -1719 -17240
rect -1685 -17274 -1651 -17240
rect -1617 -17274 -1583 -17240
rect -1549 -17274 -1515 -17240
rect -1481 -17274 -1447 -17240
rect -1413 -17274 -1379 -17240
rect -1345 -17274 -1311 -17240
rect -1277 -17257 -1052 -17240
rect -994 -17240 -34 -17202
rect -994 -17257 -769 -17240
rect -1277 -17274 -1238 -17257
rect -1826 -17290 -1238 -17274
rect -808 -17274 -769 -17257
rect -735 -17274 -701 -17240
rect -667 -17274 -633 -17240
rect -599 -17274 -565 -17240
rect -531 -17274 -497 -17240
rect -463 -17274 -429 -17240
rect -395 -17274 -361 -17240
rect -327 -17274 -293 -17240
rect -259 -17257 -34 -17240
rect -259 -17274 -220 -17257
rect -808 -17290 -220 -17274
rect -8952 -17348 -8364 -17332
rect -8952 -17365 -8913 -17348
rect -9138 -17382 -8913 -17365
rect -8879 -17382 -8845 -17348
rect -8811 -17382 -8777 -17348
rect -8743 -17382 -8709 -17348
rect -8675 -17382 -8641 -17348
rect -8607 -17382 -8573 -17348
rect -8539 -17382 -8505 -17348
rect -8471 -17382 -8437 -17348
rect -8403 -17365 -8364 -17348
rect -7934 -17348 -7346 -17332
rect -7934 -17365 -7895 -17348
rect -8403 -17382 -8178 -17365
rect -9138 -17420 -8178 -17382
rect -8120 -17382 -7895 -17365
rect -7861 -17382 -7827 -17348
rect -7793 -17382 -7759 -17348
rect -7725 -17382 -7691 -17348
rect -7657 -17382 -7623 -17348
rect -7589 -17382 -7555 -17348
rect -7521 -17382 -7487 -17348
rect -7453 -17382 -7419 -17348
rect -7385 -17365 -7346 -17348
rect -6916 -17348 -6328 -17332
rect -6916 -17365 -6877 -17348
rect -7385 -17382 -7160 -17365
rect -8120 -17420 -7160 -17382
rect -7102 -17382 -6877 -17365
rect -6843 -17382 -6809 -17348
rect -6775 -17382 -6741 -17348
rect -6707 -17382 -6673 -17348
rect -6639 -17382 -6605 -17348
rect -6571 -17382 -6537 -17348
rect -6503 -17382 -6469 -17348
rect -6435 -17382 -6401 -17348
rect -6367 -17365 -6328 -17348
rect -5898 -17348 -5310 -17332
rect -5898 -17365 -5859 -17348
rect -6367 -17382 -6142 -17365
rect -7102 -17420 -6142 -17382
rect -6084 -17382 -5859 -17365
rect -5825 -17382 -5791 -17348
rect -5757 -17382 -5723 -17348
rect -5689 -17382 -5655 -17348
rect -5621 -17382 -5587 -17348
rect -5553 -17382 -5519 -17348
rect -5485 -17382 -5451 -17348
rect -5417 -17382 -5383 -17348
rect -5349 -17365 -5310 -17348
rect -4880 -17348 -4292 -17332
rect -4880 -17365 -4841 -17348
rect -5349 -17382 -5124 -17365
rect -6084 -17420 -5124 -17382
rect -5066 -17382 -4841 -17365
rect -4807 -17382 -4773 -17348
rect -4739 -17382 -4705 -17348
rect -4671 -17382 -4637 -17348
rect -4603 -17382 -4569 -17348
rect -4535 -17382 -4501 -17348
rect -4467 -17382 -4433 -17348
rect -4399 -17382 -4365 -17348
rect -4331 -17365 -4292 -17348
rect -3862 -17348 -3274 -17332
rect -3862 -17365 -3823 -17348
rect -4331 -17382 -4106 -17365
rect -5066 -17420 -4106 -17382
rect -4048 -17382 -3823 -17365
rect -3789 -17382 -3755 -17348
rect -3721 -17382 -3687 -17348
rect -3653 -17382 -3619 -17348
rect -3585 -17382 -3551 -17348
rect -3517 -17382 -3483 -17348
rect -3449 -17382 -3415 -17348
rect -3381 -17382 -3347 -17348
rect -3313 -17365 -3274 -17348
rect -2844 -17348 -2256 -17332
rect -2844 -17365 -2805 -17348
rect -3313 -17382 -3088 -17365
rect -4048 -17420 -3088 -17382
rect -3030 -17382 -2805 -17365
rect -2771 -17382 -2737 -17348
rect -2703 -17382 -2669 -17348
rect -2635 -17382 -2601 -17348
rect -2567 -17382 -2533 -17348
rect -2499 -17382 -2465 -17348
rect -2431 -17382 -2397 -17348
rect -2363 -17382 -2329 -17348
rect -2295 -17365 -2256 -17348
rect -1826 -17348 -1238 -17332
rect -1826 -17365 -1787 -17348
rect -2295 -17382 -2070 -17365
rect -3030 -17420 -2070 -17382
rect -2012 -17382 -1787 -17365
rect -1753 -17382 -1719 -17348
rect -1685 -17382 -1651 -17348
rect -1617 -17382 -1583 -17348
rect -1549 -17382 -1515 -17348
rect -1481 -17382 -1447 -17348
rect -1413 -17382 -1379 -17348
rect -1345 -17382 -1311 -17348
rect -1277 -17365 -1238 -17348
rect -808 -17348 -220 -17332
rect -808 -17365 -769 -17348
rect -1277 -17382 -1052 -17365
rect -2012 -17420 -1052 -17382
rect -994 -17382 -769 -17365
rect -735 -17382 -701 -17348
rect -667 -17382 -633 -17348
rect -599 -17382 -565 -17348
rect -531 -17382 -497 -17348
rect -463 -17382 -429 -17348
rect -395 -17382 -361 -17348
rect -327 -17382 -293 -17348
rect -259 -17365 -220 -17348
rect 2626 -17336 3586 -17298
rect 2626 -17353 2851 -17336
rect -259 -17382 -34 -17365
rect -994 -17420 -34 -17382
rect 2812 -17370 2851 -17353
rect 2885 -17370 2919 -17336
rect 2953 -17370 2987 -17336
rect 3021 -17370 3055 -17336
rect 3089 -17370 3123 -17336
rect 3157 -17370 3191 -17336
rect 3225 -17370 3259 -17336
rect 3293 -17370 3327 -17336
rect 3361 -17353 3586 -17336
rect 3644 -17336 4604 -17298
rect 3644 -17353 3869 -17336
rect 3361 -17370 3400 -17353
rect 2812 -17386 3400 -17370
rect 3830 -17370 3869 -17353
rect 3903 -17370 3937 -17336
rect 3971 -17370 4005 -17336
rect 4039 -17370 4073 -17336
rect 4107 -17370 4141 -17336
rect 4175 -17370 4209 -17336
rect 4243 -17370 4277 -17336
rect 4311 -17370 4345 -17336
rect 4379 -17353 4604 -17336
rect 4662 -17336 5622 -17298
rect 4662 -17353 4887 -17336
rect 4379 -17370 4418 -17353
rect 3830 -17386 4418 -17370
rect 4848 -17370 4887 -17353
rect 4921 -17370 4955 -17336
rect 4989 -17370 5023 -17336
rect 5057 -17370 5091 -17336
rect 5125 -17370 5159 -17336
rect 5193 -17370 5227 -17336
rect 5261 -17370 5295 -17336
rect 5329 -17370 5363 -17336
rect 5397 -17353 5622 -17336
rect 5680 -17336 6640 -17298
rect 5680 -17353 5905 -17336
rect 5397 -17370 5436 -17353
rect 4848 -17386 5436 -17370
rect 5866 -17370 5905 -17353
rect 5939 -17370 5973 -17336
rect 6007 -17370 6041 -17336
rect 6075 -17370 6109 -17336
rect 6143 -17370 6177 -17336
rect 6211 -17370 6245 -17336
rect 6279 -17370 6313 -17336
rect 6347 -17370 6381 -17336
rect 6415 -17353 6640 -17336
rect 6698 -17336 7658 -17298
rect 6698 -17353 6923 -17336
rect 6415 -17370 6454 -17353
rect 5866 -17386 6454 -17370
rect 6884 -17370 6923 -17353
rect 6957 -17370 6991 -17336
rect 7025 -17370 7059 -17336
rect 7093 -17370 7127 -17336
rect 7161 -17370 7195 -17336
rect 7229 -17370 7263 -17336
rect 7297 -17370 7331 -17336
rect 7365 -17370 7399 -17336
rect 7433 -17353 7658 -17336
rect 7716 -17336 8676 -17298
rect 7716 -17353 7941 -17336
rect 7433 -17370 7472 -17353
rect 6884 -17386 7472 -17370
rect 7902 -17370 7941 -17353
rect 7975 -17370 8009 -17336
rect 8043 -17370 8077 -17336
rect 8111 -17370 8145 -17336
rect 8179 -17370 8213 -17336
rect 8247 -17370 8281 -17336
rect 8315 -17370 8349 -17336
rect 8383 -17370 8417 -17336
rect 8451 -17353 8676 -17336
rect 8734 -17336 9694 -17298
rect 8734 -17353 8959 -17336
rect 8451 -17370 8490 -17353
rect 7902 -17386 8490 -17370
rect 8920 -17370 8959 -17353
rect 8993 -17370 9027 -17336
rect 9061 -17370 9095 -17336
rect 9129 -17370 9163 -17336
rect 9197 -17370 9231 -17336
rect 9265 -17370 9299 -17336
rect 9333 -17370 9367 -17336
rect 9401 -17370 9435 -17336
rect 9469 -17353 9694 -17336
rect 9752 -17336 10712 -17298
rect 9752 -17353 9977 -17336
rect 9469 -17370 9508 -17353
rect 8920 -17386 9508 -17370
rect 9938 -17370 9977 -17353
rect 10011 -17370 10045 -17336
rect 10079 -17370 10113 -17336
rect 10147 -17370 10181 -17336
rect 10215 -17370 10249 -17336
rect 10283 -17370 10317 -17336
rect 10351 -17370 10385 -17336
rect 10419 -17370 10453 -17336
rect 10487 -17353 10712 -17336
rect 10770 -17336 11730 -17298
rect 10770 -17353 10995 -17336
rect 10487 -17370 10526 -17353
rect 9938 -17386 10526 -17370
rect 10956 -17370 10995 -17353
rect 11029 -17370 11063 -17336
rect 11097 -17370 11131 -17336
rect 11165 -17370 11199 -17336
rect 11233 -17370 11267 -17336
rect 11301 -17370 11335 -17336
rect 11369 -17370 11403 -17336
rect 11437 -17370 11471 -17336
rect 11505 -17353 11730 -17336
rect 11788 -17336 12748 -17298
rect 11788 -17353 12013 -17336
rect 11505 -17370 11544 -17353
rect 10956 -17386 11544 -17370
rect 11974 -17370 12013 -17353
rect 12047 -17370 12081 -17336
rect 12115 -17370 12149 -17336
rect 12183 -17370 12217 -17336
rect 12251 -17370 12285 -17336
rect 12319 -17370 12353 -17336
rect 12387 -17370 12421 -17336
rect 12455 -17370 12489 -17336
rect 12523 -17353 12748 -17336
rect 12806 -17336 13766 -17298
rect 12806 -17353 13031 -17336
rect 12523 -17370 12562 -17353
rect 11974 -17386 12562 -17370
rect 12992 -17370 13031 -17353
rect 13065 -17370 13099 -17336
rect 13133 -17370 13167 -17336
rect 13201 -17370 13235 -17336
rect 13269 -17370 13303 -17336
rect 13337 -17370 13371 -17336
rect 13405 -17370 13439 -17336
rect 13473 -17370 13507 -17336
rect 13541 -17353 13766 -17336
rect 13824 -17336 14784 -17298
rect 13824 -17353 14049 -17336
rect 13541 -17370 13580 -17353
rect 12992 -17386 13580 -17370
rect 14010 -17370 14049 -17353
rect 14083 -17370 14117 -17336
rect 14151 -17370 14185 -17336
rect 14219 -17370 14253 -17336
rect 14287 -17370 14321 -17336
rect 14355 -17370 14389 -17336
rect 14423 -17370 14457 -17336
rect 14491 -17370 14525 -17336
rect 14559 -17353 14784 -17336
rect 14842 -17336 15802 -17298
rect 14842 -17353 15067 -17336
rect 14559 -17370 14598 -17353
rect 14010 -17386 14598 -17370
rect 15028 -17370 15067 -17353
rect 15101 -17370 15135 -17336
rect 15169 -17370 15203 -17336
rect 15237 -17370 15271 -17336
rect 15305 -17370 15339 -17336
rect 15373 -17370 15407 -17336
rect 15441 -17370 15475 -17336
rect 15509 -17370 15543 -17336
rect 15577 -17353 15802 -17336
rect 15860 -17336 16820 -17298
rect 15860 -17353 16085 -17336
rect 15577 -17370 15616 -17353
rect 15028 -17386 15616 -17370
rect 16046 -17370 16085 -17353
rect 16119 -17370 16153 -17336
rect 16187 -17370 16221 -17336
rect 16255 -17370 16289 -17336
rect 16323 -17370 16357 -17336
rect 16391 -17370 16425 -17336
rect 16459 -17370 16493 -17336
rect 16527 -17370 16561 -17336
rect 16595 -17353 16820 -17336
rect 16878 -17336 17838 -17298
rect 16878 -17353 17103 -17336
rect 16595 -17370 16634 -17353
rect 16046 -17386 16634 -17370
rect 17064 -17370 17103 -17353
rect 17137 -17370 17171 -17336
rect 17205 -17370 17239 -17336
rect 17273 -17370 17307 -17336
rect 17341 -17370 17375 -17336
rect 17409 -17370 17443 -17336
rect 17477 -17370 17511 -17336
rect 17545 -17370 17579 -17336
rect 17613 -17353 17838 -17336
rect 17896 -17336 18856 -17298
rect 17896 -17353 18121 -17336
rect 17613 -17370 17652 -17353
rect 17064 -17386 17652 -17370
rect 18082 -17370 18121 -17353
rect 18155 -17370 18189 -17336
rect 18223 -17370 18257 -17336
rect 18291 -17370 18325 -17336
rect 18359 -17370 18393 -17336
rect 18427 -17370 18461 -17336
rect 18495 -17370 18529 -17336
rect 18563 -17370 18597 -17336
rect 18631 -17353 18856 -17336
rect 18914 -17336 19874 -17298
rect 18914 -17353 19139 -17336
rect 18631 -17370 18670 -17353
rect 18082 -17386 18670 -17370
rect 19100 -17370 19139 -17353
rect 19173 -17370 19207 -17336
rect 19241 -17370 19275 -17336
rect 19309 -17370 19343 -17336
rect 19377 -17370 19411 -17336
rect 19445 -17370 19479 -17336
rect 19513 -17370 19547 -17336
rect 19581 -17370 19615 -17336
rect 19649 -17353 19874 -17336
rect 19932 -17336 20892 -17298
rect 19932 -17353 20157 -17336
rect 19649 -17370 19688 -17353
rect 19100 -17386 19688 -17370
rect 20118 -17370 20157 -17353
rect 20191 -17370 20225 -17336
rect 20259 -17370 20293 -17336
rect 20327 -17370 20361 -17336
rect 20395 -17370 20429 -17336
rect 20463 -17370 20497 -17336
rect 20531 -17370 20565 -17336
rect 20599 -17370 20633 -17336
rect 20667 -17353 20892 -17336
rect 20950 -17336 21910 -17298
rect 20950 -17353 21175 -17336
rect 20667 -17370 20706 -17353
rect 20118 -17386 20706 -17370
rect 21136 -17370 21175 -17353
rect 21209 -17370 21243 -17336
rect 21277 -17370 21311 -17336
rect 21345 -17370 21379 -17336
rect 21413 -17370 21447 -17336
rect 21481 -17370 21515 -17336
rect 21549 -17370 21583 -17336
rect 21617 -17370 21651 -17336
rect 21685 -17353 21910 -17336
rect 21968 -17336 22928 -17298
rect 21968 -17353 22193 -17336
rect 21685 -17370 21724 -17353
rect 21136 -17386 21724 -17370
rect 22154 -17370 22193 -17353
rect 22227 -17370 22261 -17336
rect 22295 -17370 22329 -17336
rect 22363 -17370 22397 -17336
rect 22431 -17370 22465 -17336
rect 22499 -17370 22533 -17336
rect 22567 -17370 22601 -17336
rect 22635 -17370 22669 -17336
rect 22703 -17353 22928 -17336
rect 22703 -17370 22742 -17353
rect 22154 -17386 22742 -17370
rect 2812 -17860 3400 -17844
rect 2812 -17877 2851 -17860
rect 2626 -17894 2851 -17877
rect 2885 -17894 2919 -17860
rect 2953 -17894 2987 -17860
rect 3021 -17894 3055 -17860
rect 3089 -17894 3123 -17860
rect 3157 -17894 3191 -17860
rect 3225 -17894 3259 -17860
rect 3293 -17894 3327 -17860
rect 3361 -17877 3400 -17860
rect 3830 -17860 4418 -17844
rect 3830 -17877 3869 -17860
rect 3361 -17894 3586 -17877
rect 2626 -17932 3586 -17894
rect 3644 -17894 3869 -17877
rect 3903 -17894 3937 -17860
rect 3971 -17894 4005 -17860
rect 4039 -17894 4073 -17860
rect 4107 -17894 4141 -17860
rect 4175 -17894 4209 -17860
rect 4243 -17894 4277 -17860
rect 4311 -17894 4345 -17860
rect 4379 -17877 4418 -17860
rect 4848 -17860 5436 -17844
rect 4848 -17877 4887 -17860
rect 4379 -17894 4604 -17877
rect 3644 -17932 4604 -17894
rect 4662 -17894 4887 -17877
rect 4921 -17894 4955 -17860
rect 4989 -17894 5023 -17860
rect 5057 -17894 5091 -17860
rect 5125 -17894 5159 -17860
rect 5193 -17894 5227 -17860
rect 5261 -17894 5295 -17860
rect 5329 -17894 5363 -17860
rect 5397 -17877 5436 -17860
rect 5866 -17860 6454 -17844
rect 5866 -17877 5905 -17860
rect 5397 -17894 5622 -17877
rect 4662 -17932 5622 -17894
rect 5680 -17894 5905 -17877
rect 5939 -17894 5973 -17860
rect 6007 -17894 6041 -17860
rect 6075 -17894 6109 -17860
rect 6143 -17894 6177 -17860
rect 6211 -17894 6245 -17860
rect 6279 -17894 6313 -17860
rect 6347 -17894 6381 -17860
rect 6415 -17877 6454 -17860
rect 6884 -17860 7472 -17844
rect 6884 -17877 6923 -17860
rect 6415 -17894 6640 -17877
rect 5680 -17932 6640 -17894
rect 6698 -17894 6923 -17877
rect 6957 -17894 6991 -17860
rect 7025 -17894 7059 -17860
rect 7093 -17894 7127 -17860
rect 7161 -17894 7195 -17860
rect 7229 -17894 7263 -17860
rect 7297 -17894 7331 -17860
rect 7365 -17894 7399 -17860
rect 7433 -17877 7472 -17860
rect 7902 -17860 8490 -17844
rect 7902 -17877 7941 -17860
rect 7433 -17894 7658 -17877
rect 6698 -17932 7658 -17894
rect 7716 -17894 7941 -17877
rect 7975 -17894 8009 -17860
rect 8043 -17894 8077 -17860
rect 8111 -17894 8145 -17860
rect 8179 -17894 8213 -17860
rect 8247 -17894 8281 -17860
rect 8315 -17894 8349 -17860
rect 8383 -17894 8417 -17860
rect 8451 -17877 8490 -17860
rect 8920 -17860 9508 -17844
rect 8920 -17877 8959 -17860
rect 8451 -17894 8676 -17877
rect 7716 -17932 8676 -17894
rect 8734 -17894 8959 -17877
rect 8993 -17894 9027 -17860
rect 9061 -17894 9095 -17860
rect 9129 -17894 9163 -17860
rect 9197 -17894 9231 -17860
rect 9265 -17894 9299 -17860
rect 9333 -17894 9367 -17860
rect 9401 -17894 9435 -17860
rect 9469 -17877 9508 -17860
rect 9938 -17860 10526 -17844
rect 9938 -17877 9977 -17860
rect 9469 -17894 9694 -17877
rect 8734 -17932 9694 -17894
rect 9752 -17894 9977 -17877
rect 10011 -17894 10045 -17860
rect 10079 -17894 10113 -17860
rect 10147 -17894 10181 -17860
rect 10215 -17894 10249 -17860
rect 10283 -17894 10317 -17860
rect 10351 -17894 10385 -17860
rect 10419 -17894 10453 -17860
rect 10487 -17877 10526 -17860
rect 10956 -17860 11544 -17844
rect 10956 -17877 10995 -17860
rect 10487 -17894 10712 -17877
rect 9752 -17932 10712 -17894
rect 10770 -17894 10995 -17877
rect 11029 -17894 11063 -17860
rect 11097 -17894 11131 -17860
rect 11165 -17894 11199 -17860
rect 11233 -17894 11267 -17860
rect 11301 -17894 11335 -17860
rect 11369 -17894 11403 -17860
rect 11437 -17894 11471 -17860
rect 11505 -17877 11544 -17860
rect 11974 -17860 12562 -17844
rect 11974 -17877 12013 -17860
rect 11505 -17894 11730 -17877
rect 10770 -17932 11730 -17894
rect 11788 -17894 12013 -17877
rect 12047 -17894 12081 -17860
rect 12115 -17894 12149 -17860
rect 12183 -17894 12217 -17860
rect 12251 -17894 12285 -17860
rect 12319 -17894 12353 -17860
rect 12387 -17894 12421 -17860
rect 12455 -17894 12489 -17860
rect 12523 -17877 12562 -17860
rect 12992 -17860 13580 -17844
rect 12992 -17877 13031 -17860
rect 12523 -17894 12748 -17877
rect 11788 -17932 12748 -17894
rect 12806 -17894 13031 -17877
rect 13065 -17894 13099 -17860
rect 13133 -17894 13167 -17860
rect 13201 -17894 13235 -17860
rect 13269 -17894 13303 -17860
rect 13337 -17894 13371 -17860
rect 13405 -17894 13439 -17860
rect 13473 -17894 13507 -17860
rect 13541 -17877 13580 -17860
rect 14010 -17860 14598 -17844
rect 14010 -17877 14049 -17860
rect 13541 -17894 13766 -17877
rect 12806 -17932 13766 -17894
rect 13824 -17894 14049 -17877
rect 14083 -17894 14117 -17860
rect 14151 -17894 14185 -17860
rect 14219 -17894 14253 -17860
rect 14287 -17894 14321 -17860
rect 14355 -17894 14389 -17860
rect 14423 -17894 14457 -17860
rect 14491 -17894 14525 -17860
rect 14559 -17877 14598 -17860
rect 15028 -17860 15616 -17844
rect 15028 -17877 15067 -17860
rect 14559 -17894 14784 -17877
rect 13824 -17932 14784 -17894
rect 14842 -17894 15067 -17877
rect 15101 -17894 15135 -17860
rect 15169 -17894 15203 -17860
rect 15237 -17894 15271 -17860
rect 15305 -17894 15339 -17860
rect 15373 -17894 15407 -17860
rect 15441 -17894 15475 -17860
rect 15509 -17894 15543 -17860
rect 15577 -17877 15616 -17860
rect 16046 -17860 16634 -17844
rect 16046 -17877 16085 -17860
rect 15577 -17894 15802 -17877
rect 14842 -17932 15802 -17894
rect 15860 -17894 16085 -17877
rect 16119 -17894 16153 -17860
rect 16187 -17894 16221 -17860
rect 16255 -17894 16289 -17860
rect 16323 -17894 16357 -17860
rect 16391 -17894 16425 -17860
rect 16459 -17894 16493 -17860
rect 16527 -17894 16561 -17860
rect 16595 -17877 16634 -17860
rect 17064 -17860 17652 -17844
rect 17064 -17877 17103 -17860
rect 16595 -17894 16820 -17877
rect 15860 -17932 16820 -17894
rect 16878 -17894 17103 -17877
rect 17137 -17894 17171 -17860
rect 17205 -17894 17239 -17860
rect 17273 -17894 17307 -17860
rect 17341 -17894 17375 -17860
rect 17409 -17894 17443 -17860
rect 17477 -17894 17511 -17860
rect 17545 -17894 17579 -17860
rect 17613 -17877 17652 -17860
rect 18082 -17860 18670 -17844
rect 18082 -17877 18121 -17860
rect 17613 -17894 17838 -17877
rect 16878 -17932 17838 -17894
rect 17896 -17894 18121 -17877
rect 18155 -17894 18189 -17860
rect 18223 -17894 18257 -17860
rect 18291 -17894 18325 -17860
rect 18359 -17894 18393 -17860
rect 18427 -17894 18461 -17860
rect 18495 -17894 18529 -17860
rect 18563 -17894 18597 -17860
rect 18631 -17877 18670 -17860
rect 19100 -17860 19688 -17844
rect 19100 -17877 19139 -17860
rect 18631 -17894 18856 -17877
rect 17896 -17932 18856 -17894
rect 18914 -17894 19139 -17877
rect 19173 -17894 19207 -17860
rect 19241 -17894 19275 -17860
rect 19309 -17894 19343 -17860
rect 19377 -17894 19411 -17860
rect 19445 -17894 19479 -17860
rect 19513 -17894 19547 -17860
rect 19581 -17894 19615 -17860
rect 19649 -17877 19688 -17860
rect 20118 -17860 20706 -17844
rect 20118 -17877 20157 -17860
rect 19649 -17894 19874 -17877
rect 18914 -17932 19874 -17894
rect 19932 -17894 20157 -17877
rect 20191 -17894 20225 -17860
rect 20259 -17894 20293 -17860
rect 20327 -17894 20361 -17860
rect 20395 -17894 20429 -17860
rect 20463 -17894 20497 -17860
rect 20531 -17894 20565 -17860
rect 20599 -17894 20633 -17860
rect 20667 -17877 20706 -17860
rect 21136 -17860 21724 -17844
rect 21136 -17877 21175 -17860
rect 20667 -17894 20892 -17877
rect 19932 -17932 20892 -17894
rect 20950 -17894 21175 -17877
rect 21209 -17894 21243 -17860
rect 21277 -17894 21311 -17860
rect 21345 -17894 21379 -17860
rect 21413 -17894 21447 -17860
rect 21481 -17894 21515 -17860
rect 21549 -17894 21583 -17860
rect 21617 -17894 21651 -17860
rect 21685 -17877 21724 -17860
rect 22154 -17860 22742 -17844
rect 22154 -17877 22193 -17860
rect 21685 -17894 21910 -17877
rect 20950 -17932 21910 -17894
rect 21968 -17894 22193 -17877
rect 22227 -17894 22261 -17860
rect 22295 -17894 22329 -17860
rect 22363 -17894 22397 -17860
rect 22431 -17894 22465 -17860
rect 22499 -17894 22533 -17860
rect 22567 -17894 22601 -17860
rect 22635 -17894 22669 -17860
rect 22703 -17877 22742 -17860
rect 22703 -17894 22928 -17877
rect 21968 -17932 22928 -17894
rect -9138 -18058 -8178 -18020
rect -9138 -18075 -8913 -18058
rect -8952 -18092 -8913 -18075
rect -8879 -18092 -8845 -18058
rect -8811 -18092 -8777 -18058
rect -8743 -18092 -8709 -18058
rect -8675 -18092 -8641 -18058
rect -8607 -18092 -8573 -18058
rect -8539 -18092 -8505 -18058
rect -8471 -18092 -8437 -18058
rect -8403 -18075 -8178 -18058
rect -8120 -18058 -7160 -18020
rect -8120 -18075 -7895 -18058
rect -8403 -18092 -8364 -18075
rect -8952 -18108 -8364 -18092
rect -7934 -18092 -7895 -18075
rect -7861 -18092 -7827 -18058
rect -7793 -18092 -7759 -18058
rect -7725 -18092 -7691 -18058
rect -7657 -18092 -7623 -18058
rect -7589 -18092 -7555 -18058
rect -7521 -18092 -7487 -18058
rect -7453 -18092 -7419 -18058
rect -7385 -18075 -7160 -18058
rect -7102 -18058 -6142 -18020
rect -7102 -18075 -6877 -18058
rect -7385 -18092 -7346 -18075
rect -7934 -18108 -7346 -18092
rect -6916 -18092 -6877 -18075
rect -6843 -18092 -6809 -18058
rect -6775 -18092 -6741 -18058
rect -6707 -18092 -6673 -18058
rect -6639 -18092 -6605 -18058
rect -6571 -18092 -6537 -18058
rect -6503 -18092 -6469 -18058
rect -6435 -18092 -6401 -18058
rect -6367 -18075 -6142 -18058
rect -6084 -18058 -5124 -18020
rect -6084 -18075 -5859 -18058
rect -6367 -18092 -6328 -18075
rect -6916 -18108 -6328 -18092
rect -5898 -18092 -5859 -18075
rect -5825 -18092 -5791 -18058
rect -5757 -18092 -5723 -18058
rect -5689 -18092 -5655 -18058
rect -5621 -18092 -5587 -18058
rect -5553 -18092 -5519 -18058
rect -5485 -18092 -5451 -18058
rect -5417 -18092 -5383 -18058
rect -5349 -18075 -5124 -18058
rect -5066 -18058 -4106 -18020
rect -5066 -18075 -4841 -18058
rect -5349 -18092 -5310 -18075
rect -5898 -18108 -5310 -18092
rect -4880 -18092 -4841 -18075
rect -4807 -18092 -4773 -18058
rect -4739 -18092 -4705 -18058
rect -4671 -18092 -4637 -18058
rect -4603 -18092 -4569 -18058
rect -4535 -18092 -4501 -18058
rect -4467 -18092 -4433 -18058
rect -4399 -18092 -4365 -18058
rect -4331 -18075 -4106 -18058
rect -4048 -18058 -3088 -18020
rect -4048 -18075 -3823 -18058
rect -4331 -18092 -4292 -18075
rect -4880 -18108 -4292 -18092
rect -3862 -18092 -3823 -18075
rect -3789 -18092 -3755 -18058
rect -3721 -18092 -3687 -18058
rect -3653 -18092 -3619 -18058
rect -3585 -18092 -3551 -18058
rect -3517 -18092 -3483 -18058
rect -3449 -18092 -3415 -18058
rect -3381 -18092 -3347 -18058
rect -3313 -18075 -3088 -18058
rect -3030 -18058 -2070 -18020
rect -3030 -18075 -2805 -18058
rect -3313 -18092 -3274 -18075
rect -3862 -18108 -3274 -18092
rect -2844 -18092 -2805 -18075
rect -2771 -18092 -2737 -18058
rect -2703 -18092 -2669 -18058
rect -2635 -18092 -2601 -18058
rect -2567 -18092 -2533 -18058
rect -2499 -18092 -2465 -18058
rect -2431 -18092 -2397 -18058
rect -2363 -18092 -2329 -18058
rect -2295 -18075 -2070 -18058
rect -2012 -18058 -1052 -18020
rect -2012 -18075 -1787 -18058
rect -2295 -18092 -2256 -18075
rect -2844 -18108 -2256 -18092
rect -1826 -18092 -1787 -18075
rect -1753 -18092 -1719 -18058
rect -1685 -18092 -1651 -18058
rect -1617 -18092 -1583 -18058
rect -1549 -18092 -1515 -18058
rect -1481 -18092 -1447 -18058
rect -1413 -18092 -1379 -18058
rect -1345 -18092 -1311 -18058
rect -1277 -18075 -1052 -18058
rect -994 -18058 -34 -18020
rect -994 -18075 -769 -18058
rect -1277 -18092 -1238 -18075
rect -1826 -18108 -1238 -18092
rect -808 -18092 -769 -18075
rect -735 -18092 -701 -18058
rect -667 -18092 -633 -18058
rect -599 -18092 -565 -18058
rect -531 -18092 -497 -18058
rect -463 -18092 -429 -18058
rect -395 -18092 -361 -18058
rect -327 -18092 -293 -18058
rect -259 -18075 -34 -18058
rect -259 -18092 -220 -18075
rect -808 -18108 -220 -18092
rect -8952 -18166 -8364 -18150
rect -8952 -18183 -8913 -18166
rect -9138 -18200 -8913 -18183
rect -8879 -18200 -8845 -18166
rect -8811 -18200 -8777 -18166
rect -8743 -18200 -8709 -18166
rect -8675 -18200 -8641 -18166
rect -8607 -18200 -8573 -18166
rect -8539 -18200 -8505 -18166
rect -8471 -18200 -8437 -18166
rect -8403 -18183 -8364 -18166
rect -7934 -18166 -7346 -18150
rect -7934 -18183 -7895 -18166
rect -8403 -18200 -8178 -18183
rect -9138 -18238 -8178 -18200
rect -8120 -18200 -7895 -18183
rect -7861 -18200 -7827 -18166
rect -7793 -18200 -7759 -18166
rect -7725 -18200 -7691 -18166
rect -7657 -18200 -7623 -18166
rect -7589 -18200 -7555 -18166
rect -7521 -18200 -7487 -18166
rect -7453 -18200 -7419 -18166
rect -7385 -18183 -7346 -18166
rect -6916 -18166 -6328 -18150
rect -6916 -18183 -6877 -18166
rect -7385 -18200 -7160 -18183
rect -8120 -18238 -7160 -18200
rect -7102 -18200 -6877 -18183
rect -6843 -18200 -6809 -18166
rect -6775 -18200 -6741 -18166
rect -6707 -18200 -6673 -18166
rect -6639 -18200 -6605 -18166
rect -6571 -18200 -6537 -18166
rect -6503 -18200 -6469 -18166
rect -6435 -18200 -6401 -18166
rect -6367 -18183 -6328 -18166
rect -5898 -18166 -5310 -18150
rect -5898 -18183 -5859 -18166
rect -6367 -18200 -6142 -18183
rect -7102 -18238 -6142 -18200
rect -6084 -18200 -5859 -18183
rect -5825 -18200 -5791 -18166
rect -5757 -18200 -5723 -18166
rect -5689 -18200 -5655 -18166
rect -5621 -18200 -5587 -18166
rect -5553 -18200 -5519 -18166
rect -5485 -18200 -5451 -18166
rect -5417 -18200 -5383 -18166
rect -5349 -18183 -5310 -18166
rect -4880 -18166 -4292 -18150
rect -4880 -18183 -4841 -18166
rect -5349 -18200 -5124 -18183
rect -6084 -18238 -5124 -18200
rect -5066 -18200 -4841 -18183
rect -4807 -18200 -4773 -18166
rect -4739 -18200 -4705 -18166
rect -4671 -18200 -4637 -18166
rect -4603 -18200 -4569 -18166
rect -4535 -18200 -4501 -18166
rect -4467 -18200 -4433 -18166
rect -4399 -18200 -4365 -18166
rect -4331 -18183 -4292 -18166
rect -3862 -18166 -3274 -18150
rect -3862 -18183 -3823 -18166
rect -4331 -18200 -4106 -18183
rect -5066 -18238 -4106 -18200
rect -4048 -18200 -3823 -18183
rect -3789 -18200 -3755 -18166
rect -3721 -18200 -3687 -18166
rect -3653 -18200 -3619 -18166
rect -3585 -18200 -3551 -18166
rect -3517 -18200 -3483 -18166
rect -3449 -18200 -3415 -18166
rect -3381 -18200 -3347 -18166
rect -3313 -18183 -3274 -18166
rect -2844 -18166 -2256 -18150
rect -2844 -18183 -2805 -18166
rect -3313 -18200 -3088 -18183
rect -4048 -18238 -3088 -18200
rect -3030 -18200 -2805 -18183
rect -2771 -18200 -2737 -18166
rect -2703 -18200 -2669 -18166
rect -2635 -18200 -2601 -18166
rect -2567 -18200 -2533 -18166
rect -2499 -18200 -2465 -18166
rect -2431 -18200 -2397 -18166
rect -2363 -18200 -2329 -18166
rect -2295 -18183 -2256 -18166
rect -1826 -18166 -1238 -18150
rect -1826 -18183 -1787 -18166
rect -2295 -18200 -2070 -18183
rect -3030 -18238 -2070 -18200
rect -2012 -18200 -1787 -18183
rect -1753 -18200 -1719 -18166
rect -1685 -18200 -1651 -18166
rect -1617 -18200 -1583 -18166
rect -1549 -18200 -1515 -18166
rect -1481 -18200 -1447 -18166
rect -1413 -18200 -1379 -18166
rect -1345 -18200 -1311 -18166
rect -1277 -18183 -1238 -18166
rect -808 -18166 -220 -18150
rect -808 -18183 -769 -18166
rect -1277 -18200 -1052 -18183
rect -2012 -18238 -1052 -18200
rect -994 -18200 -769 -18183
rect -735 -18200 -701 -18166
rect -667 -18200 -633 -18166
rect -599 -18200 -565 -18166
rect -531 -18200 -497 -18166
rect -463 -18200 -429 -18166
rect -395 -18200 -361 -18166
rect -327 -18200 -293 -18166
rect -259 -18183 -220 -18166
rect -259 -18200 -34 -18183
rect -994 -18238 -34 -18200
rect 2626 -18570 3586 -18532
rect 2626 -18587 2851 -18570
rect 2812 -18604 2851 -18587
rect 2885 -18604 2919 -18570
rect 2953 -18604 2987 -18570
rect 3021 -18604 3055 -18570
rect 3089 -18604 3123 -18570
rect 3157 -18604 3191 -18570
rect 3225 -18604 3259 -18570
rect 3293 -18604 3327 -18570
rect 3361 -18587 3586 -18570
rect 3644 -18570 4604 -18532
rect 3644 -18587 3869 -18570
rect 3361 -18604 3400 -18587
rect 2812 -18620 3400 -18604
rect 3830 -18604 3869 -18587
rect 3903 -18604 3937 -18570
rect 3971 -18604 4005 -18570
rect 4039 -18604 4073 -18570
rect 4107 -18604 4141 -18570
rect 4175 -18604 4209 -18570
rect 4243 -18604 4277 -18570
rect 4311 -18604 4345 -18570
rect 4379 -18587 4604 -18570
rect 4662 -18570 5622 -18532
rect 4662 -18587 4887 -18570
rect 4379 -18604 4418 -18587
rect 3830 -18620 4418 -18604
rect 4848 -18604 4887 -18587
rect 4921 -18604 4955 -18570
rect 4989 -18604 5023 -18570
rect 5057 -18604 5091 -18570
rect 5125 -18604 5159 -18570
rect 5193 -18604 5227 -18570
rect 5261 -18604 5295 -18570
rect 5329 -18604 5363 -18570
rect 5397 -18587 5622 -18570
rect 5680 -18570 6640 -18532
rect 5680 -18587 5905 -18570
rect 5397 -18604 5436 -18587
rect 4848 -18620 5436 -18604
rect 5866 -18604 5905 -18587
rect 5939 -18604 5973 -18570
rect 6007 -18604 6041 -18570
rect 6075 -18604 6109 -18570
rect 6143 -18604 6177 -18570
rect 6211 -18604 6245 -18570
rect 6279 -18604 6313 -18570
rect 6347 -18604 6381 -18570
rect 6415 -18587 6640 -18570
rect 6698 -18570 7658 -18532
rect 6698 -18587 6923 -18570
rect 6415 -18604 6454 -18587
rect 5866 -18620 6454 -18604
rect 6884 -18604 6923 -18587
rect 6957 -18604 6991 -18570
rect 7025 -18604 7059 -18570
rect 7093 -18604 7127 -18570
rect 7161 -18604 7195 -18570
rect 7229 -18604 7263 -18570
rect 7297 -18604 7331 -18570
rect 7365 -18604 7399 -18570
rect 7433 -18587 7658 -18570
rect 7716 -18570 8676 -18532
rect 7716 -18587 7941 -18570
rect 7433 -18604 7472 -18587
rect 6884 -18620 7472 -18604
rect 7902 -18604 7941 -18587
rect 7975 -18604 8009 -18570
rect 8043 -18604 8077 -18570
rect 8111 -18604 8145 -18570
rect 8179 -18604 8213 -18570
rect 8247 -18604 8281 -18570
rect 8315 -18604 8349 -18570
rect 8383 -18604 8417 -18570
rect 8451 -18587 8676 -18570
rect 8734 -18570 9694 -18532
rect 8734 -18587 8959 -18570
rect 8451 -18604 8490 -18587
rect 7902 -18620 8490 -18604
rect 8920 -18604 8959 -18587
rect 8993 -18604 9027 -18570
rect 9061 -18604 9095 -18570
rect 9129 -18604 9163 -18570
rect 9197 -18604 9231 -18570
rect 9265 -18604 9299 -18570
rect 9333 -18604 9367 -18570
rect 9401 -18604 9435 -18570
rect 9469 -18587 9694 -18570
rect 9752 -18570 10712 -18532
rect 9752 -18587 9977 -18570
rect 9469 -18604 9508 -18587
rect 8920 -18620 9508 -18604
rect 9938 -18604 9977 -18587
rect 10011 -18604 10045 -18570
rect 10079 -18604 10113 -18570
rect 10147 -18604 10181 -18570
rect 10215 -18604 10249 -18570
rect 10283 -18604 10317 -18570
rect 10351 -18604 10385 -18570
rect 10419 -18604 10453 -18570
rect 10487 -18587 10712 -18570
rect 10770 -18570 11730 -18532
rect 10770 -18587 10995 -18570
rect 10487 -18604 10526 -18587
rect 9938 -18620 10526 -18604
rect 10956 -18604 10995 -18587
rect 11029 -18604 11063 -18570
rect 11097 -18604 11131 -18570
rect 11165 -18604 11199 -18570
rect 11233 -18604 11267 -18570
rect 11301 -18604 11335 -18570
rect 11369 -18604 11403 -18570
rect 11437 -18604 11471 -18570
rect 11505 -18587 11730 -18570
rect 11788 -18570 12748 -18532
rect 11788 -18587 12013 -18570
rect 11505 -18604 11544 -18587
rect 10956 -18620 11544 -18604
rect 11974 -18604 12013 -18587
rect 12047 -18604 12081 -18570
rect 12115 -18604 12149 -18570
rect 12183 -18604 12217 -18570
rect 12251 -18604 12285 -18570
rect 12319 -18604 12353 -18570
rect 12387 -18604 12421 -18570
rect 12455 -18604 12489 -18570
rect 12523 -18587 12748 -18570
rect 12806 -18570 13766 -18532
rect 12806 -18587 13031 -18570
rect 12523 -18604 12562 -18587
rect 11974 -18620 12562 -18604
rect 12992 -18604 13031 -18587
rect 13065 -18604 13099 -18570
rect 13133 -18604 13167 -18570
rect 13201 -18604 13235 -18570
rect 13269 -18604 13303 -18570
rect 13337 -18604 13371 -18570
rect 13405 -18604 13439 -18570
rect 13473 -18604 13507 -18570
rect 13541 -18587 13766 -18570
rect 13824 -18570 14784 -18532
rect 13824 -18587 14049 -18570
rect 13541 -18604 13580 -18587
rect 12992 -18620 13580 -18604
rect 14010 -18604 14049 -18587
rect 14083 -18604 14117 -18570
rect 14151 -18604 14185 -18570
rect 14219 -18604 14253 -18570
rect 14287 -18604 14321 -18570
rect 14355 -18604 14389 -18570
rect 14423 -18604 14457 -18570
rect 14491 -18604 14525 -18570
rect 14559 -18587 14784 -18570
rect 14842 -18570 15802 -18532
rect 14842 -18587 15067 -18570
rect 14559 -18604 14598 -18587
rect 14010 -18620 14598 -18604
rect 15028 -18604 15067 -18587
rect 15101 -18604 15135 -18570
rect 15169 -18604 15203 -18570
rect 15237 -18604 15271 -18570
rect 15305 -18604 15339 -18570
rect 15373 -18604 15407 -18570
rect 15441 -18604 15475 -18570
rect 15509 -18604 15543 -18570
rect 15577 -18587 15802 -18570
rect 15860 -18570 16820 -18532
rect 15860 -18587 16085 -18570
rect 15577 -18604 15616 -18587
rect 15028 -18620 15616 -18604
rect 16046 -18604 16085 -18587
rect 16119 -18604 16153 -18570
rect 16187 -18604 16221 -18570
rect 16255 -18604 16289 -18570
rect 16323 -18604 16357 -18570
rect 16391 -18604 16425 -18570
rect 16459 -18604 16493 -18570
rect 16527 -18604 16561 -18570
rect 16595 -18587 16820 -18570
rect 16878 -18570 17838 -18532
rect 16878 -18587 17103 -18570
rect 16595 -18604 16634 -18587
rect 16046 -18620 16634 -18604
rect 17064 -18604 17103 -18587
rect 17137 -18604 17171 -18570
rect 17205 -18604 17239 -18570
rect 17273 -18604 17307 -18570
rect 17341 -18604 17375 -18570
rect 17409 -18604 17443 -18570
rect 17477 -18604 17511 -18570
rect 17545 -18604 17579 -18570
rect 17613 -18587 17838 -18570
rect 17896 -18570 18856 -18532
rect 17896 -18587 18121 -18570
rect 17613 -18604 17652 -18587
rect 17064 -18620 17652 -18604
rect 18082 -18604 18121 -18587
rect 18155 -18604 18189 -18570
rect 18223 -18604 18257 -18570
rect 18291 -18604 18325 -18570
rect 18359 -18604 18393 -18570
rect 18427 -18604 18461 -18570
rect 18495 -18604 18529 -18570
rect 18563 -18604 18597 -18570
rect 18631 -18587 18856 -18570
rect 18914 -18570 19874 -18532
rect 18914 -18587 19139 -18570
rect 18631 -18604 18670 -18587
rect 18082 -18620 18670 -18604
rect 19100 -18604 19139 -18587
rect 19173 -18604 19207 -18570
rect 19241 -18604 19275 -18570
rect 19309 -18604 19343 -18570
rect 19377 -18604 19411 -18570
rect 19445 -18604 19479 -18570
rect 19513 -18604 19547 -18570
rect 19581 -18604 19615 -18570
rect 19649 -18587 19874 -18570
rect 19932 -18570 20892 -18532
rect 19932 -18587 20157 -18570
rect 19649 -18604 19688 -18587
rect 19100 -18620 19688 -18604
rect 20118 -18604 20157 -18587
rect 20191 -18604 20225 -18570
rect 20259 -18604 20293 -18570
rect 20327 -18604 20361 -18570
rect 20395 -18604 20429 -18570
rect 20463 -18604 20497 -18570
rect 20531 -18604 20565 -18570
rect 20599 -18604 20633 -18570
rect 20667 -18587 20892 -18570
rect 20950 -18570 21910 -18532
rect 20950 -18587 21175 -18570
rect 20667 -18604 20706 -18587
rect 20118 -18620 20706 -18604
rect 21136 -18604 21175 -18587
rect 21209 -18604 21243 -18570
rect 21277 -18604 21311 -18570
rect 21345 -18604 21379 -18570
rect 21413 -18604 21447 -18570
rect 21481 -18604 21515 -18570
rect 21549 -18604 21583 -18570
rect 21617 -18604 21651 -18570
rect 21685 -18587 21910 -18570
rect 21968 -18570 22928 -18532
rect 21968 -18587 22193 -18570
rect 21685 -18604 21724 -18587
rect 21136 -18620 21724 -18604
rect 22154 -18604 22193 -18587
rect 22227 -18604 22261 -18570
rect 22295 -18604 22329 -18570
rect 22363 -18604 22397 -18570
rect 22431 -18604 22465 -18570
rect 22499 -18604 22533 -18570
rect 22567 -18604 22601 -18570
rect 22635 -18604 22669 -18570
rect 22703 -18587 22928 -18570
rect 22703 -18604 22742 -18587
rect 22154 -18620 22742 -18604
rect -9138 -18876 -8178 -18838
rect -9138 -18893 -8913 -18876
rect -8952 -18910 -8913 -18893
rect -8879 -18910 -8845 -18876
rect -8811 -18910 -8777 -18876
rect -8743 -18910 -8709 -18876
rect -8675 -18910 -8641 -18876
rect -8607 -18910 -8573 -18876
rect -8539 -18910 -8505 -18876
rect -8471 -18910 -8437 -18876
rect -8403 -18893 -8178 -18876
rect -8120 -18876 -7160 -18838
rect -8120 -18893 -7895 -18876
rect -8403 -18910 -8364 -18893
rect -8952 -18926 -8364 -18910
rect -7934 -18910 -7895 -18893
rect -7861 -18910 -7827 -18876
rect -7793 -18910 -7759 -18876
rect -7725 -18910 -7691 -18876
rect -7657 -18910 -7623 -18876
rect -7589 -18910 -7555 -18876
rect -7521 -18910 -7487 -18876
rect -7453 -18910 -7419 -18876
rect -7385 -18893 -7160 -18876
rect -7102 -18876 -6142 -18838
rect -7102 -18893 -6877 -18876
rect -7385 -18910 -7346 -18893
rect -7934 -18926 -7346 -18910
rect -6916 -18910 -6877 -18893
rect -6843 -18910 -6809 -18876
rect -6775 -18910 -6741 -18876
rect -6707 -18910 -6673 -18876
rect -6639 -18910 -6605 -18876
rect -6571 -18910 -6537 -18876
rect -6503 -18910 -6469 -18876
rect -6435 -18910 -6401 -18876
rect -6367 -18893 -6142 -18876
rect -6084 -18876 -5124 -18838
rect -6084 -18893 -5859 -18876
rect -6367 -18910 -6328 -18893
rect -6916 -18926 -6328 -18910
rect -5898 -18910 -5859 -18893
rect -5825 -18910 -5791 -18876
rect -5757 -18910 -5723 -18876
rect -5689 -18910 -5655 -18876
rect -5621 -18910 -5587 -18876
rect -5553 -18910 -5519 -18876
rect -5485 -18910 -5451 -18876
rect -5417 -18910 -5383 -18876
rect -5349 -18893 -5124 -18876
rect -5066 -18876 -4106 -18838
rect -5066 -18893 -4841 -18876
rect -5349 -18910 -5310 -18893
rect -5898 -18926 -5310 -18910
rect -4880 -18910 -4841 -18893
rect -4807 -18910 -4773 -18876
rect -4739 -18910 -4705 -18876
rect -4671 -18910 -4637 -18876
rect -4603 -18910 -4569 -18876
rect -4535 -18910 -4501 -18876
rect -4467 -18910 -4433 -18876
rect -4399 -18910 -4365 -18876
rect -4331 -18893 -4106 -18876
rect -4048 -18876 -3088 -18838
rect -4048 -18893 -3823 -18876
rect -4331 -18910 -4292 -18893
rect -4880 -18926 -4292 -18910
rect -3862 -18910 -3823 -18893
rect -3789 -18910 -3755 -18876
rect -3721 -18910 -3687 -18876
rect -3653 -18910 -3619 -18876
rect -3585 -18910 -3551 -18876
rect -3517 -18910 -3483 -18876
rect -3449 -18910 -3415 -18876
rect -3381 -18910 -3347 -18876
rect -3313 -18893 -3088 -18876
rect -3030 -18876 -2070 -18838
rect -3030 -18893 -2805 -18876
rect -3313 -18910 -3274 -18893
rect -3862 -18926 -3274 -18910
rect -2844 -18910 -2805 -18893
rect -2771 -18910 -2737 -18876
rect -2703 -18910 -2669 -18876
rect -2635 -18910 -2601 -18876
rect -2567 -18910 -2533 -18876
rect -2499 -18910 -2465 -18876
rect -2431 -18910 -2397 -18876
rect -2363 -18910 -2329 -18876
rect -2295 -18893 -2070 -18876
rect -2012 -18876 -1052 -18838
rect -2012 -18893 -1787 -18876
rect -2295 -18910 -2256 -18893
rect -2844 -18926 -2256 -18910
rect -1826 -18910 -1787 -18893
rect -1753 -18910 -1719 -18876
rect -1685 -18910 -1651 -18876
rect -1617 -18910 -1583 -18876
rect -1549 -18910 -1515 -18876
rect -1481 -18910 -1447 -18876
rect -1413 -18910 -1379 -18876
rect -1345 -18910 -1311 -18876
rect -1277 -18893 -1052 -18876
rect -994 -18876 -34 -18838
rect -994 -18893 -769 -18876
rect -1277 -18910 -1238 -18893
rect -1826 -18926 -1238 -18910
rect -808 -18910 -769 -18893
rect -735 -18910 -701 -18876
rect -667 -18910 -633 -18876
rect -599 -18910 -565 -18876
rect -531 -18910 -497 -18876
rect -463 -18910 -429 -18876
rect -395 -18910 -361 -18876
rect -327 -18910 -293 -18876
rect -259 -18893 -34 -18876
rect -259 -18910 -220 -18893
rect -808 -18926 -220 -18910
rect 2812 -19092 3400 -19076
rect 2812 -19109 2851 -19092
rect 2626 -19126 2851 -19109
rect 2885 -19126 2919 -19092
rect 2953 -19126 2987 -19092
rect 3021 -19126 3055 -19092
rect 3089 -19126 3123 -19092
rect 3157 -19126 3191 -19092
rect 3225 -19126 3259 -19092
rect 3293 -19126 3327 -19092
rect 3361 -19109 3400 -19092
rect 3830 -19092 4418 -19076
rect 3830 -19109 3869 -19092
rect 3361 -19126 3586 -19109
rect 2626 -19164 3586 -19126
rect 3644 -19126 3869 -19109
rect 3903 -19126 3937 -19092
rect 3971 -19126 4005 -19092
rect 4039 -19126 4073 -19092
rect 4107 -19126 4141 -19092
rect 4175 -19126 4209 -19092
rect 4243 -19126 4277 -19092
rect 4311 -19126 4345 -19092
rect 4379 -19109 4418 -19092
rect 4848 -19092 5436 -19076
rect 4848 -19109 4887 -19092
rect 4379 -19126 4604 -19109
rect 3644 -19164 4604 -19126
rect 4662 -19126 4887 -19109
rect 4921 -19126 4955 -19092
rect 4989 -19126 5023 -19092
rect 5057 -19126 5091 -19092
rect 5125 -19126 5159 -19092
rect 5193 -19126 5227 -19092
rect 5261 -19126 5295 -19092
rect 5329 -19126 5363 -19092
rect 5397 -19109 5436 -19092
rect 5866 -19092 6454 -19076
rect 5866 -19109 5905 -19092
rect 5397 -19126 5622 -19109
rect 4662 -19164 5622 -19126
rect 5680 -19126 5905 -19109
rect 5939 -19126 5973 -19092
rect 6007 -19126 6041 -19092
rect 6075 -19126 6109 -19092
rect 6143 -19126 6177 -19092
rect 6211 -19126 6245 -19092
rect 6279 -19126 6313 -19092
rect 6347 -19126 6381 -19092
rect 6415 -19109 6454 -19092
rect 6884 -19092 7472 -19076
rect 6884 -19109 6923 -19092
rect 6415 -19126 6640 -19109
rect 5680 -19164 6640 -19126
rect 6698 -19126 6923 -19109
rect 6957 -19126 6991 -19092
rect 7025 -19126 7059 -19092
rect 7093 -19126 7127 -19092
rect 7161 -19126 7195 -19092
rect 7229 -19126 7263 -19092
rect 7297 -19126 7331 -19092
rect 7365 -19126 7399 -19092
rect 7433 -19109 7472 -19092
rect 7902 -19092 8490 -19076
rect 7902 -19109 7941 -19092
rect 7433 -19126 7658 -19109
rect 6698 -19164 7658 -19126
rect 7716 -19126 7941 -19109
rect 7975 -19126 8009 -19092
rect 8043 -19126 8077 -19092
rect 8111 -19126 8145 -19092
rect 8179 -19126 8213 -19092
rect 8247 -19126 8281 -19092
rect 8315 -19126 8349 -19092
rect 8383 -19126 8417 -19092
rect 8451 -19109 8490 -19092
rect 8920 -19092 9508 -19076
rect 8920 -19109 8959 -19092
rect 8451 -19126 8676 -19109
rect 7716 -19164 8676 -19126
rect 8734 -19126 8959 -19109
rect 8993 -19126 9027 -19092
rect 9061 -19126 9095 -19092
rect 9129 -19126 9163 -19092
rect 9197 -19126 9231 -19092
rect 9265 -19126 9299 -19092
rect 9333 -19126 9367 -19092
rect 9401 -19126 9435 -19092
rect 9469 -19109 9508 -19092
rect 9938 -19092 10526 -19076
rect 9938 -19109 9977 -19092
rect 9469 -19126 9694 -19109
rect 8734 -19164 9694 -19126
rect 9752 -19126 9977 -19109
rect 10011 -19126 10045 -19092
rect 10079 -19126 10113 -19092
rect 10147 -19126 10181 -19092
rect 10215 -19126 10249 -19092
rect 10283 -19126 10317 -19092
rect 10351 -19126 10385 -19092
rect 10419 -19126 10453 -19092
rect 10487 -19109 10526 -19092
rect 10956 -19092 11544 -19076
rect 10956 -19109 10995 -19092
rect 10487 -19126 10712 -19109
rect 9752 -19164 10712 -19126
rect 10770 -19126 10995 -19109
rect 11029 -19126 11063 -19092
rect 11097 -19126 11131 -19092
rect 11165 -19126 11199 -19092
rect 11233 -19126 11267 -19092
rect 11301 -19126 11335 -19092
rect 11369 -19126 11403 -19092
rect 11437 -19126 11471 -19092
rect 11505 -19109 11544 -19092
rect 11974 -19092 12562 -19076
rect 11974 -19109 12013 -19092
rect 11505 -19126 11730 -19109
rect 10770 -19164 11730 -19126
rect 11788 -19126 12013 -19109
rect 12047 -19126 12081 -19092
rect 12115 -19126 12149 -19092
rect 12183 -19126 12217 -19092
rect 12251 -19126 12285 -19092
rect 12319 -19126 12353 -19092
rect 12387 -19126 12421 -19092
rect 12455 -19126 12489 -19092
rect 12523 -19109 12562 -19092
rect 12992 -19092 13580 -19076
rect 12992 -19109 13031 -19092
rect 12523 -19126 12748 -19109
rect 11788 -19164 12748 -19126
rect 12806 -19126 13031 -19109
rect 13065 -19126 13099 -19092
rect 13133 -19126 13167 -19092
rect 13201 -19126 13235 -19092
rect 13269 -19126 13303 -19092
rect 13337 -19126 13371 -19092
rect 13405 -19126 13439 -19092
rect 13473 -19126 13507 -19092
rect 13541 -19109 13580 -19092
rect 14010 -19092 14598 -19076
rect 14010 -19109 14049 -19092
rect 13541 -19126 13766 -19109
rect 12806 -19164 13766 -19126
rect 13824 -19126 14049 -19109
rect 14083 -19126 14117 -19092
rect 14151 -19126 14185 -19092
rect 14219 -19126 14253 -19092
rect 14287 -19126 14321 -19092
rect 14355 -19126 14389 -19092
rect 14423 -19126 14457 -19092
rect 14491 -19126 14525 -19092
rect 14559 -19109 14598 -19092
rect 15028 -19092 15616 -19076
rect 15028 -19109 15067 -19092
rect 14559 -19126 14784 -19109
rect 13824 -19164 14784 -19126
rect 14842 -19126 15067 -19109
rect 15101 -19126 15135 -19092
rect 15169 -19126 15203 -19092
rect 15237 -19126 15271 -19092
rect 15305 -19126 15339 -19092
rect 15373 -19126 15407 -19092
rect 15441 -19126 15475 -19092
rect 15509 -19126 15543 -19092
rect 15577 -19109 15616 -19092
rect 16046 -19092 16634 -19076
rect 16046 -19109 16085 -19092
rect 15577 -19126 15802 -19109
rect 14842 -19164 15802 -19126
rect 15860 -19126 16085 -19109
rect 16119 -19126 16153 -19092
rect 16187 -19126 16221 -19092
rect 16255 -19126 16289 -19092
rect 16323 -19126 16357 -19092
rect 16391 -19126 16425 -19092
rect 16459 -19126 16493 -19092
rect 16527 -19126 16561 -19092
rect 16595 -19109 16634 -19092
rect 17064 -19092 17652 -19076
rect 17064 -19109 17103 -19092
rect 16595 -19126 16820 -19109
rect 15860 -19164 16820 -19126
rect 16878 -19126 17103 -19109
rect 17137 -19126 17171 -19092
rect 17205 -19126 17239 -19092
rect 17273 -19126 17307 -19092
rect 17341 -19126 17375 -19092
rect 17409 -19126 17443 -19092
rect 17477 -19126 17511 -19092
rect 17545 -19126 17579 -19092
rect 17613 -19109 17652 -19092
rect 18082 -19092 18670 -19076
rect 18082 -19109 18121 -19092
rect 17613 -19126 17838 -19109
rect 16878 -19164 17838 -19126
rect 17896 -19126 18121 -19109
rect 18155 -19126 18189 -19092
rect 18223 -19126 18257 -19092
rect 18291 -19126 18325 -19092
rect 18359 -19126 18393 -19092
rect 18427 -19126 18461 -19092
rect 18495 -19126 18529 -19092
rect 18563 -19126 18597 -19092
rect 18631 -19109 18670 -19092
rect 19100 -19092 19688 -19076
rect 19100 -19109 19139 -19092
rect 18631 -19126 18856 -19109
rect 17896 -19164 18856 -19126
rect 18914 -19126 19139 -19109
rect 19173 -19126 19207 -19092
rect 19241 -19126 19275 -19092
rect 19309 -19126 19343 -19092
rect 19377 -19126 19411 -19092
rect 19445 -19126 19479 -19092
rect 19513 -19126 19547 -19092
rect 19581 -19126 19615 -19092
rect 19649 -19109 19688 -19092
rect 20118 -19092 20706 -19076
rect 20118 -19109 20157 -19092
rect 19649 -19126 19874 -19109
rect 18914 -19164 19874 -19126
rect 19932 -19126 20157 -19109
rect 20191 -19126 20225 -19092
rect 20259 -19126 20293 -19092
rect 20327 -19126 20361 -19092
rect 20395 -19126 20429 -19092
rect 20463 -19126 20497 -19092
rect 20531 -19126 20565 -19092
rect 20599 -19126 20633 -19092
rect 20667 -19109 20706 -19092
rect 21136 -19092 21724 -19076
rect 21136 -19109 21175 -19092
rect 20667 -19126 20892 -19109
rect 19932 -19164 20892 -19126
rect 20950 -19126 21175 -19109
rect 21209 -19126 21243 -19092
rect 21277 -19126 21311 -19092
rect 21345 -19126 21379 -19092
rect 21413 -19126 21447 -19092
rect 21481 -19126 21515 -19092
rect 21549 -19126 21583 -19092
rect 21617 -19126 21651 -19092
rect 21685 -19109 21724 -19092
rect 22154 -19092 22742 -19076
rect 22154 -19109 22193 -19092
rect 21685 -19126 21910 -19109
rect 20950 -19164 21910 -19126
rect 21968 -19126 22193 -19109
rect 22227 -19126 22261 -19092
rect 22295 -19126 22329 -19092
rect 22363 -19126 22397 -19092
rect 22431 -19126 22465 -19092
rect 22499 -19126 22533 -19092
rect 22567 -19126 22601 -19092
rect 22635 -19126 22669 -19092
rect 22703 -19109 22742 -19092
rect 22703 -19126 22928 -19109
rect 21968 -19164 22928 -19126
rect 2626 -19802 3586 -19764
rect 2626 -19819 2851 -19802
rect 2812 -19836 2851 -19819
rect 2885 -19836 2919 -19802
rect 2953 -19836 2987 -19802
rect 3021 -19836 3055 -19802
rect 3089 -19836 3123 -19802
rect 3157 -19836 3191 -19802
rect 3225 -19836 3259 -19802
rect 3293 -19836 3327 -19802
rect 3361 -19819 3586 -19802
rect 3644 -19802 4604 -19764
rect 3644 -19819 3869 -19802
rect 3361 -19836 3400 -19819
rect 2812 -19852 3400 -19836
rect 3830 -19836 3869 -19819
rect 3903 -19836 3937 -19802
rect 3971 -19836 4005 -19802
rect 4039 -19836 4073 -19802
rect 4107 -19836 4141 -19802
rect 4175 -19836 4209 -19802
rect 4243 -19836 4277 -19802
rect 4311 -19836 4345 -19802
rect 4379 -19819 4604 -19802
rect 4662 -19802 5622 -19764
rect 4662 -19819 4887 -19802
rect 4379 -19836 4418 -19819
rect 3830 -19852 4418 -19836
rect 4848 -19836 4887 -19819
rect 4921 -19836 4955 -19802
rect 4989 -19836 5023 -19802
rect 5057 -19836 5091 -19802
rect 5125 -19836 5159 -19802
rect 5193 -19836 5227 -19802
rect 5261 -19836 5295 -19802
rect 5329 -19836 5363 -19802
rect 5397 -19819 5622 -19802
rect 5680 -19802 6640 -19764
rect 5680 -19819 5905 -19802
rect 5397 -19836 5436 -19819
rect 4848 -19852 5436 -19836
rect 5866 -19836 5905 -19819
rect 5939 -19836 5973 -19802
rect 6007 -19836 6041 -19802
rect 6075 -19836 6109 -19802
rect 6143 -19836 6177 -19802
rect 6211 -19836 6245 -19802
rect 6279 -19836 6313 -19802
rect 6347 -19836 6381 -19802
rect 6415 -19819 6640 -19802
rect 6698 -19802 7658 -19764
rect 6698 -19819 6923 -19802
rect 6415 -19836 6454 -19819
rect 5866 -19852 6454 -19836
rect 6884 -19836 6923 -19819
rect 6957 -19836 6991 -19802
rect 7025 -19836 7059 -19802
rect 7093 -19836 7127 -19802
rect 7161 -19836 7195 -19802
rect 7229 -19836 7263 -19802
rect 7297 -19836 7331 -19802
rect 7365 -19836 7399 -19802
rect 7433 -19819 7658 -19802
rect 7716 -19802 8676 -19764
rect 7716 -19819 7941 -19802
rect 7433 -19836 7472 -19819
rect 6884 -19852 7472 -19836
rect 7902 -19836 7941 -19819
rect 7975 -19836 8009 -19802
rect 8043 -19836 8077 -19802
rect 8111 -19836 8145 -19802
rect 8179 -19836 8213 -19802
rect 8247 -19836 8281 -19802
rect 8315 -19836 8349 -19802
rect 8383 -19836 8417 -19802
rect 8451 -19819 8676 -19802
rect 8734 -19802 9694 -19764
rect 8734 -19819 8959 -19802
rect 8451 -19836 8490 -19819
rect 7902 -19852 8490 -19836
rect 8920 -19836 8959 -19819
rect 8993 -19836 9027 -19802
rect 9061 -19836 9095 -19802
rect 9129 -19836 9163 -19802
rect 9197 -19836 9231 -19802
rect 9265 -19836 9299 -19802
rect 9333 -19836 9367 -19802
rect 9401 -19836 9435 -19802
rect 9469 -19819 9694 -19802
rect 9752 -19802 10712 -19764
rect 9752 -19819 9977 -19802
rect 9469 -19836 9508 -19819
rect 8920 -19852 9508 -19836
rect 9938 -19836 9977 -19819
rect 10011 -19836 10045 -19802
rect 10079 -19836 10113 -19802
rect 10147 -19836 10181 -19802
rect 10215 -19836 10249 -19802
rect 10283 -19836 10317 -19802
rect 10351 -19836 10385 -19802
rect 10419 -19836 10453 -19802
rect 10487 -19819 10712 -19802
rect 10770 -19802 11730 -19764
rect 10770 -19819 10995 -19802
rect 10487 -19836 10526 -19819
rect 9938 -19852 10526 -19836
rect 10956 -19836 10995 -19819
rect 11029 -19836 11063 -19802
rect 11097 -19836 11131 -19802
rect 11165 -19836 11199 -19802
rect 11233 -19836 11267 -19802
rect 11301 -19836 11335 -19802
rect 11369 -19836 11403 -19802
rect 11437 -19836 11471 -19802
rect 11505 -19819 11730 -19802
rect 11788 -19802 12748 -19764
rect 11788 -19819 12013 -19802
rect 11505 -19836 11544 -19819
rect 10956 -19852 11544 -19836
rect 11974 -19836 12013 -19819
rect 12047 -19836 12081 -19802
rect 12115 -19836 12149 -19802
rect 12183 -19836 12217 -19802
rect 12251 -19836 12285 -19802
rect 12319 -19836 12353 -19802
rect 12387 -19836 12421 -19802
rect 12455 -19836 12489 -19802
rect 12523 -19819 12748 -19802
rect 12806 -19802 13766 -19764
rect 12806 -19819 13031 -19802
rect 12523 -19836 12562 -19819
rect 11974 -19852 12562 -19836
rect 12992 -19836 13031 -19819
rect 13065 -19836 13099 -19802
rect 13133 -19836 13167 -19802
rect 13201 -19836 13235 -19802
rect 13269 -19836 13303 -19802
rect 13337 -19836 13371 -19802
rect 13405 -19836 13439 -19802
rect 13473 -19836 13507 -19802
rect 13541 -19819 13766 -19802
rect 13824 -19802 14784 -19764
rect 13824 -19819 14049 -19802
rect 13541 -19836 13580 -19819
rect 12992 -19852 13580 -19836
rect 14010 -19836 14049 -19819
rect 14083 -19836 14117 -19802
rect 14151 -19836 14185 -19802
rect 14219 -19836 14253 -19802
rect 14287 -19836 14321 -19802
rect 14355 -19836 14389 -19802
rect 14423 -19836 14457 -19802
rect 14491 -19836 14525 -19802
rect 14559 -19819 14784 -19802
rect 14842 -19802 15802 -19764
rect 14842 -19819 15067 -19802
rect 14559 -19836 14598 -19819
rect 14010 -19852 14598 -19836
rect 15028 -19836 15067 -19819
rect 15101 -19836 15135 -19802
rect 15169 -19836 15203 -19802
rect 15237 -19836 15271 -19802
rect 15305 -19836 15339 -19802
rect 15373 -19836 15407 -19802
rect 15441 -19836 15475 -19802
rect 15509 -19836 15543 -19802
rect 15577 -19819 15802 -19802
rect 15860 -19802 16820 -19764
rect 15860 -19819 16085 -19802
rect 15577 -19836 15616 -19819
rect 15028 -19852 15616 -19836
rect 16046 -19836 16085 -19819
rect 16119 -19836 16153 -19802
rect 16187 -19836 16221 -19802
rect 16255 -19836 16289 -19802
rect 16323 -19836 16357 -19802
rect 16391 -19836 16425 -19802
rect 16459 -19836 16493 -19802
rect 16527 -19836 16561 -19802
rect 16595 -19819 16820 -19802
rect 16878 -19802 17838 -19764
rect 16878 -19819 17103 -19802
rect 16595 -19836 16634 -19819
rect 16046 -19852 16634 -19836
rect 17064 -19836 17103 -19819
rect 17137 -19836 17171 -19802
rect 17205 -19836 17239 -19802
rect 17273 -19836 17307 -19802
rect 17341 -19836 17375 -19802
rect 17409 -19836 17443 -19802
rect 17477 -19836 17511 -19802
rect 17545 -19836 17579 -19802
rect 17613 -19819 17838 -19802
rect 17896 -19802 18856 -19764
rect 17896 -19819 18121 -19802
rect 17613 -19836 17652 -19819
rect 17064 -19852 17652 -19836
rect 18082 -19836 18121 -19819
rect 18155 -19836 18189 -19802
rect 18223 -19836 18257 -19802
rect 18291 -19836 18325 -19802
rect 18359 -19836 18393 -19802
rect 18427 -19836 18461 -19802
rect 18495 -19836 18529 -19802
rect 18563 -19836 18597 -19802
rect 18631 -19819 18856 -19802
rect 18914 -19802 19874 -19764
rect 18914 -19819 19139 -19802
rect 18631 -19836 18670 -19819
rect 18082 -19852 18670 -19836
rect 19100 -19836 19139 -19819
rect 19173 -19836 19207 -19802
rect 19241 -19836 19275 -19802
rect 19309 -19836 19343 -19802
rect 19377 -19836 19411 -19802
rect 19445 -19836 19479 -19802
rect 19513 -19836 19547 -19802
rect 19581 -19836 19615 -19802
rect 19649 -19819 19874 -19802
rect 19932 -19802 20892 -19764
rect 19932 -19819 20157 -19802
rect 19649 -19836 19688 -19819
rect 19100 -19852 19688 -19836
rect 20118 -19836 20157 -19819
rect 20191 -19836 20225 -19802
rect 20259 -19836 20293 -19802
rect 20327 -19836 20361 -19802
rect 20395 -19836 20429 -19802
rect 20463 -19836 20497 -19802
rect 20531 -19836 20565 -19802
rect 20599 -19836 20633 -19802
rect 20667 -19819 20892 -19802
rect 20950 -19802 21910 -19764
rect 20950 -19819 21175 -19802
rect 20667 -19836 20706 -19819
rect 20118 -19852 20706 -19836
rect 21136 -19836 21175 -19819
rect 21209 -19836 21243 -19802
rect 21277 -19836 21311 -19802
rect 21345 -19836 21379 -19802
rect 21413 -19836 21447 -19802
rect 21481 -19836 21515 -19802
rect 21549 -19836 21583 -19802
rect 21617 -19836 21651 -19802
rect 21685 -19819 21910 -19802
rect 21968 -19802 22928 -19764
rect 21968 -19819 22193 -19802
rect 21685 -19836 21724 -19819
rect 21136 -19852 21724 -19836
rect 22154 -19836 22193 -19819
rect 22227 -19836 22261 -19802
rect 22295 -19836 22329 -19802
rect 22363 -19836 22397 -19802
rect 22431 -19836 22465 -19802
rect 22499 -19836 22533 -19802
rect 22567 -19836 22601 -19802
rect 22635 -19836 22669 -19802
rect 22703 -19819 22928 -19802
rect 22703 -19836 22742 -19819
rect 22154 -19852 22742 -19836
rect 2812 -20326 3400 -20310
rect 2812 -20343 2851 -20326
rect 2626 -20360 2851 -20343
rect 2885 -20360 2919 -20326
rect 2953 -20360 2987 -20326
rect 3021 -20360 3055 -20326
rect 3089 -20360 3123 -20326
rect 3157 -20360 3191 -20326
rect 3225 -20360 3259 -20326
rect 3293 -20360 3327 -20326
rect 3361 -20343 3400 -20326
rect 3830 -20326 4418 -20310
rect 3830 -20343 3869 -20326
rect 3361 -20360 3586 -20343
rect 2626 -20398 3586 -20360
rect 3644 -20360 3869 -20343
rect 3903 -20360 3937 -20326
rect 3971 -20360 4005 -20326
rect 4039 -20360 4073 -20326
rect 4107 -20360 4141 -20326
rect 4175 -20360 4209 -20326
rect 4243 -20360 4277 -20326
rect 4311 -20360 4345 -20326
rect 4379 -20343 4418 -20326
rect 4848 -20326 5436 -20310
rect 4848 -20343 4887 -20326
rect 4379 -20360 4604 -20343
rect 3644 -20398 4604 -20360
rect 4662 -20360 4887 -20343
rect 4921 -20360 4955 -20326
rect 4989 -20360 5023 -20326
rect 5057 -20360 5091 -20326
rect 5125 -20360 5159 -20326
rect 5193 -20360 5227 -20326
rect 5261 -20360 5295 -20326
rect 5329 -20360 5363 -20326
rect 5397 -20343 5436 -20326
rect 5866 -20326 6454 -20310
rect 5866 -20343 5905 -20326
rect 5397 -20360 5622 -20343
rect 4662 -20398 5622 -20360
rect 5680 -20360 5905 -20343
rect 5939 -20360 5973 -20326
rect 6007 -20360 6041 -20326
rect 6075 -20360 6109 -20326
rect 6143 -20360 6177 -20326
rect 6211 -20360 6245 -20326
rect 6279 -20360 6313 -20326
rect 6347 -20360 6381 -20326
rect 6415 -20343 6454 -20326
rect 6884 -20326 7472 -20310
rect 6884 -20343 6923 -20326
rect 6415 -20360 6640 -20343
rect 5680 -20398 6640 -20360
rect 6698 -20360 6923 -20343
rect 6957 -20360 6991 -20326
rect 7025 -20360 7059 -20326
rect 7093 -20360 7127 -20326
rect 7161 -20360 7195 -20326
rect 7229 -20360 7263 -20326
rect 7297 -20360 7331 -20326
rect 7365 -20360 7399 -20326
rect 7433 -20343 7472 -20326
rect 7902 -20326 8490 -20310
rect 7902 -20343 7941 -20326
rect 7433 -20360 7658 -20343
rect 6698 -20398 7658 -20360
rect 7716 -20360 7941 -20343
rect 7975 -20360 8009 -20326
rect 8043 -20360 8077 -20326
rect 8111 -20360 8145 -20326
rect 8179 -20360 8213 -20326
rect 8247 -20360 8281 -20326
rect 8315 -20360 8349 -20326
rect 8383 -20360 8417 -20326
rect 8451 -20343 8490 -20326
rect 8920 -20326 9508 -20310
rect 8920 -20343 8959 -20326
rect 8451 -20360 8676 -20343
rect 7716 -20398 8676 -20360
rect 8734 -20360 8959 -20343
rect 8993 -20360 9027 -20326
rect 9061 -20360 9095 -20326
rect 9129 -20360 9163 -20326
rect 9197 -20360 9231 -20326
rect 9265 -20360 9299 -20326
rect 9333 -20360 9367 -20326
rect 9401 -20360 9435 -20326
rect 9469 -20343 9508 -20326
rect 9938 -20326 10526 -20310
rect 9938 -20343 9977 -20326
rect 9469 -20360 9694 -20343
rect 8734 -20398 9694 -20360
rect 9752 -20360 9977 -20343
rect 10011 -20360 10045 -20326
rect 10079 -20360 10113 -20326
rect 10147 -20360 10181 -20326
rect 10215 -20360 10249 -20326
rect 10283 -20360 10317 -20326
rect 10351 -20360 10385 -20326
rect 10419 -20360 10453 -20326
rect 10487 -20343 10526 -20326
rect 10956 -20326 11544 -20310
rect 10956 -20343 10995 -20326
rect 10487 -20360 10712 -20343
rect 9752 -20398 10712 -20360
rect 10770 -20360 10995 -20343
rect 11029 -20360 11063 -20326
rect 11097 -20360 11131 -20326
rect 11165 -20360 11199 -20326
rect 11233 -20360 11267 -20326
rect 11301 -20360 11335 -20326
rect 11369 -20360 11403 -20326
rect 11437 -20360 11471 -20326
rect 11505 -20343 11544 -20326
rect 11974 -20326 12562 -20310
rect 11974 -20343 12013 -20326
rect 11505 -20360 11730 -20343
rect 10770 -20398 11730 -20360
rect 11788 -20360 12013 -20343
rect 12047 -20360 12081 -20326
rect 12115 -20360 12149 -20326
rect 12183 -20360 12217 -20326
rect 12251 -20360 12285 -20326
rect 12319 -20360 12353 -20326
rect 12387 -20360 12421 -20326
rect 12455 -20360 12489 -20326
rect 12523 -20343 12562 -20326
rect 12992 -20326 13580 -20310
rect 12992 -20343 13031 -20326
rect 12523 -20360 12748 -20343
rect 11788 -20398 12748 -20360
rect 12806 -20360 13031 -20343
rect 13065 -20360 13099 -20326
rect 13133 -20360 13167 -20326
rect 13201 -20360 13235 -20326
rect 13269 -20360 13303 -20326
rect 13337 -20360 13371 -20326
rect 13405 -20360 13439 -20326
rect 13473 -20360 13507 -20326
rect 13541 -20343 13580 -20326
rect 14010 -20326 14598 -20310
rect 14010 -20343 14049 -20326
rect 13541 -20360 13766 -20343
rect 12806 -20398 13766 -20360
rect 13824 -20360 14049 -20343
rect 14083 -20360 14117 -20326
rect 14151 -20360 14185 -20326
rect 14219 -20360 14253 -20326
rect 14287 -20360 14321 -20326
rect 14355 -20360 14389 -20326
rect 14423 -20360 14457 -20326
rect 14491 -20360 14525 -20326
rect 14559 -20343 14598 -20326
rect 15028 -20326 15616 -20310
rect 15028 -20343 15067 -20326
rect 14559 -20360 14784 -20343
rect 13824 -20398 14784 -20360
rect 14842 -20360 15067 -20343
rect 15101 -20360 15135 -20326
rect 15169 -20360 15203 -20326
rect 15237 -20360 15271 -20326
rect 15305 -20360 15339 -20326
rect 15373 -20360 15407 -20326
rect 15441 -20360 15475 -20326
rect 15509 -20360 15543 -20326
rect 15577 -20343 15616 -20326
rect 16046 -20326 16634 -20310
rect 16046 -20343 16085 -20326
rect 15577 -20360 15802 -20343
rect 14842 -20398 15802 -20360
rect 15860 -20360 16085 -20343
rect 16119 -20360 16153 -20326
rect 16187 -20360 16221 -20326
rect 16255 -20360 16289 -20326
rect 16323 -20360 16357 -20326
rect 16391 -20360 16425 -20326
rect 16459 -20360 16493 -20326
rect 16527 -20360 16561 -20326
rect 16595 -20343 16634 -20326
rect 17064 -20326 17652 -20310
rect 17064 -20343 17103 -20326
rect 16595 -20360 16820 -20343
rect 15860 -20398 16820 -20360
rect 16878 -20360 17103 -20343
rect 17137 -20360 17171 -20326
rect 17205 -20360 17239 -20326
rect 17273 -20360 17307 -20326
rect 17341 -20360 17375 -20326
rect 17409 -20360 17443 -20326
rect 17477 -20360 17511 -20326
rect 17545 -20360 17579 -20326
rect 17613 -20343 17652 -20326
rect 18082 -20326 18670 -20310
rect 18082 -20343 18121 -20326
rect 17613 -20360 17838 -20343
rect 16878 -20398 17838 -20360
rect 17896 -20360 18121 -20343
rect 18155 -20360 18189 -20326
rect 18223 -20360 18257 -20326
rect 18291 -20360 18325 -20326
rect 18359 -20360 18393 -20326
rect 18427 -20360 18461 -20326
rect 18495 -20360 18529 -20326
rect 18563 -20360 18597 -20326
rect 18631 -20343 18670 -20326
rect 19100 -20326 19688 -20310
rect 19100 -20343 19139 -20326
rect 18631 -20360 18856 -20343
rect 17896 -20398 18856 -20360
rect 18914 -20360 19139 -20343
rect 19173 -20360 19207 -20326
rect 19241 -20360 19275 -20326
rect 19309 -20360 19343 -20326
rect 19377 -20360 19411 -20326
rect 19445 -20360 19479 -20326
rect 19513 -20360 19547 -20326
rect 19581 -20360 19615 -20326
rect 19649 -20343 19688 -20326
rect 20118 -20326 20706 -20310
rect 20118 -20343 20157 -20326
rect 19649 -20360 19874 -20343
rect 18914 -20398 19874 -20360
rect 19932 -20360 20157 -20343
rect 20191 -20360 20225 -20326
rect 20259 -20360 20293 -20326
rect 20327 -20360 20361 -20326
rect 20395 -20360 20429 -20326
rect 20463 -20360 20497 -20326
rect 20531 -20360 20565 -20326
rect 20599 -20360 20633 -20326
rect 20667 -20343 20706 -20326
rect 21136 -20326 21724 -20310
rect 21136 -20343 21175 -20326
rect 20667 -20360 20892 -20343
rect 19932 -20398 20892 -20360
rect 20950 -20360 21175 -20343
rect 21209 -20360 21243 -20326
rect 21277 -20360 21311 -20326
rect 21345 -20360 21379 -20326
rect 21413 -20360 21447 -20326
rect 21481 -20360 21515 -20326
rect 21549 -20360 21583 -20326
rect 21617 -20360 21651 -20326
rect 21685 -20343 21724 -20326
rect 22154 -20326 22742 -20310
rect 22154 -20343 22193 -20326
rect 21685 -20360 21910 -20343
rect 20950 -20398 21910 -20360
rect 21968 -20360 22193 -20343
rect 22227 -20360 22261 -20326
rect 22295 -20360 22329 -20326
rect 22363 -20360 22397 -20326
rect 22431 -20360 22465 -20326
rect 22499 -20360 22533 -20326
rect 22567 -20360 22601 -20326
rect 22635 -20360 22669 -20326
rect 22703 -20343 22742 -20326
rect 22703 -20360 22928 -20343
rect 21968 -20398 22928 -20360
rect 2626 -21036 3586 -20998
rect 2626 -21053 2851 -21036
rect 2812 -21070 2851 -21053
rect 2885 -21070 2919 -21036
rect 2953 -21070 2987 -21036
rect 3021 -21070 3055 -21036
rect 3089 -21070 3123 -21036
rect 3157 -21070 3191 -21036
rect 3225 -21070 3259 -21036
rect 3293 -21070 3327 -21036
rect 3361 -21053 3586 -21036
rect 3644 -21036 4604 -20998
rect 3644 -21053 3869 -21036
rect 3361 -21070 3400 -21053
rect 2812 -21086 3400 -21070
rect 3830 -21070 3869 -21053
rect 3903 -21070 3937 -21036
rect 3971 -21070 4005 -21036
rect 4039 -21070 4073 -21036
rect 4107 -21070 4141 -21036
rect 4175 -21070 4209 -21036
rect 4243 -21070 4277 -21036
rect 4311 -21070 4345 -21036
rect 4379 -21053 4604 -21036
rect 4662 -21036 5622 -20998
rect 4662 -21053 4887 -21036
rect 4379 -21070 4418 -21053
rect 3830 -21086 4418 -21070
rect 4848 -21070 4887 -21053
rect 4921 -21070 4955 -21036
rect 4989 -21070 5023 -21036
rect 5057 -21070 5091 -21036
rect 5125 -21070 5159 -21036
rect 5193 -21070 5227 -21036
rect 5261 -21070 5295 -21036
rect 5329 -21070 5363 -21036
rect 5397 -21053 5622 -21036
rect 5680 -21036 6640 -20998
rect 5680 -21053 5905 -21036
rect 5397 -21070 5436 -21053
rect 4848 -21086 5436 -21070
rect 5866 -21070 5905 -21053
rect 5939 -21070 5973 -21036
rect 6007 -21070 6041 -21036
rect 6075 -21070 6109 -21036
rect 6143 -21070 6177 -21036
rect 6211 -21070 6245 -21036
rect 6279 -21070 6313 -21036
rect 6347 -21070 6381 -21036
rect 6415 -21053 6640 -21036
rect 6698 -21036 7658 -20998
rect 6698 -21053 6923 -21036
rect 6415 -21070 6454 -21053
rect 5866 -21086 6454 -21070
rect 6884 -21070 6923 -21053
rect 6957 -21070 6991 -21036
rect 7025 -21070 7059 -21036
rect 7093 -21070 7127 -21036
rect 7161 -21070 7195 -21036
rect 7229 -21070 7263 -21036
rect 7297 -21070 7331 -21036
rect 7365 -21070 7399 -21036
rect 7433 -21053 7658 -21036
rect 7716 -21036 8676 -20998
rect 7716 -21053 7941 -21036
rect 7433 -21070 7472 -21053
rect 6884 -21086 7472 -21070
rect 7902 -21070 7941 -21053
rect 7975 -21070 8009 -21036
rect 8043 -21070 8077 -21036
rect 8111 -21070 8145 -21036
rect 8179 -21070 8213 -21036
rect 8247 -21070 8281 -21036
rect 8315 -21070 8349 -21036
rect 8383 -21070 8417 -21036
rect 8451 -21053 8676 -21036
rect 8734 -21036 9694 -20998
rect 8734 -21053 8959 -21036
rect 8451 -21070 8490 -21053
rect 7902 -21086 8490 -21070
rect 8920 -21070 8959 -21053
rect 8993 -21070 9027 -21036
rect 9061 -21070 9095 -21036
rect 9129 -21070 9163 -21036
rect 9197 -21070 9231 -21036
rect 9265 -21070 9299 -21036
rect 9333 -21070 9367 -21036
rect 9401 -21070 9435 -21036
rect 9469 -21053 9694 -21036
rect 9752 -21036 10712 -20998
rect 9752 -21053 9977 -21036
rect 9469 -21070 9508 -21053
rect 8920 -21086 9508 -21070
rect 9938 -21070 9977 -21053
rect 10011 -21070 10045 -21036
rect 10079 -21070 10113 -21036
rect 10147 -21070 10181 -21036
rect 10215 -21070 10249 -21036
rect 10283 -21070 10317 -21036
rect 10351 -21070 10385 -21036
rect 10419 -21070 10453 -21036
rect 10487 -21053 10712 -21036
rect 10770 -21036 11730 -20998
rect 10770 -21053 10995 -21036
rect 10487 -21070 10526 -21053
rect 9938 -21086 10526 -21070
rect 10956 -21070 10995 -21053
rect 11029 -21070 11063 -21036
rect 11097 -21070 11131 -21036
rect 11165 -21070 11199 -21036
rect 11233 -21070 11267 -21036
rect 11301 -21070 11335 -21036
rect 11369 -21070 11403 -21036
rect 11437 -21070 11471 -21036
rect 11505 -21053 11730 -21036
rect 11788 -21036 12748 -20998
rect 11788 -21053 12013 -21036
rect 11505 -21070 11544 -21053
rect 10956 -21086 11544 -21070
rect 11974 -21070 12013 -21053
rect 12047 -21070 12081 -21036
rect 12115 -21070 12149 -21036
rect 12183 -21070 12217 -21036
rect 12251 -21070 12285 -21036
rect 12319 -21070 12353 -21036
rect 12387 -21070 12421 -21036
rect 12455 -21070 12489 -21036
rect 12523 -21053 12748 -21036
rect 12806 -21036 13766 -20998
rect 12806 -21053 13031 -21036
rect 12523 -21070 12562 -21053
rect 11974 -21086 12562 -21070
rect 12992 -21070 13031 -21053
rect 13065 -21070 13099 -21036
rect 13133 -21070 13167 -21036
rect 13201 -21070 13235 -21036
rect 13269 -21070 13303 -21036
rect 13337 -21070 13371 -21036
rect 13405 -21070 13439 -21036
rect 13473 -21070 13507 -21036
rect 13541 -21053 13766 -21036
rect 13824 -21036 14784 -20998
rect 13824 -21053 14049 -21036
rect 13541 -21070 13580 -21053
rect 12992 -21086 13580 -21070
rect 14010 -21070 14049 -21053
rect 14083 -21070 14117 -21036
rect 14151 -21070 14185 -21036
rect 14219 -21070 14253 -21036
rect 14287 -21070 14321 -21036
rect 14355 -21070 14389 -21036
rect 14423 -21070 14457 -21036
rect 14491 -21070 14525 -21036
rect 14559 -21053 14784 -21036
rect 14842 -21036 15802 -20998
rect 14842 -21053 15067 -21036
rect 14559 -21070 14598 -21053
rect 14010 -21086 14598 -21070
rect 15028 -21070 15067 -21053
rect 15101 -21070 15135 -21036
rect 15169 -21070 15203 -21036
rect 15237 -21070 15271 -21036
rect 15305 -21070 15339 -21036
rect 15373 -21070 15407 -21036
rect 15441 -21070 15475 -21036
rect 15509 -21070 15543 -21036
rect 15577 -21053 15802 -21036
rect 15860 -21036 16820 -20998
rect 15860 -21053 16085 -21036
rect 15577 -21070 15616 -21053
rect 15028 -21086 15616 -21070
rect 16046 -21070 16085 -21053
rect 16119 -21070 16153 -21036
rect 16187 -21070 16221 -21036
rect 16255 -21070 16289 -21036
rect 16323 -21070 16357 -21036
rect 16391 -21070 16425 -21036
rect 16459 -21070 16493 -21036
rect 16527 -21070 16561 -21036
rect 16595 -21053 16820 -21036
rect 16878 -21036 17838 -20998
rect 16878 -21053 17103 -21036
rect 16595 -21070 16634 -21053
rect 16046 -21086 16634 -21070
rect 17064 -21070 17103 -21053
rect 17137 -21070 17171 -21036
rect 17205 -21070 17239 -21036
rect 17273 -21070 17307 -21036
rect 17341 -21070 17375 -21036
rect 17409 -21070 17443 -21036
rect 17477 -21070 17511 -21036
rect 17545 -21070 17579 -21036
rect 17613 -21053 17838 -21036
rect 17896 -21036 18856 -20998
rect 17896 -21053 18121 -21036
rect 17613 -21070 17652 -21053
rect 17064 -21086 17652 -21070
rect 18082 -21070 18121 -21053
rect 18155 -21070 18189 -21036
rect 18223 -21070 18257 -21036
rect 18291 -21070 18325 -21036
rect 18359 -21070 18393 -21036
rect 18427 -21070 18461 -21036
rect 18495 -21070 18529 -21036
rect 18563 -21070 18597 -21036
rect 18631 -21053 18856 -21036
rect 18914 -21036 19874 -20998
rect 18914 -21053 19139 -21036
rect 18631 -21070 18670 -21053
rect 18082 -21086 18670 -21070
rect 19100 -21070 19139 -21053
rect 19173 -21070 19207 -21036
rect 19241 -21070 19275 -21036
rect 19309 -21070 19343 -21036
rect 19377 -21070 19411 -21036
rect 19445 -21070 19479 -21036
rect 19513 -21070 19547 -21036
rect 19581 -21070 19615 -21036
rect 19649 -21053 19874 -21036
rect 19932 -21036 20892 -20998
rect 19932 -21053 20157 -21036
rect 19649 -21070 19688 -21053
rect 19100 -21086 19688 -21070
rect 20118 -21070 20157 -21053
rect 20191 -21070 20225 -21036
rect 20259 -21070 20293 -21036
rect 20327 -21070 20361 -21036
rect 20395 -21070 20429 -21036
rect 20463 -21070 20497 -21036
rect 20531 -21070 20565 -21036
rect 20599 -21070 20633 -21036
rect 20667 -21053 20892 -21036
rect 20950 -21036 21910 -20998
rect 20950 -21053 21175 -21036
rect 20667 -21070 20706 -21053
rect 20118 -21086 20706 -21070
rect 21136 -21070 21175 -21053
rect 21209 -21070 21243 -21036
rect 21277 -21070 21311 -21036
rect 21345 -21070 21379 -21036
rect 21413 -21070 21447 -21036
rect 21481 -21070 21515 -21036
rect 21549 -21070 21583 -21036
rect 21617 -21070 21651 -21036
rect 21685 -21053 21910 -21036
rect 21968 -21036 22928 -20998
rect 21968 -21053 22193 -21036
rect 21685 -21070 21724 -21053
rect 21136 -21086 21724 -21070
rect 22154 -21070 22193 -21053
rect 22227 -21070 22261 -21036
rect 22295 -21070 22329 -21036
rect 22363 -21070 22397 -21036
rect 22431 -21070 22465 -21036
rect 22499 -21070 22533 -21036
rect 22567 -21070 22601 -21036
rect 22635 -21070 22669 -21036
rect 22703 -21053 22928 -21036
rect 22703 -21070 22742 -21053
rect 22154 -21086 22742 -21070
rect 2812 -21560 3400 -21544
rect 2812 -21577 2851 -21560
rect 2626 -21594 2851 -21577
rect 2885 -21594 2919 -21560
rect 2953 -21594 2987 -21560
rect 3021 -21594 3055 -21560
rect 3089 -21594 3123 -21560
rect 3157 -21594 3191 -21560
rect 3225 -21594 3259 -21560
rect 3293 -21594 3327 -21560
rect 3361 -21577 3400 -21560
rect 3830 -21560 4418 -21544
rect 3830 -21577 3869 -21560
rect 3361 -21594 3586 -21577
rect 2626 -21632 3586 -21594
rect 3644 -21594 3869 -21577
rect 3903 -21594 3937 -21560
rect 3971 -21594 4005 -21560
rect 4039 -21594 4073 -21560
rect 4107 -21594 4141 -21560
rect 4175 -21594 4209 -21560
rect 4243 -21594 4277 -21560
rect 4311 -21594 4345 -21560
rect 4379 -21577 4418 -21560
rect 4848 -21560 5436 -21544
rect 4848 -21577 4887 -21560
rect 4379 -21594 4604 -21577
rect 3644 -21632 4604 -21594
rect 4662 -21594 4887 -21577
rect 4921 -21594 4955 -21560
rect 4989 -21594 5023 -21560
rect 5057 -21594 5091 -21560
rect 5125 -21594 5159 -21560
rect 5193 -21594 5227 -21560
rect 5261 -21594 5295 -21560
rect 5329 -21594 5363 -21560
rect 5397 -21577 5436 -21560
rect 5866 -21560 6454 -21544
rect 5866 -21577 5905 -21560
rect 5397 -21594 5622 -21577
rect 4662 -21632 5622 -21594
rect 5680 -21594 5905 -21577
rect 5939 -21594 5973 -21560
rect 6007 -21594 6041 -21560
rect 6075 -21594 6109 -21560
rect 6143 -21594 6177 -21560
rect 6211 -21594 6245 -21560
rect 6279 -21594 6313 -21560
rect 6347 -21594 6381 -21560
rect 6415 -21577 6454 -21560
rect 6884 -21560 7472 -21544
rect 6884 -21577 6923 -21560
rect 6415 -21594 6640 -21577
rect 5680 -21632 6640 -21594
rect 6698 -21594 6923 -21577
rect 6957 -21594 6991 -21560
rect 7025 -21594 7059 -21560
rect 7093 -21594 7127 -21560
rect 7161 -21594 7195 -21560
rect 7229 -21594 7263 -21560
rect 7297 -21594 7331 -21560
rect 7365 -21594 7399 -21560
rect 7433 -21577 7472 -21560
rect 7902 -21560 8490 -21544
rect 7902 -21577 7941 -21560
rect 7433 -21594 7658 -21577
rect 6698 -21632 7658 -21594
rect 7716 -21594 7941 -21577
rect 7975 -21594 8009 -21560
rect 8043 -21594 8077 -21560
rect 8111 -21594 8145 -21560
rect 8179 -21594 8213 -21560
rect 8247 -21594 8281 -21560
rect 8315 -21594 8349 -21560
rect 8383 -21594 8417 -21560
rect 8451 -21577 8490 -21560
rect 8920 -21560 9508 -21544
rect 8920 -21577 8959 -21560
rect 8451 -21594 8676 -21577
rect 7716 -21632 8676 -21594
rect 8734 -21594 8959 -21577
rect 8993 -21594 9027 -21560
rect 9061 -21594 9095 -21560
rect 9129 -21594 9163 -21560
rect 9197 -21594 9231 -21560
rect 9265 -21594 9299 -21560
rect 9333 -21594 9367 -21560
rect 9401 -21594 9435 -21560
rect 9469 -21577 9508 -21560
rect 9938 -21560 10526 -21544
rect 9938 -21577 9977 -21560
rect 9469 -21594 9694 -21577
rect 8734 -21632 9694 -21594
rect 9752 -21594 9977 -21577
rect 10011 -21594 10045 -21560
rect 10079 -21594 10113 -21560
rect 10147 -21594 10181 -21560
rect 10215 -21594 10249 -21560
rect 10283 -21594 10317 -21560
rect 10351 -21594 10385 -21560
rect 10419 -21594 10453 -21560
rect 10487 -21577 10526 -21560
rect 10956 -21560 11544 -21544
rect 10956 -21577 10995 -21560
rect 10487 -21594 10712 -21577
rect 9752 -21632 10712 -21594
rect 10770 -21594 10995 -21577
rect 11029 -21594 11063 -21560
rect 11097 -21594 11131 -21560
rect 11165 -21594 11199 -21560
rect 11233 -21594 11267 -21560
rect 11301 -21594 11335 -21560
rect 11369 -21594 11403 -21560
rect 11437 -21594 11471 -21560
rect 11505 -21577 11544 -21560
rect 11974 -21560 12562 -21544
rect 11974 -21577 12013 -21560
rect 11505 -21594 11730 -21577
rect 10770 -21632 11730 -21594
rect 11788 -21594 12013 -21577
rect 12047 -21594 12081 -21560
rect 12115 -21594 12149 -21560
rect 12183 -21594 12217 -21560
rect 12251 -21594 12285 -21560
rect 12319 -21594 12353 -21560
rect 12387 -21594 12421 -21560
rect 12455 -21594 12489 -21560
rect 12523 -21577 12562 -21560
rect 12992 -21560 13580 -21544
rect 12992 -21577 13031 -21560
rect 12523 -21594 12748 -21577
rect 11788 -21632 12748 -21594
rect 12806 -21594 13031 -21577
rect 13065 -21594 13099 -21560
rect 13133 -21594 13167 -21560
rect 13201 -21594 13235 -21560
rect 13269 -21594 13303 -21560
rect 13337 -21594 13371 -21560
rect 13405 -21594 13439 -21560
rect 13473 -21594 13507 -21560
rect 13541 -21577 13580 -21560
rect 14010 -21560 14598 -21544
rect 14010 -21577 14049 -21560
rect 13541 -21594 13766 -21577
rect 12806 -21632 13766 -21594
rect 13824 -21594 14049 -21577
rect 14083 -21594 14117 -21560
rect 14151 -21594 14185 -21560
rect 14219 -21594 14253 -21560
rect 14287 -21594 14321 -21560
rect 14355 -21594 14389 -21560
rect 14423 -21594 14457 -21560
rect 14491 -21594 14525 -21560
rect 14559 -21577 14598 -21560
rect 15028 -21560 15616 -21544
rect 15028 -21577 15067 -21560
rect 14559 -21594 14784 -21577
rect 13824 -21632 14784 -21594
rect 14842 -21594 15067 -21577
rect 15101 -21594 15135 -21560
rect 15169 -21594 15203 -21560
rect 15237 -21594 15271 -21560
rect 15305 -21594 15339 -21560
rect 15373 -21594 15407 -21560
rect 15441 -21594 15475 -21560
rect 15509 -21594 15543 -21560
rect 15577 -21577 15616 -21560
rect 16046 -21560 16634 -21544
rect 16046 -21577 16085 -21560
rect 15577 -21594 15802 -21577
rect 14842 -21632 15802 -21594
rect 15860 -21594 16085 -21577
rect 16119 -21594 16153 -21560
rect 16187 -21594 16221 -21560
rect 16255 -21594 16289 -21560
rect 16323 -21594 16357 -21560
rect 16391 -21594 16425 -21560
rect 16459 -21594 16493 -21560
rect 16527 -21594 16561 -21560
rect 16595 -21577 16634 -21560
rect 17064 -21560 17652 -21544
rect 17064 -21577 17103 -21560
rect 16595 -21594 16820 -21577
rect 15860 -21632 16820 -21594
rect 16878 -21594 17103 -21577
rect 17137 -21594 17171 -21560
rect 17205 -21594 17239 -21560
rect 17273 -21594 17307 -21560
rect 17341 -21594 17375 -21560
rect 17409 -21594 17443 -21560
rect 17477 -21594 17511 -21560
rect 17545 -21594 17579 -21560
rect 17613 -21577 17652 -21560
rect 18082 -21560 18670 -21544
rect 18082 -21577 18121 -21560
rect 17613 -21594 17838 -21577
rect 16878 -21632 17838 -21594
rect 17896 -21594 18121 -21577
rect 18155 -21594 18189 -21560
rect 18223 -21594 18257 -21560
rect 18291 -21594 18325 -21560
rect 18359 -21594 18393 -21560
rect 18427 -21594 18461 -21560
rect 18495 -21594 18529 -21560
rect 18563 -21594 18597 -21560
rect 18631 -21577 18670 -21560
rect 19100 -21560 19688 -21544
rect 19100 -21577 19139 -21560
rect 18631 -21594 18856 -21577
rect 17896 -21632 18856 -21594
rect 18914 -21594 19139 -21577
rect 19173 -21594 19207 -21560
rect 19241 -21594 19275 -21560
rect 19309 -21594 19343 -21560
rect 19377 -21594 19411 -21560
rect 19445 -21594 19479 -21560
rect 19513 -21594 19547 -21560
rect 19581 -21594 19615 -21560
rect 19649 -21577 19688 -21560
rect 20118 -21560 20706 -21544
rect 20118 -21577 20157 -21560
rect 19649 -21594 19874 -21577
rect 18914 -21632 19874 -21594
rect 19932 -21594 20157 -21577
rect 20191 -21594 20225 -21560
rect 20259 -21594 20293 -21560
rect 20327 -21594 20361 -21560
rect 20395 -21594 20429 -21560
rect 20463 -21594 20497 -21560
rect 20531 -21594 20565 -21560
rect 20599 -21594 20633 -21560
rect 20667 -21577 20706 -21560
rect 21136 -21560 21724 -21544
rect 21136 -21577 21175 -21560
rect 20667 -21594 20892 -21577
rect 19932 -21632 20892 -21594
rect 20950 -21594 21175 -21577
rect 21209 -21594 21243 -21560
rect 21277 -21594 21311 -21560
rect 21345 -21594 21379 -21560
rect 21413 -21594 21447 -21560
rect 21481 -21594 21515 -21560
rect 21549 -21594 21583 -21560
rect 21617 -21594 21651 -21560
rect 21685 -21577 21724 -21560
rect 22154 -21560 22742 -21544
rect 22154 -21577 22193 -21560
rect 21685 -21594 21910 -21577
rect 20950 -21632 21910 -21594
rect 21968 -21594 22193 -21577
rect 22227 -21594 22261 -21560
rect 22295 -21594 22329 -21560
rect 22363 -21594 22397 -21560
rect 22431 -21594 22465 -21560
rect 22499 -21594 22533 -21560
rect 22567 -21594 22601 -21560
rect 22635 -21594 22669 -21560
rect 22703 -21577 22742 -21560
rect 22703 -21594 22928 -21577
rect 21968 -21632 22928 -21594
rect 2626 -22270 3586 -22232
rect 2626 -22287 2851 -22270
rect 2812 -22304 2851 -22287
rect 2885 -22304 2919 -22270
rect 2953 -22304 2987 -22270
rect 3021 -22304 3055 -22270
rect 3089 -22304 3123 -22270
rect 3157 -22304 3191 -22270
rect 3225 -22304 3259 -22270
rect 3293 -22304 3327 -22270
rect 3361 -22287 3586 -22270
rect 3644 -22270 4604 -22232
rect 3644 -22287 3869 -22270
rect 3361 -22304 3400 -22287
rect 2812 -22320 3400 -22304
rect 3830 -22304 3869 -22287
rect 3903 -22304 3937 -22270
rect 3971 -22304 4005 -22270
rect 4039 -22304 4073 -22270
rect 4107 -22304 4141 -22270
rect 4175 -22304 4209 -22270
rect 4243 -22304 4277 -22270
rect 4311 -22304 4345 -22270
rect 4379 -22287 4604 -22270
rect 4662 -22270 5622 -22232
rect 4662 -22287 4887 -22270
rect 4379 -22304 4418 -22287
rect 3830 -22320 4418 -22304
rect 4848 -22304 4887 -22287
rect 4921 -22304 4955 -22270
rect 4989 -22304 5023 -22270
rect 5057 -22304 5091 -22270
rect 5125 -22304 5159 -22270
rect 5193 -22304 5227 -22270
rect 5261 -22304 5295 -22270
rect 5329 -22304 5363 -22270
rect 5397 -22287 5622 -22270
rect 5680 -22270 6640 -22232
rect 5680 -22287 5905 -22270
rect 5397 -22304 5436 -22287
rect 4848 -22320 5436 -22304
rect 5866 -22304 5905 -22287
rect 5939 -22304 5973 -22270
rect 6007 -22304 6041 -22270
rect 6075 -22304 6109 -22270
rect 6143 -22304 6177 -22270
rect 6211 -22304 6245 -22270
rect 6279 -22304 6313 -22270
rect 6347 -22304 6381 -22270
rect 6415 -22287 6640 -22270
rect 6698 -22270 7658 -22232
rect 6698 -22287 6923 -22270
rect 6415 -22304 6454 -22287
rect 5866 -22320 6454 -22304
rect 6884 -22304 6923 -22287
rect 6957 -22304 6991 -22270
rect 7025 -22304 7059 -22270
rect 7093 -22304 7127 -22270
rect 7161 -22304 7195 -22270
rect 7229 -22304 7263 -22270
rect 7297 -22304 7331 -22270
rect 7365 -22304 7399 -22270
rect 7433 -22287 7658 -22270
rect 7716 -22270 8676 -22232
rect 7716 -22287 7941 -22270
rect 7433 -22304 7472 -22287
rect 6884 -22320 7472 -22304
rect 7902 -22304 7941 -22287
rect 7975 -22304 8009 -22270
rect 8043 -22304 8077 -22270
rect 8111 -22304 8145 -22270
rect 8179 -22304 8213 -22270
rect 8247 -22304 8281 -22270
rect 8315 -22304 8349 -22270
rect 8383 -22304 8417 -22270
rect 8451 -22287 8676 -22270
rect 8734 -22270 9694 -22232
rect 8734 -22287 8959 -22270
rect 8451 -22304 8490 -22287
rect 7902 -22320 8490 -22304
rect 8920 -22304 8959 -22287
rect 8993 -22304 9027 -22270
rect 9061 -22304 9095 -22270
rect 9129 -22304 9163 -22270
rect 9197 -22304 9231 -22270
rect 9265 -22304 9299 -22270
rect 9333 -22304 9367 -22270
rect 9401 -22304 9435 -22270
rect 9469 -22287 9694 -22270
rect 9752 -22270 10712 -22232
rect 9752 -22287 9977 -22270
rect 9469 -22304 9508 -22287
rect 8920 -22320 9508 -22304
rect 9938 -22304 9977 -22287
rect 10011 -22304 10045 -22270
rect 10079 -22304 10113 -22270
rect 10147 -22304 10181 -22270
rect 10215 -22304 10249 -22270
rect 10283 -22304 10317 -22270
rect 10351 -22304 10385 -22270
rect 10419 -22304 10453 -22270
rect 10487 -22287 10712 -22270
rect 10770 -22270 11730 -22232
rect 10770 -22287 10995 -22270
rect 10487 -22304 10526 -22287
rect 9938 -22320 10526 -22304
rect 10956 -22304 10995 -22287
rect 11029 -22304 11063 -22270
rect 11097 -22304 11131 -22270
rect 11165 -22304 11199 -22270
rect 11233 -22304 11267 -22270
rect 11301 -22304 11335 -22270
rect 11369 -22304 11403 -22270
rect 11437 -22304 11471 -22270
rect 11505 -22287 11730 -22270
rect 11788 -22270 12748 -22232
rect 11788 -22287 12013 -22270
rect 11505 -22304 11544 -22287
rect 10956 -22320 11544 -22304
rect 11974 -22304 12013 -22287
rect 12047 -22304 12081 -22270
rect 12115 -22304 12149 -22270
rect 12183 -22304 12217 -22270
rect 12251 -22304 12285 -22270
rect 12319 -22304 12353 -22270
rect 12387 -22304 12421 -22270
rect 12455 -22304 12489 -22270
rect 12523 -22287 12748 -22270
rect 12806 -22270 13766 -22232
rect 12806 -22287 13031 -22270
rect 12523 -22304 12562 -22287
rect 11974 -22320 12562 -22304
rect 12992 -22304 13031 -22287
rect 13065 -22304 13099 -22270
rect 13133 -22304 13167 -22270
rect 13201 -22304 13235 -22270
rect 13269 -22304 13303 -22270
rect 13337 -22304 13371 -22270
rect 13405 -22304 13439 -22270
rect 13473 -22304 13507 -22270
rect 13541 -22287 13766 -22270
rect 13824 -22270 14784 -22232
rect 13824 -22287 14049 -22270
rect 13541 -22304 13580 -22287
rect 12992 -22320 13580 -22304
rect 14010 -22304 14049 -22287
rect 14083 -22304 14117 -22270
rect 14151 -22304 14185 -22270
rect 14219 -22304 14253 -22270
rect 14287 -22304 14321 -22270
rect 14355 -22304 14389 -22270
rect 14423 -22304 14457 -22270
rect 14491 -22304 14525 -22270
rect 14559 -22287 14784 -22270
rect 14842 -22270 15802 -22232
rect 14842 -22287 15067 -22270
rect 14559 -22304 14598 -22287
rect 14010 -22320 14598 -22304
rect 15028 -22304 15067 -22287
rect 15101 -22304 15135 -22270
rect 15169 -22304 15203 -22270
rect 15237 -22304 15271 -22270
rect 15305 -22304 15339 -22270
rect 15373 -22304 15407 -22270
rect 15441 -22304 15475 -22270
rect 15509 -22304 15543 -22270
rect 15577 -22287 15802 -22270
rect 15860 -22270 16820 -22232
rect 15860 -22287 16085 -22270
rect 15577 -22304 15616 -22287
rect 15028 -22320 15616 -22304
rect 16046 -22304 16085 -22287
rect 16119 -22304 16153 -22270
rect 16187 -22304 16221 -22270
rect 16255 -22304 16289 -22270
rect 16323 -22304 16357 -22270
rect 16391 -22304 16425 -22270
rect 16459 -22304 16493 -22270
rect 16527 -22304 16561 -22270
rect 16595 -22287 16820 -22270
rect 16878 -22270 17838 -22232
rect 16878 -22287 17103 -22270
rect 16595 -22304 16634 -22287
rect 16046 -22320 16634 -22304
rect 17064 -22304 17103 -22287
rect 17137 -22304 17171 -22270
rect 17205 -22304 17239 -22270
rect 17273 -22304 17307 -22270
rect 17341 -22304 17375 -22270
rect 17409 -22304 17443 -22270
rect 17477 -22304 17511 -22270
rect 17545 -22304 17579 -22270
rect 17613 -22287 17838 -22270
rect 17896 -22270 18856 -22232
rect 17896 -22287 18121 -22270
rect 17613 -22304 17652 -22287
rect 17064 -22320 17652 -22304
rect 18082 -22304 18121 -22287
rect 18155 -22304 18189 -22270
rect 18223 -22304 18257 -22270
rect 18291 -22304 18325 -22270
rect 18359 -22304 18393 -22270
rect 18427 -22304 18461 -22270
rect 18495 -22304 18529 -22270
rect 18563 -22304 18597 -22270
rect 18631 -22287 18856 -22270
rect 18914 -22270 19874 -22232
rect 18914 -22287 19139 -22270
rect 18631 -22304 18670 -22287
rect 18082 -22320 18670 -22304
rect 19100 -22304 19139 -22287
rect 19173 -22304 19207 -22270
rect 19241 -22304 19275 -22270
rect 19309 -22304 19343 -22270
rect 19377 -22304 19411 -22270
rect 19445 -22304 19479 -22270
rect 19513 -22304 19547 -22270
rect 19581 -22304 19615 -22270
rect 19649 -22287 19874 -22270
rect 19932 -22270 20892 -22232
rect 19932 -22287 20157 -22270
rect 19649 -22304 19688 -22287
rect 19100 -22320 19688 -22304
rect 20118 -22304 20157 -22287
rect 20191 -22304 20225 -22270
rect 20259 -22304 20293 -22270
rect 20327 -22304 20361 -22270
rect 20395 -22304 20429 -22270
rect 20463 -22304 20497 -22270
rect 20531 -22304 20565 -22270
rect 20599 -22304 20633 -22270
rect 20667 -22287 20892 -22270
rect 20950 -22270 21910 -22232
rect 20950 -22287 21175 -22270
rect 20667 -22304 20706 -22287
rect 20118 -22320 20706 -22304
rect 21136 -22304 21175 -22287
rect 21209 -22304 21243 -22270
rect 21277 -22304 21311 -22270
rect 21345 -22304 21379 -22270
rect 21413 -22304 21447 -22270
rect 21481 -22304 21515 -22270
rect 21549 -22304 21583 -22270
rect 21617 -22304 21651 -22270
rect 21685 -22287 21910 -22270
rect 21968 -22270 22928 -22232
rect 21968 -22287 22193 -22270
rect 21685 -22304 21724 -22287
rect 21136 -22320 21724 -22304
rect 22154 -22304 22193 -22287
rect 22227 -22304 22261 -22270
rect 22295 -22304 22329 -22270
rect 22363 -22304 22397 -22270
rect 22431 -22304 22465 -22270
rect 22499 -22304 22533 -22270
rect 22567 -22304 22601 -22270
rect 22635 -22304 22669 -22270
rect 22703 -22287 22928 -22270
rect 22703 -22304 22742 -22287
rect 22154 -22320 22742 -22304
rect 2812 -22792 3400 -22776
rect 2812 -22809 2851 -22792
rect 2626 -22826 2851 -22809
rect 2885 -22826 2919 -22792
rect 2953 -22826 2987 -22792
rect 3021 -22826 3055 -22792
rect 3089 -22826 3123 -22792
rect 3157 -22826 3191 -22792
rect 3225 -22826 3259 -22792
rect 3293 -22826 3327 -22792
rect 3361 -22809 3400 -22792
rect 3830 -22792 4418 -22776
rect 3830 -22809 3869 -22792
rect 3361 -22826 3586 -22809
rect 2626 -22864 3586 -22826
rect 3644 -22826 3869 -22809
rect 3903 -22826 3937 -22792
rect 3971 -22826 4005 -22792
rect 4039 -22826 4073 -22792
rect 4107 -22826 4141 -22792
rect 4175 -22826 4209 -22792
rect 4243 -22826 4277 -22792
rect 4311 -22826 4345 -22792
rect 4379 -22809 4418 -22792
rect 4848 -22792 5436 -22776
rect 4848 -22809 4887 -22792
rect 4379 -22826 4604 -22809
rect 3644 -22864 4604 -22826
rect 4662 -22826 4887 -22809
rect 4921 -22826 4955 -22792
rect 4989 -22826 5023 -22792
rect 5057 -22826 5091 -22792
rect 5125 -22826 5159 -22792
rect 5193 -22826 5227 -22792
rect 5261 -22826 5295 -22792
rect 5329 -22826 5363 -22792
rect 5397 -22809 5436 -22792
rect 5866 -22792 6454 -22776
rect 5866 -22809 5905 -22792
rect 5397 -22826 5622 -22809
rect 4662 -22864 5622 -22826
rect 5680 -22826 5905 -22809
rect 5939 -22826 5973 -22792
rect 6007 -22826 6041 -22792
rect 6075 -22826 6109 -22792
rect 6143 -22826 6177 -22792
rect 6211 -22826 6245 -22792
rect 6279 -22826 6313 -22792
rect 6347 -22826 6381 -22792
rect 6415 -22809 6454 -22792
rect 6884 -22792 7472 -22776
rect 6884 -22809 6923 -22792
rect 6415 -22826 6640 -22809
rect 5680 -22864 6640 -22826
rect 6698 -22826 6923 -22809
rect 6957 -22826 6991 -22792
rect 7025 -22826 7059 -22792
rect 7093 -22826 7127 -22792
rect 7161 -22826 7195 -22792
rect 7229 -22826 7263 -22792
rect 7297 -22826 7331 -22792
rect 7365 -22826 7399 -22792
rect 7433 -22809 7472 -22792
rect 7902 -22792 8490 -22776
rect 7902 -22809 7941 -22792
rect 7433 -22826 7658 -22809
rect 6698 -22864 7658 -22826
rect 7716 -22826 7941 -22809
rect 7975 -22826 8009 -22792
rect 8043 -22826 8077 -22792
rect 8111 -22826 8145 -22792
rect 8179 -22826 8213 -22792
rect 8247 -22826 8281 -22792
rect 8315 -22826 8349 -22792
rect 8383 -22826 8417 -22792
rect 8451 -22809 8490 -22792
rect 8920 -22792 9508 -22776
rect 8920 -22809 8959 -22792
rect 8451 -22826 8676 -22809
rect 7716 -22864 8676 -22826
rect 8734 -22826 8959 -22809
rect 8993 -22826 9027 -22792
rect 9061 -22826 9095 -22792
rect 9129 -22826 9163 -22792
rect 9197 -22826 9231 -22792
rect 9265 -22826 9299 -22792
rect 9333 -22826 9367 -22792
rect 9401 -22826 9435 -22792
rect 9469 -22809 9508 -22792
rect 9938 -22792 10526 -22776
rect 9938 -22809 9977 -22792
rect 9469 -22826 9694 -22809
rect 8734 -22864 9694 -22826
rect 9752 -22826 9977 -22809
rect 10011 -22826 10045 -22792
rect 10079 -22826 10113 -22792
rect 10147 -22826 10181 -22792
rect 10215 -22826 10249 -22792
rect 10283 -22826 10317 -22792
rect 10351 -22826 10385 -22792
rect 10419 -22826 10453 -22792
rect 10487 -22809 10526 -22792
rect 10956 -22792 11544 -22776
rect 10956 -22809 10995 -22792
rect 10487 -22826 10712 -22809
rect 9752 -22864 10712 -22826
rect 10770 -22826 10995 -22809
rect 11029 -22826 11063 -22792
rect 11097 -22826 11131 -22792
rect 11165 -22826 11199 -22792
rect 11233 -22826 11267 -22792
rect 11301 -22826 11335 -22792
rect 11369 -22826 11403 -22792
rect 11437 -22826 11471 -22792
rect 11505 -22809 11544 -22792
rect 11974 -22792 12562 -22776
rect 11974 -22809 12013 -22792
rect 11505 -22826 11730 -22809
rect 10770 -22864 11730 -22826
rect 11788 -22826 12013 -22809
rect 12047 -22826 12081 -22792
rect 12115 -22826 12149 -22792
rect 12183 -22826 12217 -22792
rect 12251 -22826 12285 -22792
rect 12319 -22826 12353 -22792
rect 12387 -22826 12421 -22792
rect 12455 -22826 12489 -22792
rect 12523 -22809 12562 -22792
rect 12992 -22792 13580 -22776
rect 12992 -22809 13031 -22792
rect 12523 -22826 12748 -22809
rect 11788 -22864 12748 -22826
rect 12806 -22826 13031 -22809
rect 13065 -22826 13099 -22792
rect 13133 -22826 13167 -22792
rect 13201 -22826 13235 -22792
rect 13269 -22826 13303 -22792
rect 13337 -22826 13371 -22792
rect 13405 -22826 13439 -22792
rect 13473 -22826 13507 -22792
rect 13541 -22809 13580 -22792
rect 14010 -22792 14598 -22776
rect 14010 -22809 14049 -22792
rect 13541 -22826 13766 -22809
rect 12806 -22864 13766 -22826
rect 13824 -22826 14049 -22809
rect 14083 -22826 14117 -22792
rect 14151 -22826 14185 -22792
rect 14219 -22826 14253 -22792
rect 14287 -22826 14321 -22792
rect 14355 -22826 14389 -22792
rect 14423 -22826 14457 -22792
rect 14491 -22826 14525 -22792
rect 14559 -22809 14598 -22792
rect 15028 -22792 15616 -22776
rect 15028 -22809 15067 -22792
rect 14559 -22826 14784 -22809
rect 13824 -22864 14784 -22826
rect 14842 -22826 15067 -22809
rect 15101 -22826 15135 -22792
rect 15169 -22826 15203 -22792
rect 15237 -22826 15271 -22792
rect 15305 -22826 15339 -22792
rect 15373 -22826 15407 -22792
rect 15441 -22826 15475 -22792
rect 15509 -22826 15543 -22792
rect 15577 -22809 15616 -22792
rect 16046 -22792 16634 -22776
rect 16046 -22809 16085 -22792
rect 15577 -22826 15802 -22809
rect 14842 -22864 15802 -22826
rect 15860 -22826 16085 -22809
rect 16119 -22826 16153 -22792
rect 16187 -22826 16221 -22792
rect 16255 -22826 16289 -22792
rect 16323 -22826 16357 -22792
rect 16391 -22826 16425 -22792
rect 16459 -22826 16493 -22792
rect 16527 -22826 16561 -22792
rect 16595 -22809 16634 -22792
rect 17064 -22792 17652 -22776
rect 17064 -22809 17103 -22792
rect 16595 -22826 16820 -22809
rect 15860 -22864 16820 -22826
rect 16878 -22826 17103 -22809
rect 17137 -22826 17171 -22792
rect 17205 -22826 17239 -22792
rect 17273 -22826 17307 -22792
rect 17341 -22826 17375 -22792
rect 17409 -22826 17443 -22792
rect 17477 -22826 17511 -22792
rect 17545 -22826 17579 -22792
rect 17613 -22809 17652 -22792
rect 18082 -22792 18670 -22776
rect 18082 -22809 18121 -22792
rect 17613 -22826 17838 -22809
rect 16878 -22864 17838 -22826
rect 17896 -22826 18121 -22809
rect 18155 -22826 18189 -22792
rect 18223 -22826 18257 -22792
rect 18291 -22826 18325 -22792
rect 18359 -22826 18393 -22792
rect 18427 -22826 18461 -22792
rect 18495 -22826 18529 -22792
rect 18563 -22826 18597 -22792
rect 18631 -22809 18670 -22792
rect 19100 -22792 19688 -22776
rect 19100 -22809 19139 -22792
rect 18631 -22826 18856 -22809
rect 17896 -22864 18856 -22826
rect 18914 -22826 19139 -22809
rect 19173 -22826 19207 -22792
rect 19241 -22826 19275 -22792
rect 19309 -22826 19343 -22792
rect 19377 -22826 19411 -22792
rect 19445 -22826 19479 -22792
rect 19513 -22826 19547 -22792
rect 19581 -22826 19615 -22792
rect 19649 -22809 19688 -22792
rect 20118 -22792 20706 -22776
rect 20118 -22809 20157 -22792
rect 19649 -22826 19874 -22809
rect 18914 -22864 19874 -22826
rect 19932 -22826 20157 -22809
rect 20191 -22826 20225 -22792
rect 20259 -22826 20293 -22792
rect 20327 -22826 20361 -22792
rect 20395 -22826 20429 -22792
rect 20463 -22826 20497 -22792
rect 20531 -22826 20565 -22792
rect 20599 -22826 20633 -22792
rect 20667 -22809 20706 -22792
rect 21136 -22792 21724 -22776
rect 21136 -22809 21175 -22792
rect 20667 -22826 20892 -22809
rect 19932 -22864 20892 -22826
rect 20950 -22826 21175 -22809
rect 21209 -22826 21243 -22792
rect 21277 -22826 21311 -22792
rect 21345 -22826 21379 -22792
rect 21413 -22826 21447 -22792
rect 21481 -22826 21515 -22792
rect 21549 -22826 21583 -22792
rect 21617 -22826 21651 -22792
rect 21685 -22809 21724 -22792
rect 22154 -22792 22742 -22776
rect 22154 -22809 22193 -22792
rect 21685 -22826 21910 -22809
rect 20950 -22864 21910 -22826
rect 21968 -22826 22193 -22809
rect 22227 -22826 22261 -22792
rect 22295 -22826 22329 -22792
rect 22363 -22826 22397 -22792
rect 22431 -22826 22465 -22792
rect 22499 -22826 22533 -22792
rect 22567 -22826 22601 -22792
rect 22635 -22826 22669 -22792
rect 22703 -22809 22742 -22792
rect 22703 -22826 22928 -22809
rect 21968 -22864 22928 -22826
rect 2626 -23502 3586 -23464
rect 2626 -23519 2851 -23502
rect 2812 -23536 2851 -23519
rect 2885 -23536 2919 -23502
rect 2953 -23536 2987 -23502
rect 3021 -23536 3055 -23502
rect 3089 -23536 3123 -23502
rect 3157 -23536 3191 -23502
rect 3225 -23536 3259 -23502
rect 3293 -23536 3327 -23502
rect 3361 -23519 3586 -23502
rect 3644 -23502 4604 -23464
rect 3644 -23519 3869 -23502
rect 3361 -23536 3400 -23519
rect 2812 -23552 3400 -23536
rect 3830 -23536 3869 -23519
rect 3903 -23536 3937 -23502
rect 3971 -23536 4005 -23502
rect 4039 -23536 4073 -23502
rect 4107 -23536 4141 -23502
rect 4175 -23536 4209 -23502
rect 4243 -23536 4277 -23502
rect 4311 -23536 4345 -23502
rect 4379 -23519 4604 -23502
rect 4662 -23502 5622 -23464
rect 4662 -23519 4887 -23502
rect 4379 -23536 4418 -23519
rect 3830 -23552 4418 -23536
rect 4848 -23536 4887 -23519
rect 4921 -23536 4955 -23502
rect 4989 -23536 5023 -23502
rect 5057 -23536 5091 -23502
rect 5125 -23536 5159 -23502
rect 5193 -23536 5227 -23502
rect 5261 -23536 5295 -23502
rect 5329 -23536 5363 -23502
rect 5397 -23519 5622 -23502
rect 5680 -23502 6640 -23464
rect 5680 -23519 5905 -23502
rect 5397 -23536 5436 -23519
rect 4848 -23552 5436 -23536
rect 5866 -23536 5905 -23519
rect 5939 -23536 5973 -23502
rect 6007 -23536 6041 -23502
rect 6075 -23536 6109 -23502
rect 6143 -23536 6177 -23502
rect 6211 -23536 6245 -23502
rect 6279 -23536 6313 -23502
rect 6347 -23536 6381 -23502
rect 6415 -23519 6640 -23502
rect 6698 -23502 7658 -23464
rect 6698 -23519 6923 -23502
rect 6415 -23536 6454 -23519
rect 5866 -23552 6454 -23536
rect 6884 -23536 6923 -23519
rect 6957 -23536 6991 -23502
rect 7025 -23536 7059 -23502
rect 7093 -23536 7127 -23502
rect 7161 -23536 7195 -23502
rect 7229 -23536 7263 -23502
rect 7297 -23536 7331 -23502
rect 7365 -23536 7399 -23502
rect 7433 -23519 7658 -23502
rect 7716 -23502 8676 -23464
rect 7716 -23519 7941 -23502
rect 7433 -23536 7472 -23519
rect 6884 -23552 7472 -23536
rect 7902 -23536 7941 -23519
rect 7975 -23536 8009 -23502
rect 8043 -23536 8077 -23502
rect 8111 -23536 8145 -23502
rect 8179 -23536 8213 -23502
rect 8247 -23536 8281 -23502
rect 8315 -23536 8349 -23502
rect 8383 -23536 8417 -23502
rect 8451 -23519 8676 -23502
rect 8734 -23502 9694 -23464
rect 8734 -23519 8959 -23502
rect 8451 -23536 8490 -23519
rect 7902 -23552 8490 -23536
rect 8920 -23536 8959 -23519
rect 8993 -23536 9027 -23502
rect 9061 -23536 9095 -23502
rect 9129 -23536 9163 -23502
rect 9197 -23536 9231 -23502
rect 9265 -23536 9299 -23502
rect 9333 -23536 9367 -23502
rect 9401 -23536 9435 -23502
rect 9469 -23519 9694 -23502
rect 9752 -23502 10712 -23464
rect 9752 -23519 9977 -23502
rect 9469 -23536 9508 -23519
rect 8920 -23552 9508 -23536
rect 9938 -23536 9977 -23519
rect 10011 -23536 10045 -23502
rect 10079 -23536 10113 -23502
rect 10147 -23536 10181 -23502
rect 10215 -23536 10249 -23502
rect 10283 -23536 10317 -23502
rect 10351 -23536 10385 -23502
rect 10419 -23536 10453 -23502
rect 10487 -23519 10712 -23502
rect 10770 -23502 11730 -23464
rect 10770 -23519 10995 -23502
rect 10487 -23536 10526 -23519
rect 9938 -23552 10526 -23536
rect 10956 -23536 10995 -23519
rect 11029 -23536 11063 -23502
rect 11097 -23536 11131 -23502
rect 11165 -23536 11199 -23502
rect 11233 -23536 11267 -23502
rect 11301 -23536 11335 -23502
rect 11369 -23536 11403 -23502
rect 11437 -23536 11471 -23502
rect 11505 -23519 11730 -23502
rect 11788 -23502 12748 -23464
rect 11788 -23519 12013 -23502
rect 11505 -23536 11544 -23519
rect 10956 -23552 11544 -23536
rect 11974 -23536 12013 -23519
rect 12047 -23536 12081 -23502
rect 12115 -23536 12149 -23502
rect 12183 -23536 12217 -23502
rect 12251 -23536 12285 -23502
rect 12319 -23536 12353 -23502
rect 12387 -23536 12421 -23502
rect 12455 -23536 12489 -23502
rect 12523 -23519 12748 -23502
rect 12806 -23502 13766 -23464
rect 12806 -23519 13031 -23502
rect 12523 -23536 12562 -23519
rect 11974 -23552 12562 -23536
rect 12992 -23536 13031 -23519
rect 13065 -23536 13099 -23502
rect 13133 -23536 13167 -23502
rect 13201 -23536 13235 -23502
rect 13269 -23536 13303 -23502
rect 13337 -23536 13371 -23502
rect 13405 -23536 13439 -23502
rect 13473 -23536 13507 -23502
rect 13541 -23519 13766 -23502
rect 13824 -23502 14784 -23464
rect 13824 -23519 14049 -23502
rect 13541 -23536 13580 -23519
rect 12992 -23552 13580 -23536
rect 14010 -23536 14049 -23519
rect 14083 -23536 14117 -23502
rect 14151 -23536 14185 -23502
rect 14219 -23536 14253 -23502
rect 14287 -23536 14321 -23502
rect 14355 -23536 14389 -23502
rect 14423 -23536 14457 -23502
rect 14491 -23536 14525 -23502
rect 14559 -23519 14784 -23502
rect 14842 -23502 15802 -23464
rect 14842 -23519 15067 -23502
rect 14559 -23536 14598 -23519
rect 14010 -23552 14598 -23536
rect 15028 -23536 15067 -23519
rect 15101 -23536 15135 -23502
rect 15169 -23536 15203 -23502
rect 15237 -23536 15271 -23502
rect 15305 -23536 15339 -23502
rect 15373 -23536 15407 -23502
rect 15441 -23536 15475 -23502
rect 15509 -23536 15543 -23502
rect 15577 -23519 15802 -23502
rect 15860 -23502 16820 -23464
rect 15860 -23519 16085 -23502
rect 15577 -23536 15616 -23519
rect 15028 -23552 15616 -23536
rect 16046 -23536 16085 -23519
rect 16119 -23536 16153 -23502
rect 16187 -23536 16221 -23502
rect 16255 -23536 16289 -23502
rect 16323 -23536 16357 -23502
rect 16391 -23536 16425 -23502
rect 16459 -23536 16493 -23502
rect 16527 -23536 16561 -23502
rect 16595 -23519 16820 -23502
rect 16878 -23502 17838 -23464
rect 16878 -23519 17103 -23502
rect 16595 -23536 16634 -23519
rect 16046 -23552 16634 -23536
rect 17064 -23536 17103 -23519
rect 17137 -23536 17171 -23502
rect 17205 -23536 17239 -23502
rect 17273 -23536 17307 -23502
rect 17341 -23536 17375 -23502
rect 17409 -23536 17443 -23502
rect 17477 -23536 17511 -23502
rect 17545 -23536 17579 -23502
rect 17613 -23519 17838 -23502
rect 17896 -23502 18856 -23464
rect 17896 -23519 18121 -23502
rect 17613 -23536 17652 -23519
rect 17064 -23552 17652 -23536
rect 18082 -23536 18121 -23519
rect 18155 -23536 18189 -23502
rect 18223 -23536 18257 -23502
rect 18291 -23536 18325 -23502
rect 18359 -23536 18393 -23502
rect 18427 -23536 18461 -23502
rect 18495 -23536 18529 -23502
rect 18563 -23536 18597 -23502
rect 18631 -23519 18856 -23502
rect 18914 -23502 19874 -23464
rect 18914 -23519 19139 -23502
rect 18631 -23536 18670 -23519
rect 18082 -23552 18670 -23536
rect 19100 -23536 19139 -23519
rect 19173 -23536 19207 -23502
rect 19241 -23536 19275 -23502
rect 19309 -23536 19343 -23502
rect 19377 -23536 19411 -23502
rect 19445 -23536 19479 -23502
rect 19513 -23536 19547 -23502
rect 19581 -23536 19615 -23502
rect 19649 -23519 19874 -23502
rect 19932 -23502 20892 -23464
rect 19932 -23519 20157 -23502
rect 19649 -23536 19688 -23519
rect 19100 -23552 19688 -23536
rect 20118 -23536 20157 -23519
rect 20191 -23536 20225 -23502
rect 20259 -23536 20293 -23502
rect 20327 -23536 20361 -23502
rect 20395 -23536 20429 -23502
rect 20463 -23536 20497 -23502
rect 20531 -23536 20565 -23502
rect 20599 -23536 20633 -23502
rect 20667 -23519 20892 -23502
rect 20950 -23502 21910 -23464
rect 20950 -23519 21175 -23502
rect 20667 -23536 20706 -23519
rect 20118 -23552 20706 -23536
rect 21136 -23536 21175 -23519
rect 21209 -23536 21243 -23502
rect 21277 -23536 21311 -23502
rect 21345 -23536 21379 -23502
rect 21413 -23536 21447 -23502
rect 21481 -23536 21515 -23502
rect 21549 -23536 21583 -23502
rect 21617 -23536 21651 -23502
rect 21685 -23519 21910 -23502
rect 21968 -23502 22928 -23464
rect 21968 -23519 22193 -23502
rect 21685 -23536 21724 -23519
rect 21136 -23552 21724 -23536
rect 22154 -23536 22193 -23519
rect 22227 -23536 22261 -23502
rect 22295 -23536 22329 -23502
rect 22363 -23536 22397 -23502
rect 22431 -23536 22465 -23502
rect 22499 -23536 22533 -23502
rect 22567 -23536 22601 -23502
rect 22635 -23536 22669 -23502
rect 22703 -23519 22928 -23502
rect 22703 -23536 22742 -23519
rect 22154 -23552 22742 -23536
rect 2812 -24026 3400 -24010
rect 2812 -24043 2851 -24026
rect 2626 -24060 2851 -24043
rect 2885 -24060 2919 -24026
rect 2953 -24060 2987 -24026
rect 3021 -24060 3055 -24026
rect 3089 -24060 3123 -24026
rect 3157 -24060 3191 -24026
rect 3225 -24060 3259 -24026
rect 3293 -24060 3327 -24026
rect 3361 -24043 3400 -24026
rect 3830 -24026 4418 -24010
rect 3830 -24043 3869 -24026
rect 3361 -24060 3586 -24043
rect 2626 -24098 3586 -24060
rect 3644 -24060 3869 -24043
rect 3903 -24060 3937 -24026
rect 3971 -24060 4005 -24026
rect 4039 -24060 4073 -24026
rect 4107 -24060 4141 -24026
rect 4175 -24060 4209 -24026
rect 4243 -24060 4277 -24026
rect 4311 -24060 4345 -24026
rect 4379 -24043 4418 -24026
rect 4848 -24026 5436 -24010
rect 4848 -24043 4887 -24026
rect 4379 -24060 4604 -24043
rect 3644 -24098 4604 -24060
rect 4662 -24060 4887 -24043
rect 4921 -24060 4955 -24026
rect 4989 -24060 5023 -24026
rect 5057 -24060 5091 -24026
rect 5125 -24060 5159 -24026
rect 5193 -24060 5227 -24026
rect 5261 -24060 5295 -24026
rect 5329 -24060 5363 -24026
rect 5397 -24043 5436 -24026
rect 5866 -24026 6454 -24010
rect 5866 -24043 5905 -24026
rect 5397 -24060 5622 -24043
rect 4662 -24098 5622 -24060
rect 5680 -24060 5905 -24043
rect 5939 -24060 5973 -24026
rect 6007 -24060 6041 -24026
rect 6075 -24060 6109 -24026
rect 6143 -24060 6177 -24026
rect 6211 -24060 6245 -24026
rect 6279 -24060 6313 -24026
rect 6347 -24060 6381 -24026
rect 6415 -24043 6454 -24026
rect 6884 -24026 7472 -24010
rect 6884 -24043 6923 -24026
rect 6415 -24060 6640 -24043
rect 5680 -24098 6640 -24060
rect 6698 -24060 6923 -24043
rect 6957 -24060 6991 -24026
rect 7025 -24060 7059 -24026
rect 7093 -24060 7127 -24026
rect 7161 -24060 7195 -24026
rect 7229 -24060 7263 -24026
rect 7297 -24060 7331 -24026
rect 7365 -24060 7399 -24026
rect 7433 -24043 7472 -24026
rect 7902 -24026 8490 -24010
rect 7902 -24043 7941 -24026
rect 7433 -24060 7658 -24043
rect 6698 -24098 7658 -24060
rect 7716 -24060 7941 -24043
rect 7975 -24060 8009 -24026
rect 8043 -24060 8077 -24026
rect 8111 -24060 8145 -24026
rect 8179 -24060 8213 -24026
rect 8247 -24060 8281 -24026
rect 8315 -24060 8349 -24026
rect 8383 -24060 8417 -24026
rect 8451 -24043 8490 -24026
rect 8920 -24026 9508 -24010
rect 8920 -24043 8959 -24026
rect 8451 -24060 8676 -24043
rect 7716 -24098 8676 -24060
rect 8734 -24060 8959 -24043
rect 8993 -24060 9027 -24026
rect 9061 -24060 9095 -24026
rect 9129 -24060 9163 -24026
rect 9197 -24060 9231 -24026
rect 9265 -24060 9299 -24026
rect 9333 -24060 9367 -24026
rect 9401 -24060 9435 -24026
rect 9469 -24043 9508 -24026
rect 9938 -24026 10526 -24010
rect 9938 -24043 9977 -24026
rect 9469 -24060 9694 -24043
rect 8734 -24098 9694 -24060
rect 9752 -24060 9977 -24043
rect 10011 -24060 10045 -24026
rect 10079 -24060 10113 -24026
rect 10147 -24060 10181 -24026
rect 10215 -24060 10249 -24026
rect 10283 -24060 10317 -24026
rect 10351 -24060 10385 -24026
rect 10419 -24060 10453 -24026
rect 10487 -24043 10526 -24026
rect 10956 -24026 11544 -24010
rect 10956 -24043 10995 -24026
rect 10487 -24060 10712 -24043
rect 9752 -24098 10712 -24060
rect 10770 -24060 10995 -24043
rect 11029 -24060 11063 -24026
rect 11097 -24060 11131 -24026
rect 11165 -24060 11199 -24026
rect 11233 -24060 11267 -24026
rect 11301 -24060 11335 -24026
rect 11369 -24060 11403 -24026
rect 11437 -24060 11471 -24026
rect 11505 -24043 11544 -24026
rect 11974 -24026 12562 -24010
rect 11974 -24043 12013 -24026
rect 11505 -24060 11730 -24043
rect 10770 -24098 11730 -24060
rect 11788 -24060 12013 -24043
rect 12047 -24060 12081 -24026
rect 12115 -24060 12149 -24026
rect 12183 -24060 12217 -24026
rect 12251 -24060 12285 -24026
rect 12319 -24060 12353 -24026
rect 12387 -24060 12421 -24026
rect 12455 -24060 12489 -24026
rect 12523 -24043 12562 -24026
rect 12992 -24026 13580 -24010
rect 12992 -24043 13031 -24026
rect 12523 -24060 12748 -24043
rect 11788 -24098 12748 -24060
rect 12806 -24060 13031 -24043
rect 13065 -24060 13099 -24026
rect 13133 -24060 13167 -24026
rect 13201 -24060 13235 -24026
rect 13269 -24060 13303 -24026
rect 13337 -24060 13371 -24026
rect 13405 -24060 13439 -24026
rect 13473 -24060 13507 -24026
rect 13541 -24043 13580 -24026
rect 14010 -24026 14598 -24010
rect 14010 -24043 14049 -24026
rect 13541 -24060 13766 -24043
rect 12806 -24098 13766 -24060
rect 13824 -24060 14049 -24043
rect 14083 -24060 14117 -24026
rect 14151 -24060 14185 -24026
rect 14219 -24060 14253 -24026
rect 14287 -24060 14321 -24026
rect 14355 -24060 14389 -24026
rect 14423 -24060 14457 -24026
rect 14491 -24060 14525 -24026
rect 14559 -24043 14598 -24026
rect 15028 -24026 15616 -24010
rect 15028 -24043 15067 -24026
rect 14559 -24060 14784 -24043
rect 13824 -24098 14784 -24060
rect 14842 -24060 15067 -24043
rect 15101 -24060 15135 -24026
rect 15169 -24060 15203 -24026
rect 15237 -24060 15271 -24026
rect 15305 -24060 15339 -24026
rect 15373 -24060 15407 -24026
rect 15441 -24060 15475 -24026
rect 15509 -24060 15543 -24026
rect 15577 -24043 15616 -24026
rect 16046 -24026 16634 -24010
rect 16046 -24043 16085 -24026
rect 15577 -24060 15802 -24043
rect 14842 -24098 15802 -24060
rect 15860 -24060 16085 -24043
rect 16119 -24060 16153 -24026
rect 16187 -24060 16221 -24026
rect 16255 -24060 16289 -24026
rect 16323 -24060 16357 -24026
rect 16391 -24060 16425 -24026
rect 16459 -24060 16493 -24026
rect 16527 -24060 16561 -24026
rect 16595 -24043 16634 -24026
rect 17064 -24026 17652 -24010
rect 17064 -24043 17103 -24026
rect 16595 -24060 16820 -24043
rect 15860 -24098 16820 -24060
rect 16878 -24060 17103 -24043
rect 17137 -24060 17171 -24026
rect 17205 -24060 17239 -24026
rect 17273 -24060 17307 -24026
rect 17341 -24060 17375 -24026
rect 17409 -24060 17443 -24026
rect 17477 -24060 17511 -24026
rect 17545 -24060 17579 -24026
rect 17613 -24043 17652 -24026
rect 18082 -24026 18670 -24010
rect 18082 -24043 18121 -24026
rect 17613 -24060 17838 -24043
rect 16878 -24098 17838 -24060
rect 17896 -24060 18121 -24043
rect 18155 -24060 18189 -24026
rect 18223 -24060 18257 -24026
rect 18291 -24060 18325 -24026
rect 18359 -24060 18393 -24026
rect 18427 -24060 18461 -24026
rect 18495 -24060 18529 -24026
rect 18563 -24060 18597 -24026
rect 18631 -24043 18670 -24026
rect 19100 -24026 19688 -24010
rect 19100 -24043 19139 -24026
rect 18631 -24060 18856 -24043
rect 17896 -24098 18856 -24060
rect 18914 -24060 19139 -24043
rect 19173 -24060 19207 -24026
rect 19241 -24060 19275 -24026
rect 19309 -24060 19343 -24026
rect 19377 -24060 19411 -24026
rect 19445 -24060 19479 -24026
rect 19513 -24060 19547 -24026
rect 19581 -24060 19615 -24026
rect 19649 -24043 19688 -24026
rect 20118 -24026 20706 -24010
rect 20118 -24043 20157 -24026
rect 19649 -24060 19874 -24043
rect 18914 -24098 19874 -24060
rect 19932 -24060 20157 -24043
rect 20191 -24060 20225 -24026
rect 20259 -24060 20293 -24026
rect 20327 -24060 20361 -24026
rect 20395 -24060 20429 -24026
rect 20463 -24060 20497 -24026
rect 20531 -24060 20565 -24026
rect 20599 -24060 20633 -24026
rect 20667 -24043 20706 -24026
rect 21136 -24026 21724 -24010
rect 21136 -24043 21175 -24026
rect 20667 -24060 20892 -24043
rect 19932 -24098 20892 -24060
rect 20950 -24060 21175 -24043
rect 21209 -24060 21243 -24026
rect 21277 -24060 21311 -24026
rect 21345 -24060 21379 -24026
rect 21413 -24060 21447 -24026
rect 21481 -24060 21515 -24026
rect 21549 -24060 21583 -24026
rect 21617 -24060 21651 -24026
rect 21685 -24043 21724 -24026
rect 22154 -24026 22742 -24010
rect 22154 -24043 22193 -24026
rect 21685 -24060 21910 -24043
rect 20950 -24098 21910 -24060
rect 21968 -24060 22193 -24043
rect 22227 -24060 22261 -24026
rect 22295 -24060 22329 -24026
rect 22363 -24060 22397 -24026
rect 22431 -24060 22465 -24026
rect 22499 -24060 22533 -24026
rect 22567 -24060 22601 -24026
rect 22635 -24060 22669 -24026
rect 22703 -24043 22742 -24026
rect 22703 -24060 22928 -24043
rect 21968 -24098 22928 -24060
rect 2626 -24736 3586 -24698
rect 2626 -24753 2851 -24736
rect 2812 -24770 2851 -24753
rect 2885 -24770 2919 -24736
rect 2953 -24770 2987 -24736
rect 3021 -24770 3055 -24736
rect 3089 -24770 3123 -24736
rect 3157 -24770 3191 -24736
rect 3225 -24770 3259 -24736
rect 3293 -24770 3327 -24736
rect 3361 -24753 3586 -24736
rect 3644 -24736 4604 -24698
rect 3644 -24753 3869 -24736
rect 3361 -24770 3400 -24753
rect 2812 -24786 3400 -24770
rect 3830 -24770 3869 -24753
rect 3903 -24770 3937 -24736
rect 3971 -24770 4005 -24736
rect 4039 -24770 4073 -24736
rect 4107 -24770 4141 -24736
rect 4175 -24770 4209 -24736
rect 4243 -24770 4277 -24736
rect 4311 -24770 4345 -24736
rect 4379 -24753 4604 -24736
rect 4662 -24736 5622 -24698
rect 4662 -24753 4887 -24736
rect 4379 -24770 4418 -24753
rect 3830 -24786 4418 -24770
rect 4848 -24770 4887 -24753
rect 4921 -24770 4955 -24736
rect 4989 -24770 5023 -24736
rect 5057 -24770 5091 -24736
rect 5125 -24770 5159 -24736
rect 5193 -24770 5227 -24736
rect 5261 -24770 5295 -24736
rect 5329 -24770 5363 -24736
rect 5397 -24753 5622 -24736
rect 5680 -24736 6640 -24698
rect 5680 -24753 5905 -24736
rect 5397 -24770 5436 -24753
rect 4848 -24786 5436 -24770
rect 5866 -24770 5905 -24753
rect 5939 -24770 5973 -24736
rect 6007 -24770 6041 -24736
rect 6075 -24770 6109 -24736
rect 6143 -24770 6177 -24736
rect 6211 -24770 6245 -24736
rect 6279 -24770 6313 -24736
rect 6347 -24770 6381 -24736
rect 6415 -24753 6640 -24736
rect 6698 -24736 7658 -24698
rect 6698 -24753 6923 -24736
rect 6415 -24770 6454 -24753
rect 5866 -24786 6454 -24770
rect 6884 -24770 6923 -24753
rect 6957 -24770 6991 -24736
rect 7025 -24770 7059 -24736
rect 7093 -24770 7127 -24736
rect 7161 -24770 7195 -24736
rect 7229 -24770 7263 -24736
rect 7297 -24770 7331 -24736
rect 7365 -24770 7399 -24736
rect 7433 -24753 7658 -24736
rect 7716 -24736 8676 -24698
rect 7716 -24753 7941 -24736
rect 7433 -24770 7472 -24753
rect 6884 -24786 7472 -24770
rect 7902 -24770 7941 -24753
rect 7975 -24770 8009 -24736
rect 8043 -24770 8077 -24736
rect 8111 -24770 8145 -24736
rect 8179 -24770 8213 -24736
rect 8247 -24770 8281 -24736
rect 8315 -24770 8349 -24736
rect 8383 -24770 8417 -24736
rect 8451 -24753 8676 -24736
rect 8734 -24736 9694 -24698
rect 8734 -24753 8959 -24736
rect 8451 -24770 8490 -24753
rect 7902 -24786 8490 -24770
rect 8920 -24770 8959 -24753
rect 8993 -24770 9027 -24736
rect 9061 -24770 9095 -24736
rect 9129 -24770 9163 -24736
rect 9197 -24770 9231 -24736
rect 9265 -24770 9299 -24736
rect 9333 -24770 9367 -24736
rect 9401 -24770 9435 -24736
rect 9469 -24753 9694 -24736
rect 9752 -24736 10712 -24698
rect 9752 -24753 9977 -24736
rect 9469 -24770 9508 -24753
rect 8920 -24786 9508 -24770
rect 9938 -24770 9977 -24753
rect 10011 -24770 10045 -24736
rect 10079 -24770 10113 -24736
rect 10147 -24770 10181 -24736
rect 10215 -24770 10249 -24736
rect 10283 -24770 10317 -24736
rect 10351 -24770 10385 -24736
rect 10419 -24770 10453 -24736
rect 10487 -24753 10712 -24736
rect 10770 -24736 11730 -24698
rect 10770 -24753 10995 -24736
rect 10487 -24770 10526 -24753
rect 9938 -24786 10526 -24770
rect 10956 -24770 10995 -24753
rect 11029 -24770 11063 -24736
rect 11097 -24770 11131 -24736
rect 11165 -24770 11199 -24736
rect 11233 -24770 11267 -24736
rect 11301 -24770 11335 -24736
rect 11369 -24770 11403 -24736
rect 11437 -24770 11471 -24736
rect 11505 -24753 11730 -24736
rect 11788 -24736 12748 -24698
rect 11788 -24753 12013 -24736
rect 11505 -24770 11544 -24753
rect 10956 -24786 11544 -24770
rect 11974 -24770 12013 -24753
rect 12047 -24770 12081 -24736
rect 12115 -24770 12149 -24736
rect 12183 -24770 12217 -24736
rect 12251 -24770 12285 -24736
rect 12319 -24770 12353 -24736
rect 12387 -24770 12421 -24736
rect 12455 -24770 12489 -24736
rect 12523 -24753 12748 -24736
rect 12806 -24736 13766 -24698
rect 12806 -24753 13031 -24736
rect 12523 -24770 12562 -24753
rect 11974 -24786 12562 -24770
rect 12992 -24770 13031 -24753
rect 13065 -24770 13099 -24736
rect 13133 -24770 13167 -24736
rect 13201 -24770 13235 -24736
rect 13269 -24770 13303 -24736
rect 13337 -24770 13371 -24736
rect 13405 -24770 13439 -24736
rect 13473 -24770 13507 -24736
rect 13541 -24753 13766 -24736
rect 13824 -24736 14784 -24698
rect 13824 -24753 14049 -24736
rect 13541 -24770 13580 -24753
rect 12992 -24786 13580 -24770
rect 14010 -24770 14049 -24753
rect 14083 -24770 14117 -24736
rect 14151 -24770 14185 -24736
rect 14219 -24770 14253 -24736
rect 14287 -24770 14321 -24736
rect 14355 -24770 14389 -24736
rect 14423 -24770 14457 -24736
rect 14491 -24770 14525 -24736
rect 14559 -24753 14784 -24736
rect 14842 -24736 15802 -24698
rect 14842 -24753 15067 -24736
rect 14559 -24770 14598 -24753
rect 14010 -24786 14598 -24770
rect 15028 -24770 15067 -24753
rect 15101 -24770 15135 -24736
rect 15169 -24770 15203 -24736
rect 15237 -24770 15271 -24736
rect 15305 -24770 15339 -24736
rect 15373 -24770 15407 -24736
rect 15441 -24770 15475 -24736
rect 15509 -24770 15543 -24736
rect 15577 -24753 15802 -24736
rect 15860 -24736 16820 -24698
rect 15860 -24753 16085 -24736
rect 15577 -24770 15616 -24753
rect 15028 -24786 15616 -24770
rect 16046 -24770 16085 -24753
rect 16119 -24770 16153 -24736
rect 16187 -24770 16221 -24736
rect 16255 -24770 16289 -24736
rect 16323 -24770 16357 -24736
rect 16391 -24770 16425 -24736
rect 16459 -24770 16493 -24736
rect 16527 -24770 16561 -24736
rect 16595 -24753 16820 -24736
rect 16878 -24736 17838 -24698
rect 16878 -24753 17103 -24736
rect 16595 -24770 16634 -24753
rect 16046 -24786 16634 -24770
rect 17064 -24770 17103 -24753
rect 17137 -24770 17171 -24736
rect 17205 -24770 17239 -24736
rect 17273 -24770 17307 -24736
rect 17341 -24770 17375 -24736
rect 17409 -24770 17443 -24736
rect 17477 -24770 17511 -24736
rect 17545 -24770 17579 -24736
rect 17613 -24753 17838 -24736
rect 17896 -24736 18856 -24698
rect 17896 -24753 18121 -24736
rect 17613 -24770 17652 -24753
rect 17064 -24786 17652 -24770
rect 18082 -24770 18121 -24753
rect 18155 -24770 18189 -24736
rect 18223 -24770 18257 -24736
rect 18291 -24770 18325 -24736
rect 18359 -24770 18393 -24736
rect 18427 -24770 18461 -24736
rect 18495 -24770 18529 -24736
rect 18563 -24770 18597 -24736
rect 18631 -24753 18856 -24736
rect 18914 -24736 19874 -24698
rect 18914 -24753 19139 -24736
rect 18631 -24770 18670 -24753
rect 18082 -24786 18670 -24770
rect 19100 -24770 19139 -24753
rect 19173 -24770 19207 -24736
rect 19241 -24770 19275 -24736
rect 19309 -24770 19343 -24736
rect 19377 -24770 19411 -24736
rect 19445 -24770 19479 -24736
rect 19513 -24770 19547 -24736
rect 19581 -24770 19615 -24736
rect 19649 -24753 19874 -24736
rect 19932 -24736 20892 -24698
rect 19932 -24753 20157 -24736
rect 19649 -24770 19688 -24753
rect 19100 -24786 19688 -24770
rect 20118 -24770 20157 -24753
rect 20191 -24770 20225 -24736
rect 20259 -24770 20293 -24736
rect 20327 -24770 20361 -24736
rect 20395 -24770 20429 -24736
rect 20463 -24770 20497 -24736
rect 20531 -24770 20565 -24736
rect 20599 -24770 20633 -24736
rect 20667 -24753 20892 -24736
rect 20950 -24736 21910 -24698
rect 20950 -24753 21175 -24736
rect 20667 -24770 20706 -24753
rect 20118 -24786 20706 -24770
rect 21136 -24770 21175 -24753
rect 21209 -24770 21243 -24736
rect 21277 -24770 21311 -24736
rect 21345 -24770 21379 -24736
rect 21413 -24770 21447 -24736
rect 21481 -24770 21515 -24736
rect 21549 -24770 21583 -24736
rect 21617 -24770 21651 -24736
rect 21685 -24753 21910 -24736
rect 21968 -24736 22928 -24698
rect 21968 -24753 22193 -24736
rect 21685 -24770 21724 -24753
rect 21136 -24786 21724 -24770
rect 22154 -24770 22193 -24753
rect 22227 -24770 22261 -24736
rect 22295 -24770 22329 -24736
rect 22363 -24770 22397 -24736
rect 22431 -24770 22465 -24736
rect 22499 -24770 22533 -24736
rect 22567 -24770 22601 -24736
rect 22635 -24770 22669 -24736
rect 22703 -24753 22928 -24736
rect 22703 -24770 22742 -24753
rect 22154 -24786 22742 -24770
<< polycont >>
rect -8913 -12474 -8879 -12440
rect -8845 -12474 -8811 -12440
rect -8777 -12474 -8743 -12440
rect -8709 -12474 -8675 -12440
rect -8641 -12474 -8607 -12440
rect -8573 -12474 -8539 -12440
rect -8505 -12474 -8471 -12440
rect -8437 -12474 -8403 -12440
rect -7895 -12474 -7861 -12440
rect -7827 -12474 -7793 -12440
rect -7759 -12474 -7725 -12440
rect -7691 -12474 -7657 -12440
rect -7623 -12474 -7589 -12440
rect -7555 -12474 -7521 -12440
rect -7487 -12474 -7453 -12440
rect -7419 -12474 -7385 -12440
rect -6877 -12474 -6843 -12440
rect -6809 -12474 -6775 -12440
rect -6741 -12474 -6707 -12440
rect -6673 -12474 -6639 -12440
rect -6605 -12474 -6571 -12440
rect -6537 -12474 -6503 -12440
rect -6469 -12474 -6435 -12440
rect -6401 -12474 -6367 -12440
rect -5859 -12474 -5825 -12440
rect -5791 -12474 -5757 -12440
rect -5723 -12474 -5689 -12440
rect -5655 -12474 -5621 -12440
rect -5587 -12474 -5553 -12440
rect -5519 -12474 -5485 -12440
rect -5451 -12474 -5417 -12440
rect -5383 -12474 -5349 -12440
rect -4841 -12474 -4807 -12440
rect -4773 -12474 -4739 -12440
rect -4705 -12474 -4671 -12440
rect -4637 -12474 -4603 -12440
rect -4569 -12474 -4535 -12440
rect -4501 -12474 -4467 -12440
rect -4433 -12474 -4399 -12440
rect -4365 -12474 -4331 -12440
rect -3823 -12474 -3789 -12440
rect -3755 -12474 -3721 -12440
rect -3687 -12474 -3653 -12440
rect -3619 -12474 -3585 -12440
rect -3551 -12474 -3517 -12440
rect -3483 -12474 -3449 -12440
rect -3415 -12474 -3381 -12440
rect -3347 -12474 -3313 -12440
rect -2805 -12474 -2771 -12440
rect -2737 -12474 -2703 -12440
rect -2669 -12474 -2635 -12440
rect -2601 -12474 -2567 -12440
rect -2533 -12474 -2499 -12440
rect -2465 -12474 -2431 -12440
rect -2397 -12474 -2363 -12440
rect -2329 -12474 -2295 -12440
rect -1787 -12474 -1753 -12440
rect -1719 -12474 -1685 -12440
rect -1651 -12474 -1617 -12440
rect -1583 -12474 -1549 -12440
rect -1515 -12474 -1481 -12440
rect -1447 -12474 -1413 -12440
rect -1379 -12474 -1345 -12440
rect -1311 -12474 -1277 -12440
rect -769 -12474 -735 -12440
rect -701 -12474 -667 -12440
rect -633 -12474 -599 -12440
rect -565 -12474 -531 -12440
rect -497 -12474 -463 -12440
rect -429 -12474 -395 -12440
rect -361 -12474 -327 -12440
rect -293 -12474 -259 -12440
rect -8913 -13184 -8879 -13150
rect -8845 -13184 -8811 -13150
rect -8777 -13184 -8743 -13150
rect -8709 -13184 -8675 -13150
rect -8641 -13184 -8607 -13150
rect -8573 -13184 -8539 -13150
rect -8505 -13184 -8471 -13150
rect -8437 -13184 -8403 -13150
rect -7895 -13184 -7861 -13150
rect -7827 -13184 -7793 -13150
rect -7759 -13184 -7725 -13150
rect -7691 -13184 -7657 -13150
rect -7623 -13184 -7589 -13150
rect -7555 -13184 -7521 -13150
rect -7487 -13184 -7453 -13150
rect -7419 -13184 -7385 -13150
rect -6877 -13184 -6843 -13150
rect -6809 -13184 -6775 -13150
rect -6741 -13184 -6707 -13150
rect -6673 -13184 -6639 -13150
rect -6605 -13184 -6571 -13150
rect -6537 -13184 -6503 -13150
rect -6469 -13184 -6435 -13150
rect -6401 -13184 -6367 -13150
rect -5859 -13184 -5825 -13150
rect -5791 -13184 -5757 -13150
rect -5723 -13184 -5689 -13150
rect -5655 -13184 -5621 -13150
rect -5587 -13184 -5553 -13150
rect -5519 -13184 -5485 -13150
rect -5451 -13184 -5417 -13150
rect -5383 -13184 -5349 -13150
rect -4841 -13184 -4807 -13150
rect -4773 -13184 -4739 -13150
rect -4705 -13184 -4671 -13150
rect -4637 -13184 -4603 -13150
rect -4569 -13184 -4535 -13150
rect -4501 -13184 -4467 -13150
rect -4433 -13184 -4399 -13150
rect -4365 -13184 -4331 -13150
rect -3823 -13184 -3789 -13150
rect -3755 -13184 -3721 -13150
rect -3687 -13184 -3653 -13150
rect -3619 -13184 -3585 -13150
rect -3551 -13184 -3517 -13150
rect -3483 -13184 -3449 -13150
rect -3415 -13184 -3381 -13150
rect -3347 -13184 -3313 -13150
rect -2805 -13184 -2771 -13150
rect -2737 -13184 -2703 -13150
rect -2669 -13184 -2635 -13150
rect -2601 -13184 -2567 -13150
rect -2533 -13184 -2499 -13150
rect -2465 -13184 -2431 -13150
rect -2397 -13184 -2363 -13150
rect -2329 -13184 -2295 -13150
rect -1787 -13184 -1753 -13150
rect -1719 -13184 -1685 -13150
rect -1651 -13184 -1617 -13150
rect -1583 -13184 -1549 -13150
rect -1515 -13184 -1481 -13150
rect -1447 -13184 -1413 -13150
rect -1379 -13184 -1345 -13150
rect -1311 -13184 -1277 -13150
rect -769 -13184 -735 -13150
rect -701 -13184 -667 -13150
rect -633 -13184 -599 -13150
rect -565 -13184 -531 -13150
rect -497 -13184 -463 -13150
rect -429 -13184 -395 -13150
rect -361 -13184 -327 -13150
rect -293 -13184 -259 -13150
rect -8913 -13292 -8879 -13258
rect -8845 -13292 -8811 -13258
rect -8777 -13292 -8743 -13258
rect -8709 -13292 -8675 -13258
rect -8641 -13292 -8607 -13258
rect -8573 -13292 -8539 -13258
rect -8505 -13292 -8471 -13258
rect -8437 -13292 -8403 -13258
rect -7895 -13292 -7861 -13258
rect -7827 -13292 -7793 -13258
rect -7759 -13292 -7725 -13258
rect -7691 -13292 -7657 -13258
rect -7623 -13292 -7589 -13258
rect -7555 -13292 -7521 -13258
rect -7487 -13292 -7453 -13258
rect -7419 -13292 -7385 -13258
rect -6877 -13292 -6843 -13258
rect -6809 -13292 -6775 -13258
rect -6741 -13292 -6707 -13258
rect -6673 -13292 -6639 -13258
rect -6605 -13292 -6571 -13258
rect -6537 -13292 -6503 -13258
rect -6469 -13292 -6435 -13258
rect -6401 -13292 -6367 -13258
rect -5859 -13292 -5825 -13258
rect -5791 -13292 -5757 -13258
rect -5723 -13292 -5689 -13258
rect -5655 -13292 -5621 -13258
rect -5587 -13292 -5553 -13258
rect -5519 -13292 -5485 -13258
rect -5451 -13292 -5417 -13258
rect -5383 -13292 -5349 -13258
rect -4841 -13292 -4807 -13258
rect -4773 -13292 -4739 -13258
rect -4705 -13292 -4671 -13258
rect -4637 -13292 -4603 -13258
rect -4569 -13292 -4535 -13258
rect -4501 -13292 -4467 -13258
rect -4433 -13292 -4399 -13258
rect -4365 -13292 -4331 -13258
rect -3823 -13292 -3789 -13258
rect -3755 -13292 -3721 -13258
rect -3687 -13292 -3653 -13258
rect -3619 -13292 -3585 -13258
rect -3551 -13292 -3517 -13258
rect -3483 -13292 -3449 -13258
rect -3415 -13292 -3381 -13258
rect -3347 -13292 -3313 -13258
rect -2805 -13292 -2771 -13258
rect -2737 -13292 -2703 -13258
rect -2669 -13292 -2635 -13258
rect -2601 -13292 -2567 -13258
rect -2533 -13292 -2499 -13258
rect -2465 -13292 -2431 -13258
rect -2397 -13292 -2363 -13258
rect -2329 -13292 -2295 -13258
rect -1787 -13292 -1753 -13258
rect -1719 -13292 -1685 -13258
rect -1651 -13292 -1617 -13258
rect -1583 -13292 -1549 -13258
rect -1515 -13292 -1481 -13258
rect -1447 -13292 -1413 -13258
rect -1379 -13292 -1345 -13258
rect -1311 -13292 -1277 -13258
rect -769 -13292 -735 -13258
rect -701 -13292 -667 -13258
rect -633 -13292 -599 -13258
rect -565 -13292 -531 -13258
rect -497 -13292 -463 -13258
rect -429 -13292 -395 -13258
rect -361 -13292 -327 -13258
rect -293 -13292 -259 -13258
rect -8913 -14002 -8879 -13968
rect -8845 -14002 -8811 -13968
rect -8777 -14002 -8743 -13968
rect -8709 -14002 -8675 -13968
rect -8641 -14002 -8607 -13968
rect -8573 -14002 -8539 -13968
rect -8505 -14002 -8471 -13968
rect -8437 -14002 -8403 -13968
rect -7895 -14002 -7861 -13968
rect -7827 -14002 -7793 -13968
rect -7759 -14002 -7725 -13968
rect -7691 -14002 -7657 -13968
rect -7623 -14002 -7589 -13968
rect -7555 -14002 -7521 -13968
rect -7487 -14002 -7453 -13968
rect -7419 -14002 -7385 -13968
rect -6877 -14002 -6843 -13968
rect -6809 -14002 -6775 -13968
rect -6741 -14002 -6707 -13968
rect -6673 -14002 -6639 -13968
rect -6605 -14002 -6571 -13968
rect -6537 -14002 -6503 -13968
rect -6469 -14002 -6435 -13968
rect -6401 -14002 -6367 -13968
rect -5859 -14002 -5825 -13968
rect -5791 -14002 -5757 -13968
rect -5723 -14002 -5689 -13968
rect -5655 -14002 -5621 -13968
rect -5587 -14002 -5553 -13968
rect -5519 -14002 -5485 -13968
rect -5451 -14002 -5417 -13968
rect -5383 -14002 -5349 -13968
rect -4841 -14002 -4807 -13968
rect -4773 -14002 -4739 -13968
rect -4705 -14002 -4671 -13968
rect -4637 -14002 -4603 -13968
rect -4569 -14002 -4535 -13968
rect -4501 -14002 -4467 -13968
rect -4433 -14002 -4399 -13968
rect -4365 -14002 -4331 -13968
rect -3823 -14002 -3789 -13968
rect -3755 -14002 -3721 -13968
rect -3687 -14002 -3653 -13968
rect -3619 -14002 -3585 -13968
rect -3551 -14002 -3517 -13968
rect -3483 -14002 -3449 -13968
rect -3415 -14002 -3381 -13968
rect -3347 -14002 -3313 -13968
rect -2805 -14002 -2771 -13968
rect -2737 -14002 -2703 -13968
rect -2669 -14002 -2635 -13968
rect -2601 -14002 -2567 -13968
rect -2533 -14002 -2499 -13968
rect -2465 -14002 -2431 -13968
rect -2397 -14002 -2363 -13968
rect -2329 -14002 -2295 -13968
rect -1787 -14002 -1753 -13968
rect -1719 -14002 -1685 -13968
rect -1651 -14002 -1617 -13968
rect -1583 -14002 -1549 -13968
rect -1515 -14002 -1481 -13968
rect -1447 -14002 -1413 -13968
rect -1379 -14002 -1345 -13968
rect -1311 -14002 -1277 -13968
rect -769 -14002 -735 -13968
rect -701 -14002 -667 -13968
rect -633 -14002 -599 -13968
rect -565 -14002 -531 -13968
rect -497 -14002 -463 -13968
rect -429 -14002 -395 -13968
rect -361 -14002 -327 -13968
rect -293 -14002 -259 -13968
rect -8913 -14110 -8879 -14076
rect -8845 -14110 -8811 -14076
rect -8777 -14110 -8743 -14076
rect -8709 -14110 -8675 -14076
rect -8641 -14110 -8607 -14076
rect -8573 -14110 -8539 -14076
rect -8505 -14110 -8471 -14076
rect -8437 -14110 -8403 -14076
rect -7895 -14110 -7861 -14076
rect -7827 -14110 -7793 -14076
rect -7759 -14110 -7725 -14076
rect -7691 -14110 -7657 -14076
rect -7623 -14110 -7589 -14076
rect -7555 -14110 -7521 -14076
rect -7487 -14110 -7453 -14076
rect -7419 -14110 -7385 -14076
rect -6877 -14110 -6843 -14076
rect -6809 -14110 -6775 -14076
rect -6741 -14110 -6707 -14076
rect -6673 -14110 -6639 -14076
rect -6605 -14110 -6571 -14076
rect -6537 -14110 -6503 -14076
rect -6469 -14110 -6435 -14076
rect -6401 -14110 -6367 -14076
rect -5859 -14110 -5825 -14076
rect -5791 -14110 -5757 -14076
rect -5723 -14110 -5689 -14076
rect -5655 -14110 -5621 -14076
rect -5587 -14110 -5553 -14076
rect -5519 -14110 -5485 -14076
rect -5451 -14110 -5417 -14076
rect -5383 -14110 -5349 -14076
rect -4841 -14110 -4807 -14076
rect -4773 -14110 -4739 -14076
rect -4705 -14110 -4671 -14076
rect -4637 -14110 -4603 -14076
rect -4569 -14110 -4535 -14076
rect -4501 -14110 -4467 -14076
rect -4433 -14110 -4399 -14076
rect -4365 -14110 -4331 -14076
rect -3823 -14110 -3789 -14076
rect -3755 -14110 -3721 -14076
rect -3687 -14110 -3653 -14076
rect -3619 -14110 -3585 -14076
rect -3551 -14110 -3517 -14076
rect -3483 -14110 -3449 -14076
rect -3415 -14110 -3381 -14076
rect -3347 -14110 -3313 -14076
rect -2805 -14110 -2771 -14076
rect -2737 -14110 -2703 -14076
rect -2669 -14110 -2635 -14076
rect -2601 -14110 -2567 -14076
rect -2533 -14110 -2499 -14076
rect -2465 -14110 -2431 -14076
rect -2397 -14110 -2363 -14076
rect -2329 -14110 -2295 -14076
rect -1787 -14110 -1753 -14076
rect -1719 -14110 -1685 -14076
rect -1651 -14110 -1617 -14076
rect -1583 -14110 -1549 -14076
rect -1515 -14110 -1481 -14076
rect -1447 -14110 -1413 -14076
rect -1379 -14110 -1345 -14076
rect -1311 -14110 -1277 -14076
rect -769 -14110 -735 -14076
rect -701 -14110 -667 -14076
rect -633 -14110 -599 -14076
rect -565 -14110 -531 -14076
rect -497 -14110 -463 -14076
rect -429 -14110 -395 -14076
rect -361 -14110 -327 -14076
rect -293 -14110 -259 -14076
rect 2853 -14194 2887 -14160
rect 2921 -14194 2955 -14160
rect 2989 -14194 3023 -14160
rect 3057 -14194 3091 -14160
rect 3125 -14194 3159 -14160
rect 3193 -14194 3227 -14160
rect 3261 -14194 3295 -14160
rect 3329 -14194 3363 -14160
rect 3871 -14194 3905 -14160
rect 3939 -14194 3973 -14160
rect 4007 -14194 4041 -14160
rect 4075 -14194 4109 -14160
rect 4143 -14194 4177 -14160
rect 4211 -14194 4245 -14160
rect 4279 -14194 4313 -14160
rect 4347 -14194 4381 -14160
rect 4889 -14194 4923 -14160
rect 4957 -14194 4991 -14160
rect 5025 -14194 5059 -14160
rect 5093 -14194 5127 -14160
rect 5161 -14194 5195 -14160
rect 5229 -14194 5263 -14160
rect 5297 -14194 5331 -14160
rect 5365 -14194 5399 -14160
rect 5907 -14194 5941 -14160
rect 5975 -14194 6009 -14160
rect 6043 -14194 6077 -14160
rect 6111 -14194 6145 -14160
rect 6179 -14194 6213 -14160
rect 6247 -14194 6281 -14160
rect 6315 -14194 6349 -14160
rect 6383 -14194 6417 -14160
rect 6925 -14194 6959 -14160
rect 6993 -14194 7027 -14160
rect 7061 -14194 7095 -14160
rect 7129 -14194 7163 -14160
rect 7197 -14194 7231 -14160
rect 7265 -14194 7299 -14160
rect 7333 -14194 7367 -14160
rect 7401 -14194 7435 -14160
rect 7943 -14194 7977 -14160
rect 8011 -14194 8045 -14160
rect 8079 -14194 8113 -14160
rect 8147 -14194 8181 -14160
rect 8215 -14194 8249 -14160
rect 8283 -14194 8317 -14160
rect 8351 -14194 8385 -14160
rect 8419 -14194 8453 -14160
rect 8961 -14194 8995 -14160
rect 9029 -14194 9063 -14160
rect 9097 -14194 9131 -14160
rect 9165 -14194 9199 -14160
rect 9233 -14194 9267 -14160
rect 9301 -14194 9335 -14160
rect 9369 -14194 9403 -14160
rect 9437 -14194 9471 -14160
rect 9979 -14194 10013 -14160
rect 10047 -14194 10081 -14160
rect 10115 -14194 10149 -14160
rect 10183 -14194 10217 -14160
rect 10251 -14194 10285 -14160
rect 10319 -14194 10353 -14160
rect 10387 -14194 10421 -14160
rect 10455 -14194 10489 -14160
rect 10997 -14194 11031 -14160
rect 11065 -14194 11099 -14160
rect 11133 -14194 11167 -14160
rect 11201 -14194 11235 -14160
rect 11269 -14194 11303 -14160
rect 11337 -14194 11371 -14160
rect 11405 -14194 11439 -14160
rect 11473 -14194 11507 -14160
rect 12015 -14194 12049 -14160
rect 12083 -14194 12117 -14160
rect 12151 -14194 12185 -14160
rect 12219 -14194 12253 -14160
rect 12287 -14194 12321 -14160
rect 12355 -14194 12389 -14160
rect 12423 -14194 12457 -14160
rect 12491 -14194 12525 -14160
rect 13033 -14194 13067 -14160
rect 13101 -14194 13135 -14160
rect 13169 -14194 13203 -14160
rect 13237 -14194 13271 -14160
rect 13305 -14194 13339 -14160
rect 13373 -14194 13407 -14160
rect 13441 -14194 13475 -14160
rect 13509 -14194 13543 -14160
rect 14051 -14194 14085 -14160
rect 14119 -14194 14153 -14160
rect 14187 -14194 14221 -14160
rect 14255 -14194 14289 -14160
rect 14323 -14194 14357 -14160
rect 14391 -14194 14425 -14160
rect 14459 -14194 14493 -14160
rect 14527 -14194 14561 -14160
rect 15069 -14194 15103 -14160
rect 15137 -14194 15171 -14160
rect 15205 -14194 15239 -14160
rect 15273 -14194 15307 -14160
rect 15341 -14194 15375 -14160
rect 15409 -14194 15443 -14160
rect 15477 -14194 15511 -14160
rect 15545 -14194 15579 -14160
rect 16087 -14194 16121 -14160
rect 16155 -14194 16189 -14160
rect 16223 -14194 16257 -14160
rect 16291 -14194 16325 -14160
rect 16359 -14194 16393 -14160
rect 16427 -14194 16461 -14160
rect 16495 -14194 16529 -14160
rect 16563 -14194 16597 -14160
rect 17105 -14194 17139 -14160
rect 17173 -14194 17207 -14160
rect 17241 -14194 17275 -14160
rect 17309 -14194 17343 -14160
rect 17377 -14194 17411 -14160
rect 17445 -14194 17479 -14160
rect 17513 -14194 17547 -14160
rect 17581 -14194 17615 -14160
rect 18123 -14194 18157 -14160
rect 18191 -14194 18225 -14160
rect 18259 -14194 18293 -14160
rect 18327 -14194 18361 -14160
rect 18395 -14194 18429 -14160
rect 18463 -14194 18497 -14160
rect 18531 -14194 18565 -14160
rect 18599 -14194 18633 -14160
rect 19141 -14194 19175 -14160
rect 19209 -14194 19243 -14160
rect 19277 -14194 19311 -14160
rect 19345 -14194 19379 -14160
rect 19413 -14194 19447 -14160
rect 19481 -14194 19515 -14160
rect 19549 -14194 19583 -14160
rect 19617 -14194 19651 -14160
rect 20159 -14194 20193 -14160
rect 20227 -14194 20261 -14160
rect 20295 -14194 20329 -14160
rect 20363 -14194 20397 -14160
rect 20431 -14194 20465 -14160
rect 20499 -14194 20533 -14160
rect 20567 -14194 20601 -14160
rect 20635 -14194 20669 -14160
rect 21177 -14194 21211 -14160
rect 21245 -14194 21279 -14160
rect 21313 -14194 21347 -14160
rect 21381 -14194 21415 -14160
rect 21449 -14194 21483 -14160
rect 21517 -14194 21551 -14160
rect 21585 -14194 21619 -14160
rect 21653 -14194 21687 -14160
rect 22195 -14194 22229 -14160
rect 22263 -14194 22297 -14160
rect 22331 -14194 22365 -14160
rect 22399 -14194 22433 -14160
rect 22467 -14194 22501 -14160
rect 22535 -14194 22569 -14160
rect 22603 -14194 22637 -14160
rect 22671 -14194 22705 -14160
rect -8913 -14820 -8879 -14786
rect -8845 -14820 -8811 -14786
rect -8777 -14820 -8743 -14786
rect -8709 -14820 -8675 -14786
rect -8641 -14820 -8607 -14786
rect -8573 -14820 -8539 -14786
rect -8505 -14820 -8471 -14786
rect -8437 -14820 -8403 -14786
rect -7895 -14820 -7861 -14786
rect -7827 -14820 -7793 -14786
rect -7759 -14820 -7725 -14786
rect -7691 -14820 -7657 -14786
rect -7623 -14820 -7589 -14786
rect -7555 -14820 -7521 -14786
rect -7487 -14820 -7453 -14786
rect -7419 -14820 -7385 -14786
rect -6877 -14820 -6843 -14786
rect -6809 -14820 -6775 -14786
rect -6741 -14820 -6707 -14786
rect -6673 -14820 -6639 -14786
rect -6605 -14820 -6571 -14786
rect -6537 -14820 -6503 -14786
rect -6469 -14820 -6435 -14786
rect -6401 -14820 -6367 -14786
rect -5859 -14820 -5825 -14786
rect -5791 -14820 -5757 -14786
rect -5723 -14820 -5689 -14786
rect -5655 -14820 -5621 -14786
rect -5587 -14820 -5553 -14786
rect -5519 -14820 -5485 -14786
rect -5451 -14820 -5417 -14786
rect -5383 -14820 -5349 -14786
rect -4841 -14820 -4807 -14786
rect -4773 -14820 -4739 -14786
rect -4705 -14820 -4671 -14786
rect -4637 -14820 -4603 -14786
rect -4569 -14820 -4535 -14786
rect -4501 -14820 -4467 -14786
rect -4433 -14820 -4399 -14786
rect -4365 -14820 -4331 -14786
rect -3823 -14820 -3789 -14786
rect -3755 -14820 -3721 -14786
rect -3687 -14820 -3653 -14786
rect -3619 -14820 -3585 -14786
rect -3551 -14820 -3517 -14786
rect -3483 -14820 -3449 -14786
rect -3415 -14820 -3381 -14786
rect -3347 -14820 -3313 -14786
rect -2805 -14820 -2771 -14786
rect -2737 -14820 -2703 -14786
rect -2669 -14820 -2635 -14786
rect -2601 -14820 -2567 -14786
rect -2533 -14820 -2499 -14786
rect -2465 -14820 -2431 -14786
rect -2397 -14820 -2363 -14786
rect -2329 -14820 -2295 -14786
rect -1787 -14820 -1753 -14786
rect -1719 -14820 -1685 -14786
rect -1651 -14820 -1617 -14786
rect -1583 -14820 -1549 -14786
rect -1515 -14820 -1481 -14786
rect -1447 -14820 -1413 -14786
rect -1379 -14820 -1345 -14786
rect -1311 -14820 -1277 -14786
rect -769 -14820 -735 -14786
rect -701 -14820 -667 -14786
rect -633 -14820 -599 -14786
rect -565 -14820 -531 -14786
rect -497 -14820 -463 -14786
rect -429 -14820 -395 -14786
rect -361 -14820 -327 -14786
rect -293 -14820 -259 -14786
rect -8913 -14928 -8879 -14894
rect -8845 -14928 -8811 -14894
rect -8777 -14928 -8743 -14894
rect -8709 -14928 -8675 -14894
rect -8641 -14928 -8607 -14894
rect -8573 -14928 -8539 -14894
rect -8505 -14928 -8471 -14894
rect -8437 -14928 -8403 -14894
rect -7895 -14928 -7861 -14894
rect -7827 -14928 -7793 -14894
rect -7759 -14928 -7725 -14894
rect -7691 -14928 -7657 -14894
rect -7623 -14928 -7589 -14894
rect -7555 -14928 -7521 -14894
rect -7487 -14928 -7453 -14894
rect -7419 -14928 -7385 -14894
rect -6877 -14928 -6843 -14894
rect -6809 -14928 -6775 -14894
rect -6741 -14928 -6707 -14894
rect -6673 -14928 -6639 -14894
rect -6605 -14928 -6571 -14894
rect -6537 -14928 -6503 -14894
rect -6469 -14928 -6435 -14894
rect -6401 -14928 -6367 -14894
rect -5859 -14928 -5825 -14894
rect -5791 -14928 -5757 -14894
rect -5723 -14928 -5689 -14894
rect -5655 -14928 -5621 -14894
rect -5587 -14928 -5553 -14894
rect -5519 -14928 -5485 -14894
rect -5451 -14928 -5417 -14894
rect -5383 -14928 -5349 -14894
rect -4841 -14928 -4807 -14894
rect -4773 -14928 -4739 -14894
rect -4705 -14928 -4671 -14894
rect -4637 -14928 -4603 -14894
rect -4569 -14928 -4535 -14894
rect -4501 -14928 -4467 -14894
rect -4433 -14928 -4399 -14894
rect -4365 -14928 -4331 -14894
rect -3823 -14928 -3789 -14894
rect -3755 -14928 -3721 -14894
rect -3687 -14928 -3653 -14894
rect -3619 -14928 -3585 -14894
rect -3551 -14928 -3517 -14894
rect -3483 -14928 -3449 -14894
rect -3415 -14928 -3381 -14894
rect -3347 -14928 -3313 -14894
rect -2805 -14928 -2771 -14894
rect -2737 -14928 -2703 -14894
rect -2669 -14928 -2635 -14894
rect -2601 -14928 -2567 -14894
rect -2533 -14928 -2499 -14894
rect -2465 -14928 -2431 -14894
rect -2397 -14928 -2363 -14894
rect -2329 -14928 -2295 -14894
rect -1787 -14928 -1753 -14894
rect -1719 -14928 -1685 -14894
rect -1651 -14928 -1617 -14894
rect -1583 -14928 -1549 -14894
rect -1515 -14928 -1481 -14894
rect -1447 -14928 -1413 -14894
rect -1379 -14928 -1345 -14894
rect -1311 -14928 -1277 -14894
rect -769 -14928 -735 -14894
rect -701 -14928 -667 -14894
rect -633 -14928 -599 -14894
rect -565 -14928 -531 -14894
rect -497 -14928 -463 -14894
rect -429 -14928 -395 -14894
rect -361 -14928 -327 -14894
rect -293 -14928 -259 -14894
rect 2853 -14904 2887 -14870
rect 2921 -14904 2955 -14870
rect 2989 -14904 3023 -14870
rect 3057 -14904 3091 -14870
rect 3125 -14904 3159 -14870
rect 3193 -14904 3227 -14870
rect 3261 -14904 3295 -14870
rect 3329 -14904 3363 -14870
rect 3871 -14904 3905 -14870
rect 3939 -14904 3973 -14870
rect 4007 -14904 4041 -14870
rect 4075 -14904 4109 -14870
rect 4143 -14904 4177 -14870
rect 4211 -14904 4245 -14870
rect 4279 -14904 4313 -14870
rect 4347 -14904 4381 -14870
rect 4889 -14904 4923 -14870
rect 4957 -14904 4991 -14870
rect 5025 -14904 5059 -14870
rect 5093 -14904 5127 -14870
rect 5161 -14904 5195 -14870
rect 5229 -14904 5263 -14870
rect 5297 -14904 5331 -14870
rect 5365 -14904 5399 -14870
rect 5907 -14904 5941 -14870
rect 5975 -14904 6009 -14870
rect 6043 -14904 6077 -14870
rect 6111 -14904 6145 -14870
rect 6179 -14904 6213 -14870
rect 6247 -14904 6281 -14870
rect 6315 -14904 6349 -14870
rect 6383 -14904 6417 -14870
rect 6925 -14904 6959 -14870
rect 6993 -14904 7027 -14870
rect 7061 -14904 7095 -14870
rect 7129 -14904 7163 -14870
rect 7197 -14904 7231 -14870
rect 7265 -14904 7299 -14870
rect 7333 -14904 7367 -14870
rect 7401 -14904 7435 -14870
rect 7943 -14904 7977 -14870
rect 8011 -14904 8045 -14870
rect 8079 -14904 8113 -14870
rect 8147 -14904 8181 -14870
rect 8215 -14904 8249 -14870
rect 8283 -14904 8317 -14870
rect 8351 -14904 8385 -14870
rect 8419 -14904 8453 -14870
rect 8961 -14904 8995 -14870
rect 9029 -14904 9063 -14870
rect 9097 -14904 9131 -14870
rect 9165 -14904 9199 -14870
rect 9233 -14904 9267 -14870
rect 9301 -14904 9335 -14870
rect 9369 -14904 9403 -14870
rect 9437 -14904 9471 -14870
rect 9979 -14904 10013 -14870
rect 10047 -14904 10081 -14870
rect 10115 -14904 10149 -14870
rect 10183 -14904 10217 -14870
rect 10251 -14904 10285 -14870
rect 10319 -14904 10353 -14870
rect 10387 -14904 10421 -14870
rect 10455 -14904 10489 -14870
rect 10997 -14904 11031 -14870
rect 11065 -14904 11099 -14870
rect 11133 -14904 11167 -14870
rect 11201 -14904 11235 -14870
rect 11269 -14904 11303 -14870
rect 11337 -14904 11371 -14870
rect 11405 -14904 11439 -14870
rect 11473 -14904 11507 -14870
rect 12015 -14904 12049 -14870
rect 12083 -14904 12117 -14870
rect 12151 -14904 12185 -14870
rect 12219 -14904 12253 -14870
rect 12287 -14904 12321 -14870
rect 12355 -14904 12389 -14870
rect 12423 -14904 12457 -14870
rect 12491 -14904 12525 -14870
rect 13033 -14904 13067 -14870
rect 13101 -14904 13135 -14870
rect 13169 -14904 13203 -14870
rect 13237 -14904 13271 -14870
rect 13305 -14904 13339 -14870
rect 13373 -14904 13407 -14870
rect 13441 -14904 13475 -14870
rect 13509 -14904 13543 -14870
rect 14051 -14904 14085 -14870
rect 14119 -14904 14153 -14870
rect 14187 -14904 14221 -14870
rect 14255 -14904 14289 -14870
rect 14323 -14904 14357 -14870
rect 14391 -14904 14425 -14870
rect 14459 -14904 14493 -14870
rect 14527 -14904 14561 -14870
rect 15069 -14904 15103 -14870
rect 15137 -14904 15171 -14870
rect 15205 -14904 15239 -14870
rect 15273 -14904 15307 -14870
rect 15341 -14904 15375 -14870
rect 15409 -14904 15443 -14870
rect 15477 -14904 15511 -14870
rect 15545 -14904 15579 -14870
rect 16087 -14904 16121 -14870
rect 16155 -14904 16189 -14870
rect 16223 -14904 16257 -14870
rect 16291 -14904 16325 -14870
rect 16359 -14904 16393 -14870
rect 16427 -14904 16461 -14870
rect 16495 -14904 16529 -14870
rect 16563 -14904 16597 -14870
rect 17105 -14904 17139 -14870
rect 17173 -14904 17207 -14870
rect 17241 -14904 17275 -14870
rect 17309 -14904 17343 -14870
rect 17377 -14904 17411 -14870
rect 17445 -14904 17479 -14870
rect 17513 -14904 17547 -14870
rect 17581 -14904 17615 -14870
rect 18123 -14904 18157 -14870
rect 18191 -14904 18225 -14870
rect 18259 -14904 18293 -14870
rect 18327 -14904 18361 -14870
rect 18395 -14904 18429 -14870
rect 18463 -14904 18497 -14870
rect 18531 -14904 18565 -14870
rect 18599 -14904 18633 -14870
rect 19141 -14904 19175 -14870
rect 19209 -14904 19243 -14870
rect 19277 -14904 19311 -14870
rect 19345 -14904 19379 -14870
rect 19413 -14904 19447 -14870
rect 19481 -14904 19515 -14870
rect 19549 -14904 19583 -14870
rect 19617 -14904 19651 -14870
rect 20159 -14904 20193 -14870
rect 20227 -14904 20261 -14870
rect 20295 -14904 20329 -14870
rect 20363 -14904 20397 -14870
rect 20431 -14904 20465 -14870
rect 20499 -14904 20533 -14870
rect 20567 -14904 20601 -14870
rect 20635 -14904 20669 -14870
rect 21177 -14904 21211 -14870
rect 21245 -14904 21279 -14870
rect 21313 -14904 21347 -14870
rect 21381 -14904 21415 -14870
rect 21449 -14904 21483 -14870
rect 21517 -14904 21551 -14870
rect 21585 -14904 21619 -14870
rect 21653 -14904 21687 -14870
rect 22195 -14904 22229 -14870
rect 22263 -14904 22297 -14870
rect 22331 -14904 22365 -14870
rect 22399 -14904 22433 -14870
rect 22467 -14904 22501 -14870
rect 22535 -14904 22569 -14870
rect 22603 -14904 22637 -14870
rect 22671 -14904 22705 -14870
rect 2853 -15426 2887 -15392
rect 2921 -15426 2955 -15392
rect 2989 -15426 3023 -15392
rect 3057 -15426 3091 -15392
rect 3125 -15426 3159 -15392
rect 3193 -15426 3227 -15392
rect 3261 -15426 3295 -15392
rect 3329 -15426 3363 -15392
rect 3871 -15426 3905 -15392
rect 3939 -15426 3973 -15392
rect 4007 -15426 4041 -15392
rect 4075 -15426 4109 -15392
rect 4143 -15426 4177 -15392
rect 4211 -15426 4245 -15392
rect 4279 -15426 4313 -15392
rect 4347 -15426 4381 -15392
rect 4889 -15426 4923 -15392
rect 4957 -15426 4991 -15392
rect 5025 -15426 5059 -15392
rect 5093 -15426 5127 -15392
rect 5161 -15426 5195 -15392
rect 5229 -15426 5263 -15392
rect 5297 -15426 5331 -15392
rect 5365 -15426 5399 -15392
rect 5907 -15426 5941 -15392
rect 5975 -15426 6009 -15392
rect 6043 -15426 6077 -15392
rect 6111 -15426 6145 -15392
rect 6179 -15426 6213 -15392
rect 6247 -15426 6281 -15392
rect 6315 -15426 6349 -15392
rect 6383 -15426 6417 -15392
rect 6925 -15426 6959 -15392
rect 6993 -15426 7027 -15392
rect 7061 -15426 7095 -15392
rect 7129 -15426 7163 -15392
rect 7197 -15426 7231 -15392
rect 7265 -15426 7299 -15392
rect 7333 -15426 7367 -15392
rect 7401 -15426 7435 -15392
rect 7943 -15426 7977 -15392
rect 8011 -15426 8045 -15392
rect 8079 -15426 8113 -15392
rect 8147 -15426 8181 -15392
rect 8215 -15426 8249 -15392
rect 8283 -15426 8317 -15392
rect 8351 -15426 8385 -15392
rect 8419 -15426 8453 -15392
rect 8961 -15426 8995 -15392
rect 9029 -15426 9063 -15392
rect 9097 -15426 9131 -15392
rect 9165 -15426 9199 -15392
rect 9233 -15426 9267 -15392
rect 9301 -15426 9335 -15392
rect 9369 -15426 9403 -15392
rect 9437 -15426 9471 -15392
rect 9979 -15426 10013 -15392
rect 10047 -15426 10081 -15392
rect 10115 -15426 10149 -15392
rect 10183 -15426 10217 -15392
rect 10251 -15426 10285 -15392
rect 10319 -15426 10353 -15392
rect 10387 -15426 10421 -15392
rect 10455 -15426 10489 -15392
rect 10997 -15426 11031 -15392
rect 11065 -15426 11099 -15392
rect 11133 -15426 11167 -15392
rect 11201 -15426 11235 -15392
rect 11269 -15426 11303 -15392
rect 11337 -15426 11371 -15392
rect 11405 -15426 11439 -15392
rect 11473 -15426 11507 -15392
rect 12015 -15426 12049 -15392
rect 12083 -15426 12117 -15392
rect 12151 -15426 12185 -15392
rect 12219 -15426 12253 -15392
rect 12287 -15426 12321 -15392
rect 12355 -15426 12389 -15392
rect 12423 -15426 12457 -15392
rect 12491 -15426 12525 -15392
rect 13033 -15426 13067 -15392
rect 13101 -15426 13135 -15392
rect 13169 -15426 13203 -15392
rect 13237 -15426 13271 -15392
rect 13305 -15426 13339 -15392
rect 13373 -15426 13407 -15392
rect 13441 -15426 13475 -15392
rect 13509 -15426 13543 -15392
rect 14051 -15426 14085 -15392
rect 14119 -15426 14153 -15392
rect 14187 -15426 14221 -15392
rect 14255 -15426 14289 -15392
rect 14323 -15426 14357 -15392
rect 14391 -15426 14425 -15392
rect 14459 -15426 14493 -15392
rect 14527 -15426 14561 -15392
rect 15069 -15426 15103 -15392
rect 15137 -15426 15171 -15392
rect 15205 -15426 15239 -15392
rect 15273 -15426 15307 -15392
rect 15341 -15426 15375 -15392
rect 15409 -15426 15443 -15392
rect 15477 -15426 15511 -15392
rect 15545 -15426 15579 -15392
rect 16087 -15426 16121 -15392
rect 16155 -15426 16189 -15392
rect 16223 -15426 16257 -15392
rect 16291 -15426 16325 -15392
rect 16359 -15426 16393 -15392
rect 16427 -15426 16461 -15392
rect 16495 -15426 16529 -15392
rect 16563 -15426 16597 -15392
rect 17105 -15426 17139 -15392
rect 17173 -15426 17207 -15392
rect 17241 -15426 17275 -15392
rect 17309 -15426 17343 -15392
rect 17377 -15426 17411 -15392
rect 17445 -15426 17479 -15392
rect 17513 -15426 17547 -15392
rect 17581 -15426 17615 -15392
rect 18123 -15426 18157 -15392
rect 18191 -15426 18225 -15392
rect 18259 -15426 18293 -15392
rect 18327 -15426 18361 -15392
rect 18395 -15426 18429 -15392
rect 18463 -15426 18497 -15392
rect 18531 -15426 18565 -15392
rect 18599 -15426 18633 -15392
rect 19141 -15426 19175 -15392
rect 19209 -15426 19243 -15392
rect 19277 -15426 19311 -15392
rect 19345 -15426 19379 -15392
rect 19413 -15426 19447 -15392
rect 19481 -15426 19515 -15392
rect 19549 -15426 19583 -15392
rect 19617 -15426 19651 -15392
rect 20159 -15426 20193 -15392
rect 20227 -15426 20261 -15392
rect 20295 -15426 20329 -15392
rect 20363 -15426 20397 -15392
rect 20431 -15426 20465 -15392
rect 20499 -15426 20533 -15392
rect 20567 -15426 20601 -15392
rect 20635 -15426 20669 -15392
rect 21177 -15426 21211 -15392
rect 21245 -15426 21279 -15392
rect 21313 -15426 21347 -15392
rect 21381 -15426 21415 -15392
rect 21449 -15426 21483 -15392
rect 21517 -15426 21551 -15392
rect 21585 -15426 21619 -15392
rect 21653 -15426 21687 -15392
rect 22195 -15426 22229 -15392
rect 22263 -15426 22297 -15392
rect 22331 -15426 22365 -15392
rect 22399 -15426 22433 -15392
rect 22467 -15426 22501 -15392
rect 22535 -15426 22569 -15392
rect 22603 -15426 22637 -15392
rect 22671 -15426 22705 -15392
rect -8913 -15638 -8879 -15604
rect -8845 -15638 -8811 -15604
rect -8777 -15638 -8743 -15604
rect -8709 -15638 -8675 -15604
rect -8641 -15638 -8607 -15604
rect -8573 -15638 -8539 -15604
rect -8505 -15638 -8471 -15604
rect -8437 -15638 -8403 -15604
rect -7895 -15638 -7861 -15604
rect -7827 -15638 -7793 -15604
rect -7759 -15638 -7725 -15604
rect -7691 -15638 -7657 -15604
rect -7623 -15638 -7589 -15604
rect -7555 -15638 -7521 -15604
rect -7487 -15638 -7453 -15604
rect -7419 -15638 -7385 -15604
rect -6877 -15638 -6843 -15604
rect -6809 -15638 -6775 -15604
rect -6741 -15638 -6707 -15604
rect -6673 -15638 -6639 -15604
rect -6605 -15638 -6571 -15604
rect -6537 -15638 -6503 -15604
rect -6469 -15638 -6435 -15604
rect -6401 -15638 -6367 -15604
rect -5859 -15638 -5825 -15604
rect -5791 -15638 -5757 -15604
rect -5723 -15638 -5689 -15604
rect -5655 -15638 -5621 -15604
rect -5587 -15638 -5553 -15604
rect -5519 -15638 -5485 -15604
rect -5451 -15638 -5417 -15604
rect -5383 -15638 -5349 -15604
rect -4841 -15638 -4807 -15604
rect -4773 -15638 -4739 -15604
rect -4705 -15638 -4671 -15604
rect -4637 -15638 -4603 -15604
rect -4569 -15638 -4535 -15604
rect -4501 -15638 -4467 -15604
rect -4433 -15638 -4399 -15604
rect -4365 -15638 -4331 -15604
rect -3823 -15638 -3789 -15604
rect -3755 -15638 -3721 -15604
rect -3687 -15638 -3653 -15604
rect -3619 -15638 -3585 -15604
rect -3551 -15638 -3517 -15604
rect -3483 -15638 -3449 -15604
rect -3415 -15638 -3381 -15604
rect -3347 -15638 -3313 -15604
rect -2805 -15638 -2771 -15604
rect -2737 -15638 -2703 -15604
rect -2669 -15638 -2635 -15604
rect -2601 -15638 -2567 -15604
rect -2533 -15638 -2499 -15604
rect -2465 -15638 -2431 -15604
rect -2397 -15638 -2363 -15604
rect -2329 -15638 -2295 -15604
rect -1787 -15638 -1753 -15604
rect -1719 -15638 -1685 -15604
rect -1651 -15638 -1617 -15604
rect -1583 -15638 -1549 -15604
rect -1515 -15638 -1481 -15604
rect -1447 -15638 -1413 -15604
rect -1379 -15638 -1345 -15604
rect -1311 -15638 -1277 -15604
rect -769 -15638 -735 -15604
rect -701 -15638 -667 -15604
rect -633 -15638 -599 -15604
rect -565 -15638 -531 -15604
rect -497 -15638 -463 -15604
rect -429 -15638 -395 -15604
rect -361 -15638 -327 -15604
rect -293 -15638 -259 -15604
rect -8913 -15746 -8879 -15712
rect -8845 -15746 -8811 -15712
rect -8777 -15746 -8743 -15712
rect -8709 -15746 -8675 -15712
rect -8641 -15746 -8607 -15712
rect -8573 -15746 -8539 -15712
rect -8505 -15746 -8471 -15712
rect -8437 -15746 -8403 -15712
rect -7895 -15746 -7861 -15712
rect -7827 -15746 -7793 -15712
rect -7759 -15746 -7725 -15712
rect -7691 -15746 -7657 -15712
rect -7623 -15746 -7589 -15712
rect -7555 -15746 -7521 -15712
rect -7487 -15746 -7453 -15712
rect -7419 -15746 -7385 -15712
rect -6877 -15746 -6843 -15712
rect -6809 -15746 -6775 -15712
rect -6741 -15746 -6707 -15712
rect -6673 -15746 -6639 -15712
rect -6605 -15746 -6571 -15712
rect -6537 -15746 -6503 -15712
rect -6469 -15746 -6435 -15712
rect -6401 -15746 -6367 -15712
rect -5859 -15746 -5825 -15712
rect -5791 -15746 -5757 -15712
rect -5723 -15746 -5689 -15712
rect -5655 -15746 -5621 -15712
rect -5587 -15746 -5553 -15712
rect -5519 -15746 -5485 -15712
rect -5451 -15746 -5417 -15712
rect -5383 -15746 -5349 -15712
rect -4841 -15746 -4807 -15712
rect -4773 -15746 -4739 -15712
rect -4705 -15746 -4671 -15712
rect -4637 -15746 -4603 -15712
rect -4569 -15746 -4535 -15712
rect -4501 -15746 -4467 -15712
rect -4433 -15746 -4399 -15712
rect -4365 -15746 -4331 -15712
rect -3823 -15746 -3789 -15712
rect -3755 -15746 -3721 -15712
rect -3687 -15746 -3653 -15712
rect -3619 -15746 -3585 -15712
rect -3551 -15746 -3517 -15712
rect -3483 -15746 -3449 -15712
rect -3415 -15746 -3381 -15712
rect -3347 -15746 -3313 -15712
rect -2805 -15746 -2771 -15712
rect -2737 -15746 -2703 -15712
rect -2669 -15746 -2635 -15712
rect -2601 -15746 -2567 -15712
rect -2533 -15746 -2499 -15712
rect -2465 -15746 -2431 -15712
rect -2397 -15746 -2363 -15712
rect -2329 -15746 -2295 -15712
rect -1787 -15746 -1753 -15712
rect -1719 -15746 -1685 -15712
rect -1651 -15746 -1617 -15712
rect -1583 -15746 -1549 -15712
rect -1515 -15746 -1481 -15712
rect -1447 -15746 -1413 -15712
rect -1379 -15746 -1345 -15712
rect -1311 -15746 -1277 -15712
rect -769 -15746 -735 -15712
rect -701 -15746 -667 -15712
rect -633 -15746 -599 -15712
rect -565 -15746 -531 -15712
rect -497 -15746 -463 -15712
rect -429 -15746 -395 -15712
rect -361 -15746 -327 -15712
rect -293 -15746 -259 -15712
rect 2853 -16136 2887 -16102
rect 2921 -16136 2955 -16102
rect 2989 -16136 3023 -16102
rect 3057 -16136 3091 -16102
rect 3125 -16136 3159 -16102
rect 3193 -16136 3227 -16102
rect 3261 -16136 3295 -16102
rect 3329 -16136 3363 -16102
rect 3871 -16136 3905 -16102
rect 3939 -16136 3973 -16102
rect 4007 -16136 4041 -16102
rect 4075 -16136 4109 -16102
rect 4143 -16136 4177 -16102
rect 4211 -16136 4245 -16102
rect 4279 -16136 4313 -16102
rect 4347 -16136 4381 -16102
rect 4889 -16136 4923 -16102
rect 4957 -16136 4991 -16102
rect 5025 -16136 5059 -16102
rect 5093 -16136 5127 -16102
rect 5161 -16136 5195 -16102
rect 5229 -16136 5263 -16102
rect 5297 -16136 5331 -16102
rect 5365 -16136 5399 -16102
rect 5907 -16136 5941 -16102
rect 5975 -16136 6009 -16102
rect 6043 -16136 6077 -16102
rect 6111 -16136 6145 -16102
rect 6179 -16136 6213 -16102
rect 6247 -16136 6281 -16102
rect 6315 -16136 6349 -16102
rect 6383 -16136 6417 -16102
rect 6925 -16136 6959 -16102
rect 6993 -16136 7027 -16102
rect 7061 -16136 7095 -16102
rect 7129 -16136 7163 -16102
rect 7197 -16136 7231 -16102
rect 7265 -16136 7299 -16102
rect 7333 -16136 7367 -16102
rect 7401 -16136 7435 -16102
rect 7943 -16136 7977 -16102
rect 8011 -16136 8045 -16102
rect 8079 -16136 8113 -16102
rect 8147 -16136 8181 -16102
rect 8215 -16136 8249 -16102
rect 8283 -16136 8317 -16102
rect 8351 -16136 8385 -16102
rect 8419 -16136 8453 -16102
rect 8961 -16136 8995 -16102
rect 9029 -16136 9063 -16102
rect 9097 -16136 9131 -16102
rect 9165 -16136 9199 -16102
rect 9233 -16136 9267 -16102
rect 9301 -16136 9335 -16102
rect 9369 -16136 9403 -16102
rect 9437 -16136 9471 -16102
rect 9979 -16136 10013 -16102
rect 10047 -16136 10081 -16102
rect 10115 -16136 10149 -16102
rect 10183 -16136 10217 -16102
rect 10251 -16136 10285 -16102
rect 10319 -16136 10353 -16102
rect 10387 -16136 10421 -16102
rect 10455 -16136 10489 -16102
rect 10997 -16136 11031 -16102
rect 11065 -16136 11099 -16102
rect 11133 -16136 11167 -16102
rect 11201 -16136 11235 -16102
rect 11269 -16136 11303 -16102
rect 11337 -16136 11371 -16102
rect 11405 -16136 11439 -16102
rect 11473 -16136 11507 -16102
rect 12015 -16136 12049 -16102
rect 12083 -16136 12117 -16102
rect 12151 -16136 12185 -16102
rect 12219 -16136 12253 -16102
rect 12287 -16136 12321 -16102
rect 12355 -16136 12389 -16102
rect 12423 -16136 12457 -16102
rect 12491 -16136 12525 -16102
rect 13033 -16136 13067 -16102
rect 13101 -16136 13135 -16102
rect 13169 -16136 13203 -16102
rect 13237 -16136 13271 -16102
rect 13305 -16136 13339 -16102
rect 13373 -16136 13407 -16102
rect 13441 -16136 13475 -16102
rect 13509 -16136 13543 -16102
rect 14051 -16136 14085 -16102
rect 14119 -16136 14153 -16102
rect 14187 -16136 14221 -16102
rect 14255 -16136 14289 -16102
rect 14323 -16136 14357 -16102
rect 14391 -16136 14425 -16102
rect 14459 -16136 14493 -16102
rect 14527 -16136 14561 -16102
rect 15069 -16136 15103 -16102
rect 15137 -16136 15171 -16102
rect 15205 -16136 15239 -16102
rect 15273 -16136 15307 -16102
rect 15341 -16136 15375 -16102
rect 15409 -16136 15443 -16102
rect 15477 -16136 15511 -16102
rect 15545 -16136 15579 -16102
rect 16087 -16136 16121 -16102
rect 16155 -16136 16189 -16102
rect 16223 -16136 16257 -16102
rect 16291 -16136 16325 -16102
rect 16359 -16136 16393 -16102
rect 16427 -16136 16461 -16102
rect 16495 -16136 16529 -16102
rect 16563 -16136 16597 -16102
rect 17105 -16136 17139 -16102
rect 17173 -16136 17207 -16102
rect 17241 -16136 17275 -16102
rect 17309 -16136 17343 -16102
rect 17377 -16136 17411 -16102
rect 17445 -16136 17479 -16102
rect 17513 -16136 17547 -16102
rect 17581 -16136 17615 -16102
rect 18123 -16136 18157 -16102
rect 18191 -16136 18225 -16102
rect 18259 -16136 18293 -16102
rect 18327 -16136 18361 -16102
rect 18395 -16136 18429 -16102
rect 18463 -16136 18497 -16102
rect 18531 -16136 18565 -16102
rect 18599 -16136 18633 -16102
rect 19141 -16136 19175 -16102
rect 19209 -16136 19243 -16102
rect 19277 -16136 19311 -16102
rect 19345 -16136 19379 -16102
rect 19413 -16136 19447 -16102
rect 19481 -16136 19515 -16102
rect 19549 -16136 19583 -16102
rect 19617 -16136 19651 -16102
rect 20159 -16136 20193 -16102
rect 20227 -16136 20261 -16102
rect 20295 -16136 20329 -16102
rect 20363 -16136 20397 -16102
rect 20431 -16136 20465 -16102
rect 20499 -16136 20533 -16102
rect 20567 -16136 20601 -16102
rect 20635 -16136 20669 -16102
rect 21177 -16136 21211 -16102
rect 21245 -16136 21279 -16102
rect 21313 -16136 21347 -16102
rect 21381 -16136 21415 -16102
rect 21449 -16136 21483 -16102
rect 21517 -16136 21551 -16102
rect 21585 -16136 21619 -16102
rect 21653 -16136 21687 -16102
rect 22195 -16136 22229 -16102
rect 22263 -16136 22297 -16102
rect 22331 -16136 22365 -16102
rect 22399 -16136 22433 -16102
rect 22467 -16136 22501 -16102
rect 22535 -16136 22569 -16102
rect 22603 -16136 22637 -16102
rect 22671 -16136 22705 -16102
rect -8913 -16456 -8879 -16422
rect -8845 -16456 -8811 -16422
rect -8777 -16456 -8743 -16422
rect -8709 -16456 -8675 -16422
rect -8641 -16456 -8607 -16422
rect -8573 -16456 -8539 -16422
rect -8505 -16456 -8471 -16422
rect -8437 -16456 -8403 -16422
rect -7895 -16456 -7861 -16422
rect -7827 -16456 -7793 -16422
rect -7759 -16456 -7725 -16422
rect -7691 -16456 -7657 -16422
rect -7623 -16456 -7589 -16422
rect -7555 -16456 -7521 -16422
rect -7487 -16456 -7453 -16422
rect -7419 -16456 -7385 -16422
rect -6877 -16456 -6843 -16422
rect -6809 -16456 -6775 -16422
rect -6741 -16456 -6707 -16422
rect -6673 -16456 -6639 -16422
rect -6605 -16456 -6571 -16422
rect -6537 -16456 -6503 -16422
rect -6469 -16456 -6435 -16422
rect -6401 -16456 -6367 -16422
rect -5859 -16456 -5825 -16422
rect -5791 -16456 -5757 -16422
rect -5723 -16456 -5689 -16422
rect -5655 -16456 -5621 -16422
rect -5587 -16456 -5553 -16422
rect -5519 -16456 -5485 -16422
rect -5451 -16456 -5417 -16422
rect -5383 -16456 -5349 -16422
rect -4841 -16456 -4807 -16422
rect -4773 -16456 -4739 -16422
rect -4705 -16456 -4671 -16422
rect -4637 -16456 -4603 -16422
rect -4569 -16456 -4535 -16422
rect -4501 -16456 -4467 -16422
rect -4433 -16456 -4399 -16422
rect -4365 -16456 -4331 -16422
rect -3823 -16456 -3789 -16422
rect -3755 -16456 -3721 -16422
rect -3687 -16456 -3653 -16422
rect -3619 -16456 -3585 -16422
rect -3551 -16456 -3517 -16422
rect -3483 -16456 -3449 -16422
rect -3415 -16456 -3381 -16422
rect -3347 -16456 -3313 -16422
rect -2805 -16456 -2771 -16422
rect -2737 -16456 -2703 -16422
rect -2669 -16456 -2635 -16422
rect -2601 -16456 -2567 -16422
rect -2533 -16456 -2499 -16422
rect -2465 -16456 -2431 -16422
rect -2397 -16456 -2363 -16422
rect -2329 -16456 -2295 -16422
rect -1787 -16456 -1753 -16422
rect -1719 -16456 -1685 -16422
rect -1651 -16456 -1617 -16422
rect -1583 -16456 -1549 -16422
rect -1515 -16456 -1481 -16422
rect -1447 -16456 -1413 -16422
rect -1379 -16456 -1345 -16422
rect -1311 -16456 -1277 -16422
rect -769 -16456 -735 -16422
rect -701 -16456 -667 -16422
rect -633 -16456 -599 -16422
rect -565 -16456 -531 -16422
rect -497 -16456 -463 -16422
rect -429 -16456 -395 -16422
rect -361 -16456 -327 -16422
rect -293 -16456 -259 -16422
rect -8913 -16564 -8879 -16530
rect -8845 -16564 -8811 -16530
rect -8777 -16564 -8743 -16530
rect -8709 -16564 -8675 -16530
rect -8641 -16564 -8607 -16530
rect -8573 -16564 -8539 -16530
rect -8505 -16564 -8471 -16530
rect -8437 -16564 -8403 -16530
rect -7895 -16564 -7861 -16530
rect -7827 -16564 -7793 -16530
rect -7759 -16564 -7725 -16530
rect -7691 -16564 -7657 -16530
rect -7623 -16564 -7589 -16530
rect -7555 -16564 -7521 -16530
rect -7487 -16564 -7453 -16530
rect -7419 -16564 -7385 -16530
rect -6877 -16564 -6843 -16530
rect -6809 -16564 -6775 -16530
rect -6741 -16564 -6707 -16530
rect -6673 -16564 -6639 -16530
rect -6605 -16564 -6571 -16530
rect -6537 -16564 -6503 -16530
rect -6469 -16564 -6435 -16530
rect -6401 -16564 -6367 -16530
rect -5859 -16564 -5825 -16530
rect -5791 -16564 -5757 -16530
rect -5723 -16564 -5689 -16530
rect -5655 -16564 -5621 -16530
rect -5587 -16564 -5553 -16530
rect -5519 -16564 -5485 -16530
rect -5451 -16564 -5417 -16530
rect -5383 -16564 -5349 -16530
rect -4841 -16564 -4807 -16530
rect -4773 -16564 -4739 -16530
rect -4705 -16564 -4671 -16530
rect -4637 -16564 -4603 -16530
rect -4569 -16564 -4535 -16530
rect -4501 -16564 -4467 -16530
rect -4433 -16564 -4399 -16530
rect -4365 -16564 -4331 -16530
rect -3823 -16564 -3789 -16530
rect -3755 -16564 -3721 -16530
rect -3687 -16564 -3653 -16530
rect -3619 -16564 -3585 -16530
rect -3551 -16564 -3517 -16530
rect -3483 -16564 -3449 -16530
rect -3415 -16564 -3381 -16530
rect -3347 -16564 -3313 -16530
rect -2805 -16564 -2771 -16530
rect -2737 -16564 -2703 -16530
rect -2669 -16564 -2635 -16530
rect -2601 -16564 -2567 -16530
rect -2533 -16564 -2499 -16530
rect -2465 -16564 -2431 -16530
rect -2397 -16564 -2363 -16530
rect -2329 -16564 -2295 -16530
rect -1787 -16564 -1753 -16530
rect -1719 -16564 -1685 -16530
rect -1651 -16564 -1617 -16530
rect -1583 -16564 -1549 -16530
rect -1515 -16564 -1481 -16530
rect -1447 -16564 -1413 -16530
rect -1379 -16564 -1345 -16530
rect -1311 -16564 -1277 -16530
rect -769 -16564 -735 -16530
rect -701 -16564 -667 -16530
rect -633 -16564 -599 -16530
rect -565 -16564 -531 -16530
rect -497 -16564 -463 -16530
rect -429 -16564 -395 -16530
rect -361 -16564 -327 -16530
rect -293 -16564 -259 -16530
rect 2851 -16660 2885 -16626
rect 2919 -16660 2953 -16626
rect 2987 -16660 3021 -16626
rect 3055 -16660 3089 -16626
rect 3123 -16660 3157 -16626
rect 3191 -16660 3225 -16626
rect 3259 -16660 3293 -16626
rect 3327 -16660 3361 -16626
rect 3869 -16660 3903 -16626
rect 3937 -16660 3971 -16626
rect 4005 -16660 4039 -16626
rect 4073 -16660 4107 -16626
rect 4141 -16660 4175 -16626
rect 4209 -16660 4243 -16626
rect 4277 -16660 4311 -16626
rect 4345 -16660 4379 -16626
rect 4887 -16660 4921 -16626
rect 4955 -16660 4989 -16626
rect 5023 -16660 5057 -16626
rect 5091 -16660 5125 -16626
rect 5159 -16660 5193 -16626
rect 5227 -16660 5261 -16626
rect 5295 -16660 5329 -16626
rect 5363 -16660 5397 -16626
rect 5905 -16660 5939 -16626
rect 5973 -16660 6007 -16626
rect 6041 -16660 6075 -16626
rect 6109 -16660 6143 -16626
rect 6177 -16660 6211 -16626
rect 6245 -16660 6279 -16626
rect 6313 -16660 6347 -16626
rect 6381 -16660 6415 -16626
rect 6923 -16660 6957 -16626
rect 6991 -16660 7025 -16626
rect 7059 -16660 7093 -16626
rect 7127 -16660 7161 -16626
rect 7195 -16660 7229 -16626
rect 7263 -16660 7297 -16626
rect 7331 -16660 7365 -16626
rect 7399 -16660 7433 -16626
rect 7941 -16660 7975 -16626
rect 8009 -16660 8043 -16626
rect 8077 -16660 8111 -16626
rect 8145 -16660 8179 -16626
rect 8213 -16660 8247 -16626
rect 8281 -16660 8315 -16626
rect 8349 -16660 8383 -16626
rect 8417 -16660 8451 -16626
rect 8959 -16660 8993 -16626
rect 9027 -16660 9061 -16626
rect 9095 -16660 9129 -16626
rect 9163 -16660 9197 -16626
rect 9231 -16660 9265 -16626
rect 9299 -16660 9333 -16626
rect 9367 -16660 9401 -16626
rect 9435 -16660 9469 -16626
rect 9977 -16660 10011 -16626
rect 10045 -16660 10079 -16626
rect 10113 -16660 10147 -16626
rect 10181 -16660 10215 -16626
rect 10249 -16660 10283 -16626
rect 10317 -16660 10351 -16626
rect 10385 -16660 10419 -16626
rect 10453 -16660 10487 -16626
rect 10995 -16660 11029 -16626
rect 11063 -16660 11097 -16626
rect 11131 -16660 11165 -16626
rect 11199 -16660 11233 -16626
rect 11267 -16660 11301 -16626
rect 11335 -16660 11369 -16626
rect 11403 -16660 11437 -16626
rect 11471 -16660 11505 -16626
rect 12013 -16660 12047 -16626
rect 12081 -16660 12115 -16626
rect 12149 -16660 12183 -16626
rect 12217 -16660 12251 -16626
rect 12285 -16660 12319 -16626
rect 12353 -16660 12387 -16626
rect 12421 -16660 12455 -16626
rect 12489 -16660 12523 -16626
rect 13031 -16660 13065 -16626
rect 13099 -16660 13133 -16626
rect 13167 -16660 13201 -16626
rect 13235 -16660 13269 -16626
rect 13303 -16660 13337 -16626
rect 13371 -16660 13405 -16626
rect 13439 -16660 13473 -16626
rect 13507 -16660 13541 -16626
rect 14049 -16660 14083 -16626
rect 14117 -16660 14151 -16626
rect 14185 -16660 14219 -16626
rect 14253 -16660 14287 -16626
rect 14321 -16660 14355 -16626
rect 14389 -16660 14423 -16626
rect 14457 -16660 14491 -16626
rect 14525 -16660 14559 -16626
rect 15067 -16660 15101 -16626
rect 15135 -16660 15169 -16626
rect 15203 -16660 15237 -16626
rect 15271 -16660 15305 -16626
rect 15339 -16660 15373 -16626
rect 15407 -16660 15441 -16626
rect 15475 -16660 15509 -16626
rect 15543 -16660 15577 -16626
rect 16085 -16660 16119 -16626
rect 16153 -16660 16187 -16626
rect 16221 -16660 16255 -16626
rect 16289 -16660 16323 -16626
rect 16357 -16660 16391 -16626
rect 16425 -16660 16459 -16626
rect 16493 -16660 16527 -16626
rect 16561 -16660 16595 -16626
rect 17103 -16660 17137 -16626
rect 17171 -16660 17205 -16626
rect 17239 -16660 17273 -16626
rect 17307 -16660 17341 -16626
rect 17375 -16660 17409 -16626
rect 17443 -16660 17477 -16626
rect 17511 -16660 17545 -16626
rect 17579 -16660 17613 -16626
rect 18121 -16660 18155 -16626
rect 18189 -16660 18223 -16626
rect 18257 -16660 18291 -16626
rect 18325 -16660 18359 -16626
rect 18393 -16660 18427 -16626
rect 18461 -16660 18495 -16626
rect 18529 -16660 18563 -16626
rect 18597 -16660 18631 -16626
rect 19139 -16660 19173 -16626
rect 19207 -16660 19241 -16626
rect 19275 -16660 19309 -16626
rect 19343 -16660 19377 -16626
rect 19411 -16660 19445 -16626
rect 19479 -16660 19513 -16626
rect 19547 -16660 19581 -16626
rect 19615 -16660 19649 -16626
rect 20157 -16660 20191 -16626
rect 20225 -16660 20259 -16626
rect 20293 -16660 20327 -16626
rect 20361 -16660 20395 -16626
rect 20429 -16660 20463 -16626
rect 20497 -16660 20531 -16626
rect 20565 -16660 20599 -16626
rect 20633 -16660 20667 -16626
rect 21175 -16660 21209 -16626
rect 21243 -16660 21277 -16626
rect 21311 -16660 21345 -16626
rect 21379 -16660 21413 -16626
rect 21447 -16660 21481 -16626
rect 21515 -16660 21549 -16626
rect 21583 -16660 21617 -16626
rect 21651 -16660 21685 -16626
rect 22193 -16660 22227 -16626
rect 22261 -16660 22295 -16626
rect 22329 -16660 22363 -16626
rect 22397 -16660 22431 -16626
rect 22465 -16660 22499 -16626
rect 22533 -16660 22567 -16626
rect 22601 -16660 22635 -16626
rect 22669 -16660 22703 -16626
rect -8913 -17274 -8879 -17240
rect -8845 -17274 -8811 -17240
rect -8777 -17274 -8743 -17240
rect -8709 -17274 -8675 -17240
rect -8641 -17274 -8607 -17240
rect -8573 -17274 -8539 -17240
rect -8505 -17274 -8471 -17240
rect -8437 -17274 -8403 -17240
rect -7895 -17274 -7861 -17240
rect -7827 -17274 -7793 -17240
rect -7759 -17274 -7725 -17240
rect -7691 -17274 -7657 -17240
rect -7623 -17274 -7589 -17240
rect -7555 -17274 -7521 -17240
rect -7487 -17274 -7453 -17240
rect -7419 -17274 -7385 -17240
rect -6877 -17274 -6843 -17240
rect -6809 -17274 -6775 -17240
rect -6741 -17274 -6707 -17240
rect -6673 -17274 -6639 -17240
rect -6605 -17274 -6571 -17240
rect -6537 -17274 -6503 -17240
rect -6469 -17274 -6435 -17240
rect -6401 -17274 -6367 -17240
rect -5859 -17274 -5825 -17240
rect -5791 -17274 -5757 -17240
rect -5723 -17274 -5689 -17240
rect -5655 -17274 -5621 -17240
rect -5587 -17274 -5553 -17240
rect -5519 -17274 -5485 -17240
rect -5451 -17274 -5417 -17240
rect -5383 -17274 -5349 -17240
rect -4841 -17274 -4807 -17240
rect -4773 -17274 -4739 -17240
rect -4705 -17274 -4671 -17240
rect -4637 -17274 -4603 -17240
rect -4569 -17274 -4535 -17240
rect -4501 -17274 -4467 -17240
rect -4433 -17274 -4399 -17240
rect -4365 -17274 -4331 -17240
rect -3823 -17274 -3789 -17240
rect -3755 -17274 -3721 -17240
rect -3687 -17274 -3653 -17240
rect -3619 -17274 -3585 -17240
rect -3551 -17274 -3517 -17240
rect -3483 -17274 -3449 -17240
rect -3415 -17274 -3381 -17240
rect -3347 -17274 -3313 -17240
rect -2805 -17274 -2771 -17240
rect -2737 -17274 -2703 -17240
rect -2669 -17274 -2635 -17240
rect -2601 -17274 -2567 -17240
rect -2533 -17274 -2499 -17240
rect -2465 -17274 -2431 -17240
rect -2397 -17274 -2363 -17240
rect -2329 -17274 -2295 -17240
rect -1787 -17274 -1753 -17240
rect -1719 -17274 -1685 -17240
rect -1651 -17274 -1617 -17240
rect -1583 -17274 -1549 -17240
rect -1515 -17274 -1481 -17240
rect -1447 -17274 -1413 -17240
rect -1379 -17274 -1345 -17240
rect -1311 -17274 -1277 -17240
rect -769 -17274 -735 -17240
rect -701 -17274 -667 -17240
rect -633 -17274 -599 -17240
rect -565 -17274 -531 -17240
rect -497 -17274 -463 -17240
rect -429 -17274 -395 -17240
rect -361 -17274 -327 -17240
rect -293 -17274 -259 -17240
rect -8913 -17382 -8879 -17348
rect -8845 -17382 -8811 -17348
rect -8777 -17382 -8743 -17348
rect -8709 -17382 -8675 -17348
rect -8641 -17382 -8607 -17348
rect -8573 -17382 -8539 -17348
rect -8505 -17382 -8471 -17348
rect -8437 -17382 -8403 -17348
rect -7895 -17382 -7861 -17348
rect -7827 -17382 -7793 -17348
rect -7759 -17382 -7725 -17348
rect -7691 -17382 -7657 -17348
rect -7623 -17382 -7589 -17348
rect -7555 -17382 -7521 -17348
rect -7487 -17382 -7453 -17348
rect -7419 -17382 -7385 -17348
rect -6877 -17382 -6843 -17348
rect -6809 -17382 -6775 -17348
rect -6741 -17382 -6707 -17348
rect -6673 -17382 -6639 -17348
rect -6605 -17382 -6571 -17348
rect -6537 -17382 -6503 -17348
rect -6469 -17382 -6435 -17348
rect -6401 -17382 -6367 -17348
rect -5859 -17382 -5825 -17348
rect -5791 -17382 -5757 -17348
rect -5723 -17382 -5689 -17348
rect -5655 -17382 -5621 -17348
rect -5587 -17382 -5553 -17348
rect -5519 -17382 -5485 -17348
rect -5451 -17382 -5417 -17348
rect -5383 -17382 -5349 -17348
rect -4841 -17382 -4807 -17348
rect -4773 -17382 -4739 -17348
rect -4705 -17382 -4671 -17348
rect -4637 -17382 -4603 -17348
rect -4569 -17382 -4535 -17348
rect -4501 -17382 -4467 -17348
rect -4433 -17382 -4399 -17348
rect -4365 -17382 -4331 -17348
rect -3823 -17382 -3789 -17348
rect -3755 -17382 -3721 -17348
rect -3687 -17382 -3653 -17348
rect -3619 -17382 -3585 -17348
rect -3551 -17382 -3517 -17348
rect -3483 -17382 -3449 -17348
rect -3415 -17382 -3381 -17348
rect -3347 -17382 -3313 -17348
rect -2805 -17382 -2771 -17348
rect -2737 -17382 -2703 -17348
rect -2669 -17382 -2635 -17348
rect -2601 -17382 -2567 -17348
rect -2533 -17382 -2499 -17348
rect -2465 -17382 -2431 -17348
rect -2397 -17382 -2363 -17348
rect -2329 -17382 -2295 -17348
rect -1787 -17382 -1753 -17348
rect -1719 -17382 -1685 -17348
rect -1651 -17382 -1617 -17348
rect -1583 -17382 -1549 -17348
rect -1515 -17382 -1481 -17348
rect -1447 -17382 -1413 -17348
rect -1379 -17382 -1345 -17348
rect -1311 -17382 -1277 -17348
rect -769 -17382 -735 -17348
rect -701 -17382 -667 -17348
rect -633 -17382 -599 -17348
rect -565 -17382 -531 -17348
rect -497 -17382 -463 -17348
rect -429 -17382 -395 -17348
rect -361 -17382 -327 -17348
rect -293 -17382 -259 -17348
rect 2851 -17370 2885 -17336
rect 2919 -17370 2953 -17336
rect 2987 -17370 3021 -17336
rect 3055 -17370 3089 -17336
rect 3123 -17370 3157 -17336
rect 3191 -17370 3225 -17336
rect 3259 -17370 3293 -17336
rect 3327 -17370 3361 -17336
rect 3869 -17370 3903 -17336
rect 3937 -17370 3971 -17336
rect 4005 -17370 4039 -17336
rect 4073 -17370 4107 -17336
rect 4141 -17370 4175 -17336
rect 4209 -17370 4243 -17336
rect 4277 -17370 4311 -17336
rect 4345 -17370 4379 -17336
rect 4887 -17370 4921 -17336
rect 4955 -17370 4989 -17336
rect 5023 -17370 5057 -17336
rect 5091 -17370 5125 -17336
rect 5159 -17370 5193 -17336
rect 5227 -17370 5261 -17336
rect 5295 -17370 5329 -17336
rect 5363 -17370 5397 -17336
rect 5905 -17370 5939 -17336
rect 5973 -17370 6007 -17336
rect 6041 -17370 6075 -17336
rect 6109 -17370 6143 -17336
rect 6177 -17370 6211 -17336
rect 6245 -17370 6279 -17336
rect 6313 -17370 6347 -17336
rect 6381 -17370 6415 -17336
rect 6923 -17370 6957 -17336
rect 6991 -17370 7025 -17336
rect 7059 -17370 7093 -17336
rect 7127 -17370 7161 -17336
rect 7195 -17370 7229 -17336
rect 7263 -17370 7297 -17336
rect 7331 -17370 7365 -17336
rect 7399 -17370 7433 -17336
rect 7941 -17370 7975 -17336
rect 8009 -17370 8043 -17336
rect 8077 -17370 8111 -17336
rect 8145 -17370 8179 -17336
rect 8213 -17370 8247 -17336
rect 8281 -17370 8315 -17336
rect 8349 -17370 8383 -17336
rect 8417 -17370 8451 -17336
rect 8959 -17370 8993 -17336
rect 9027 -17370 9061 -17336
rect 9095 -17370 9129 -17336
rect 9163 -17370 9197 -17336
rect 9231 -17370 9265 -17336
rect 9299 -17370 9333 -17336
rect 9367 -17370 9401 -17336
rect 9435 -17370 9469 -17336
rect 9977 -17370 10011 -17336
rect 10045 -17370 10079 -17336
rect 10113 -17370 10147 -17336
rect 10181 -17370 10215 -17336
rect 10249 -17370 10283 -17336
rect 10317 -17370 10351 -17336
rect 10385 -17370 10419 -17336
rect 10453 -17370 10487 -17336
rect 10995 -17370 11029 -17336
rect 11063 -17370 11097 -17336
rect 11131 -17370 11165 -17336
rect 11199 -17370 11233 -17336
rect 11267 -17370 11301 -17336
rect 11335 -17370 11369 -17336
rect 11403 -17370 11437 -17336
rect 11471 -17370 11505 -17336
rect 12013 -17370 12047 -17336
rect 12081 -17370 12115 -17336
rect 12149 -17370 12183 -17336
rect 12217 -17370 12251 -17336
rect 12285 -17370 12319 -17336
rect 12353 -17370 12387 -17336
rect 12421 -17370 12455 -17336
rect 12489 -17370 12523 -17336
rect 13031 -17370 13065 -17336
rect 13099 -17370 13133 -17336
rect 13167 -17370 13201 -17336
rect 13235 -17370 13269 -17336
rect 13303 -17370 13337 -17336
rect 13371 -17370 13405 -17336
rect 13439 -17370 13473 -17336
rect 13507 -17370 13541 -17336
rect 14049 -17370 14083 -17336
rect 14117 -17370 14151 -17336
rect 14185 -17370 14219 -17336
rect 14253 -17370 14287 -17336
rect 14321 -17370 14355 -17336
rect 14389 -17370 14423 -17336
rect 14457 -17370 14491 -17336
rect 14525 -17370 14559 -17336
rect 15067 -17370 15101 -17336
rect 15135 -17370 15169 -17336
rect 15203 -17370 15237 -17336
rect 15271 -17370 15305 -17336
rect 15339 -17370 15373 -17336
rect 15407 -17370 15441 -17336
rect 15475 -17370 15509 -17336
rect 15543 -17370 15577 -17336
rect 16085 -17370 16119 -17336
rect 16153 -17370 16187 -17336
rect 16221 -17370 16255 -17336
rect 16289 -17370 16323 -17336
rect 16357 -17370 16391 -17336
rect 16425 -17370 16459 -17336
rect 16493 -17370 16527 -17336
rect 16561 -17370 16595 -17336
rect 17103 -17370 17137 -17336
rect 17171 -17370 17205 -17336
rect 17239 -17370 17273 -17336
rect 17307 -17370 17341 -17336
rect 17375 -17370 17409 -17336
rect 17443 -17370 17477 -17336
rect 17511 -17370 17545 -17336
rect 17579 -17370 17613 -17336
rect 18121 -17370 18155 -17336
rect 18189 -17370 18223 -17336
rect 18257 -17370 18291 -17336
rect 18325 -17370 18359 -17336
rect 18393 -17370 18427 -17336
rect 18461 -17370 18495 -17336
rect 18529 -17370 18563 -17336
rect 18597 -17370 18631 -17336
rect 19139 -17370 19173 -17336
rect 19207 -17370 19241 -17336
rect 19275 -17370 19309 -17336
rect 19343 -17370 19377 -17336
rect 19411 -17370 19445 -17336
rect 19479 -17370 19513 -17336
rect 19547 -17370 19581 -17336
rect 19615 -17370 19649 -17336
rect 20157 -17370 20191 -17336
rect 20225 -17370 20259 -17336
rect 20293 -17370 20327 -17336
rect 20361 -17370 20395 -17336
rect 20429 -17370 20463 -17336
rect 20497 -17370 20531 -17336
rect 20565 -17370 20599 -17336
rect 20633 -17370 20667 -17336
rect 21175 -17370 21209 -17336
rect 21243 -17370 21277 -17336
rect 21311 -17370 21345 -17336
rect 21379 -17370 21413 -17336
rect 21447 -17370 21481 -17336
rect 21515 -17370 21549 -17336
rect 21583 -17370 21617 -17336
rect 21651 -17370 21685 -17336
rect 22193 -17370 22227 -17336
rect 22261 -17370 22295 -17336
rect 22329 -17370 22363 -17336
rect 22397 -17370 22431 -17336
rect 22465 -17370 22499 -17336
rect 22533 -17370 22567 -17336
rect 22601 -17370 22635 -17336
rect 22669 -17370 22703 -17336
rect 2851 -17894 2885 -17860
rect 2919 -17894 2953 -17860
rect 2987 -17894 3021 -17860
rect 3055 -17894 3089 -17860
rect 3123 -17894 3157 -17860
rect 3191 -17894 3225 -17860
rect 3259 -17894 3293 -17860
rect 3327 -17894 3361 -17860
rect 3869 -17894 3903 -17860
rect 3937 -17894 3971 -17860
rect 4005 -17894 4039 -17860
rect 4073 -17894 4107 -17860
rect 4141 -17894 4175 -17860
rect 4209 -17894 4243 -17860
rect 4277 -17894 4311 -17860
rect 4345 -17894 4379 -17860
rect 4887 -17894 4921 -17860
rect 4955 -17894 4989 -17860
rect 5023 -17894 5057 -17860
rect 5091 -17894 5125 -17860
rect 5159 -17894 5193 -17860
rect 5227 -17894 5261 -17860
rect 5295 -17894 5329 -17860
rect 5363 -17894 5397 -17860
rect 5905 -17894 5939 -17860
rect 5973 -17894 6007 -17860
rect 6041 -17894 6075 -17860
rect 6109 -17894 6143 -17860
rect 6177 -17894 6211 -17860
rect 6245 -17894 6279 -17860
rect 6313 -17894 6347 -17860
rect 6381 -17894 6415 -17860
rect 6923 -17894 6957 -17860
rect 6991 -17894 7025 -17860
rect 7059 -17894 7093 -17860
rect 7127 -17894 7161 -17860
rect 7195 -17894 7229 -17860
rect 7263 -17894 7297 -17860
rect 7331 -17894 7365 -17860
rect 7399 -17894 7433 -17860
rect 7941 -17894 7975 -17860
rect 8009 -17894 8043 -17860
rect 8077 -17894 8111 -17860
rect 8145 -17894 8179 -17860
rect 8213 -17894 8247 -17860
rect 8281 -17894 8315 -17860
rect 8349 -17894 8383 -17860
rect 8417 -17894 8451 -17860
rect 8959 -17894 8993 -17860
rect 9027 -17894 9061 -17860
rect 9095 -17894 9129 -17860
rect 9163 -17894 9197 -17860
rect 9231 -17894 9265 -17860
rect 9299 -17894 9333 -17860
rect 9367 -17894 9401 -17860
rect 9435 -17894 9469 -17860
rect 9977 -17894 10011 -17860
rect 10045 -17894 10079 -17860
rect 10113 -17894 10147 -17860
rect 10181 -17894 10215 -17860
rect 10249 -17894 10283 -17860
rect 10317 -17894 10351 -17860
rect 10385 -17894 10419 -17860
rect 10453 -17894 10487 -17860
rect 10995 -17894 11029 -17860
rect 11063 -17894 11097 -17860
rect 11131 -17894 11165 -17860
rect 11199 -17894 11233 -17860
rect 11267 -17894 11301 -17860
rect 11335 -17894 11369 -17860
rect 11403 -17894 11437 -17860
rect 11471 -17894 11505 -17860
rect 12013 -17894 12047 -17860
rect 12081 -17894 12115 -17860
rect 12149 -17894 12183 -17860
rect 12217 -17894 12251 -17860
rect 12285 -17894 12319 -17860
rect 12353 -17894 12387 -17860
rect 12421 -17894 12455 -17860
rect 12489 -17894 12523 -17860
rect 13031 -17894 13065 -17860
rect 13099 -17894 13133 -17860
rect 13167 -17894 13201 -17860
rect 13235 -17894 13269 -17860
rect 13303 -17894 13337 -17860
rect 13371 -17894 13405 -17860
rect 13439 -17894 13473 -17860
rect 13507 -17894 13541 -17860
rect 14049 -17894 14083 -17860
rect 14117 -17894 14151 -17860
rect 14185 -17894 14219 -17860
rect 14253 -17894 14287 -17860
rect 14321 -17894 14355 -17860
rect 14389 -17894 14423 -17860
rect 14457 -17894 14491 -17860
rect 14525 -17894 14559 -17860
rect 15067 -17894 15101 -17860
rect 15135 -17894 15169 -17860
rect 15203 -17894 15237 -17860
rect 15271 -17894 15305 -17860
rect 15339 -17894 15373 -17860
rect 15407 -17894 15441 -17860
rect 15475 -17894 15509 -17860
rect 15543 -17894 15577 -17860
rect 16085 -17894 16119 -17860
rect 16153 -17894 16187 -17860
rect 16221 -17894 16255 -17860
rect 16289 -17894 16323 -17860
rect 16357 -17894 16391 -17860
rect 16425 -17894 16459 -17860
rect 16493 -17894 16527 -17860
rect 16561 -17894 16595 -17860
rect 17103 -17894 17137 -17860
rect 17171 -17894 17205 -17860
rect 17239 -17894 17273 -17860
rect 17307 -17894 17341 -17860
rect 17375 -17894 17409 -17860
rect 17443 -17894 17477 -17860
rect 17511 -17894 17545 -17860
rect 17579 -17894 17613 -17860
rect 18121 -17894 18155 -17860
rect 18189 -17894 18223 -17860
rect 18257 -17894 18291 -17860
rect 18325 -17894 18359 -17860
rect 18393 -17894 18427 -17860
rect 18461 -17894 18495 -17860
rect 18529 -17894 18563 -17860
rect 18597 -17894 18631 -17860
rect 19139 -17894 19173 -17860
rect 19207 -17894 19241 -17860
rect 19275 -17894 19309 -17860
rect 19343 -17894 19377 -17860
rect 19411 -17894 19445 -17860
rect 19479 -17894 19513 -17860
rect 19547 -17894 19581 -17860
rect 19615 -17894 19649 -17860
rect 20157 -17894 20191 -17860
rect 20225 -17894 20259 -17860
rect 20293 -17894 20327 -17860
rect 20361 -17894 20395 -17860
rect 20429 -17894 20463 -17860
rect 20497 -17894 20531 -17860
rect 20565 -17894 20599 -17860
rect 20633 -17894 20667 -17860
rect 21175 -17894 21209 -17860
rect 21243 -17894 21277 -17860
rect 21311 -17894 21345 -17860
rect 21379 -17894 21413 -17860
rect 21447 -17894 21481 -17860
rect 21515 -17894 21549 -17860
rect 21583 -17894 21617 -17860
rect 21651 -17894 21685 -17860
rect 22193 -17894 22227 -17860
rect 22261 -17894 22295 -17860
rect 22329 -17894 22363 -17860
rect 22397 -17894 22431 -17860
rect 22465 -17894 22499 -17860
rect 22533 -17894 22567 -17860
rect 22601 -17894 22635 -17860
rect 22669 -17894 22703 -17860
rect -8913 -18092 -8879 -18058
rect -8845 -18092 -8811 -18058
rect -8777 -18092 -8743 -18058
rect -8709 -18092 -8675 -18058
rect -8641 -18092 -8607 -18058
rect -8573 -18092 -8539 -18058
rect -8505 -18092 -8471 -18058
rect -8437 -18092 -8403 -18058
rect -7895 -18092 -7861 -18058
rect -7827 -18092 -7793 -18058
rect -7759 -18092 -7725 -18058
rect -7691 -18092 -7657 -18058
rect -7623 -18092 -7589 -18058
rect -7555 -18092 -7521 -18058
rect -7487 -18092 -7453 -18058
rect -7419 -18092 -7385 -18058
rect -6877 -18092 -6843 -18058
rect -6809 -18092 -6775 -18058
rect -6741 -18092 -6707 -18058
rect -6673 -18092 -6639 -18058
rect -6605 -18092 -6571 -18058
rect -6537 -18092 -6503 -18058
rect -6469 -18092 -6435 -18058
rect -6401 -18092 -6367 -18058
rect -5859 -18092 -5825 -18058
rect -5791 -18092 -5757 -18058
rect -5723 -18092 -5689 -18058
rect -5655 -18092 -5621 -18058
rect -5587 -18092 -5553 -18058
rect -5519 -18092 -5485 -18058
rect -5451 -18092 -5417 -18058
rect -5383 -18092 -5349 -18058
rect -4841 -18092 -4807 -18058
rect -4773 -18092 -4739 -18058
rect -4705 -18092 -4671 -18058
rect -4637 -18092 -4603 -18058
rect -4569 -18092 -4535 -18058
rect -4501 -18092 -4467 -18058
rect -4433 -18092 -4399 -18058
rect -4365 -18092 -4331 -18058
rect -3823 -18092 -3789 -18058
rect -3755 -18092 -3721 -18058
rect -3687 -18092 -3653 -18058
rect -3619 -18092 -3585 -18058
rect -3551 -18092 -3517 -18058
rect -3483 -18092 -3449 -18058
rect -3415 -18092 -3381 -18058
rect -3347 -18092 -3313 -18058
rect -2805 -18092 -2771 -18058
rect -2737 -18092 -2703 -18058
rect -2669 -18092 -2635 -18058
rect -2601 -18092 -2567 -18058
rect -2533 -18092 -2499 -18058
rect -2465 -18092 -2431 -18058
rect -2397 -18092 -2363 -18058
rect -2329 -18092 -2295 -18058
rect -1787 -18092 -1753 -18058
rect -1719 -18092 -1685 -18058
rect -1651 -18092 -1617 -18058
rect -1583 -18092 -1549 -18058
rect -1515 -18092 -1481 -18058
rect -1447 -18092 -1413 -18058
rect -1379 -18092 -1345 -18058
rect -1311 -18092 -1277 -18058
rect -769 -18092 -735 -18058
rect -701 -18092 -667 -18058
rect -633 -18092 -599 -18058
rect -565 -18092 -531 -18058
rect -497 -18092 -463 -18058
rect -429 -18092 -395 -18058
rect -361 -18092 -327 -18058
rect -293 -18092 -259 -18058
rect -8913 -18200 -8879 -18166
rect -8845 -18200 -8811 -18166
rect -8777 -18200 -8743 -18166
rect -8709 -18200 -8675 -18166
rect -8641 -18200 -8607 -18166
rect -8573 -18200 -8539 -18166
rect -8505 -18200 -8471 -18166
rect -8437 -18200 -8403 -18166
rect -7895 -18200 -7861 -18166
rect -7827 -18200 -7793 -18166
rect -7759 -18200 -7725 -18166
rect -7691 -18200 -7657 -18166
rect -7623 -18200 -7589 -18166
rect -7555 -18200 -7521 -18166
rect -7487 -18200 -7453 -18166
rect -7419 -18200 -7385 -18166
rect -6877 -18200 -6843 -18166
rect -6809 -18200 -6775 -18166
rect -6741 -18200 -6707 -18166
rect -6673 -18200 -6639 -18166
rect -6605 -18200 -6571 -18166
rect -6537 -18200 -6503 -18166
rect -6469 -18200 -6435 -18166
rect -6401 -18200 -6367 -18166
rect -5859 -18200 -5825 -18166
rect -5791 -18200 -5757 -18166
rect -5723 -18200 -5689 -18166
rect -5655 -18200 -5621 -18166
rect -5587 -18200 -5553 -18166
rect -5519 -18200 -5485 -18166
rect -5451 -18200 -5417 -18166
rect -5383 -18200 -5349 -18166
rect -4841 -18200 -4807 -18166
rect -4773 -18200 -4739 -18166
rect -4705 -18200 -4671 -18166
rect -4637 -18200 -4603 -18166
rect -4569 -18200 -4535 -18166
rect -4501 -18200 -4467 -18166
rect -4433 -18200 -4399 -18166
rect -4365 -18200 -4331 -18166
rect -3823 -18200 -3789 -18166
rect -3755 -18200 -3721 -18166
rect -3687 -18200 -3653 -18166
rect -3619 -18200 -3585 -18166
rect -3551 -18200 -3517 -18166
rect -3483 -18200 -3449 -18166
rect -3415 -18200 -3381 -18166
rect -3347 -18200 -3313 -18166
rect -2805 -18200 -2771 -18166
rect -2737 -18200 -2703 -18166
rect -2669 -18200 -2635 -18166
rect -2601 -18200 -2567 -18166
rect -2533 -18200 -2499 -18166
rect -2465 -18200 -2431 -18166
rect -2397 -18200 -2363 -18166
rect -2329 -18200 -2295 -18166
rect -1787 -18200 -1753 -18166
rect -1719 -18200 -1685 -18166
rect -1651 -18200 -1617 -18166
rect -1583 -18200 -1549 -18166
rect -1515 -18200 -1481 -18166
rect -1447 -18200 -1413 -18166
rect -1379 -18200 -1345 -18166
rect -1311 -18200 -1277 -18166
rect -769 -18200 -735 -18166
rect -701 -18200 -667 -18166
rect -633 -18200 -599 -18166
rect -565 -18200 -531 -18166
rect -497 -18200 -463 -18166
rect -429 -18200 -395 -18166
rect -361 -18200 -327 -18166
rect -293 -18200 -259 -18166
rect 2851 -18604 2885 -18570
rect 2919 -18604 2953 -18570
rect 2987 -18604 3021 -18570
rect 3055 -18604 3089 -18570
rect 3123 -18604 3157 -18570
rect 3191 -18604 3225 -18570
rect 3259 -18604 3293 -18570
rect 3327 -18604 3361 -18570
rect 3869 -18604 3903 -18570
rect 3937 -18604 3971 -18570
rect 4005 -18604 4039 -18570
rect 4073 -18604 4107 -18570
rect 4141 -18604 4175 -18570
rect 4209 -18604 4243 -18570
rect 4277 -18604 4311 -18570
rect 4345 -18604 4379 -18570
rect 4887 -18604 4921 -18570
rect 4955 -18604 4989 -18570
rect 5023 -18604 5057 -18570
rect 5091 -18604 5125 -18570
rect 5159 -18604 5193 -18570
rect 5227 -18604 5261 -18570
rect 5295 -18604 5329 -18570
rect 5363 -18604 5397 -18570
rect 5905 -18604 5939 -18570
rect 5973 -18604 6007 -18570
rect 6041 -18604 6075 -18570
rect 6109 -18604 6143 -18570
rect 6177 -18604 6211 -18570
rect 6245 -18604 6279 -18570
rect 6313 -18604 6347 -18570
rect 6381 -18604 6415 -18570
rect 6923 -18604 6957 -18570
rect 6991 -18604 7025 -18570
rect 7059 -18604 7093 -18570
rect 7127 -18604 7161 -18570
rect 7195 -18604 7229 -18570
rect 7263 -18604 7297 -18570
rect 7331 -18604 7365 -18570
rect 7399 -18604 7433 -18570
rect 7941 -18604 7975 -18570
rect 8009 -18604 8043 -18570
rect 8077 -18604 8111 -18570
rect 8145 -18604 8179 -18570
rect 8213 -18604 8247 -18570
rect 8281 -18604 8315 -18570
rect 8349 -18604 8383 -18570
rect 8417 -18604 8451 -18570
rect 8959 -18604 8993 -18570
rect 9027 -18604 9061 -18570
rect 9095 -18604 9129 -18570
rect 9163 -18604 9197 -18570
rect 9231 -18604 9265 -18570
rect 9299 -18604 9333 -18570
rect 9367 -18604 9401 -18570
rect 9435 -18604 9469 -18570
rect 9977 -18604 10011 -18570
rect 10045 -18604 10079 -18570
rect 10113 -18604 10147 -18570
rect 10181 -18604 10215 -18570
rect 10249 -18604 10283 -18570
rect 10317 -18604 10351 -18570
rect 10385 -18604 10419 -18570
rect 10453 -18604 10487 -18570
rect 10995 -18604 11029 -18570
rect 11063 -18604 11097 -18570
rect 11131 -18604 11165 -18570
rect 11199 -18604 11233 -18570
rect 11267 -18604 11301 -18570
rect 11335 -18604 11369 -18570
rect 11403 -18604 11437 -18570
rect 11471 -18604 11505 -18570
rect 12013 -18604 12047 -18570
rect 12081 -18604 12115 -18570
rect 12149 -18604 12183 -18570
rect 12217 -18604 12251 -18570
rect 12285 -18604 12319 -18570
rect 12353 -18604 12387 -18570
rect 12421 -18604 12455 -18570
rect 12489 -18604 12523 -18570
rect 13031 -18604 13065 -18570
rect 13099 -18604 13133 -18570
rect 13167 -18604 13201 -18570
rect 13235 -18604 13269 -18570
rect 13303 -18604 13337 -18570
rect 13371 -18604 13405 -18570
rect 13439 -18604 13473 -18570
rect 13507 -18604 13541 -18570
rect 14049 -18604 14083 -18570
rect 14117 -18604 14151 -18570
rect 14185 -18604 14219 -18570
rect 14253 -18604 14287 -18570
rect 14321 -18604 14355 -18570
rect 14389 -18604 14423 -18570
rect 14457 -18604 14491 -18570
rect 14525 -18604 14559 -18570
rect 15067 -18604 15101 -18570
rect 15135 -18604 15169 -18570
rect 15203 -18604 15237 -18570
rect 15271 -18604 15305 -18570
rect 15339 -18604 15373 -18570
rect 15407 -18604 15441 -18570
rect 15475 -18604 15509 -18570
rect 15543 -18604 15577 -18570
rect 16085 -18604 16119 -18570
rect 16153 -18604 16187 -18570
rect 16221 -18604 16255 -18570
rect 16289 -18604 16323 -18570
rect 16357 -18604 16391 -18570
rect 16425 -18604 16459 -18570
rect 16493 -18604 16527 -18570
rect 16561 -18604 16595 -18570
rect 17103 -18604 17137 -18570
rect 17171 -18604 17205 -18570
rect 17239 -18604 17273 -18570
rect 17307 -18604 17341 -18570
rect 17375 -18604 17409 -18570
rect 17443 -18604 17477 -18570
rect 17511 -18604 17545 -18570
rect 17579 -18604 17613 -18570
rect 18121 -18604 18155 -18570
rect 18189 -18604 18223 -18570
rect 18257 -18604 18291 -18570
rect 18325 -18604 18359 -18570
rect 18393 -18604 18427 -18570
rect 18461 -18604 18495 -18570
rect 18529 -18604 18563 -18570
rect 18597 -18604 18631 -18570
rect 19139 -18604 19173 -18570
rect 19207 -18604 19241 -18570
rect 19275 -18604 19309 -18570
rect 19343 -18604 19377 -18570
rect 19411 -18604 19445 -18570
rect 19479 -18604 19513 -18570
rect 19547 -18604 19581 -18570
rect 19615 -18604 19649 -18570
rect 20157 -18604 20191 -18570
rect 20225 -18604 20259 -18570
rect 20293 -18604 20327 -18570
rect 20361 -18604 20395 -18570
rect 20429 -18604 20463 -18570
rect 20497 -18604 20531 -18570
rect 20565 -18604 20599 -18570
rect 20633 -18604 20667 -18570
rect 21175 -18604 21209 -18570
rect 21243 -18604 21277 -18570
rect 21311 -18604 21345 -18570
rect 21379 -18604 21413 -18570
rect 21447 -18604 21481 -18570
rect 21515 -18604 21549 -18570
rect 21583 -18604 21617 -18570
rect 21651 -18604 21685 -18570
rect 22193 -18604 22227 -18570
rect 22261 -18604 22295 -18570
rect 22329 -18604 22363 -18570
rect 22397 -18604 22431 -18570
rect 22465 -18604 22499 -18570
rect 22533 -18604 22567 -18570
rect 22601 -18604 22635 -18570
rect 22669 -18604 22703 -18570
rect -8913 -18910 -8879 -18876
rect -8845 -18910 -8811 -18876
rect -8777 -18910 -8743 -18876
rect -8709 -18910 -8675 -18876
rect -8641 -18910 -8607 -18876
rect -8573 -18910 -8539 -18876
rect -8505 -18910 -8471 -18876
rect -8437 -18910 -8403 -18876
rect -7895 -18910 -7861 -18876
rect -7827 -18910 -7793 -18876
rect -7759 -18910 -7725 -18876
rect -7691 -18910 -7657 -18876
rect -7623 -18910 -7589 -18876
rect -7555 -18910 -7521 -18876
rect -7487 -18910 -7453 -18876
rect -7419 -18910 -7385 -18876
rect -6877 -18910 -6843 -18876
rect -6809 -18910 -6775 -18876
rect -6741 -18910 -6707 -18876
rect -6673 -18910 -6639 -18876
rect -6605 -18910 -6571 -18876
rect -6537 -18910 -6503 -18876
rect -6469 -18910 -6435 -18876
rect -6401 -18910 -6367 -18876
rect -5859 -18910 -5825 -18876
rect -5791 -18910 -5757 -18876
rect -5723 -18910 -5689 -18876
rect -5655 -18910 -5621 -18876
rect -5587 -18910 -5553 -18876
rect -5519 -18910 -5485 -18876
rect -5451 -18910 -5417 -18876
rect -5383 -18910 -5349 -18876
rect -4841 -18910 -4807 -18876
rect -4773 -18910 -4739 -18876
rect -4705 -18910 -4671 -18876
rect -4637 -18910 -4603 -18876
rect -4569 -18910 -4535 -18876
rect -4501 -18910 -4467 -18876
rect -4433 -18910 -4399 -18876
rect -4365 -18910 -4331 -18876
rect -3823 -18910 -3789 -18876
rect -3755 -18910 -3721 -18876
rect -3687 -18910 -3653 -18876
rect -3619 -18910 -3585 -18876
rect -3551 -18910 -3517 -18876
rect -3483 -18910 -3449 -18876
rect -3415 -18910 -3381 -18876
rect -3347 -18910 -3313 -18876
rect -2805 -18910 -2771 -18876
rect -2737 -18910 -2703 -18876
rect -2669 -18910 -2635 -18876
rect -2601 -18910 -2567 -18876
rect -2533 -18910 -2499 -18876
rect -2465 -18910 -2431 -18876
rect -2397 -18910 -2363 -18876
rect -2329 -18910 -2295 -18876
rect -1787 -18910 -1753 -18876
rect -1719 -18910 -1685 -18876
rect -1651 -18910 -1617 -18876
rect -1583 -18910 -1549 -18876
rect -1515 -18910 -1481 -18876
rect -1447 -18910 -1413 -18876
rect -1379 -18910 -1345 -18876
rect -1311 -18910 -1277 -18876
rect -769 -18910 -735 -18876
rect -701 -18910 -667 -18876
rect -633 -18910 -599 -18876
rect -565 -18910 -531 -18876
rect -497 -18910 -463 -18876
rect -429 -18910 -395 -18876
rect -361 -18910 -327 -18876
rect -293 -18910 -259 -18876
rect 2851 -19126 2885 -19092
rect 2919 -19126 2953 -19092
rect 2987 -19126 3021 -19092
rect 3055 -19126 3089 -19092
rect 3123 -19126 3157 -19092
rect 3191 -19126 3225 -19092
rect 3259 -19126 3293 -19092
rect 3327 -19126 3361 -19092
rect 3869 -19126 3903 -19092
rect 3937 -19126 3971 -19092
rect 4005 -19126 4039 -19092
rect 4073 -19126 4107 -19092
rect 4141 -19126 4175 -19092
rect 4209 -19126 4243 -19092
rect 4277 -19126 4311 -19092
rect 4345 -19126 4379 -19092
rect 4887 -19126 4921 -19092
rect 4955 -19126 4989 -19092
rect 5023 -19126 5057 -19092
rect 5091 -19126 5125 -19092
rect 5159 -19126 5193 -19092
rect 5227 -19126 5261 -19092
rect 5295 -19126 5329 -19092
rect 5363 -19126 5397 -19092
rect 5905 -19126 5939 -19092
rect 5973 -19126 6007 -19092
rect 6041 -19126 6075 -19092
rect 6109 -19126 6143 -19092
rect 6177 -19126 6211 -19092
rect 6245 -19126 6279 -19092
rect 6313 -19126 6347 -19092
rect 6381 -19126 6415 -19092
rect 6923 -19126 6957 -19092
rect 6991 -19126 7025 -19092
rect 7059 -19126 7093 -19092
rect 7127 -19126 7161 -19092
rect 7195 -19126 7229 -19092
rect 7263 -19126 7297 -19092
rect 7331 -19126 7365 -19092
rect 7399 -19126 7433 -19092
rect 7941 -19126 7975 -19092
rect 8009 -19126 8043 -19092
rect 8077 -19126 8111 -19092
rect 8145 -19126 8179 -19092
rect 8213 -19126 8247 -19092
rect 8281 -19126 8315 -19092
rect 8349 -19126 8383 -19092
rect 8417 -19126 8451 -19092
rect 8959 -19126 8993 -19092
rect 9027 -19126 9061 -19092
rect 9095 -19126 9129 -19092
rect 9163 -19126 9197 -19092
rect 9231 -19126 9265 -19092
rect 9299 -19126 9333 -19092
rect 9367 -19126 9401 -19092
rect 9435 -19126 9469 -19092
rect 9977 -19126 10011 -19092
rect 10045 -19126 10079 -19092
rect 10113 -19126 10147 -19092
rect 10181 -19126 10215 -19092
rect 10249 -19126 10283 -19092
rect 10317 -19126 10351 -19092
rect 10385 -19126 10419 -19092
rect 10453 -19126 10487 -19092
rect 10995 -19126 11029 -19092
rect 11063 -19126 11097 -19092
rect 11131 -19126 11165 -19092
rect 11199 -19126 11233 -19092
rect 11267 -19126 11301 -19092
rect 11335 -19126 11369 -19092
rect 11403 -19126 11437 -19092
rect 11471 -19126 11505 -19092
rect 12013 -19126 12047 -19092
rect 12081 -19126 12115 -19092
rect 12149 -19126 12183 -19092
rect 12217 -19126 12251 -19092
rect 12285 -19126 12319 -19092
rect 12353 -19126 12387 -19092
rect 12421 -19126 12455 -19092
rect 12489 -19126 12523 -19092
rect 13031 -19126 13065 -19092
rect 13099 -19126 13133 -19092
rect 13167 -19126 13201 -19092
rect 13235 -19126 13269 -19092
rect 13303 -19126 13337 -19092
rect 13371 -19126 13405 -19092
rect 13439 -19126 13473 -19092
rect 13507 -19126 13541 -19092
rect 14049 -19126 14083 -19092
rect 14117 -19126 14151 -19092
rect 14185 -19126 14219 -19092
rect 14253 -19126 14287 -19092
rect 14321 -19126 14355 -19092
rect 14389 -19126 14423 -19092
rect 14457 -19126 14491 -19092
rect 14525 -19126 14559 -19092
rect 15067 -19126 15101 -19092
rect 15135 -19126 15169 -19092
rect 15203 -19126 15237 -19092
rect 15271 -19126 15305 -19092
rect 15339 -19126 15373 -19092
rect 15407 -19126 15441 -19092
rect 15475 -19126 15509 -19092
rect 15543 -19126 15577 -19092
rect 16085 -19126 16119 -19092
rect 16153 -19126 16187 -19092
rect 16221 -19126 16255 -19092
rect 16289 -19126 16323 -19092
rect 16357 -19126 16391 -19092
rect 16425 -19126 16459 -19092
rect 16493 -19126 16527 -19092
rect 16561 -19126 16595 -19092
rect 17103 -19126 17137 -19092
rect 17171 -19126 17205 -19092
rect 17239 -19126 17273 -19092
rect 17307 -19126 17341 -19092
rect 17375 -19126 17409 -19092
rect 17443 -19126 17477 -19092
rect 17511 -19126 17545 -19092
rect 17579 -19126 17613 -19092
rect 18121 -19126 18155 -19092
rect 18189 -19126 18223 -19092
rect 18257 -19126 18291 -19092
rect 18325 -19126 18359 -19092
rect 18393 -19126 18427 -19092
rect 18461 -19126 18495 -19092
rect 18529 -19126 18563 -19092
rect 18597 -19126 18631 -19092
rect 19139 -19126 19173 -19092
rect 19207 -19126 19241 -19092
rect 19275 -19126 19309 -19092
rect 19343 -19126 19377 -19092
rect 19411 -19126 19445 -19092
rect 19479 -19126 19513 -19092
rect 19547 -19126 19581 -19092
rect 19615 -19126 19649 -19092
rect 20157 -19126 20191 -19092
rect 20225 -19126 20259 -19092
rect 20293 -19126 20327 -19092
rect 20361 -19126 20395 -19092
rect 20429 -19126 20463 -19092
rect 20497 -19126 20531 -19092
rect 20565 -19126 20599 -19092
rect 20633 -19126 20667 -19092
rect 21175 -19126 21209 -19092
rect 21243 -19126 21277 -19092
rect 21311 -19126 21345 -19092
rect 21379 -19126 21413 -19092
rect 21447 -19126 21481 -19092
rect 21515 -19126 21549 -19092
rect 21583 -19126 21617 -19092
rect 21651 -19126 21685 -19092
rect 22193 -19126 22227 -19092
rect 22261 -19126 22295 -19092
rect 22329 -19126 22363 -19092
rect 22397 -19126 22431 -19092
rect 22465 -19126 22499 -19092
rect 22533 -19126 22567 -19092
rect 22601 -19126 22635 -19092
rect 22669 -19126 22703 -19092
rect 2851 -19836 2885 -19802
rect 2919 -19836 2953 -19802
rect 2987 -19836 3021 -19802
rect 3055 -19836 3089 -19802
rect 3123 -19836 3157 -19802
rect 3191 -19836 3225 -19802
rect 3259 -19836 3293 -19802
rect 3327 -19836 3361 -19802
rect 3869 -19836 3903 -19802
rect 3937 -19836 3971 -19802
rect 4005 -19836 4039 -19802
rect 4073 -19836 4107 -19802
rect 4141 -19836 4175 -19802
rect 4209 -19836 4243 -19802
rect 4277 -19836 4311 -19802
rect 4345 -19836 4379 -19802
rect 4887 -19836 4921 -19802
rect 4955 -19836 4989 -19802
rect 5023 -19836 5057 -19802
rect 5091 -19836 5125 -19802
rect 5159 -19836 5193 -19802
rect 5227 -19836 5261 -19802
rect 5295 -19836 5329 -19802
rect 5363 -19836 5397 -19802
rect 5905 -19836 5939 -19802
rect 5973 -19836 6007 -19802
rect 6041 -19836 6075 -19802
rect 6109 -19836 6143 -19802
rect 6177 -19836 6211 -19802
rect 6245 -19836 6279 -19802
rect 6313 -19836 6347 -19802
rect 6381 -19836 6415 -19802
rect 6923 -19836 6957 -19802
rect 6991 -19836 7025 -19802
rect 7059 -19836 7093 -19802
rect 7127 -19836 7161 -19802
rect 7195 -19836 7229 -19802
rect 7263 -19836 7297 -19802
rect 7331 -19836 7365 -19802
rect 7399 -19836 7433 -19802
rect 7941 -19836 7975 -19802
rect 8009 -19836 8043 -19802
rect 8077 -19836 8111 -19802
rect 8145 -19836 8179 -19802
rect 8213 -19836 8247 -19802
rect 8281 -19836 8315 -19802
rect 8349 -19836 8383 -19802
rect 8417 -19836 8451 -19802
rect 8959 -19836 8993 -19802
rect 9027 -19836 9061 -19802
rect 9095 -19836 9129 -19802
rect 9163 -19836 9197 -19802
rect 9231 -19836 9265 -19802
rect 9299 -19836 9333 -19802
rect 9367 -19836 9401 -19802
rect 9435 -19836 9469 -19802
rect 9977 -19836 10011 -19802
rect 10045 -19836 10079 -19802
rect 10113 -19836 10147 -19802
rect 10181 -19836 10215 -19802
rect 10249 -19836 10283 -19802
rect 10317 -19836 10351 -19802
rect 10385 -19836 10419 -19802
rect 10453 -19836 10487 -19802
rect 10995 -19836 11029 -19802
rect 11063 -19836 11097 -19802
rect 11131 -19836 11165 -19802
rect 11199 -19836 11233 -19802
rect 11267 -19836 11301 -19802
rect 11335 -19836 11369 -19802
rect 11403 -19836 11437 -19802
rect 11471 -19836 11505 -19802
rect 12013 -19836 12047 -19802
rect 12081 -19836 12115 -19802
rect 12149 -19836 12183 -19802
rect 12217 -19836 12251 -19802
rect 12285 -19836 12319 -19802
rect 12353 -19836 12387 -19802
rect 12421 -19836 12455 -19802
rect 12489 -19836 12523 -19802
rect 13031 -19836 13065 -19802
rect 13099 -19836 13133 -19802
rect 13167 -19836 13201 -19802
rect 13235 -19836 13269 -19802
rect 13303 -19836 13337 -19802
rect 13371 -19836 13405 -19802
rect 13439 -19836 13473 -19802
rect 13507 -19836 13541 -19802
rect 14049 -19836 14083 -19802
rect 14117 -19836 14151 -19802
rect 14185 -19836 14219 -19802
rect 14253 -19836 14287 -19802
rect 14321 -19836 14355 -19802
rect 14389 -19836 14423 -19802
rect 14457 -19836 14491 -19802
rect 14525 -19836 14559 -19802
rect 15067 -19836 15101 -19802
rect 15135 -19836 15169 -19802
rect 15203 -19836 15237 -19802
rect 15271 -19836 15305 -19802
rect 15339 -19836 15373 -19802
rect 15407 -19836 15441 -19802
rect 15475 -19836 15509 -19802
rect 15543 -19836 15577 -19802
rect 16085 -19836 16119 -19802
rect 16153 -19836 16187 -19802
rect 16221 -19836 16255 -19802
rect 16289 -19836 16323 -19802
rect 16357 -19836 16391 -19802
rect 16425 -19836 16459 -19802
rect 16493 -19836 16527 -19802
rect 16561 -19836 16595 -19802
rect 17103 -19836 17137 -19802
rect 17171 -19836 17205 -19802
rect 17239 -19836 17273 -19802
rect 17307 -19836 17341 -19802
rect 17375 -19836 17409 -19802
rect 17443 -19836 17477 -19802
rect 17511 -19836 17545 -19802
rect 17579 -19836 17613 -19802
rect 18121 -19836 18155 -19802
rect 18189 -19836 18223 -19802
rect 18257 -19836 18291 -19802
rect 18325 -19836 18359 -19802
rect 18393 -19836 18427 -19802
rect 18461 -19836 18495 -19802
rect 18529 -19836 18563 -19802
rect 18597 -19836 18631 -19802
rect 19139 -19836 19173 -19802
rect 19207 -19836 19241 -19802
rect 19275 -19836 19309 -19802
rect 19343 -19836 19377 -19802
rect 19411 -19836 19445 -19802
rect 19479 -19836 19513 -19802
rect 19547 -19836 19581 -19802
rect 19615 -19836 19649 -19802
rect 20157 -19836 20191 -19802
rect 20225 -19836 20259 -19802
rect 20293 -19836 20327 -19802
rect 20361 -19836 20395 -19802
rect 20429 -19836 20463 -19802
rect 20497 -19836 20531 -19802
rect 20565 -19836 20599 -19802
rect 20633 -19836 20667 -19802
rect 21175 -19836 21209 -19802
rect 21243 -19836 21277 -19802
rect 21311 -19836 21345 -19802
rect 21379 -19836 21413 -19802
rect 21447 -19836 21481 -19802
rect 21515 -19836 21549 -19802
rect 21583 -19836 21617 -19802
rect 21651 -19836 21685 -19802
rect 22193 -19836 22227 -19802
rect 22261 -19836 22295 -19802
rect 22329 -19836 22363 -19802
rect 22397 -19836 22431 -19802
rect 22465 -19836 22499 -19802
rect 22533 -19836 22567 -19802
rect 22601 -19836 22635 -19802
rect 22669 -19836 22703 -19802
rect 2851 -20360 2885 -20326
rect 2919 -20360 2953 -20326
rect 2987 -20360 3021 -20326
rect 3055 -20360 3089 -20326
rect 3123 -20360 3157 -20326
rect 3191 -20360 3225 -20326
rect 3259 -20360 3293 -20326
rect 3327 -20360 3361 -20326
rect 3869 -20360 3903 -20326
rect 3937 -20360 3971 -20326
rect 4005 -20360 4039 -20326
rect 4073 -20360 4107 -20326
rect 4141 -20360 4175 -20326
rect 4209 -20360 4243 -20326
rect 4277 -20360 4311 -20326
rect 4345 -20360 4379 -20326
rect 4887 -20360 4921 -20326
rect 4955 -20360 4989 -20326
rect 5023 -20360 5057 -20326
rect 5091 -20360 5125 -20326
rect 5159 -20360 5193 -20326
rect 5227 -20360 5261 -20326
rect 5295 -20360 5329 -20326
rect 5363 -20360 5397 -20326
rect 5905 -20360 5939 -20326
rect 5973 -20360 6007 -20326
rect 6041 -20360 6075 -20326
rect 6109 -20360 6143 -20326
rect 6177 -20360 6211 -20326
rect 6245 -20360 6279 -20326
rect 6313 -20360 6347 -20326
rect 6381 -20360 6415 -20326
rect 6923 -20360 6957 -20326
rect 6991 -20360 7025 -20326
rect 7059 -20360 7093 -20326
rect 7127 -20360 7161 -20326
rect 7195 -20360 7229 -20326
rect 7263 -20360 7297 -20326
rect 7331 -20360 7365 -20326
rect 7399 -20360 7433 -20326
rect 7941 -20360 7975 -20326
rect 8009 -20360 8043 -20326
rect 8077 -20360 8111 -20326
rect 8145 -20360 8179 -20326
rect 8213 -20360 8247 -20326
rect 8281 -20360 8315 -20326
rect 8349 -20360 8383 -20326
rect 8417 -20360 8451 -20326
rect 8959 -20360 8993 -20326
rect 9027 -20360 9061 -20326
rect 9095 -20360 9129 -20326
rect 9163 -20360 9197 -20326
rect 9231 -20360 9265 -20326
rect 9299 -20360 9333 -20326
rect 9367 -20360 9401 -20326
rect 9435 -20360 9469 -20326
rect 9977 -20360 10011 -20326
rect 10045 -20360 10079 -20326
rect 10113 -20360 10147 -20326
rect 10181 -20360 10215 -20326
rect 10249 -20360 10283 -20326
rect 10317 -20360 10351 -20326
rect 10385 -20360 10419 -20326
rect 10453 -20360 10487 -20326
rect 10995 -20360 11029 -20326
rect 11063 -20360 11097 -20326
rect 11131 -20360 11165 -20326
rect 11199 -20360 11233 -20326
rect 11267 -20360 11301 -20326
rect 11335 -20360 11369 -20326
rect 11403 -20360 11437 -20326
rect 11471 -20360 11505 -20326
rect 12013 -20360 12047 -20326
rect 12081 -20360 12115 -20326
rect 12149 -20360 12183 -20326
rect 12217 -20360 12251 -20326
rect 12285 -20360 12319 -20326
rect 12353 -20360 12387 -20326
rect 12421 -20360 12455 -20326
rect 12489 -20360 12523 -20326
rect 13031 -20360 13065 -20326
rect 13099 -20360 13133 -20326
rect 13167 -20360 13201 -20326
rect 13235 -20360 13269 -20326
rect 13303 -20360 13337 -20326
rect 13371 -20360 13405 -20326
rect 13439 -20360 13473 -20326
rect 13507 -20360 13541 -20326
rect 14049 -20360 14083 -20326
rect 14117 -20360 14151 -20326
rect 14185 -20360 14219 -20326
rect 14253 -20360 14287 -20326
rect 14321 -20360 14355 -20326
rect 14389 -20360 14423 -20326
rect 14457 -20360 14491 -20326
rect 14525 -20360 14559 -20326
rect 15067 -20360 15101 -20326
rect 15135 -20360 15169 -20326
rect 15203 -20360 15237 -20326
rect 15271 -20360 15305 -20326
rect 15339 -20360 15373 -20326
rect 15407 -20360 15441 -20326
rect 15475 -20360 15509 -20326
rect 15543 -20360 15577 -20326
rect 16085 -20360 16119 -20326
rect 16153 -20360 16187 -20326
rect 16221 -20360 16255 -20326
rect 16289 -20360 16323 -20326
rect 16357 -20360 16391 -20326
rect 16425 -20360 16459 -20326
rect 16493 -20360 16527 -20326
rect 16561 -20360 16595 -20326
rect 17103 -20360 17137 -20326
rect 17171 -20360 17205 -20326
rect 17239 -20360 17273 -20326
rect 17307 -20360 17341 -20326
rect 17375 -20360 17409 -20326
rect 17443 -20360 17477 -20326
rect 17511 -20360 17545 -20326
rect 17579 -20360 17613 -20326
rect 18121 -20360 18155 -20326
rect 18189 -20360 18223 -20326
rect 18257 -20360 18291 -20326
rect 18325 -20360 18359 -20326
rect 18393 -20360 18427 -20326
rect 18461 -20360 18495 -20326
rect 18529 -20360 18563 -20326
rect 18597 -20360 18631 -20326
rect 19139 -20360 19173 -20326
rect 19207 -20360 19241 -20326
rect 19275 -20360 19309 -20326
rect 19343 -20360 19377 -20326
rect 19411 -20360 19445 -20326
rect 19479 -20360 19513 -20326
rect 19547 -20360 19581 -20326
rect 19615 -20360 19649 -20326
rect 20157 -20360 20191 -20326
rect 20225 -20360 20259 -20326
rect 20293 -20360 20327 -20326
rect 20361 -20360 20395 -20326
rect 20429 -20360 20463 -20326
rect 20497 -20360 20531 -20326
rect 20565 -20360 20599 -20326
rect 20633 -20360 20667 -20326
rect 21175 -20360 21209 -20326
rect 21243 -20360 21277 -20326
rect 21311 -20360 21345 -20326
rect 21379 -20360 21413 -20326
rect 21447 -20360 21481 -20326
rect 21515 -20360 21549 -20326
rect 21583 -20360 21617 -20326
rect 21651 -20360 21685 -20326
rect 22193 -20360 22227 -20326
rect 22261 -20360 22295 -20326
rect 22329 -20360 22363 -20326
rect 22397 -20360 22431 -20326
rect 22465 -20360 22499 -20326
rect 22533 -20360 22567 -20326
rect 22601 -20360 22635 -20326
rect 22669 -20360 22703 -20326
rect 2851 -21070 2885 -21036
rect 2919 -21070 2953 -21036
rect 2987 -21070 3021 -21036
rect 3055 -21070 3089 -21036
rect 3123 -21070 3157 -21036
rect 3191 -21070 3225 -21036
rect 3259 -21070 3293 -21036
rect 3327 -21070 3361 -21036
rect 3869 -21070 3903 -21036
rect 3937 -21070 3971 -21036
rect 4005 -21070 4039 -21036
rect 4073 -21070 4107 -21036
rect 4141 -21070 4175 -21036
rect 4209 -21070 4243 -21036
rect 4277 -21070 4311 -21036
rect 4345 -21070 4379 -21036
rect 4887 -21070 4921 -21036
rect 4955 -21070 4989 -21036
rect 5023 -21070 5057 -21036
rect 5091 -21070 5125 -21036
rect 5159 -21070 5193 -21036
rect 5227 -21070 5261 -21036
rect 5295 -21070 5329 -21036
rect 5363 -21070 5397 -21036
rect 5905 -21070 5939 -21036
rect 5973 -21070 6007 -21036
rect 6041 -21070 6075 -21036
rect 6109 -21070 6143 -21036
rect 6177 -21070 6211 -21036
rect 6245 -21070 6279 -21036
rect 6313 -21070 6347 -21036
rect 6381 -21070 6415 -21036
rect 6923 -21070 6957 -21036
rect 6991 -21070 7025 -21036
rect 7059 -21070 7093 -21036
rect 7127 -21070 7161 -21036
rect 7195 -21070 7229 -21036
rect 7263 -21070 7297 -21036
rect 7331 -21070 7365 -21036
rect 7399 -21070 7433 -21036
rect 7941 -21070 7975 -21036
rect 8009 -21070 8043 -21036
rect 8077 -21070 8111 -21036
rect 8145 -21070 8179 -21036
rect 8213 -21070 8247 -21036
rect 8281 -21070 8315 -21036
rect 8349 -21070 8383 -21036
rect 8417 -21070 8451 -21036
rect 8959 -21070 8993 -21036
rect 9027 -21070 9061 -21036
rect 9095 -21070 9129 -21036
rect 9163 -21070 9197 -21036
rect 9231 -21070 9265 -21036
rect 9299 -21070 9333 -21036
rect 9367 -21070 9401 -21036
rect 9435 -21070 9469 -21036
rect 9977 -21070 10011 -21036
rect 10045 -21070 10079 -21036
rect 10113 -21070 10147 -21036
rect 10181 -21070 10215 -21036
rect 10249 -21070 10283 -21036
rect 10317 -21070 10351 -21036
rect 10385 -21070 10419 -21036
rect 10453 -21070 10487 -21036
rect 10995 -21070 11029 -21036
rect 11063 -21070 11097 -21036
rect 11131 -21070 11165 -21036
rect 11199 -21070 11233 -21036
rect 11267 -21070 11301 -21036
rect 11335 -21070 11369 -21036
rect 11403 -21070 11437 -21036
rect 11471 -21070 11505 -21036
rect 12013 -21070 12047 -21036
rect 12081 -21070 12115 -21036
rect 12149 -21070 12183 -21036
rect 12217 -21070 12251 -21036
rect 12285 -21070 12319 -21036
rect 12353 -21070 12387 -21036
rect 12421 -21070 12455 -21036
rect 12489 -21070 12523 -21036
rect 13031 -21070 13065 -21036
rect 13099 -21070 13133 -21036
rect 13167 -21070 13201 -21036
rect 13235 -21070 13269 -21036
rect 13303 -21070 13337 -21036
rect 13371 -21070 13405 -21036
rect 13439 -21070 13473 -21036
rect 13507 -21070 13541 -21036
rect 14049 -21070 14083 -21036
rect 14117 -21070 14151 -21036
rect 14185 -21070 14219 -21036
rect 14253 -21070 14287 -21036
rect 14321 -21070 14355 -21036
rect 14389 -21070 14423 -21036
rect 14457 -21070 14491 -21036
rect 14525 -21070 14559 -21036
rect 15067 -21070 15101 -21036
rect 15135 -21070 15169 -21036
rect 15203 -21070 15237 -21036
rect 15271 -21070 15305 -21036
rect 15339 -21070 15373 -21036
rect 15407 -21070 15441 -21036
rect 15475 -21070 15509 -21036
rect 15543 -21070 15577 -21036
rect 16085 -21070 16119 -21036
rect 16153 -21070 16187 -21036
rect 16221 -21070 16255 -21036
rect 16289 -21070 16323 -21036
rect 16357 -21070 16391 -21036
rect 16425 -21070 16459 -21036
rect 16493 -21070 16527 -21036
rect 16561 -21070 16595 -21036
rect 17103 -21070 17137 -21036
rect 17171 -21070 17205 -21036
rect 17239 -21070 17273 -21036
rect 17307 -21070 17341 -21036
rect 17375 -21070 17409 -21036
rect 17443 -21070 17477 -21036
rect 17511 -21070 17545 -21036
rect 17579 -21070 17613 -21036
rect 18121 -21070 18155 -21036
rect 18189 -21070 18223 -21036
rect 18257 -21070 18291 -21036
rect 18325 -21070 18359 -21036
rect 18393 -21070 18427 -21036
rect 18461 -21070 18495 -21036
rect 18529 -21070 18563 -21036
rect 18597 -21070 18631 -21036
rect 19139 -21070 19173 -21036
rect 19207 -21070 19241 -21036
rect 19275 -21070 19309 -21036
rect 19343 -21070 19377 -21036
rect 19411 -21070 19445 -21036
rect 19479 -21070 19513 -21036
rect 19547 -21070 19581 -21036
rect 19615 -21070 19649 -21036
rect 20157 -21070 20191 -21036
rect 20225 -21070 20259 -21036
rect 20293 -21070 20327 -21036
rect 20361 -21070 20395 -21036
rect 20429 -21070 20463 -21036
rect 20497 -21070 20531 -21036
rect 20565 -21070 20599 -21036
rect 20633 -21070 20667 -21036
rect 21175 -21070 21209 -21036
rect 21243 -21070 21277 -21036
rect 21311 -21070 21345 -21036
rect 21379 -21070 21413 -21036
rect 21447 -21070 21481 -21036
rect 21515 -21070 21549 -21036
rect 21583 -21070 21617 -21036
rect 21651 -21070 21685 -21036
rect 22193 -21070 22227 -21036
rect 22261 -21070 22295 -21036
rect 22329 -21070 22363 -21036
rect 22397 -21070 22431 -21036
rect 22465 -21070 22499 -21036
rect 22533 -21070 22567 -21036
rect 22601 -21070 22635 -21036
rect 22669 -21070 22703 -21036
rect 2851 -21594 2885 -21560
rect 2919 -21594 2953 -21560
rect 2987 -21594 3021 -21560
rect 3055 -21594 3089 -21560
rect 3123 -21594 3157 -21560
rect 3191 -21594 3225 -21560
rect 3259 -21594 3293 -21560
rect 3327 -21594 3361 -21560
rect 3869 -21594 3903 -21560
rect 3937 -21594 3971 -21560
rect 4005 -21594 4039 -21560
rect 4073 -21594 4107 -21560
rect 4141 -21594 4175 -21560
rect 4209 -21594 4243 -21560
rect 4277 -21594 4311 -21560
rect 4345 -21594 4379 -21560
rect 4887 -21594 4921 -21560
rect 4955 -21594 4989 -21560
rect 5023 -21594 5057 -21560
rect 5091 -21594 5125 -21560
rect 5159 -21594 5193 -21560
rect 5227 -21594 5261 -21560
rect 5295 -21594 5329 -21560
rect 5363 -21594 5397 -21560
rect 5905 -21594 5939 -21560
rect 5973 -21594 6007 -21560
rect 6041 -21594 6075 -21560
rect 6109 -21594 6143 -21560
rect 6177 -21594 6211 -21560
rect 6245 -21594 6279 -21560
rect 6313 -21594 6347 -21560
rect 6381 -21594 6415 -21560
rect 6923 -21594 6957 -21560
rect 6991 -21594 7025 -21560
rect 7059 -21594 7093 -21560
rect 7127 -21594 7161 -21560
rect 7195 -21594 7229 -21560
rect 7263 -21594 7297 -21560
rect 7331 -21594 7365 -21560
rect 7399 -21594 7433 -21560
rect 7941 -21594 7975 -21560
rect 8009 -21594 8043 -21560
rect 8077 -21594 8111 -21560
rect 8145 -21594 8179 -21560
rect 8213 -21594 8247 -21560
rect 8281 -21594 8315 -21560
rect 8349 -21594 8383 -21560
rect 8417 -21594 8451 -21560
rect 8959 -21594 8993 -21560
rect 9027 -21594 9061 -21560
rect 9095 -21594 9129 -21560
rect 9163 -21594 9197 -21560
rect 9231 -21594 9265 -21560
rect 9299 -21594 9333 -21560
rect 9367 -21594 9401 -21560
rect 9435 -21594 9469 -21560
rect 9977 -21594 10011 -21560
rect 10045 -21594 10079 -21560
rect 10113 -21594 10147 -21560
rect 10181 -21594 10215 -21560
rect 10249 -21594 10283 -21560
rect 10317 -21594 10351 -21560
rect 10385 -21594 10419 -21560
rect 10453 -21594 10487 -21560
rect 10995 -21594 11029 -21560
rect 11063 -21594 11097 -21560
rect 11131 -21594 11165 -21560
rect 11199 -21594 11233 -21560
rect 11267 -21594 11301 -21560
rect 11335 -21594 11369 -21560
rect 11403 -21594 11437 -21560
rect 11471 -21594 11505 -21560
rect 12013 -21594 12047 -21560
rect 12081 -21594 12115 -21560
rect 12149 -21594 12183 -21560
rect 12217 -21594 12251 -21560
rect 12285 -21594 12319 -21560
rect 12353 -21594 12387 -21560
rect 12421 -21594 12455 -21560
rect 12489 -21594 12523 -21560
rect 13031 -21594 13065 -21560
rect 13099 -21594 13133 -21560
rect 13167 -21594 13201 -21560
rect 13235 -21594 13269 -21560
rect 13303 -21594 13337 -21560
rect 13371 -21594 13405 -21560
rect 13439 -21594 13473 -21560
rect 13507 -21594 13541 -21560
rect 14049 -21594 14083 -21560
rect 14117 -21594 14151 -21560
rect 14185 -21594 14219 -21560
rect 14253 -21594 14287 -21560
rect 14321 -21594 14355 -21560
rect 14389 -21594 14423 -21560
rect 14457 -21594 14491 -21560
rect 14525 -21594 14559 -21560
rect 15067 -21594 15101 -21560
rect 15135 -21594 15169 -21560
rect 15203 -21594 15237 -21560
rect 15271 -21594 15305 -21560
rect 15339 -21594 15373 -21560
rect 15407 -21594 15441 -21560
rect 15475 -21594 15509 -21560
rect 15543 -21594 15577 -21560
rect 16085 -21594 16119 -21560
rect 16153 -21594 16187 -21560
rect 16221 -21594 16255 -21560
rect 16289 -21594 16323 -21560
rect 16357 -21594 16391 -21560
rect 16425 -21594 16459 -21560
rect 16493 -21594 16527 -21560
rect 16561 -21594 16595 -21560
rect 17103 -21594 17137 -21560
rect 17171 -21594 17205 -21560
rect 17239 -21594 17273 -21560
rect 17307 -21594 17341 -21560
rect 17375 -21594 17409 -21560
rect 17443 -21594 17477 -21560
rect 17511 -21594 17545 -21560
rect 17579 -21594 17613 -21560
rect 18121 -21594 18155 -21560
rect 18189 -21594 18223 -21560
rect 18257 -21594 18291 -21560
rect 18325 -21594 18359 -21560
rect 18393 -21594 18427 -21560
rect 18461 -21594 18495 -21560
rect 18529 -21594 18563 -21560
rect 18597 -21594 18631 -21560
rect 19139 -21594 19173 -21560
rect 19207 -21594 19241 -21560
rect 19275 -21594 19309 -21560
rect 19343 -21594 19377 -21560
rect 19411 -21594 19445 -21560
rect 19479 -21594 19513 -21560
rect 19547 -21594 19581 -21560
rect 19615 -21594 19649 -21560
rect 20157 -21594 20191 -21560
rect 20225 -21594 20259 -21560
rect 20293 -21594 20327 -21560
rect 20361 -21594 20395 -21560
rect 20429 -21594 20463 -21560
rect 20497 -21594 20531 -21560
rect 20565 -21594 20599 -21560
rect 20633 -21594 20667 -21560
rect 21175 -21594 21209 -21560
rect 21243 -21594 21277 -21560
rect 21311 -21594 21345 -21560
rect 21379 -21594 21413 -21560
rect 21447 -21594 21481 -21560
rect 21515 -21594 21549 -21560
rect 21583 -21594 21617 -21560
rect 21651 -21594 21685 -21560
rect 22193 -21594 22227 -21560
rect 22261 -21594 22295 -21560
rect 22329 -21594 22363 -21560
rect 22397 -21594 22431 -21560
rect 22465 -21594 22499 -21560
rect 22533 -21594 22567 -21560
rect 22601 -21594 22635 -21560
rect 22669 -21594 22703 -21560
rect 2851 -22304 2885 -22270
rect 2919 -22304 2953 -22270
rect 2987 -22304 3021 -22270
rect 3055 -22304 3089 -22270
rect 3123 -22304 3157 -22270
rect 3191 -22304 3225 -22270
rect 3259 -22304 3293 -22270
rect 3327 -22304 3361 -22270
rect 3869 -22304 3903 -22270
rect 3937 -22304 3971 -22270
rect 4005 -22304 4039 -22270
rect 4073 -22304 4107 -22270
rect 4141 -22304 4175 -22270
rect 4209 -22304 4243 -22270
rect 4277 -22304 4311 -22270
rect 4345 -22304 4379 -22270
rect 4887 -22304 4921 -22270
rect 4955 -22304 4989 -22270
rect 5023 -22304 5057 -22270
rect 5091 -22304 5125 -22270
rect 5159 -22304 5193 -22270
rect 5227 -22304 5261 -22270
rect 5295 -22304 5329 -22270
rect 5363 -22304 5397 -22270
rect 5905 -22304 5939 -22270
rect 5973 -22304 6007 -22270
rect 6041 -22304 6075 -22270
rect 6109 -22304 6143 -22270
rect 6177 -22304 6211 -22270
rect 6245 -22304 6279 -22270
rect 6313 -22304 6347 -22270
rect 6381 -22304 6415 -22270
rect 6923 -22304 6957 -22270
rect 6991 -22304 7025 -22270
rect 7059 -22304 7093 -22270
rect 7127 -22304 7161 -22270
rect 7195 -22304 7229 -22270
rect 7263 -22304 7297 -22270
rect 7331 -22304 7365 -22270
rect 7399 -22304 7433 -22270
rect 7941 -22304 7975 -22270
rect 8009 -22304 8043 -22270
rect 8077 -22304 8111 -22270
rect 8145 -22304 8179 -22270
rect 8213 -22304 8247 -22270
rect 8281 -22304 8315 -22270
rect 8349 -22304 8383 -22270
rect 8417 -22304 8451 -22270
rect 8959 -22304 8993 -22270
rect 9027 -22304 9061 -22270
rect 9095 -22304 9129 -22270
rect 9163 -22304 9197 -22270
rect 9231 -22304 9265 -22270
rect 9299 -22304 9333 -22270
rect 9367 -22304 9401 -22270
rect 9435 -22304 9469 -22270
rect 9977 -22304 10011 -22270
rect 10045 -22304 10079 -22270
rect 10113 -22304 10147 -22270
rect 10181 -22304 10215 -22270
rect 10249 -22304 10283 -22270
rect 10317 -22304 10351 -22270
rect 10385 -22304 10419 -22270
rect 10453 -22304 10487 -22270
rect 10995 -22304 11029 -22270
rect 11063 -22304 11097 -22270
rect 11131 -22304 11165 -22270
rect 11199 -22304 11233 -22270
rect 11267 -22304 11301 -22270
rect 11335 -22304 11369 -22270
rect 11403 -22304 11437 -22270
rect 11471 -22304 11505 -22270
rect 12013 -22304 12047 -22270
rect 12081 -22304 12115 -22270
rect 12149 -22304 12183 -22270
rect 12217 -22304 12251 -22270
rect 12285 -22304 12319 -22270
rect 12353 -22304 12387 -22270
rect 12421 -22304 12455 -22270
rect 12489 -22304 12523 -22270
rect 13031 -22304 13065 -22270
rect 13099 -22304 13133 -22270
rect 13167 -22304 13201 -22270
rect 13235 -22304 13269 -22270
rect 13303 -22304 13337 -22270
rect 13371 -22304 13405 -22270
rect 13439 -22304 13473 -22270
rect 13507 -22304 13541 -22270
rect 14049 -22304 14083 -22270
rect 14117 -22304 14151 -22270
rect 14185 -22304 14219 -22270
rect 14253 -22304 14287 -22270
rect 14321 -22304 14355 -22270
rect 14389 -22304 14423 -22270
rect 14457 -22304 14491 -22270
rect 14525 -22304 14559 -22270
rect 15067 -22304 15101 -22270
rect 15135 -22304 15169 -22270
rect 15203 -22304 15237 -22270
rect 15271 -22304 15305 -22270
rect 15339 -22304 15373 -22270
rect 15407 -22304 15441 -22270
rect 15475 -22304 15509 -22270
rect 15543 -22304 15577 -22270
rect 16085 -22304 16119 -22270
rect 16153 -22304 16187 -22270
rect 16221 -22304 16255 -22270
rect 16289 -22304 16323 -22270
rect 16357 -22304 16391 -22270
rect 16425 -22304 16459 -22270
rect 16493 -22304 16527 -22270
rect 16561 -22304 16595 -22270
rect 17103 -22304 17137 -22270
rect 17171 -22304 17205 -22270
rect 17239 -22304 17273 -22270
rect 17307 -22304 17341 -22270
rect 17375 -22304 17409 -22270
rect 17443 -22304 17477 -22270
rect 17511 -22304 17545 -22270
rect 17579 -22304 17613 -22270
rect 18121 -22304 18155 -22270
rect 18189 -22304 18223 -22270
rect 18257 -22304 18291 -22270
rect 18325 -22304 18359 -22270
rect 18393 -22304 18427 -22270
rect 18461 -22304 18495 -22270
rect 18529 -22304 18563 -22270
rect 18597 -22304 18631 -22270
rect 19139 -22304 19173 -22270
rect 19207 -22304 19241 -22270
rect 19275 -22304 19309 -22270
rect 19343 -22304 19377 -22270
rect 19411 -22304 19445 -22270
rect 19479 -22304 19513 -22270
rect 19547 -22304 19581 -22270
rect 19615 -22304 19649 -22270
rect 20157 -22304 20191 -22270
rect 20225 -22304 20259 -22270
rect 20293 -22304 20327 -22270
rect 20361 -22304 20395 -22270
rect 20429 -22304 20463 -22270
rect 20497 -22304 20531 -22270
rect 20565 -22304 20599 -22270
rect 20633 -22304 20667 -22270
rect 21175 -22304 21209 -22270
rect 21243 -22304 21277 -22270
rect 21311 -22304 21345 -22270
rect 21379 -22304 21413 -22270
rect 21447 -22304 21481 -22270
rect 21515 -22304 21549 -22270
rect 21583 -22304 21617 -22270
rect 21651 -22304 21685 -22270
rect 22193 -22304 22227 -22270
rect 22261 -22304 22295 -22270
rect 22329 -22304 22363 -22270
rect 22397 -22304 22431 -22270
rect 22465 -22304 22499 -22270
rect 22533 -22304 22567 -22270
rect 22601 -22304 22635 -22270
rect 22669 -22304 22703 -22270
rect 2851 -22826 2885 -22792
rect 2919 -22826 2953 -22792
rect 2987 -22826 3021 -22792
rect 3055 -22826 3089 -22792
rect 3123 -22826 3157 -22792
rect 3191 -22826 3225 -22792
rect 3259 -22826 3293 -22792
rect 3327 -22826 3361 -22792
rect 3869 -22826 3903 -22792
rect 3937 -22826 3971 -22792
rect 4005 -22826 4039 -22792
rect 4073 -22826 4107 -22792
rect 4141 -22826 4175 -22792
rect 4209 -22826 4243 -22792
rect 4277 -22826 4311 -22792
rect 4345 -22826 4379 -22792
rect 4887 -22826 4921 -22792
rect 4955 -22826 4989 -22792
rect 5023 -22826 5057 -22792
rect 5091 -22826 5125 -22792
rect 5159 -22826 5193 -22792
rect 5227 -22826 5261 -22792
rect 5295 -22826 5329 -22792
rect 5363 -22826 5397 -22792
rect 5905 -22826 5939 -22792
rect 5973 -22826 6007 -22792
rect 6041 -22826 6075 -22792
rect 6109 -22826 6143 -22792
rect 6177 -22826 6211 -22792
rect 6245 -22826 6279 -22792
rect 6313 -22826 6347 -22792
rect 6381 -22826 6415 -22792
rect 6923 -22826 6957 -22792
rect 6991 -22826 7025 -22792
rect 7059 -22826 7093 -22792
rect 7127 -22826 7161 -22792
rect 7195 -22826 7229 -22792
rect 7263 -22826 7297 -22792
rect 7331 -22826 7365 -22792
rect 7399 -22826 7433 -22792
rect 7941 -22826 7975 -22792
rect 8009 -22826 8043 -22792
rect 8077 -22826 8111 -22792
rect 8145 -22826 8179 -22792
rect 8213 -22826 8247 -22792
rect 8281 -22826 8315 -22792
rect 8349 -22826 8383 -22792
rect 8417 -22826 8451 -22792
rect 8959 -22826 8993 -22792
rect 9027 -22826 9061 -22792
rect 9095 -22826 9129 -22792
rect 9163 -22826 9197 -22792
rect 9231 -22826 9265 -22792
rect 9299 -22826 9333 -22792
rect 9367 -22826 9401 -22792
rect 9435 -22826 9469 -22792
rect 9977 -22826 10011 -22792
rect 10045 -22826 10079 -22792
rect 10113 -22826 10147 -22792
rect 10181 -22826 10215 -22792
rect 10249 -22826 10283 -22792
rect 10317 -22826 10351 -22792
rect 10385 -22826 10419 -22792
rect 10453 -22826 10487 -22792
rect 10995 -22826 11029 -22792
rect 11063 -22826 11097 -22792
rect 11131 -22826 11165 -22792
rect 11199 -22826 11233 -22792
rect 11267 -22826 11301 -22792
rect 11335 -22826 11369 -22792
rect 11403 -22826 11437 -22792
rect 11471 -22826 11505 -22792
rect 12013 -22826 12047 -22792
rect 12081 -22826 12115 -22792
rect 12149 -22826 12183 -22792
rect 12217 -22826 12251 -22792
rect 12285 -22826 12319 -22792
rect 12353 -22826 12387 -22792
rect 12421 -22826 12455 -22792
rect 12489 -22826 12523 -22792
rect 13031 -22826 13065 -22792
rect 13099 -22826 13133 -22792
rect 13167 -22826 13201 -22792
rect 13235 -22826 13269 -22792
rect 13303 -22826 13337 -22792
rect 13371 -22826 13405 -22792
rect 13439 -22826 13473 -22792
rect 13507 -22826 13541 -22792
rect 14049 -22826 14083 -22792
rect 14117 -22826 14151 -22792
rect 14185 -22826 14219 -22792
rect 14253 -22826 14287 -22792
rect 14321 -22826 14355 -22792
rect 14389 -22826 14423 -22792
rect 14457 -22826 14491 -22792
rect 14525 -22826 14559 -22792
rect 15067 -22826 15101 -22792
rect 15135 -22826 15169 -22792
rect 15203 -22826 15237 -22792
rect 15271 -22826 15305 -22792
rect 15339 -22826 15373 -22792
rect 15407 -22826 15441 -22792
rect 15475 -22826 15509 -22792
rect 15543 -22826 15577 -22792
rect 16085 -22826 16119 -22792
rect 16153 -22826 16187 -22792
rect 16221 -22826 16255 -22792
rect 16289 -22826 16323 -22792
rect 16357 -22826 16391 -22792
rect 16425 -22826 16459 -22792
rect 16493 -22826 16527 -22792
rect 16561 -22826 16595 -22792
rect 17103 -22826 17137 -22792
rect 17171 -22826 17205 -22792
rect 17239 -22826 17273 -22792
rect 17307 -22826 17341 -22792
rect 17375 -22826 17409 -22792
rect 17443 -22826 17477 -22792
rect 17511 -22826 17545 -22792
rect 17579 -22826 17613 -22792
rect 18121 -22826 18155 -22792
rect 18189 -22826 18223 -22792
rect 18257 -22826 18291 -22792
rect 18325 -22826 18359 -22792
rect 18393 -22826 18427 -22792
rect 18461 -22826 18495 -22792
rect 18529 -22826 18563 -22792
rect 18597 -22826 18631 -22792
rect 19139 -22826 19173 -22792
rect 19207 -22826 19241 -22792
rect 19275 -22826 19309 -22792
rect 19343 -22826 19377 -22792
rect 19411 -22826 19445 -22792
rect 19479 -22826 19513 -22792
rect 19547 -22826 19581 -22792
rect 19615 -22826 19649 -22792
rect 20157 -22826 20191 -22792
rect 20225 -22826 20259 -22792
rect 20293 -22826 20327 -22792
rect 20361 -22826 20395 -22792
rect 20429 -22826 20463 -22792
rect 20497 -22826 20531 -22792
rect 20565 -22826 20599 -22792
rect 20633 -22826 20667 -22792
rect 21175 -22826 21209 -22792
rect 21243 -22826 21277 -22792
rect 21311 -22826 21345 -22792
rect 21379 -22826 21413 -22792
rect 21447 -22826 21481 -22792
rect 21515 -22826 21549 -22792
rect 21583 -22826 21617 -22792
rect 21651 -22826 21685 -22792
rect 22193 -22826 22227 -22792
rect 22261 -22826 22295 -22792
rect 22329 -22826 22363 -22792
rect 22397 -22826 22431 -22792
rect 22465 -22826 22499 -22792
rect 22533 -22826 22567 -22792
rect 22601 -22826 22635 -22792
rect 22669 -22826 22703 -22792
rect 2851 -23536 2885 -23502
rect 2919 -23536 2953 -23502
rect 2987 -23536 3021 -23502
rect 3055 -23536 3089 -23502
rect 3123 -23536 3157 -23502
rect 3191 -23536 3225 -23502
rect 3259 -23536 3293 -23502
rect 3327 -23536 3361 -23502
rect 3869 -23536 3903 -23502
rect 3937 -23536 3971 -23502
rect 4005 -23536 4039 -23502
rect 4073 -23536 4107 -23502
rect 4141 -23536 4175 -23502
rect 4209 -23536 4243 -23502
rect 4277 -23536 4311 -23502
rect 4345 -23536 4379 -23502
rect 4887 -23536 4921 -23502
rect 4955 -23536 4989 -23502
rect 5023 -23536 5057 -23502
rect 5091 -23536 5125 -23502
rect 5159 -23536 5193 -23502
rect 5227 -23536 5261 -23502
rect 5295 -23536 5329 -23502
rect 5363 -23536 5397 -23502
rect 5905 -23536 5939 -23502
rect 5973 -23536 6007 -23502
rect 6041 -23536 6075 -23502
rect 6109 -23536 6143 -23502
rect 6177 -23536 6211 -23502
rect 6245 -23536 6279 -23502
rect 6313 -23536 6347 -23502
rect 6381 -23536 6415 -23502
rect 6923 -23536 6957 -23502
rect 6991 -23536 7025 -23502
rect 7059 -23536 7093 -23502
rect 7127 -23536 7161 -23502
rect 7195 -23536 7229 -23502
rect 7263 -23536 7297 -23502
rect 7331 -23536 7365 -23502
rect 7399 -23536 7433 -23502
rect 7941 -23536 7975 -23502
rect 8009 -23536 8043 -23502
rect 8077 -23536 8111 -23502
rect 8145 -23536 8179 -23502
rect 8213 -23536 8247 -23502
rect 8281 -23536 8315 -23502
rect 8349 -23536 8383 -23502
rect 8417 -23536 8451 -23502
rect 8959 -23536 8993 -23502
rect 9027 -23536 9061 -23502
rect 9095 -23536 9129 -23502
rect 9163 -23536 9197 -23502
rect 9231 -23536 9265 -23502
rect 9299 -23536 9333 -23502
rect 9367 -23536 9401 -23502
rect 9435 -23536 9469 -23502
rect 9977 -23536 10011 -23502
rect 10045 -23536 10079 -23502
rect 10113 -23536 10147 -23502
rect 10181 -23536 10215 -23502
rect 10249 -23536 10283 -23502
rect 10317 -23536 10351 -23502
rect 10385 -23536 10419 -23502
rect 10453 -23536 10487 -23502
rect 10995 -23536 11029 -23502
rect 11063 -23536 11097 -23502
rect 11131 -23536 11165 -23502
rect 11199 -23536 11233 -23502
rect 11267 -23536 11301 -23502
rect 11335 -23536 11369 -23502
rect 11403 -23536 11437 -23502
rect 11471 -23536 11505 -23502
rect 12013 -23536 12047 -23502
rect 12081 -23536 12115 -23502
rect 12149 -23536 12183 -23502
rect 12217 -23536 12251 -23502
rect 12285 -23536 12319 -23502
rect 12353 -23536 12387 -23502
rect 12421 -23536 12455 -23502
rect 12489 -23536 12523 -23502
rect 13031 -23536 13065 -23502
rect 13099 -23536 13133 -23502
rect 13167 -23536 13201 -23502
rect 13235 -23536 13269 -23502
rect 13303 -23536 13337 -23502
rect 13371 -23536 13405 -23502
rect 13439 -23536 13473 -23502
rect 13507 -23536 13541 -23502
rect 14049 -23536 14083 -23502
rect 14117 -23536 14151 -23502
rect 14185 -23536 14219 -23502
rect 14253 -23536 14287 -23502
rect 14321 -23536 14355 -23502
rect 14389 -23536 14423 -23502
rect 14457 -23536 14491 -23502
rect 14525 -23536 14559 -23502
rect 15067 -23536 15101 -23502
rect 15135 -23536 15169 -23502
rect 15203 -23536 15237 -23502
rect 15271 -23536 15305 -23502
rect 15339 -23536 15373 -23502
rect 15407 -23536 15441 -23502
rect 15475 -23536 15509 -23502
rect 15543 -23536 15577 -23502
rect 16085 -23536 16119 -23502
rect 16153 -23536 16187 -23502
rect 16221 -23536 16255 -23502
rect 16289 -23536 16323 -23502
rect 16357 -23536 16391 -23502
rect 16425 -23536 16459 -23502
rect 16493 -23536 16527 -23502
rect 16561 -23536 16595 -23502
rect 17103 -23536 17137 -23502
rect 17171 -23536 17205 -23502
rect 17239 -23536 17273 -23502
rect 17307 -23536 17341 -23502
rect 17375 -23536 17409 -23502
rect 17443 -23536 17477 -23502
rect 17511 -23536 17545 -23502
rect 17579 -23536 17613 -23502
rect 18121 -23536 18155 -23502
rect 18189 -23536 18223 -23502
rect 18257 -23536 18291 -23502
rect 18325 -23536 18359 -23502
rect 18393 -23536 18427 -23502
rect 18461 -23536 18495 -23502
rect 18529 -23536 18563 -23502
rect 18597 -23536 18631 -23502
rect 19139 -23536 19173 -23502
rect 19207 -23536 19241 -23502
rect 19275 -23536 19309 -23502
rect 19343 -23536 19377 -23502
rect 19411 -23536 19445 -23502
rect 19479 -23536 19513 -23502
rect 19547 -23536 19581 -23502
rect 19615 -23536 19649 -23502
rect 20157 -23536 20191 -23502
rect 20225 -23536 20259 -23502
rect 20293 -23536 20327 -23502
rect 20361 -23536 20395 -23502
rect 20429 -23536 20463 -23502
rect 20497 -23536 20531 -23502
rect 20565 -23536 20599 -23502
rect 20633 -23536 20667 -23502
rect 21175 -23536 21209 -23502
rect 21243 -23536 21277 -23502
rect 21311 -23536 21345 -23502
rect 21379 -23536 21413 -23502
rect 21447 -23536 21481 -23502
rect 21515 -23536 21549 -23502
rect 21583 -23536 21617 -23502
rect 21651 -23536 21685 -23502
rect 22193 -23536 22227 -23502
rect 22261 -23536 22295 -23502
rect 22329 -23536 22363 -23502
rect 22397 -23536 22431 -23502
rect 22465 -23536 22499 -23502
rect 22533 -23536 22567 -23502
rect 22601 -23536 22635 -23502
rect 22669 -23536 22703 -23502
rect 2851 -24060 2885 -24026
rect 2919 -24060 2953 -24026
rect 2987 -24060 3021 -24026
rect 3055 -24060 3089 -24026
rect 3123 -24060 3157 -24026
rect 3191 -24060 3225 -24026
rect 3259 -24060 3293 -24026
rect 3327 -24060 3361 -24026
rect 3869 -24060 3903 -24026
rect 3937 -24060 3971 -24026
rect 4005 -24060 4039 -24026
rect 4073 -24060 4107 -24026
rect 4141 -24060 4175 -24026
rect 4209 -24060 4243 -24026
rect 4277 -24060 4311 -24026
rect 4345 -24060 4379 -24026
rect 4887 -24060 4921 -24026
rect 4955 -24060 4989 -24026
rect 5023 -24060 5057 -24026
rect 5091 -24060 5125 -24026
rect 5159 -24060 5193 -24026
rect 5227 -24060 5261 -24026
rect 5295 -24060 5329 -24026
rect 5363 -24060 5397 -24026
rect 5905 -24060 5939 -24026
rect 5973 -24060 6007 -24026
rect 6041 -24060 6075 -24026
rect 6109 -24060 6143 -24026
rect 6177 -24060 6211 -24026
rect 6245 -24060 6279 -24026
rect 6313 -24060 6347 -24026
rect 6381 -24060 6415 -24026
rect 6923 -24060 6957 -24026
rect 6991 -24060 7025 -24026
rect 7059 -24060 7093 -24026
rect 7127 -24060 7161 -24026
rect 7195 -24060 7229 -24026
rect 7263 -24060 7297 -24026
rect 7331 -24060 7365 -24026
rect 7399 -24060 7433 -24026
rect 7941 -24060 7975 -24026
rect 8009 -24060 8043 -24026
rect 8077 -24060 8111 -24026
rect 8145 -24060 8179 -24026
rect 8213 -24060 8247 -24026
rect 8281 -24060 8315 -24026
rect 8349 -24060 8383 -24026
rect 8417 -24060 8451 -24026
rect 8959 -24060 8993 -24026
rect 9027 -24060 9061 -24026
rect 9095 -24060 9129 -24026
rect 9163 -24060 9197 -24026
rect 9231 -24060 9265 -24026
rect 9299 -24060 9333 -24026
rect 9367 -24060 9401 -24026
rect 9435 -24060 9469 -24026
rect 9977 -24060 10011 -24026
rect 10045 -24060 10079 -24026
rect 10113 -24060 10147 -24026
rect 10181 -24060 10215 -24026
rect 10249 -24060 10283 -24026
rect 10317 -24060 10351 -24026
rect 10385 -24060 10419 -24026
rect 10453 -24060 10487 -24026
rect 10995 -24060 11029 -24026
rect 11063 -24060 11097 -24026
rect 11131 -24060 11165 -24026
rect 11199 -24060 11233 -24026
rect 11267 -24060 11301 -24026
rect 11335 -24060 11369 -24026
rect 11403 -24060 11437 -24026
rect 11471 -24060 11505 -24026
rect 12013 -24060 12047 -24026
rect 12081 -24060 12115 -24026
rect 12149 -24060 12183 -24026
rect 12217 -24060 12251 -24026
rect 12285 -24060 12319 -24026
rect 12353 -24060 12387 -24026
rect 12421 -24060 12455 -24026
rect 12489 -24060 12523 -24026
rect 13031 -24060 13065 -24026
rect 13099 -24060 13133 -24026
rect 13167 -24060 13201 -24026
rect 13235 -24060 13269 -24026
rect 13303 -24060 13337 -24026
rect 13371 -24060 13405 -24026
rect 13439 -24060 13473 -24026
rect 13507 -24060 13541 -24026
rect 14049 -24060 14083 -24026
rect 14117 -24060 14151 -24026
rect 14185 -24060 14219 -24026
rect 14253 -24060 14287 -24026
rect 14321 -24060 14355 -24026
rect 14389 -24060 14423 -24026
rect 14457 -24060 14491 -24026
rect 14525 -24060 14559 -24026
rect 15067 -24060 15101 -24026
rect 15135 -24060 15169 -24026
rect 15203 -24060 15237 -24026
rect 15271 -24060 15305 -24026
rect 15339 -24060 15373 -24026
rect 15407 -24060 15441 -24026
rect 15475 -24060 15509 -24026
rect 15543 -24060 15577 -24026
rect 16085 -24060 16119 -24026
rect 16153 -24060 16187 -24026
rect 16221 -24060 16255 -24026
rect 16289 -24060 16323 -24026
rect 16357 -24060 16391 -24026
rect 16425 -24060 16459 -24026
rect 16493 -24060 16527 -24026
rect 16561 -24060 16595 -24026
rect 17103 -24060 17137 -24026
rect 17171 -24060 17205 -24026
rect 17239 -24060 17273 -24026
rect 17307 -24060 17341 -24026
rect 17375 -24060 17409 -24026
rect 17443 -24060 17477 -24026
rect 17511 -24060 17545 -24026
rect 17579 -24060 17613 -24026
rect 18121 -24060 18155 -24026
rect 18189 -24060 18223 -24026
rect 18257 -24060 18291 -24026
rect 18325 -24060 18359 -24026
rect 18393 -24060 18427 -24026
rect 18461 -24060 18495 -24026
rect 18529 -24060 18563 -24026
rect 18597 -24060 18631 -24026
rect 19139 -24060 19173 -24026
rect 19207 -24060 19241 -24026
rect 19275 -24060 19309 -24026
rect 19343 -24060 19377 -24026
rect 19411 -24060 19445 -24026
rect 19479 -24060 19513 -24026
rect 19547 -24060 19581 -24026
rect 19615 -24060 19649 -24026
rect 20157 -24060 20191 -24026
rect 20225 -24060 20259 -24026
rect 20293 -24060 20327 -24026
rect 20361 -24060 20395 -24026
rect 20429 -24060 20463 -24026
rect 20497 -24060 20531 -24026
rect 20565 -24060 20599 -24026
rect 20633 -24060 20667 -24026
rect 21175 -24060 21209 -24026
rect 21243 -24060 21277 -24026
rect 21311 -24060 21345 -24026
rect 21379 -24060 21413 -24026
rect 21447 -24060 21481 -24026
rect 21515 -24060 21549 -24026
rect 21583 -24060 21617 -24026
rect 21651 -24060 21685 -24026
rect 22193 -24060 22227 -24026
rect 22261 -24060 22295 -24026
rect 22329 -24060 22363 -24026
rect 22397 -24060 22431 -24026
rect 22465 -24060 22499 -24026
rect 22533 -24060 22567 -24026
rect 22601 -24060 22635 -24026
rect 22669 -24060 22703 -24026
rect 2851 -24770 2885 -24736
rect 2919 -24770 2953 -24736
rect 2987 -24770 3021 -24736
rect 3055 -24770 3089 -24736
rect 3123 -24770 3157 -24736
rect 3191 -24770 3225 -24736
rect 3259 -24770 3293 -24736
rect 3327 -24770 3361 -24736
rect 3869 -24770 3903 -24736
rect 3937 -24770 3971 -24736
rect 4005 -24770 4039 -24736
rect 4073 -24770 4107 -24736
rect 4141 -24770 4175 -24736
rect 4209 -24770 4243 -24736
rect 4277 -24770 4311 -24736
rect 4345 -24770 4379 -24736
rect 4887 -24770 4921 -24736
rect 4955 -24770 4989 -24736
rect 5023 -24770 5057 -24736
rect 5091 -24770 5125 -24736
rect 5159 -24770 5193 -24736
rect 5227 -24770 5261 -24736
rect 5295 -24770 5329 -24736
rect 5363 -24770 5397 -24736
rect 5905 -24770 5939 -24736
rect 5973 -24770 6007 -24736
rect 6041 -24770 6075 -24736
rect 6109 -24770 6143 -24736
rect 6177 -24770 6211 -24736
rect 6245 -24770 6279 -24736
rect 6313 -24770 6347 -24736
rect 6381 -24770 6415 -24736
rect 6923 -24770 6957 -24736
rect 6991 -24770 7025 -24736
rect 7059 -24770 7093 -24736
rect 7127 -24770 7161 -24736
rect 7195 -24770 7229 -24736
rect 7263 -24770 7297 -24736
rect 7331 -24770 7365 -24736
rect 7399 -24770 7433 -24736
rect 7941 -24770 7975 -24736
rect 8009 -24770 8043 -24736
rect 8077 -24770 8111 -24736
rect 8145 -24770 8179 -24736
rect 8213 -24770 8247 -24736
rect 8281 -24770 8315 -24736
rect 8349 -24770 8383 -24736
rect 8417 -24770 8451 -24736
rect 8959 -24770 8993 -24736
rect 9027 -24770 9061 -24736
rect 9095 -24770 9129 -24736
rect 9163 -24770 9197 -24736
rect 9231 -24770 9265 -24736
rect 9299 -24770 9333 -24736
rect 9367 -24770 9401 -24736
rect 9435 -24770 9469 -24736
rect 9977 -24770 10011 -24736
rect 10045 -24770 10079 -24736
rect 10113 -24770 10147 -24736
rect 10181 -24770 10215 -24736
rect 10249 -24770 10283 -24736
rect 10317 -24770 10351 -24736
rect 10385 -24770 10419 -24736
rect 10453 -24770 10487 -24736
rect 10995 -24770 11029 -24736
rect 11063 -24770 11097 -24736
rect 11131 -24770 11165 -24736
rect 11199 -24770 11233 -24736
rect 11267 -24770 11301 -24736
rect 11335 -24770 11369 -24736
rect 11403 -24770 11437 -24736
rect 11471 -24770 11505 -24736
rect 12013 -24770 12047 -24736
rect 12081 -24770 12115 -24736
rect 12149 -24770 12183 -24736
rect 12217 -24770 12251 -24736
rect 12285 -24770 12319 -24736
rect 12353 -24770 12387 -24736
rect 12421 -24770 12455 -24736
rect 12489 -24770 12523 -24736
rect 13031 -24770 13065 -24736
rect 13099 -24770 13133 -24736
rect 13167 -24770 13201 -24736
rect 13235 -24770 13269 -24736
rect 13303 -24770 13337 -24736
rect 13371 -24770 13405 -24736
rect 13439 -24770 13473 -24736
rect 13507 -24770 13541 -24736
rect 14049 -24770 14083 -24736
rect 14117 -24770 14151 -24736
rect 14185 -24770 14219 -24736
rect 14253 -24770 14287 -24736
rect 14321 -24770 14355 -24736
rect 14389 -24770 14423 -24736
rect 14457 -24770 14491 -24736
rect 14525 -24770 14559 -24736
rect 15067 -24770 15101 -24736
rect 15135 -24770 15169 -24736
rect 15203 -24770 15237 -24736
rect 15271 -24770 15305 -24736
rect 15339 -24770 15373 -24736
rect 15407 -24770 15441 -24736
rect 15475 -24770 15509 -24736
rect 15543 -24770 15577 -24736
rect 16085 -24770 16119 -24736
rect 16153 -24770 16187 -24736
rect 16221 -24770 16255 -24736
rect 16289 -24770 16323 -24736
rect 16357 -24770 16391 -24736
rect 16425 -24770 16459 -24736
rect 16493 -24770 16527 -24736
rect 16561 -24770 16595 -24736
rect 17103 -24770 17137 -24736
rect 17171 -24770 17205 -24736
rect 17239 -24770 17273 -24736
rect 17307 -24770 17341 -24736
rect 17375 -24770 17409 -24736
rect 17443 -24770 17477 -24736
rect 17511 -24770 17545 -24736
rect 17579 -24770 17613 -24736
rect 18121 -24770 18155 -24736
rect 18189 -24770 18223 -24736
rect 18257 -24770 18291 -24736
rect 18325 -24770 18359 -24736
rect 18393 -24770 18427 -24736
rect 18461 -24770 18495 -24736
rect 18529 -24770 18563 -24736
rect 18597 -24770 18631 -24736
rect 19139 -24770 19173 -24736
rect 19207 -24770 19241 -24736
rect 19275 -24770 19309 -24736
rect 19343 -24770 19377 -24736
rect 19411 -24770 19445 -24736
rect 19479 -24770 19513 -24736
rect 19547 -24770 19581 -24736
rect 19615 -24770 19649 -24736
rect 20157 -24770 20191 -24736
rect 20225 -24770 20259 -24736
rect 20293 -24770 20327 -24736
rect 20361 -24770 20395 -24736
rect 20429 -24770 20463 -24736
rect 20497 -24770 20531 -24736
rect 20565 -24770 20599 -24736
rect 20633 -24770 20667 -24736
rect 21175 -24770 21209 -24736
rect 21243 -24770 21277 -24736
rect 21311 -24770 21345 -24736
rect 21379 -24770 21413 -24736
rect 21447 -24770 21481 -24736
rect 21515 -24770 21549 -24736
rect 21583 -24770 21617 -24736
rect 21651 -24770 21685 -24736
rect 22193 -24770 22227 -24736
rect 22261 -24770 22295 -24736
rect 22329 -24770 22363 -24736
rect 22397 -24770 22431 -24736
rect 22465 -24770 22499 -24736
rect 22533 -24770 22567 -24736
rect 22601 -24770 22635 -24736
rect 22669 -24770 22703 -24736
<< locali >>
rect 378 4289 24822 4322
rect 378 4255 487 4289
rect 521 4255 547 4289
rect 593 4255 615 4289
rect 665 4255 683 4289
rect 737 4255 751 4289
rect 809 4255 819 4289
rect 881 4255 887 4289
rect 953 4255 955 4289
rect 989 4255 991 4289
rect 1057 4255 1063 4289
rect 1125 4255 1135 4289
rect 1193 4255 1207 4289
rect 1261 4255 1279 4289
rect 1329 4255 1351 4289
rect 1397 4255 1423 4289
rect 1465 4255 1495 4289
rect 1533 4255 1567 4289
rect 1601 4255 1635 4289
rect 1673 4255 1703 4289
rect 1745 4255 1771 4289
rect 1817 4255 1839 4289
rect 1889 4255 1907 4289
rect 1961 4255 1975 4289
rect 2033 4255 2043 4289
rect 2105 4255 2111 4289
rect 2177 4255 2179 4289
rect 2213 4255 2215 4289
rect 2281 4255 2287 4289
rect 2349 4255 2359 4289
rect 2417 4255 2431 4289
rect 2485 4255 2503 4289
rect 2553 4255 2575 4289
rect 2621 4255 2647 4289
rect 2689 4255 2719 4289
rect 2757 4255 2791 4289
rect 2825 4255 2859 4289
rect 2897 4255 2927 4289
rect 2969 4255 2995 4289
rect 3041 4255 3063 4289
rect 3113 4255 3131 4289
rect 3185 4255 3199 4289
rect 3257 4255 3267 4289
rect 3329 4255 3335 4289
rect 3401 4255 3403 4289
rect 3437 4255 3439 4289
rect 3505 4255 3511 4289
rect 3573 4255 3583 4289
rect 3641 4255 3655 4289
rect 3709 4255 3727 4289
rect 3777 4255 3799 4289
rect 3845 4255 3871 4289
rect 3913 4255 3943 4289
rect 3981 4255 4015 4289
rect 4049 4255 4083 4289
rect 4121 4255 4151 4289
rect 4193 4255 4219 4289
rect 4265 4255 4287 4289
rect 4337 4255 4355 4289
rect 4409 4255 4423 4289
rect 4481 4255 4491 4289
rect 4553 4255 4559 4289
rect 4625 4255 4627 4289
rect 4661 4255 4663 4289
rect 4729 4255 4735 4289
rect 4797 4255 4807 4289
rect 4865 4255 4879 4289
rect 4933 4255 4951 4289
rect 5001 4255 5023 4289
rect 5069 4255 5095 4289
rect 5137 4255 5167 4289
rect 5205 4255 5239 4289
rect 5273 4255 5307 4289
rect 5345 4255 5375 4289
rect 5417 4255 5443 4289
rect 5489 4255 5511 4289
rect 5561 4255 5579 4289
rect 5633 4255 5647 4289
rect 5705 4255 5715 4289
rect 5777 4255 5783 4289
rect 5849 4255 5851 4289
rect 5885 4255 5887 4289
rect 5953 4255 5959 4289
rect 6021 4255 6031 4289
rect 6089 4255 6103 4289
rect 6157 4255 6175 4289
rect 6225 4255 6247 4289
rect 6293 4255 6319 4289
rect 6361 4255 6391 4289
rect 6429 4255 6463 4289
rect 6497 4255 6531 4289
rect 6569 4255 6599 4289
rect 6641 4255 6667 4289
rect 6713 4255 6735 4289
rect 6785 4255 6803 4289
rect 6857 4255 6871 4289
rect 6929 4255 6939 4289
rect 7001 4255 7007 4289
rect 7073 4255 7075 4289
rect 7109 4255 7111 4289
rect 7177 4255 7183 4289
rect 7245 4255 7255 4289
rect 7313 4255 7327 4289
rect 7381 4255 7399 4289
rect 7449 4255 7471 4289
rect 7517 4255 7543 4289
rect 7585 4255 7615 4289
rect 7653 4255 7687 4289
rect 7721 4255 7755 4289
rect 7793 4255 7823 4289
rect 7865 4255 7891 4289
rect 7937 4255 7959 4289
rect 8009 4255 8027 4289
rect 8081 4255 8095 4289
rect 8153 4255 8163 4289
rect 8225 4255 8231 4289
rect 8297 4255 8299 4289
rect 8333 4255 8335 4289
rect 8401 4255 8407 4289
rect 8469 4255 8479 4289
rect 8537 4255 8551 4289
rect 8605 4255 8623 4289
rect 8673 4255 8695 4289
rect 8741 4255 8767 4289
rect 8809 4255 8839 4289
rect 8877 4255 8911 4289
rect 8945 4255 8979 4289
rect 9017 4255 9047 4289
rect 9089 4255 9115 4289
rect 9161 4255 9183 4289
rect 9233 4255 9251 4289
rect 9305 4255 9319 4289
rect 9377 4255 9387 4289
rect 9449 4255 9455 4289
rect 9521 4255 9523 4289
rect 9557 4255 9559 4289
rect 9625 4255 9631 4289
rect 9693 4255 9703 4289
rect 9761 4255 9775 4289
rect 9829 4255 9847 4289
rect 9897 4255 9919 4289
rect 9965 4255 9991 4289
rect 10033 4255 10063 4289
rect 10101 4255 10135 4289
rect 10169 4255 10203 4289
rect 10241 4255 10271 4289
rect 10313 4255 10339 4289
rect 10385 4255 10407 4289
rect 10457 4255 10475 4289
rect 10529 4255 10543 4289
rect 10601 4255 10611 4289
rect 10673 4255 10679 4289
rect 10745 4255 10747 4289
rect 10781 4255 10783 4289
rect 10849 4255 10855 4289
rect 10917 4255 10927 4289
rect 10985 4255 10999 4289
rect 11053 4255 11071 4289
rect 11121 4255 11143 4289
rect 11189 4255 11215 4289
rect 11257 4255 11287 4289
rect 11325 4255 11359 4289
rect 11393 4255 11427 4289
rect 11465 4255 11495 4289
rect 11537 4255 11563 4289
rect 11609 4255 11631 4289
rect 11681 4255 11699 4289
rect 11753 4255 11767 4289
rect 11825 4255 11835 4289
rect 11897 4255 11903 4289
rect 11969 4255 11971 4289
rect 12005 4255 12007 4289
rect 12073 4255 12079 4289
rect 12141 4255 12151 4289
rect 12209 4255 12223 4289
rect 12277 4255 12295 4289
rect 12345 4255 12367 4289
rect 12413 4255 12439 4289
rect 12481 4255 12511 4289
rect 12549 4255 12583 4289
rect 12617 4255 12651 4289
rect 12689 4255 12719 4289
rect 12761 4255 12787 4289
rect 12833 4255 12855 4289
rect 12905 4255 12923 4289
rect 12977 4255 12991 4289
rect 13049 4255 13059 4289
rect 13121 4255 13127 4289
rect 13193 4255 13195 4289
rect 13229 4255 13231 4289
rect 13297 4255 13303 4289
rect 13365 4255 13375 4289
rect 13433 4255 13447 4289
rect 13501 4255 13519 4289
rect 13569 4255 13591 4289
rect 13637 4255 13663 4289
rect 13705 4255 13735 4289
rect 13773 4255 13807 4289
rect 13841 4255 13875 4289
rect 13913 4255 13943 4289
rect 13985 4255 14011 4289
rect 14057 4255 14079 4289
rect 14129 4255 14147 4289
rect 14201 4255 14215 4289
rect 14273 4255 14283 4289
rect 14345 4255 14351 4289
rect 14417 4255 14419 4289
rect 14453 4255 14455 4289
rect 14521 4255 14527 4289
rect 14589 4255 14599 4289
rect 14657 4255 14671 4289
rect 14725 4255 14743 4289
rect 14793 4255 14815 4289
rect 14861 4255 14887 4289
rect 14929 4255 14959 4289
rect 14997 4255 15031 4289
rect 15065 4255 15099 4289
rect 15137 4255 15167 4289
rect 15209 4255 15235 4289
rect 15281 4255 15303 4289
rect 15353 4255 15371 4289
rect 15425 4255 15439 4289
rect 15497 4255 15507 4289
rect 15569 4255 15575 4289
rect 15641 4255 15643 4289
rect 15677 4255 15679 4289
rect 15745 4255 15751 4289
rect 15813 4255 15823 4289
rect 15881 4255 15895 4289
rect 15949 4255 15967 4289
rect 16017 4255 16039 4289
rect 16085 4255 16111 4289
rect 16153 4255 16183 4289
rect 16221 4255 16255 4289
rect 16289 4255 16323 4289
rect 16361 4255 16391 4289
rect 16433 4255 16459 4289
rect 16505 4255 16527 4289
rect 16577 4255 16595 4289
rect 16649 4255 16663 4289
rect 16721 4255 16731 4289
rect 16793 4255 16799 4289
rect 16865 4255 16867 4289
rect 16901 4255 16903 4289
rect 16969 4255 16975 4289
rect 17037 4255 17047 4289
rect 17105 4255 17119 4289
rect 17173 4255 17191 4289
rect 17241 4255 17263 4289
rect 17309 4255 17335 4289
rect 17377 4255 17407 4289
rect 17445 4255 17479 4289
rect 17513 4255 17547 4289
rect 17585 4255 17615 4289
rect 17657 4255 17683 4289
rect 17729 4255 17751 4289
rect 17801 4255 17819 4289
rect 17873 4255 17887 4289
rect 17945 4255 17955 4289
rect 18017 4255 18023 4289
rect 18089 4255 18091 4289
rect 18125 4255 18127 4289
rect 18193 4255 18199 4289
rect 18261 4255 18271 4289
rect 18329 4255 18343 4289
rect 18397 4255 18415 4289
rect 18465 4255 18487 4289
rect 18533 4255 18559 4289
rect 18601 4255 18631 4289
rect 18669 4255 18703 4289
rect 18737 4255 18771 4289
rect 18809 4255 18839 4289
rect 18881 4255 18907 4289
rect 18953 4255 18975 4289
rect 19025 4255 19043 4289
rect 19097 4255 19111 4289
rect 19169 4255 19179 4289
rect 19241 4255 19247 4289
rect 19313 4255 19315 4289
rect 19349 4255 19351 4289
rect 19417 4255 19423 4289
rect 19485 4255 19495 4289
rect 19553 4255 19567 4289
rect 19621 4255 19639 4289
rect 19689 4255 19711 4289
rect 19757 4255 19783 4289
rect 19825 4255 19855 4289
rect 19893 4255 19927 4289
rect 19961 4255 19995 4289
rect 20033 4255 20063 4289
rect 20105 4255 20131 4289
rect 20177 4255 20199 4289
rect 20249 4255 20267 4289
rect 20321 4255 20335 4289
rect 20393 4255 20403 4289
rect 20465 4255 20471 4289
rect 20537 4255 20539 4289
rect 20573 4255 20575 4289
rect 20641 4255 20647 4289
rect 20709 4255 20719 4289
rect 20777 4255 20791 4289
rect 20845 4255 20863 4289
rect 20913 4255 20935 4289
rect 20981 4255 21007 4289
rect 21049 4255 21079 4289
rect 21117 4255 21151 4289
rect 21185 4255 21219 4289
rect 21257 4255 21287 4289
rect 21329 4255 21355 4289
rect 21401 4255 21423 4289
rect 21473 4255 21491 4289
rect 21545 4255 21559 4289
rect 21617 4255 21627 4289
rect 21689 4255 21695 4289
rect 21761 4255 21763 4289
rect 21797 4255 21799 4289
rect 21865 4255 21871 4289
rect 21933 4255 21943 4289
rect 22001 4255 22015 4289
rect 22069 4255 22087 4289
rect 22137 4255 22159 4289
rect 22205 4255 22231 4289
rect 22273 4255 22303 4289
rect 22341 4255 22375 4289
rect 22409 4255 22443 4289
rect 22481 4255 22511 4289
rect 22553 4255 22579 4289
rect 22625 4255 22647 4289
rect 22697 4255 22715 4289
rect 22769 4255 22783 4289
rect 22841 4255 22851 4289
rect 22913 4255 22919 4289
rect 22985 4255 22987 4289
rect 23021 4255 23023 4289
rect 23089 4255 23095 4289
rect 23157 4255 23167 4289
rect 23225 4255 23239 4289
rect 23293 4255 23311 4289
rect 23361 4255 23383 4289
rect 23429 4255 23455 4289
rect 23497 4255 23527 4289
rect 23565 4255 23599 4289
rect 23633 4255 23667 4289
rect 23705 4255 23735 4289
rect 23777 4255 23803 4289
rect 23849 4255 23871 4289
rect 23921 4255 23939 4289
rect 23993 4255 24007 4289
rect 24065 4255 24075 4289
rect 24137 4255 24143 4289
rect 24209 4255 24211 4289
rect 24245 4255 24247 4289
rect 24313 4255 24319 4289
rect 24381 4255 24391 4289
rect 24449 4255 24463 4289
rect 24517 4255 24535 4289
rect 24585 4255 24607 4289
rect 24653 4255 24679 4289
rect 24713 4255 24822 4289
rect 378 4222 24822 4255
rect 378 4144 478 4222
rect 378 4110 411 4144
rect 445 4110 478 4144
rect 378 4076 478 4110
rect 378 4042 411 4076
rect 445 4042 478 4076
rect 378 4008 478 4042
rect 378 3974 411 4008
rect 445 3974 478 4008
rect 378 3940 478 3974
rect 378 3906 411 3940
rect 445 3906 478 3940
rect 378 3872 478 3906
rect 378 3838 411 3872
rect 445 3838 478 3872
rect 378 3804 478 3838
rect 378 3770 411 3804
rect 445 3770 478 3804
rect 378 3736 478 3770
rect 378 3702 411 3736
rect 445 3702 478 3736
rect 378 3700 478 3702
rect 378 3634 411 3700
rect 445 3634 478 3700
rect 378 3628 478 3634
rect 378 3566 411 3628
rect 445 3566 478 3628
rect 378 3556 478 3566
rect 378 3498 411 3556
rect 445 3498 478 3556
rect 378 3484 478 3498
rect 378 3430 411 3484
rect 445 3430 478 3484
rect 378 3412 478 3430
rect 378 3362 411 3412
rect 445 3362 478 3412
rect 378 3340 478 3362
rect 378 3294 411 3340
rect 445 3294 478 3340
rect 378 3268 478 3294
rect 378 3226 411 3268
rect 445 3226 478 3268
rect 378 3196 478 3226
rect 378 3158 411 3196
rect 445 3158 478 3196
rect 378 3124 478 3158
rect 378 3090 411 3124
rect 445 3090 478 3124
rect 378 3056 478 3090
rect 378 3018 411 3056
rect 445 3018 478 3056
rect 378 2988 478 3018
rect 378 2946 411 2988
rect 445 2946 478 2988
rect 378 2920 478 2946
rect 378 2874 411 2920
rect 445 2874 478 2920
rect 378 2852 478 2874
rect 378 2802 411 2852
rect 445 2802 478 2852
rect 378 2784 478 2802
rect 378 2730 411 2784
rect 445 2730 478 2784
rect 378 2716 478 2730
rect 378 2658 411 2716
rect 445 2658 478 2716
rect 378 2648 478 2658
rect 378 2586 411 2648
rect 445 2586 478 2648
rect 378 2580 478 2586
rect 378 2514 411 2580
rect 445 2514 478 2580
rect 378 2512 478 2514
rect 378 2478 411 2512
rect 445 2478 478 2512
rect 378 2476 478 2478
rect 378 2410 411 2476
rect 445 2410 478 2476
rect 378 2404 478 2410
rect 378 2342 411 2404
rect 445 2342 478 2404
rect 378 2332 478 2342
rect 378 2274 411 2332
rect 445 2274 478 2332
rect 378 2260 478 2274
rect 378 2206 411 2260
rect 445 2206 478 2260
rect 378 2188 478 2206
rect 378 2138 411 2188
rect 445 2138 478 2188
rect 378 2116 478 2138
rect 378 2070 411 2116
rect 445 2070 478 2116
rect 378 2044 478 2070
rect 378 2002 411 2044
rect 445 2002 478 2044
rect 378 1972 478 2002
rect 378 1934 411 1972
rect 445 1934 478 1972
rect 378 1900 478 1934
rect 378 1866 411 1900
rect 445 1866 478 1900
rect 378 1832 478 1866
rect 378 1794 411 1832
rect 445 1794 478 1832
rect 378 1764 478 1794
rect 378 1722 411 1764
rect 445 1722 478 1764
rect 378 1696 478 1722
rect 378 1650 411 1696
rect 445 1650 478 1696
rect 378 1628 478 1650
rect 378 1578 411 1628
rect 445 1578 478 1628
rect 378 1560 478 1578
rect 378 1506 411 1560
rect 445 1506 478 1560
rect 378 1492 478 1506
rect 378 1434 411 1492
rect 445 1434 478 1492
rect 378 1424 478 1434
rect 378 1362 411 1424
rect 445 1362 478 1424
rect 378 1356 478 1362
rect 378 1290 411 1356
rect 445 1290 478 1356
rect 378 1288 478 1290
rect 378 1254 411 1288
rect 445 1254 478 1288
rect 378 1252 478 1254
rect 378 1186 411 1252
rect 445 1186 478 1252
rect 378 1180 478 1186
rect 378 1118 411 1180
rect 445 1118 478 1180
rect 378 1108 478 1118
rect 378 1050 411 1108
rect 445 1050 478 1108
rect 378 1036 478 1050
rect 378 982 411 1036
rect 445 982 478 1036
rect 378 964 478 982
rect 378 914 411 964
rect 445 914 478 964
rect 378 892 478 914
rect 378 846 411 892
rect 445 846 478 892
rect 378 820 478 846
rect 378 778 411 820
rect 445 778 478 820
rect 378 748 478 778
rect 378 710 411 748
rect 445 710 478 748
rect 378 676 478 710
rect 378 642 411 676
rect 445 642 478 676
rect 378 608 478 642
rect 378 570 411 608
rect 445 570 478 608
rect 378 540 478 570
rect 378 498 411 540
rect 445 498 478 540
rect 378 472 478 498
rect 378 426 411 472
rect 445 426 478 472
rect 378 404 478 426
rect 378 354 411 404
rect 445 354 478 404
rect 378 336 478 354
rect 378 282 411 336
rect 445 282 478 336
rect 378 268 478 282
rect 378 210 411 268
rect 445 210 478 268
rect 378 200 478 210
rect 378 138 411 200
rect 445 138 478 200
rect 378 132 478 138
rect 378 66 411 132
rect 445 66 478 132
rect 378 64 478 66
rect 378 30 411 64
rect 445 30 478 64
rect 378 28 478 30
rect 378 -38 411 28
rect 445 -38 478 28
rect 378 -44 478 -38
rect 378 -106 411 -44
rect 445 -106 478 -44
rect 378 -116 478 -106
rect 378 -174 411 -116
rect 445 -174 478 -116
rect 378 -188 478 -174
rect 378 -242 411 -188
rect 445 -242 478 -188
rect 378 -260 478 -242
rect 378 -310 411 -260
rect 445 -310 478 -260
rect 378 -332 478 -310
rect 378 -378 411 -332
rect 445 -378 478 -332
rect 378 -404 478 -378
rect 378 -446 411 -404
rect 445 -446 478 -404
rect 378 -476 478 -446
rect 378 -514 411 -476
rect 445 -514 478 -476
rect 378 -548 478 -514
rect 378 -582 411 -548
rect 445 -582 478 -548
rect 378 -616 478 -582
rect 378 -654 411 -616
rect 445 -654 478 -616
rect 378 -684 478 -654
rect 378 -726 411 -684
rect 445 -726 478 -684
rect 378 -752 478 -726
rect 378 -798 411 -752
rect 445 -798 478 -752
rect 378 -820 478 -798
rect 378 -870 411 -820
rect 445 -870 478 -820
rect 378 -888 478 -870
rect 378 -942 411 -888
rect 445 -942 478 -888
rect 378 -956 478 -942
rect 378 -1014 411 -956
rect 445 -1014 478 -956
rect 378 -1024 478 -1014
rect 378 -1086 411 -1024
rect 445 -1086 478 -1024
rect 378 -1092 478 -1086
rect 378 -1158 411 -1092
rect 445 -1158 478 -1092
rect 378 -1160 478 -1158
rect 378 -1194 411 -1160
rect 445 -1194 478 -1160
rect 378 -1196 478 -1194
rect 378 -1262 411 -1196
rect 445 -1262 478 -1196
rect 378 -1268 478 -1262
rect 378 -1330 411 -1268
rect 445 -1330 478 -1268
rect 378 -1340 478 -1330
rect 378 -1398 411 -1340
rect 445 -1398 478 -1340
rect 378 -1412 478 -1398
rect 378 -1466 411 -1412
rect 445 -1466 478 -1412
rect 378 -1484 478 -1466
rect 378 -1534 411 -1484
rect 445 -1534 478 -1484
rect 378 -1556 478 -1534
rect 378 -1602 411 -1556
rect 445 -1602 478 -1556
rect 378 -1628 478 -1602
rect 378 -1670 411 -1628
rect 445 -1670 478 -1628
rect 378 -1700 478 -1670
rect 378 -1738 411 -1700
rect 445 -1738 478 -1700
rect 378 -1772 478 -1738
rect 378 -1806 411 -1772
rect 445 -1806 478 -1772
rect 378 -1840 478 -1806
rect 378 -1878 411 -1840
rect 445 -1878 478 -1840
rect 378 -1908 478 -1878
rect 378 -1950 411 -1908
rect 445 -1950 478 -1908
rect 378 -1976 478 -1950
rect 378 -2022 411 -1976
rect 445 -2022 478 -1976
rect 378 -2044 478 -2022
rect 378 -2094 411 -2044
rect 445 -2094 478 -2044
rect 378 -2112 478 -2094
rect 378 -2166 411 -2112
rect 445 -2166 478 -2112
rect 378 -2180 478 -2166
rect 378 -2238 411 -2180
rect 445 -2238 478 -2180
rect 378 -2248 478 -2238
rect 378 -2310 411 -2248
rect 445 -2310 478 -2248
rect 378 -2316 478 -2310
rect 378 -2382 411 -2316
rect 445 -2382 478 -2316
rect 378 -2384 478 -2382
rect 378 -2418 411 -2384
rect 445 -2418 478 -2384
rect 378 -2420 478 -2418
rect 378 -2486 411 -2420
rect 445 -2486 478 -2420
rect 378 -2492 478 -2486
rect 378 -2554 411 -2492
rect 445 -2554 478 -2492
rect 378 -2564 478 -2554
rect 378 -2622 411 -2564
rect 445 -2622 478 -2564
rect 378 -2636 478 -2622
rect 378 -2690 411 -2636
rect 445 -2690 478 -2636
rect 378 -2708 478 -2690
rect 378 -2758 411 -2708
rect 445 -2758 478 -2708
rect 378 -2780 478 -2758
rect 378 -2826 411 -2780
rect 445 -2826 478 -2780
rect 378 -2852 478 -2826
rect 378 -2894 411 -2852
rect 445 -2894 478 -2852
rect 378 -2924 478 -2894
rect 378 -2962 411 -2924
rect 445 -2962 478 -2924
rect 378 -2996 478 -2962
rect 378 -3030 411 -2996
rect 445 -3030 478 -2996
rect 378 -3064 478 -3030
rect 378 -3102 411 -3064
rect 445 -3102 478 -3064
rect 378 -3132 478 -3102
rect 378 -3174 411 -3132
rect 445 -3174 478 -3132
rect 378 -3200 478 -3174
rect 378 -3246 411 -3200
rect 445 -3246 478 -3200
rect 378 -3268 478 -3246
rect 378 -3318 411 -3268
rect 445 -3318 478 -3268
rect 378 -3336 478 -3318
rect 378 -3390 411 -3336
rect 445 -3390 478 -3336
rect 378 -3404 478 -3390
rect 378 -3462 411 -3404
rect 445 -3462 478 -3404
rect 378 -3472 478 -3462
rect 378 -3534 411 -3472
rect 445 -3534 478 -3472
rect 378 -3540 478 -3534
rect 378 -3606 411 -3540
rect 445 -3606 478 -3540
rect 378 -3608 478 -3606
rect 378 -3642 411 -3608
rect 445 -3642 478 -3608
rect 378 -3644 478 -3642
rect 378 -3710 411 -3644
rect 445 -3710 478 -3644
rect 378 -3716 478 -3710
rect 378 -3778 411 -3716
rect 445 -3778 478 -3716
rect 378 -3788 478 -3778
rect 378 -3846 411 -3788
rect 445 -3846 478 -3788
rect 378 -3860 478 -3846
rect 378 -3914 411 -3860
rect 445 -3914 478 -3860
rect 378 -3932 478 -3914
rect 378 -3982 411 -3932
rect 445 -3982 478 -3932
rect 378 -4004 478 -3982
rect 378 -4050 411 -4004
rect 445 -4050 478 -4004
rect 378 -4076 478 -4050
rect 378 -4118 411 -4076
rect 445 -4118 478 -4076
rect 378 -4148 478 -4118
rect 378 -4186 411 -4148
rect 445 -4186 478 -4148
rect 378 -4220 478 -4186
rect 378 -4254 411 -4220
rect 445 -4254 478 -4220
rect 378 -4288 478 -4254
rect 378 -4326 411 -4288
rect 445 -4326 478 -4288
rect 378 -4356 478 -4326
rect 378 -4398 411 -4356
rect 445 -4398 478 -4356
rect 378 -4424 478 -4398
rect 378 -4470 411 -4424
rect 445 -4470 478 -4424
rect 378 -4492 478 -4470
rect 378 -4542 411 -4492
rect 445 -4542 478 -4492
rect 378 -4560 478 -4542
rect 378 -4614 411 -4560
rect 445 -4614 478 -4560
rect 378 -4628 478 -4614
rect 378 -4686 411 -4628
rect 445 -4686 478 -4628
rect 378 -4696 478 -4686
rect 378 -4758 411 -4696
rect 445 -4758 478 -4696
rect 378 -4764 478 -4758
rect 378 -4830 411 -4764
rect 445 -4830 478 -4764
rect 378 -4832 478 -4830
rect 378 -4866 411 -4832
rect 445 -4866 478 -4832
rect 378 -4868 478 -4866
rect 378 -4934 411 -4868
rect 445 -4934 478 -4868
rect 378 -4940 478 -4934
rect 378 -5002 411 -4940
rect 445 -5002 478 -4940
rect 378 -5012 478 -5002
rect 378 -5070 411 -5012
rect 445 -5070 478 -5012
rect 378 -5084 478 -5070
rect 378 -5138 411 -5084
rect 445 -5138 478 -5084
rect 378 -5156 478 -5138
rect 378 -5206 411 -5156
rect 445 -5206 478 -5156
rect 378 -5228 478 -5206
rect 378 -5274 411 -5228
rect 445 -5274 478 -5228
rect 378 -5300 478 -5274
rect 378 -5342 411 -5300
rect 445 -5342 478 -5300
rect 378 -5372 478 -5342
rect 378 -5410 411 -5372
rect 445 -5410 478 -5372
rect 378 -5444 478 -5410
rect 378 -5478 411 -5444
rect 445 -5478 478 -5444
rect 378 -5512 478 -5478
rect 378 -5550 411 -5512
rect 445 -5550 478 -5512
rect 378 -5580 478 -5550
rect 378 -5622 411 -5580
rect 445 -5622 478 -5580
rect 378 -5648 478 -5622
rect 378 -5694 411 -5648
rect 445 -5694 478 -5648
rect 378 -5716 478 -5694
rect 378 -5766 411 -5716
rect 445 -5766 478 -5716
rect 378 -5784 478 -5766
rect 378 -5838 411 -5784
rect 445 -5838 478 -5784
rect 378 -5852 478 -5838
rect 378 -5910 411 -5852
rect 445 -5910 478 -5852
rect 378 -5920 478 -5910
rect 378 -5982 411 -5920
rect 445 -5982 478 -5920
rect 378 -5988 478 -5982
rect 378 -6054 411 -5988
rect 445 -6054 478 -5988
rect 378 -6056 478 -6054
rect 378 -6090 411 -6056
rect 445 -6090 478 -6056
rect 378 -6092 478 -6090
rect 378 -6158 411 -6092
rect 445 -6158 478 -6092
rect 378 -6164 478 -6158
rect 378 -6226 411 -6164
rect 445 -6226 478 -6164
rect 378 -6236 478 -6226
rect 378 -6294 411 -6236
rect 445 -6294 478 -6236
rect 378 -6308 478 -6294
rect 378 -6362 411 -6308
rect 445 -6362 478 -6308
rect 378 -6380 478 -6362
rect 378 -6430 411 -6380
rect 445 -6430 478 -6380
rect 378 -6452 478 -6430
rect 378 -6498 411 -6452
rect 445 -6498 478 -6452
rect 378 -6524 478 -6498
rect 378 -6566 411 -6524
rect 445 -6566 478 -6524
rect 378 -6596 478 -6566
rect 378 -6634 411 -6596
rect 445 -6634 478 -6596
rect 378 -6668 478 -6634
rect 378 -6702 411 -6668
rect 445 -6702 478 -6668
rect 378 -6736 478 -6702
rect 378 -6774 411 -6736
rect 445 -6774 478 -6736
rect 378 -6804 478 -6774
rect 378 -6846 411 -6804
rect 445 -6846 478 -6804
rect 378 -6872 478 -6846
rect 378 -6918 411 -6872
rect 445 -6918 478 -6872
rect 378 -6940 478 -6918
rect 378 -6990 411 -6940
rect 445 -6990 478 -6940
rect 378 -7008 478 -6990
rect 378 -7062 411 -7008
rect 445 -7062 478 -7008
rect 378 -7076 478 -7062
rect 378 -7134 411 -7076
rect 445 -7134 478 -7076
rect 378 -7144 478 -7134
rect 378 -7206 411 -7144
rect 445 -7206 478 -7144
rect 378 -7212 478 -7206
rect 378 -7278 411 -7212
rect 445 -7278 478 -7212
rect 378 -7280 478 -7278
rect 378 -7314 411 -7280
rect 445 -7314 478 -7280
rect 378 -7316 478 -7314
rect 378 -7382 411 -7316
rect 445 -7382 478 -7316
rect 378 -7388 478 -7382
rect 378 -7450 411 -7388
rect 445 -7450 478 -7388
rect 378 -7460 478 -7450
rect 378 -7518 411 -7460
rect 445 -7518 478 -7460
rect 378 -7532 478 -7518
rect 378 -7586 411 -7532
rect 445 -7586 478 -7532
rect 378 -7604 478 -7586
rect 378 -7654 411 -7604
rect 445 -7654 478 -7604
rect 378 -7676 478 -7654
rect 378 -7722 411 -7676
rect 445 -7722 478 -7676
rect 378 -7748 478 -7722
rect 378 -7790 411 -7748
rect 445 -7790 478 -7748
rect 378 -7820 478 -7790
rect 378 -7858 411 -7820
rect 445 -7858 478 -7820
rect 378 -7892 478 -7858
rect 378 -7926 411 -7892
rect 445 -7926 478 -7892
rect 378 -7960 478 -7926
rect 378 -7998 411 -7960
rect 445 -7998 478 -7960
rect 378 -8028 478 -7998
rect 378 -8070 411 -8028
rect 445 -8070 478 -8028
rect 378 -8096 478 -8070
rect 378 -8142 411 -8096
rect 445 -8142 478 -8096
rect 378 -8164 478 -8142
rect 378 -8214 411 -8164
rect 445 -8214 478 -8164
rect 378 -8232 478 -8214
rect 378 -8286 411 -8232
rect 445 -8286 478 -8232
rect 378 -8300 478 -8286
rect 378 -8358 411 -8300
rect 445 -8358 478 -8300
rect 378 -8368 478 -8358
rect 378 -8430 411 -8368
rect 445 -8430 478 -8368
rect 378 -8436 478 -8430
rect 378 -8502 411 -8436
rect 445 -8502 478 -8436
rect 378 -8504 478 -8502
rect 378 -8538 411 -8504
rect 445 -8538 478 -8504
rect 378 -8540 478 -8538
rect 378 -8606 411 -8540
rect 445 -8606 478 -8540
rect 378 -8612 478 -8606
rect 378 -8674 411 -8612
rect 445 -8674 478 -8612
rect 378 -8684 478 -8674
rect 378 -8742 411 -8684
rect 445 -8742 478 -8684
rect 378 -8756 478 -8742
rect 378 -8810 411 -8756
rect 445 -8810 478 -8756
rect 378 -8828 478 -8810
rect 378 -8878 411 -8828
rect 445 -8878 478 -8828
rect 378 -8900 478 -8878
rect 378 -8946 411 -8900
rect 445 -8946 478 -8900
rect 378 -8972 478 -8946
rect 378 -9014 411 -8972
rect 445 -9014 478 -8972
rect 378 -9044 478 -9014
rect 378 -9082 411 -9044
rect 445 -9082 478 -9044
rect 378 -9116 478 -9082
rect 378 -9150 411 -9116
rect 445 -9150 478 -9116
rect 378 -9184 478 -9150
rect 378 -9222 411 -9184
rect 445 -9222 478 -9184
rect 378 -9252 478 -9222
rect 378 -9294 411 -9252
rect 445 -9294 478 -9252
rect 378 -9320 478 -9294
rect 378 -9366 411 -9320
rect 445 -9366 478 -9320
rect 378 -9388 478 -9366
rect 378 -9438 411 -9388
rect 445 -9438 478 -9388
rect 378 -9456 478 -9438
rect 378 -9510 411 -9456
rect 445 -9510 478 -9456
rect 378 -9524 478 -9510
rect 378 -9582 411 -9524
rect 445 -9582 478 -9524
rect 378 -9592 478 -9582
rect 378 -9654 411 -9592
rect 445 -9654 478 -9592
rect 378 -9660 478 -9654
rect 378 -9726 411 -9660
rect 445 -9726 478 -9660
rect 378 -9728 478 -9726
rect 378 -9762 411 -9728
rect 445 -9762 478 -9728
rect 378 -9796 478 -9762
rect 378 -9830 411 -9796
rect 445 -9830 478 -9796
rect 378 -9864 478 -9830
rect 378 -9898 411 -9864
rect 445 -9898 478 -9864
rect 378 -9932 478 -9898
rect 378 -9966 411 -9932
rect 445 -9966 478 -9932
rect 378 -10000 478 -9966
rect 378 -10034 411 -10000
rect 445 -10034 478 -10000
rect 378 -10068 478 -10034
rect 378 -10102 411 -10068
rect 445 -10102 478 -10068
rect 378 -10136 478 -10102
rect 378 -10170 411 -10136
rect 445 -10170 478 -10136
rect 378 -10248 478 -10170
rect 24722 4144 24822 4222
rect 24722 4110 24755 4144
rect 24789 4110 24822 4144
rect 24722 4076 24822 4110
rect 24722 4042 24755 4076
rect 24789 4042 24822 4076
rect 24722 4008 24822 4042
rect 24722 3974 24755 4008
rect 24789 3974 24822 4008
rect 24722 3940 24822 3974
rect 24722 3906 24755 3940
rect 24789 3906 24822 3940
rect 24722 3872 24822 3906
rect 24722 3838 24755 3872
rect 24789 3838 24822 3872
rect 24722 3804 24822 3838
rect 24722 3770 24755 3804
rect 24789 3770 24822 3804
rect 24722 3736 24822 3770
rect 24722 3702 24755 3736
rect 24789 3702 24822 3736
rect 24722 3700 24822 3702
rect 24722 3634 24755 3700
rect 24789 3634 24822 3700
rect 24722 3628 24822 3634
rect 24722 3566 24755 3628
rect 24789 3566 24822 3628
rect 24722 3556 24822 3566
rect 24722 3498 24755 3556
rect 24789 3498 24822 3556
rect 24722 3484 24822 3498
rect 24722 3430 24755 3484
rect 24789 3430 24822 3484
rect 24722 3412 24822 3430
rect 24722 3362 24755 3412
rect 24789 3362 24822 3412
rect 24722 3340 24822 3362
rect 24722 3294 24755 3340
rect 24789 3294 24822 3340
rect 24722 3268 24822 3294
rect 24722 3226 24755 3268
rect 24789 3226 24822 3268
rect 24722 3196 24822 3226
rect 24722 3158 24755 3196
rect 24789 3158 24822 3196
rect 24722 3124 24822 3158
rect 24722 3090 24755 3124
rect 24789 3090 24822 3124
rect 24722 3056 24822 3090
rect 24722 3018 24755 3056
rect 24789 3018 24822 3056
rect 24722 2988 24822 3018
rect 24722 2946 24755 2988
rect 24789 2946 24822 2988
rect 24722 2920 24822 2946
rect 24722 2874 24755 2920
rect 24789 2874 24822 2920
rect 24722 2852 24822 2874
rect 24722 2802 24755 2852
rect 24789 2802 24822 2852
rect 24722 2784 24822 2802
rect 24722 2730 24755 2784
rect 24789 2730 24822 2784
rect 24722 2716 24822 2730
rect 24722 2658 24755 2716
rect 24789 2658 24822 2716
rect 24722 2648 24822 2658
rect 24722 2586 24755 2648
rect 24789 2586 24822 2648
rect 24722 2580 24822 2586
rect 24722 2514 24755 2580
rect 24789 2514 24822 2580
rect 24722 2512 24822 2514
rect 24722 2478 24755 2512
rect 24789 2478 24822 2512
rect 24722 2476 24822 2478
rect 24722 2410 24755 2476
rect 24789 2410 24822 2476
rect 24722 2404 24822 2410
rect 24722 2342 24755 2404
rect 24789 2342 24822 2404
rect 24722 2332 24822 2342
rect 24722 2274 24755 2332
rect 24789 2274 24822 2332
rect 24722 2260 24822 2274
rect 24722 2206 24755 2260
rect 24789 2206 24822 2260
rect 24722 2188 24822 2206
rect 24722 2138 24755 2188
rect 24789 2138 24822 2188
rect 24722 2116 24822 2138
rect 24722 2070 24755 2116
rect 24789 2070 24822 2116
rect 24722 2044 24822 2070
rect 24722 2002 24755 2044
rect 24789 2002 24822 2044
rect 24722 1972 24822 2002
rect 24722 1934 24755 1972
rect 24789 1934 24822 1972
rect 24722 1900 24822 1934
rect 24722 1866 24755 1900
rect 24789 1866 24822 1900
rect 24722 1832 24822 1866
rect 24722 1794 24755 1832
rect 24789 1794 24822 1832
rect 24722 1764 24822 1794
rect 24722 1722 24755 1764
rect 24789 1722 24822 1764
rect 24722 1696 24822 1722
rect 24722 1650 24755 1696
rect 24789 1650 24822 1696
rect 24722 1628 24822 1650
rect 24722 1578 24755 1628
rect 24789 1578 24822 1628
rect 24722 1560 24822 1578
rect 24722 1506 24755 1560
rect 24789 1506 24822 1560
rect 24722 1492 24822 1506
rect 24722 1434 24755 1492
rect 24789 1434 24822 1492
rect 24722 1424 24822 1434
rect 24722 1362 24755 1424
rect 24789 1362 24822 1424
rect 24722 1356 24822 1362
rect 24722 1290 24755 1356
rect 24789 1290 24822 1356
rect 24722 1288 24822 1290
rect 24722 1254 24755 1288
rect 24789 1254 24822 1288
rect 24722 1252 24822 1254
rect 24722 1186 24755 1252
rect 24789 1186 24822 1252
rect 24722 1180 24822 1186
rect 24722 1118 24755 1180
rect 24789 1118 24822 1180
rect 24722 1108 24822 1118
rect 24722 1050 24755 1108
rect 24789 1050 24822 1108
rect 24722 1036 24822 1050
rect 24722 982 24755 1036
rect 24789 982 24822 1036
rect 24722 964 24822 982
rect 24722 914 24755 964
rect 24789 914 24822 964
rect 24722 892 24822 914
rect 24722 846 24755 892
rect 24789 846 24822 892
rect 24722 820 24822 846
rect 24722 778 24755 820
rect 24789 778 24822 820
rect 24722 748 24822 778
rect 24722 710 24755 748
rect 24789 710 24822 748
rect 24722 676 24822 710
rect 24722 642 24755 676
rect 24789 642 24822 676
rect 24722 608 24822 642
rect 24722 570 24755 608
rect 24789 570 24822 608
rect 24722 540 24822 570
rect 24722 498 24755 540
rect 24789 498 24822 540
rect 24722 472 24822 498
rect 24722 426 24755 472
rect 24789 426 24822 472
rect 24722 404 24822 426
rect 24722 354 24755 404
rect 24789 354 24822 404
rect 24722 336 24822 354
rect 24722 282 24755 336
rect 24789 282 24822 336
rect 24722 268 24822 282
rect 24722 210 24755 268
rect 24789 210 24822 268
rect 24722 200 24822 210
rect 24722 138 24755 200
rect 24789 138 24822 200
rect 24722 132 24822 138
rect 24722 66 24755 132
rect 24789 66 24822 132
rect 24722 64 24822 66
rect 24722 30 24755 64
rect 24789 30 24822 64
rect 24722 28 24822 30
rect 24722 -38 24755 28
rect 24789 -38 24822 28
rect 24722 -44 24822 -38
rect 24722 -106 24755 -44
rect 24789 -106 24822 -44
rect 24722 -116 24822 -106
rect 24722 -174 24755 -116
rect 24789 -174 24822 -116
rect 24722 -188 24822 -174
rect 24722 -242 24755 -188
rect 24789 -242 24822 -188
rect 24722 -260 24822 -242
rect 24722 -310 24755 -260
rect 24789 -310 24822 -260
rect 24722 -332 24822 -310
rect 24722 -378 24755 -332
rect 24789 -378 24822 -332
rect 24722 -404 24822 -378
rect 24722 -446 24755 -404
rect 24789 -446 24822 -404
rect 24722 -476 24822 -446
rect 24722 -514 24755 -476
rect 24789 -514 24822 -476
rect 24722 -548 24822 -514
rect 24722 -582 24755 -548
rect 24789 -582 24822 -548
rect 24722 -616 24822 -582
rect 24722 -654 24755 -616
rect 24789 -654 24822 -616
rect 24722 -684 24822 -654
rect 24722 -726 24755 -684
rect 24789 -726 24822 -684
rect 24722 -752 24822 -726
rect 24722 -798 24755 -752
rect 24789 -798 24822 -752
rect 24722 -820 24822 -798
rect 24722 -870 24755 -820
rect 24789 -870 24822 -820
rect 24722 -888 24822 -870
rect 24722 -942 24755 -888
rect 24789 -942 24822 -888
rect 24722 -956 24822 -942
rect 24722 -1014 24755 -956
rect 24789 -1014 24822 -956
rect 24722 -1024 24822 -1014
rect 24722 -1086 24755 -1024
rect 24789 -1086 24822 -1024
rect 24722 -1092 24822 -1086
rect 24722 -1158 24755 -1092
rect 24789 -1158 24822 -1092
rect 24722 -1160 24822 -1158
rect 24722 -1194 24755 -1160
rect 24789 -1194 24822 -1160
rect 24722 -1196 24822 -1194
rect 24722 -1262 24755 -1196
rect 24789 -1262 24822 -1196
rect 24722 -1268 24822 -1262
rect 24722 -1330 24755 -1268
rect 24789 -1330 24822 -1268
rect 24722 -1340 24822 -1330
rect 24722 -1398 24755 -1340
rect 24789 -1398 24822 -1340
rect 24722 -1412 24822 -1398
rect 24722 -1466 24755 -1412
rect 24789 -1466 24822 -1412
rect 24722 -1484 24822 -1466
rect 24722 -1534 24755 -1484
rect 24789 -1534 24822 -1484
rect 24722 -1556 24822 -1534
rect 24722 -1602 24755 -1556
rect 24789 -1602 24822 -1556
rect 24722 -1628 24822 -1602
rect 24722 -1670 24755 -1628
rect 24789 -1670 24822 -1628
rect 24722 -1700 24822 -1670
rect 24722 -1738 24755 -1700
rect 24789 -1738 24822 -1700
rect 24722 -1772 24822 -1738
rect 24722 -1806 24755 -1772
rect 24789 -1806 24822 -1772
rect 24722 -1840 24822 -1806
rect 24722 -1878 24755 -1840
rect 24789 -1878 24822 -1840
rect 24722 -1908 24822 -1878
rect 24722 -1950 24755 -1908
rect 24789 -1950 24822 -1908
rect 24722 -1976 24822 -1950
rect 24722 -2022 24755 -1976
rect 24789 -2022 24822 -1976
rect 24722 -2044 24822 -2022
rect 24722 -2094 24755 -2044
rect 24789 -2094 24822 -2044
rect 24722 -2112 24822 -2094
rect 24722 -2166 24755 -2112
rect 24789 -2166 24822 -2112
rect 24722 -2180 24822 -2166
rect 24722 -2238 24755 -2180
rect 24789 -2238 24822 -2180
rect 24722 -2248 24822 -2238
rect 24722 -2310 24755 -2248
rect 24789 -2310 24822 -2248
rect 24722 -2316 24822 -2310
rect 24722 -2382 24755 -2316
rect 24789 -2382 24822 -2316
rect 24722 -2384 24822 -2382
rect 24722 -2418 24755 -2384
rect 24789 -2418 24822 -2384
rect 24722 -2420 24822 -2418
rect 24722 -2486 24755 -2420
rect 24789 -2486 24822 -2420
rect 24722 -2492 24822 -2486
rect 24722 -2554 24755 -2492
rect 24789 -2554 24822 -2492
rect 24722 -2564 24822 -2554
rect 24722 -2622 24755 -2564
rect 24789 -2622 24822 -2564
rect 24722 -2636 24822 -2622
rect 24722 -2690 24755 -2636
rect 24789 -2690 24822 -2636
rect 24722 -2708 24822 -2690
rect 24722 -2758 24755 -2708
rect 24789 -2758 24822 -2708
rect 24722 -2780 24822 -2758
rect 24722 -2826 24755 -2780
rect 24789 -2826 24822 -2780
rect 24722 -2852 24822 -2826
rect 24722 -2894 24755 -2852
rect 24789 -2894 24822 -2852
rect 24722 -2924 24822 -2894
rect 24722 -2962 24755 -2924
rect 24789 -2962 24822 -2924
rect 24722 -2996 24822 -2962
rect 24722 -3030 24755 -2996
rect 24789 -3030 24822 -2996
rect 24722 -3064 24822 -3030
rect 24722 -3102 24755 -3064
rect 24789 -3102 24822 -3064
rect 24722 -3132 24822 -3102
rect 24722 -3174 24755 -3132
rect 24789 -3174 24822 -3132
rect 24722 -3200 24822 -3174
rect 24722 -3246 24755 -3200
rect 24789 -3246 24822 -3200
rect 24722 -3268 24822 -3246
rect 24722 -3318 24755 -3268
rect 24789 -3318 24822 -3268
rect 24722 -3336 24822 -3318
rect 24722 -3390 24755 -3336
rect 24789 -3390 24822 -3336
rect 24722 -3404 24822 -3390
rect 24722 -3462 24755 -3404
rect 24789 -3462 24822 -3404
rect 24722 -3472 24822 -3462
rect 24722 -3534 24755 -3472
rect 24789 -3534 24822 -3472
rect 24722 -3540 24822 -3534
rect 24722 -3606 24755 -3540
rect 24789 -3606 24822 -3540
rect 24722 -3608 24822 -3606
rect 24722 -3642 24755 -3608
rect 24789 -3642 24822 -3608
rect 24722 -3644 24822 -3642
rect 24722 -3710 24755 -3644
rect 24789 -3710 24822 -3644
rect 24722 -3716 24822 -3710
rect 24722 -3778 24755 -3716
rect 24789 -3778 24822 -3716
rect 24722 -3788 24822 -3778
rect 24722 -3846 24755 -3788
rect 24789 -3846 24822 -3788
rect 24722 -3860 24822 -3846
rect 24722 -3914 24755 -3860
rect 24789 -3914 24822 -3860
rect 24722 -3932 24822 -3914
rect 24722 -3982 24755 -3932
rect 24789 -3982 24822 -3932
rect 24722 -4004 24822 -3982
rect 24722 -4050 24755 -4004
rect 24789 -4050 24822 -4004
rect 24722 -4076 24822 -4050
rect 24722 -4118 24755 -4076
rect 24789 -4118 24822 -4076
rect 24722 -4148 24822 -4118
rect 24722 -4186 24755 -4148
rect 24789 -4186 24822 -4148
rect 24722 -4220 24822 -4186
rect 24722 -4254 24755 -4220
rect 24789 -4254 24822 -4220
rect 24722 -4288 24822 -4254
rect 24722 -4326 24755 -4288
rect 24789 -4326 24822 -4288
rect 24722 -4356 24822 -4326
rect 24722 -4398 24755 -4356
rect 24789 -4398 24822 -4356
rect 24722 -4424 24822 -4398
rect 24722 -4470 24755 -4424
rect 24789 -4470 24822 -4424
rect 24722 -4492 24822 -4470
rect 24722 -4542 24755 -4492
rect 24789 -4542 24822 -4492
rect 24722 -4560 24822 -4542
rect 24722 -4614 24755 -4560
rect 24789 -4614 24822 -4560
rect 24722 -4628 24822 -4614
rect 24722 -4686 24755 -4628
rect 24789 -4686 24822 -4628
rect 24722 -4696 24822 -4686
rect 24722 -4758 24755 -4696
rect 24789 -4758 24822 -4696
rect 24722 -4764 24822 -4758
rect 24722 -4830 24755 -4764
rect 24789 -4830 24822 -4764
rect 24722 -4832 24822 -4830
rect 24722 -4866 24755 -4832
rect 24789 -4866 24822 -4832
rect 24722 -4868 24822 -4866
rect 24722 -4934 24755 -4868
rect 24789 -4934 24822 -4868
rect 24722 -4940 24822 -4934
rect 24722 -5002 24755 -4940
rect 24789 -5002 24822 -4940
rect 24722 -5012 24822 -5002
rect 24722 -5070 24755 -5012
rect 24789 -5070 24822 -5012
rect 24722 -5084 24822 -5070
rect 24722 -5138 24755 -5084
rect 24789 -5138 24822 -5084
rect 24722 -5156 24822 -5138
rect 24722 -5206 24755 -5156
rect 24789 -5206 24822 -5156
rect 24722 -5228 24822 -5206
rect 24722 -5274 24755 -5228
rect 24789 -5274 24822 -5228
rect 24722 -5300 24822 -5274
rect 24722 -5342 24755 -5300
rect 24789 -5342 24822 -5300
rect 24722 -5372 24822 -5342
rect 24722 -5410 24755 -5372
rect 24789 -5410 24822 -5372
rect 24722 -5444 24822 -5410
rect 24722 -5478 24755 -5444
rect 24789 -5478 24822 -5444
rect 24722 -5512 24822 -5478
rect 24722 -5550 24755 -5512
rect 24789 -5550 24822 -5512
rect 24722 -5580 24822 -5550
rect 24722 -5622 24755 -5580
rect 24789 -5622 24822 -5580
rect 24722 -5648 24822 -5622
rect 24722 -5694 24755 -5648
rect 24789 -5694 24822 -5648
rect 24722 -5716 24822 -5694
rect 24722 -5766 24755 -5716
rect 24789 -5766 24822 -5716
rect 24722 -5784 24822 -5766
rect 24722 -5838 24755 -5784
rect 24789 -5838 24822 -5784
rect 24722 -5852 24822 -5838
rect 24722 -5910 24755 -5852
rect 24789 -5910 24822 -5852
rect 24722 -5920 24822 -5910
rect 24722 -5982 24755 -5920
rect 24789 -5982 24822 -5920
rect 24722 -5988 24822 -5982
rect 24722 -6054 24755 -5988
rect 24789 -6054 24822 -5988
rect 24722 -6056 24822 -6054
rect 24722 -6090 24755 -6056
rect 24789 -6090 24822 -6056
rect 24722 -6092 24822 -6090
rect 24722 -6158 24755 -6092
rect 24789 -6158 24822 -6092
rect 24722 -6164 24822 -6158
rect 24722 -6226 24755 -6164
rect 24789 -6226 24822 -6164
rect 24722 -6236 24822 -6226
rect 24722 -6294 24755 -6236
rect 24789 -6294 24822 -6236
rect 24722 -6308 24822 -6294
rect 24722 -6362 24755 -6308
rect 24789 -6362 24822 -6308
rect 24722 -6380 24822 -6362
rect 24722 -6430 24755 -6380
rect 24789 -6430 24822 -6380
rect 24722 -6452 24822 -6430
rect 24722 -6498 24755 -6452
rect 24789 -6498 24822 -6452
rect 24722 -6524 24822 -6498
rect 24722 -6566 24755 -6524
rect 24789 -6566 24822 -6524
rect 24722 -6596 24822 -6566
rect 24722 -6634 24755 -6596
rect 24789 -6634 24822 -6596
rect 24722 -6668 24822 -6634
rect 24722 -6702 24755 -6668
rect 24789 -6702 24822 -6668
rect 24722 -6736 24822 -6702
rect 24722 -6774 24755 -6736
rect 24789 -6774 24822 -6736
rect 24722 -6804 24822 -6774
rect 24722 -6846 24755 -6804
rect 24789 -6846 24822 -6804
rect 24722 -6872 24822 -6846
rect 24722 -6918 24755 -6872
rect 24789 -6918 24822 -6872
rect 24722 -6940 24822 -6918
rect 24722 -6990 24755 -6940
rect 24789 -6990 24822 -6940
rect 24722 -7008 24822 -6990
rect 24722 -7062 24755 -7008
rect 24789 -7062 24822 -7008
rect 24722 -7076 24822 -7062
rect 24722 -7134 24755 -7076
rect 24789 -7134 24822 -7076
rect 24722 -7144 24822 -7134
rect 24722 -7206 24755 -7144
rect 24789 -7206 24822 -7144
rect 24722 -7212 24822 -7206
rect 24722 -7278 24755 -7212
rect 24789 -7278 24822 -7212
rect 24722 -7280 24822 -7278
rect 24722 -7314 24755 -7280
rect 24789 -7314 24822 -7280
rect 24722 -7316 24822 -7314
rect 24722 -7382 24755 -7316
rect 24789 -7382 24822 -7316
rect 24722 -7388 24822 -7382
rect 24722 -7450 24755 -7388
rect 24789 -7450 24822 -7388
rect 24722 -7460 24822 -7450
rect 24722 -7518 24755 -7460
rect 24789 -7518 24822 -7460
rect 24722 -7532 24822 -7518
rect 24722 -7586 24755 -7532
rect 24789 -7586 24822 -7532
rect 24722 -7604 24822 -7586
rect 24722 -7654 24755 -7604
rect 24789 -7654 24822 -7604
rect 24722 -7676 24822 -7654
rect 24722 -7722 24755 -7676
rect 24789 -7722 24822 -7676
rect 24722 -7748 24822 -7722
rect 24722 -7790 24755 -7748
rect 24789 -7790 24822 -7748
rect 24722 -7820 24822 -7790
rect 24722 -7858 24755 -7820
rect 24789 -7858 24822 -7820
rect 24722 -7892 24822 -7858
rect 24722 -7926 24755 -7892
rect 24789 -7926 24822 -7892
rect 24722 -7960 24822 -7926
rect 24722 -7998 24755 -7960
rect 24789 -7998 24822 -7960
rect 24722 -8028 24822 -7998
rect 24722 -8070 24755 -8028
rect 24789 -8070 24822 -8028
rect 24722 -8096 24822 -8070
rect 24722 -8142 24755 -8096
rect 24789 -8142 24822 -8096
rect 24722 -8164 24822 -8142
rect 24722 -8214 24755 -8164
rect 24789 -8214 24822 -8164
rect 24722 -8232 24822 -8214
rect 24722 -8286 24755 -8232
rect 24789 -8286 24822 -8232
rect 24722 -8300 24822 -8286
rect 24722 -8358 24755 -8300
rect 24789 -8358 24822 -8300
rect 24722 -8368 24822 -8358
rect 24722 -8430 24755 -8368
rect 24789 -8430 24822 -8368
rect 24722 -8436 24822 -8430
rect 24722 -8502 24755 -8436
rect 24789 -8502 24822 -8436
rect 24722 -8504 24822 -8502
rect 24722 -8538 24755 -8504
rect 24789 -8538 24822 -8504
rect 24722 -8540 24822 -8538
rect 24722 -8606 24755 -8540
rect 24789 -8606 24822 -8540
rect 24722 -8612 24822 -8606
rect 24722 -8674 24755 -8612
rect 24789 -8674 24822 -8612
rect 24722 -8684 24822 -8674
rect 24722 -8742 24755 -8684
rect 24789 -8742 24822 -8684
rect 24722 -8756 24822 -8742
rect 24722 -8810 24755 -8756
rect 24789 -8810 24822 -8756
rect 24722 -8828 24822 -8810
rect 24722 -8878 24755 -8828
rect 24789 -8878 24822 -8828
rect 24722 -8900 24822 -8878
rect 24722 -8946 24755 -8900
rect 24789 -8946 24822 -8900
rect 24722 -8972 24822 -8946
rect 24722 -9014 24755 -8972
rect 24789 -9014 24822 -8972
rect 24722 -9044 24822 -9014
rect 24722 -9082 24755 -9044
rect 24789 -9082 24822 -9044
rect 24722 -9116 24822 -9082
rect 24722 -9150 24755 -9116
rect 24789 -9150 24822 -9116
rect 24722 -9184 24822 -9150
rect 24722 -9222 24755 -9184
rect 24789 -9222 24822 -9184
rect 24722 -9252 24822 -9222
rect 24722 -9294 24755 -9252
rect 24789 -9294 24822 -9252
rect 24722 -9320 24822 -9294
rect 24722 -9366 24755 -9320
rect 24789 -9366 24822 -9320
rect 24722 -9388 24822 -9366
rect 24722 -9438 24755 -9388
rect 24789 -9438 24822 -9388
rect 24722 -9456 24822 -9438
rect 24722 -9510 24755 -9456
rect 24789 -9510 24822 -9456
rect 24722 -9524 24822 -9510
rect 24722 -9582 24755 -9524
rect 24789 -9582 24822 -9524
rect 24722 -9592 24822 -9582
rect 24722 -9654 24755 -9592
rect 24789 -9654 24822 -9592
rect 24722 -9660 24822 -9654
rect 24722 -9726 24755 -9660
rect 24789 -9726 24822 -9660
rect 24722 -9728 24822 -9726
rect 24722 -9762 24755 -9728
rect 24789 -9762 24822 -9728
rect 24722 -9796 24822 -9762
rect 24722 -9830 24755 -9796
rect 24789 -9830 24822 -9796
rect 24722 -9864 24822 -9830
rect 24722 -9898 24755 -9864
rect 24789 -9898 24822 -9864
rect 24722 -9932 24822 -9898
rect 24722 -9966 24755 -9932
rect 24789 -9966 24822 -9932
rect 24722 -10000 24822 -9966
rect 24722 -10034 24755 -10000
rect 24789 -10034 24822 -10000
rect 24722 -10068 24822 -10034
rect 24722 -10102 24755 -10068
rect 24789 -10102 24822 -10068
rect 24722 -10136 24822 -10102
rect 24722 -10170 24755 -10136
rect 24789 -10170 24822 -10136
rect 24722 -10248 24822 -10170
rect 378 -10281 24822 -10248
rect 378 -10315 487 -10281
rect 521 -10315 547 -10281
rect 593 -10315 615 -10281
rect 665 -10315 683 -10281
rect 737 -10315 751 -10281
rect 809 -10315 819 -10281
rect 881 -10315 887 -10281
rect 953 -10315 955 -10281
rect 989 -10315 991 -10281
rect 1057 -10315 1063 -10281
rect 1125 -10315 1135 -10281
rect 1193 -10315 1207 -10281
rect 1261 -10315 1279 -10281
rect 1329 -10315 1351 -10281
rect 1397 -10315 1423 -10281
rect 1465 -10315 1495 -10281
rect 1533 -10315 1567 -10281
rect 1601 -10315 1635 -10281
rect 1673 -10315 1703 -10281
rect 1745 -10315 1771 -10281
rect 1817 -10315 1839 -10281
rect 1889 -10315 1907 -10281
rect 1961 -10315 1975 -10281
rect 2033 -10315 2043 -10281
rect 2105 -10315 2111 -10281
rect 2177 -10315 2179 -10281
rect 2213 -10315 2215 -10281
rect 2281 -10315 2287 -10281
rect 2349 -10315 2359 -10281
rect 2417 -10315 2431 -10281
rect 2485 -10315 2503 -10281
rect 2553 -10315 2575 -10281
rect 2621 -10315 2647 -10281
rect 2689 -10315 2719 -10281
rect 2757 -10315 2791 -10281
rect 2825 -10315 2859 -10281
rect 2897 -10315 2927 -10281
rect 2969 -10315 2995 -10281
rect 3041 -10315 3063 -10281
rect 3113 -10315 3131 -10281
rect 3185 -10315 3199 -10281
rect 3257 -10315 3267 -10281
rect 3329 -10315 3335 -10281
rect 3401 -10315 3403 -10281
rect 3437 -10315 3439 -10281
rect 3505 -10315 3511 -10281
rect 3573 -10315 3583 -10281
rect 3641 -10315 3655 -10281
rect 3709 -10315 3727 -10281
rect 3777 -10315 3799 -10281
rect 3845 -10315 3871 -10281
rect 3913 -10315 3943 -10281
rect 3981 -10315 4015 -10281
rect 4049 -10315 4083 -10281
rect 4121 -10315 4151 -10281
rect 4193 -10315 4219 -10281
rect 4265 -10315 4287 -10281
rect 4337 -10315 4355 -10281
rect 4409 -10315 4423 -10281
rect 4481 -10315 4491 -10281
rect 4553 -10315 4559 -10281
rect 4625 -10315 4627 -10281
rect 4661 -10315 4663 -10281
rect 4729 -10315 4735 -10281
rect 4797 -10315 4807 -10281
rect 4865 -10315 4879 -10281
rect 4933 -10315 4951 -10281
rect 5001 -10315 5023 -10281
rect 5069 -10315 5095 -10281
rect 5137 -10315 5167 -10281
rect 5205 -10315 5239 -10281
rect 5273 -10315 5307 -10281
rect 5345 -10315 5375 -10281
rect 5417 -10315 5443 -10281
rect 5489 -10315 5511 -10281
rect 5561 -10315 5579 -10281
rect 5633 -10315 5647 -10281
rect 5705 -10315 5715 -10281
rect 5777 -10315 5783 -10281
rect 5849 -10315 5851 -10281
rect 5885 -10315 5887 -10281
rect 5953 -10315 5959 -10281
rect 6021 -10315 6031 -10281
rect 6089 -10315 6103 -10281
rect 6157 -10315 6175 -10281
rect 6225 -10315 6247 -10281
rect 6293 -10315 6319 -10281
rect 6361 -10315 6391 -10281
rect 6429 -10315 6463 -10281
rect 6497 -10315 6531 -10281
rect 6569 -10315 6599 -10281
rect 6641 -10315 6667 -10281
rect 6713 -10315 6735 -10281
rect 6785 -10315 6803 -10281
rect 6857 -10315 6871 -10281
rect 6929 -10315 6939 -10281
rect 7001 -10315 7007 -10281
rect 7073 -10315 7075 -10281
rect 7109 -10315 7111 -10281
rect 7177 -10315 7183 -10281
rect 7245 -10315 7255 -10281
rect 7313 -10315 7327 -10281
rect 7381 -10315 7399 -10281
rect 7449 -10315 7471 -10281
rect 7517 -10315 7543 -10281
rect 7585 -10315 7615 -10281
rect 7653 -10315 7687 -10281
rect 7721 -10315 7755 -10281
rect 7793 -10315 7823 -10281
rect 7865 -10315 7891 -10281
rect 7937 -10315 7959 -10281
rect 8009 -10315 8027 -10281
rect 8081 -10315 8095 -10281
rect 8153 -10315 8163 -10281
rect 8225 -10315 8231 -10281
rect 8297 -10315 8299 -10281
rect 8333 -10315 8335 -10281
rect 8401 -10315 8407 -10281
rect 8469 -10315 8479 -10281
rect 8537 -10315 8551 -10281
rect 8605 -10315 8623 -10281
rect 8673 -10315 8695 -10281
rect 8741 -10315 8767 -10281
rect 8809 -10315 8839 -10281
rect 8877 -10315 8911 -10281
rect 8945 -10315 8979 -10281
rect 9017 -10315 9047 -10281
rect 9089 -10315 9115 -10281
rect 9161 -10315 9183 -10281
rect 9233 -10315 9251 -10281
rect 9305 -10315 9319 -10281
rect 9377 -10315 9387 -10281
rect 9449 -10315 9455 -10281
rect 9521 -10315 9523 -10281
rect 9557 -10315 9559 -10281
rect 9625 -10315 9631 -10281
rect 9693 -10315 9703 -10281
rect 9761 -10315 9775 -10281
rect 9829 -10315 9847 -10281
rect 9897 -10315 9919 -10281
rect 9965 -10315 9991 -10281
rect 10033 -10315 10063 -10281
rect 10101 -10315 10135 -10281
rect 10169 -10315 10203 -10281
rect 10241 -10315 10271 -10281
rect 10313 -10315 10339 -10281
rect 10385 -10315 10407 -10281
rect 10457 -10315 10475 -10281
rect 10529 -10315 10543 -10281
rect 10601 -10315 10611 -10281
rect 10673 -10315 10679 -10281
rect 10745 -10315 10747 -10281
rect 10781 -10315 10783 -10281
rect 10849 -10315 10855 -10281
rect 10917 -10315 10927 -10281
rect 10985 -10315 10999 -10281
rect 11053 -10315 11071 -10281
rect 11121 -10315 11143 -10281
rect 11189 -10315 11215 -10281
rect 11257 -10315 11287 -10281
rect 11325 -10315 11359 -10281
rect 11393 -10315 11427 -10281
rect 11465 -10315 11495 -10281
rect 11537 -10315 11563 -10281
rect 11609 -10315 11631 -10281
rect 11681 -10315 11699 -10281
rect 11753 -10315 11767 -10281
rect 11825 -10315 11835 -10281
rect 11897 -10315 11903 -10281
rect 11969 -10315 11971 -10281
rect 12005 -10315 12007 -10281
rect 12073 -10315 12079 -10281
rect 12141 -10315 12151 -10281
rect 12209 -10315 12223 -10281
rect 12277 -10315 12295 -10281
rect 12345 -10315 12367 -10281
rect 12413 -10315 12439 -10281
rect 12481 -10315 12511 -10281
rect 12549 -10315 12583 -10281
rect 12617 -10315 12651 -10281
rect 12689 -10315 12719 -10281
rect 12761 -10315 12787 -10281
rect 12833 -10315 12855 -10281
rect 12905 -10315 12923 -10281
rect 12977 -10315 12991 -10281
rect 13049 -10315 13059 -10281
rect 13121 -10315 13127 -10281
rect 13193 -10315 13195 -10281
rect 13229 -10315 13231 -10281
rect 13297 -10315 13303 -10281
rect 13365 -10315 13375 -10281
rect 13433 -10315 13447 -10281
rect 13501 -10315 13519 -10281
rect 13569 -10315 13591 -10281
rect 13637 -10315 13663 -10281
rect 13705 -10315 13735 -10281
rect 13773 -10315 13807 -10281
rect 13841 -10315 13875 -10281
rect 13913 -10315 13943 -10281
rect 13985 -10315 14011 -10281
rect 14057 -10315 14079 -10281
rect 14129 -10315 14147 -10281
rect 14201 -10315 14215 -10281
rect 14273 -10315 14283 -10281
rect 14345 -10315 14351 -10281
rect 14417 -10315 14419 -10281
rect 14453 -10315 14455 -10281
rect 14521 -10315 14527 -10281
rect 14589 -10315 14599 -10281
rect 14657 -10315 14671 -10281
rect 14725 -10315 14743 -10281
rect 14793 -10315 14815 -10281
rect 14861 -10315 14887 -10281
rect 14929 -10315 14959 -10281
rect 14997 -10315 15031 -10281
rect 15065 -10315 15099 -10281
rect 15137 -10315 15167 -10281
rect 15209 -10315 15235 -10281
rect 15281 -10315 15303 -10281
rect 15353 -10315 15371 -10281
rect 15425 -10315 15439 -10281
rect 15497 -10315 15507 -10281
rect 15569 -10315 15575 -10281
rect 15641 -10315 15643 -10281
rect 15677 -10315 15679 -10281
rect 15745 -10315 15751 -10281
rect 15813 -10315 15823 -10281
rect 15881 -10315 15895 -10281
rect 15949 -10315 15967 -10281
rect 16017 -10315 16039 -10281
rect 16085 -10315 16111 -10281
rect 16153 -10315 16183 -10281
rect 16221 -10315 16255 -10281
rect 16289 -10315 16323 -10281
rect 16361 -10315 16391 -10281
rect 16433 -10315 16459 -10281
rect 16505 -10315 16527 -10281
rect 16577 -10315 16595 -10281
rect 16649 -10315 16663 -10281
rect 16721 -10315 16731 -10281
rect 16793 -10315 16799 -10281
rect 16865 -10315 16867 -10281
rect 16901 -10315 16903 -10281
rect 16969 -10315 16975 -10281
rect 17037 -10315 17047 -10281
rect 17105 -10315 17119 -10281
rect 17173 -10315 17191 -10281
rect 17241 -10315 17263 -10281
rect 17309 -10315 17335 -10281
rect 17377 -10315 17407 -10281
rect 17445 -10315 17479 -10281
rect 17513 -10315 17547 -10281
rect 17585 -10315 17615 -10281
rect 17657 -10315 17683 -10281
rect 17729 -10315 17751 -10281
rect 17801 -10315 17819 -10281
rect 17873 -10315 17887 -10281
rect 17945 -10315 17955 -10281
rect 18017 -10315 18023 -10281
rect 18089 -10315 18091 -10281
rect 18125 -10315 18127 -10281
rect 18193 -10315 18199 -10281
rect 18261 -10315 18271 -10281
rect 18329 -10315 18343 -10281
rect 18397 -10315 18415 -10281
rect 18465 -10315 18487 -10281
rect 18533 -10315 18559 -10281
rect 18601 -10315 18631 -10281
rect 18669 -10315 18703 -10281
rect 18737 -10315 18771 -10281
rect 18809 -10315 18839 -10281
rect 18881 -10315 18907 -10281
rect 18953 -10315 18975 -10281
rect 19025 -10315 19043 -10281
rect 19097 -10315 19111 -10281
rect 19169 -10315 19179 -10281
rect 19241 -10315 19247 -10281
rect 19313 -10315 19315 -10281
rect 19349 -10315 19351 -10281
rect 19417 -10315 19423 -10281
rect 19485 -10315 19495 -10281
rect 19553 -10315 19567 -10281
rect 19621 -10315 19639 -10281
rect 19689 -10315 19711 -10281
rect 19757 -10315 19783 -10281
rect 19825 -10315 19855 -10281
rect 19893 -10315 19927 -10281
rect 19961 -10315 19995 -10281
rect 20033 -10315 20063 -10281
rect 20105 -10315 20131 -10281
rect 20177 -10315 20199 -10281
rect 20249 -10315 20267 -10281
rect 20321 -10315 20335 -10281
rect 20393 -10315 20403 -10281
rect 20465 -10315 20471 -10281
rect 20537 -10315 20539 -10281
rect 20573 -10315 20575 -10281
rect 20641 -10315 20647 -10281
rect 20709 -10315 20719 -10281
rect 20777 -10315 20791 -10281
rect 20845 -10315 20863 -10281
rect 20913 -10315 20935 -10281
rect 20981 -10315 21007 -10281
rect 21049 -10315 21079 -10281
rect 21117 -10315 21151 -10281
rect 21185 -10315 21219 -10281
rect 21257 -10315 21287 -10281
rect 21329 -10315 21355 -10281
rect 21401 -10315 21423 -10281
rect 21473 -10315 21491 -10281
rect 21545 -10315 21559 -10281
rect 21617 -10315 21627 -10281
rect 21689 -10315 21695 -10281
rect 21761 -10315 21763 -10281
rect 21797 -10315 21799 -10281
rect 21865 -10315 21871 -10281
rect 21933 -10315 21943 -10281
rect 22001 -10315 22015 -10281
rect 22069 -10315 22087 -10281
rect 22137 -10315 22159 -10281
rect 22205 -10315 22231 -10281
rect 22273 -10315 22303 -10281
rect 22341 -10315 22375 -10281
rect 22409 -10315 22443 -10281
rect 22481 -10315 22511 -10281
rect 22553 -10315 22579 -10281
rect 22625 -10315 22647 -10281
rect 22697 -10315 22715 -10281
rect 22769 -10315 22783 -10281
rect 22841 -10315 22851 -10281
rect 22913 -10315 22919 -10281
rect 22985 -10315 22987 -10281
rect 23021 -10315 23023 -10281
rect 23089 -10315 23095 -10281
rect 23157 -10315 23167 -10281
rect 23225 -10315 23239 -10281
rect 23293 -10315 23311 -10281
rect 23361 -10315 23383 -10281
rect 23429 -10315 23455 -10281
rect 23497 -10315 23527 -10281
rect 23565 -10315 23599 -10281
rect 23633 -10315 23667 -10281
rect 23705 -10315 23735 -10281
rect 23777 -10315 23803 -10281
rect 23849 -10315 23871 -10281
rect 23921 -10315 23939 -10281
rect 23993 -10315 24007 -10281
rect 24065 -10315 24075 -10281
rect 24137 -10315 24143 -10281
rect 24209 -10315 24211 -10281
rect 24245 -10315 24247 -10281
rect 24313 -10315 24319 -10281
rect 24381 -10315 24391 -10281
rect 24449 -10315 24463 -10281
rect 24517 -10315 24535 -10281
rect 24585 -10315 24607 -10281
rect 24653 -10315 24679 -10281
rect 24713 -10315 24822 -10281
rect 378 -10348 24822 -10315
rect -12322 -11211 24922 -11178
rect -12322 -11245 -12221 -11211
rect -12187 -11245 -12149 -11211
rect -12111 -11245 -12077 -11211
rect -12043 -11245 -12009 -11211
rect -11971 -11245 -11941 -11211
rect -11899 -11245 -11873 -11211
rect -11827 -11245 -11805 -11211
rect -11755 -11245 -11737 -11211
rect -11683 -11245 -11669 -11211
rect -11611 -11245 -11601 -11211
rect -11539 -11245 -11533 -11211
rect -11467 -11245 -11465 -11211
rect -11431 -11245 -11429 -11211
rect -11363 -11245 -11357 -11211
rect -11295 -11245 -11285 -11211
rect -11227 -11245 -11213 -11211
rect -11159 -11245 -11141 -11211
rect -11091 -11245 -11069 -11211
rect -11023 -11245 -10997 -11211
rect -10955 -11245 -10925 -11211
rect -10887 -11245 -10853 -11211
rect -10819 -11245 -10785 -11211
rect -10747 -11245 -10717 -11211
rect -10675 -11245 -10649 -11211
rect -10603 -11245 -10581 -11211
rect -10531 -11245 -10513 -11211
rect -10459 -11245 -10445 -11211
rect -10387 -11245 -10377 -11211
rect -10315 -11245 -10309 -11211
rect -10243 -11245 -10241 -11211
rect -10207 -11245 -10205 -11211
rect -10139 -11245 -10133 -11211
rect -10071 -11245 -10061 -11211
rect -10003 -11245 -9989 -11211
rect -9935 -11245 -9917 -11211
rect -9867 -11245 -9845 -11211
rect -9799 -11245 -9773 -11211
rect -9731 -11245 -9701 -11211
rect -9663 -11245 -9629 -11211
rect -9595 -11245 -9561 -11211
rect -9523 -11245 -9493 -11211
rect -9451 -11245 -9425 -11211
rect -9379 -11245 -9357 -11211
rect -9307 -11245 -9289 -11211
rect -9235 -11245 -9221 -11211
rect -9163 -11245 -9153 -11211
rect -9091 -11245 -9085 -11211
rect -9019 -11245 -9017 -11211
rect -8983 -11245 -8981 -11211
rect -8915 -11245 -8909 -11211
rect -8847 -11245 -8837 -11211
rect -8779 -11245 -8765 -11211
rect -8711 -11245 -8693 -11211
rect -8643 -11245 -8621 -11211
rect -8575 -11245 -8549 -11211
rect -8507 -11245 -8477 -11211
rect -8439 -11245 -8405 -11211
rect -8371 -11245 -8337 -11211
rect -8299 -11245 -8269 -11211
rect -8227 -11245 -8201 -11211
rect -8155 -11245 -8133 -11211
rect -8083 -11245 -8065 -11211
rect -8011 -11245 -7997 -11211
rect -7939 -11245 -7929 -11211
rect -7867 -11245 -7861 -11211
rect -7795 -11245 -7793 -11211
rect -7759 -11245 -7757 -11211
rect -7691 -11245 -7685 -11211
rect -7623 -11245 -7613 -11211
rect -7555 -11245 -7541 -11211
rect -7487 -11245 -7469 -11211
rect -7419 -11245 -7397 -11211
rect -7351 -11245 -7325 -11211
rect -7283 -11245 -7253 -11211
rect -7215 -11245 -7181 -11211
rect -7147 -11245 -7113 -11211
rect -7075 -11245 -7045 -11211
rect -7003 -11245 -6977 -11211
rect -6931 -11245 -6909 -11211
rect -6859 -11245 -6841 -11211
rect -6787 -11245 -6773 -11211
rect -6715 -11245 -6705 -11211
rect -6643 -11245 -6637 -11211
rect -6571 -11245 -6569 -11211
rect -6535 -11245 -6533 -11211
rect -6467 -11245 -6461 -11211
rect -6399 -11245 -6389 -11211
rect -6331 -11245 -6317 -11211
rect -6263 -11245 -6245 -11211
rect -6195 -11245 -6173 -11211
rect -6127 -11245 -6101 -11211
rect -6059 -11245 -6029 -11211
rect -5991 -11245 -5957 -11211
rect -5923 -11245 -5889 -11211
rect -5851 -11245 -5821 -11211
rect -5779 -11245 -5753 -11211
rect -5707 -11245 -5685 -11211
rect -5635 -11245 -5617 -11211
rect -5563 -11245 -5549 -11211
rect -5491 -11245 -5481 -11211
rect -5419 -11245 -5413 -11211
rect -5347 -11245 -5345 -11211
rect -5311 -11245 -5309 -11211
rect -5243 -11245 -5237 -11211
rect -5175 -11245 -5165 -11211
rect -5107 -11245 -5093 -11211
rect -5039 -11245 -5021 -11211
rect -4971 -11245 -4949 -11211
rect -4903 -11245 -4877 -11211
rect -4835 -11245 -4805 -11211
rect -4767 -11245 -4733 -11211
rect -4699 -11245 -4665 -11211
rect -4627 -11245 -4597 -11211
rect -4555 -11245 -4529 -11211
rect -4483 -11245 -4461 -11211
rect -4411 -11245 -4393 -11211
rect -4339 -11245 -4325 -11211
rect -4267 -11245 -4257 -11211
rect -4195 -11245 -4189 -11211
rect -4123 -11245 -4121 -11211
rect -4087 -11245 -4085 -11211
rect -4019 -11245 -4013 -11211
rect -3951 -11245 -3941 -11211
rect -3883 -11245 -3869 -11211
rect -3815 -11245 -3797 -11211
rect -3747 -11245 -3725 -11211
rect -3679 -11245 -3653 -11211
rect -3611 -11245 -3581 -11211
rect -3543 -11245 -3509 -11211
rect -3475 -11245 -3441 -11211
rect -3403 -11245 -3373 -11211
rect -3331 -11245 -3305 -11211
rect -3259 -11245 -3237 -11211
rect -3187 -11245 -3169 -11211
rect -3115 -11245 -3101 -11211
rect -3043 -11245 -3033 -11211
rect -2971 -11245 -2965 -11211
rect -2899 -11245 -2897 -11211
rect -2863 -11245 -2861 -11211
rect -2795 -11245 -2789 -11211
rect -2727 -11245 -2717 -11211
rect -2659 -11245 -2645 -11211
rect -2591 -11245 -2573 -11211
rect -2523 -11245 -2501 -11211
rect -2455 -11245 -2429 -11211
rect -2387 -11245 -2357 -11211
rect -2319 -11245 -2285 -11211
rect -2251 -11245 -2217 -11211
rect -2179 -11245 -2149 -11211
rect -2107 -11245 -2081 -11211
rect -2035 -11245 -2013 -11211
rect -1963 -11245 -1945 -11211
rect -1891 -11245 -1877 -11211
rect -1819 -11245 -1809 -11211
rect -1747 -11245 -1741 -11211
rect -1675 -11245 -1673 -11211
rect -1639 -11245 -1637 -11211
rect -1571 -11245 -1565 -11211
rect -1503 -11245 -1493 -11211
rect -1435 -11245 -1421 -11211
rect -1367 -11245 -1349 -11211
rect -1299 -11245 -1277 -11211
rect -1231 -11245 -1205 -11211
rect -1163 -11245 -1133 -11211
rect -1095 -11245 -1061 -11211
rect -1027 -11245 -993 -11211
rect -955 -11245 -925 -11211
rect -883 -11245 -857 -11211
rect -811 -11245 -789 -11211
rect -739 -11245 -721 -11211
rect -667 -11245 -653 -11211
rect -595 -11245 -585 -11211
rect -523 -11245 -517 -11211
rect -451 -11245 -449 -11211
rect -415 -11245 -413 -11211
rect -347 -11245 -341 -11211
rect -279 -11245 -269 -11211
rect -211 -11245 -197 -11211
rect -143 -11245 -125 -11211
rect -75 -11245 -53 -11211
rect -7 -11245 19 -11211
rect 61 -11245 91 -11211
rect 129 -11245 163 -11211
rect 197 -11245 231 -11211
rect 269 -11245 299 -11211
rect 341 -11245 367 -11211
rect 413 -11245 435 -11211
rect 485 -11245 503 -11211
rect 557 -11245 571 -11211
rect 629 -11245 639 -11211
rect 701 -11245 707 -11211
rect 773 -11245 775 -11211
rect 809 -11245 811 -11211
rect 877 -11245 883 -11211
rect 945 -11245 955 -11211
rect 1013 -11245 1027 -11211
rect 1081 -11245 1099 -11211
rect 1149 -11245 1171 -11211
rect 1217 -11245 1243 -11211
rect 1285 -11245 1315 -11211
rect 1353 -11245 1387 -11211
rect 1421 -11245 1455 -11211
rect 1493 -11245 1523 -11211
rect 1565 -11245 1591 -11211
rect 1637 -11245 1659 -11211
rect 1709 -11245 1727 -11211
rect 1781 -11245 1795 -11211
rect 1853 -11245 1863 -11211
rect 1925 -11245 1931 -11211
rect 1997 -11245 1999 -11211
rect 2033 -11245 2035 -11211
rect 2101 -11245 2107 -11211
rect 2169 -11245 2179 -11211
rect 2237 -11245 2251 -11211
rect 2305 -11245 2323 -11211
rect 2373 -11245 2395 -11211
rect 2441 -11245 2467 -11211
rect 2509 -11245 2539 -11211
rect 2577 -11245 2611 -11211
rect 2645 -11245 2679 -11211
rect 2717 -11245 2747 -11211
rect 2789 -11245 2815 -11211
rect 2861 -11245 2883 -11211
rect 2933 -11245 2951 -11211
rect 3005 -11245 3019 -11211
rect 3077 -11245 3087 -11211
rect 3149 -11245 3155 -11211
rect 3221 -11245 3223 -11211
rect 3257 -11245 3259 -11211
rect 3325 -11245 3331 -11211
rect 3393 -11245 3403 -11211
rect 3461 -11245 3475 -11211
rect 3529 -11245 3547 -11211
rect 3597 -11245 3619 -11211
rect 3665 -11245 3691 -11211
rect 3733 -11245 3763 -11211
rect 3801 -11245 3835 -11211
rect 3869 -11245 3903 -11211
rect 3941 -11245 3971 -11211
rect 4013 -11245 4039 -11211
rect 4085 -11245 4107 -11211
rect 4157 -11245 4175 -11211
rect 4229 -11245 4243 -11211
rect 4301 -11245 4311 -11211
rect 4373 -11245 4379 -11211
rect 4445 -11245 4447 -11211
rect 4481 -11245 4483 -11211
rect 4549 -11245 4555 -11211
rect 4617 -11245 4627 -11211
rect 4685 -11245 4699 -11211
rect 4753 -11245 4771 -11211
rect 4821 -11245 4843 -11211
rect 4889 -11245 4915 -11211
rect 4957 -11245 4987 -11211
rect 5025 -11245 5059 -11211
rect 5093 -11245 5127 -11211
rect 5165 -11245 5195 -11211
rect 5237 -11245 5263 -11211
rect 5309 -11245 5331 -11211
rect 5381 -11245 5399 -11211
rect 5453 -11245 5467 -11211
rect 5525 -11245 5535 -11211
rect 5597 -11245 5603 -11211
rect 5669 -11245 5671 -11211
rect 5705 -11245 5707 -11211
rect 5773 -11245 5779 -11211
rect 5841 -11245 5851 -11211
rect 5909 -11245 5923 -11211
rect 5977 -11245 5995 -11211
rect 6045 -11245 6067 -11211
rect 6113 -11245 6139 -11211
rect 6181 -11245 6211 -11211
rect 6249 -11245 6283 -11211
rect 6317 -11245 6351 -11211
rect 6389 -11245 6419 -11211
rect 6461 -11245 6487 -11211
rect 6533 -11245 6555 -11211
rect 6605 -11245 6623 -11211
rect 6677 -11245 6691 -11211
rect 6749 -11245 6759 -11211
rect 6821 -11245 6827 -11211
rect 6893 -11245 6895 -11211
rect 6929 -11245 6931 -11211
rect 6997 -11245 7003 -11211
rect 7065 -11245 7075 -11211
rect 7133 -11245 7147 -11211
rect 7201 -11245 7219 -11211
rect 7269 -11245 7291 -11211
rect 7337 -11245 7363 -11211
rect 7405 -11245 7435 -11211
rect 7473 -11245 7507 -11211
rect 7541 -11245 7575 -11211
rect 7613 -11245 7643 -11211
rect 7685 -11245 7711 -11211
rect 7757 -11245 7779 -11211
rect 7829 -11245 7847 -11211
rect 7901 -11245 7915 -11211
rect 7973 -11245 7983 -11211
rect 8045 -11245 8051 -11211
rect 8117 -11245 8119 -11211
rect 8153 -11245 8155 -11211
rect 8221 -11245 8227 -11211
rect 8289 -11245 8299 -11211
rect 8357 -11245 8371 -11211
rect 8425 -11245 8443 -11211
rect 8493 -11245 8515 -11211
rect 8561 -11245 8587 -11211
rect 8629 -11245 8659 -11211
rect 8697 -11245 8731 -11211
rect 8765 -11245 8799 -11211
rect 8837 -11245 8867 -11211
rect 8909 -11245 8935 -11211
rect 8981 -11245 9003 -11211
rect 9053 -11245 9071 -11211
rect 9125 -11245 9139 -11211
rect 9197 -11245 9207 -11211
rect 9269 -11245 9275 -11211
rect 9341 -11245 9343 -11211
rect 9377 -11245 9379 -11211
rect 9445 -11245 9451 -11211
rect 9513 -11245 9523 -11211
rect 9581 -11245 9595 -11211
rect 9649 -11245 9667 -11211
rect 9717 -11245 9739 -11211
rect 9785 -11245 9811 -11211
rect 9853 -11245 9883 -11211
rect 9921 -11245 9955 -11211
rect 9989 -11245 10023 -11211
rect 10061 -11245 10091 -11211
rect 10133 -11245 10159 -11211
rect 10205 -11245 10227 -11211
rect 10277 -11245 10295 -11211
rect 10349 -11245 10363 -11211
rect 10421 -11245 10431 -11211
rect 10493 -11245 10499 -11211
rect 10565 -11245 10567 -11211
rect 10601 -11245 10603 -11211
rect 10669 -11245 10675 -11211
rect 10737 -11245 10747 -11211
rect 10805 -11245 10819 -11211
rect 10873 -11245 10891 -11211
rect 10941 -11245 10963 -11211
rect 11009 -11245 11035 -11211
rect 11077 -11245 11107 -11211
rect 11145 -11245 11179 -11211
rect 11213 -11245 11247 -11211
rect 11285 -11245 11315 -11211
rect 11357 -11245 11383 -11211
rect 11429 -11245 11451 -11211
rect 11501 -11245 11519 -11211
rect 11573 -11245 11587 -11211
rect 11645 -11245 11655 -11211
rect 11717 -11245 11723 -11211
rect 11789 -11245 11791 -11211
rect 11825 -11245 11827 -11211
rect 11893 -11245 11899 -11211
rect 11961 -11245 11971 -11211
rect 12029 -11245 12043 -11211
rect 12097 -11245 12115 -11211
rect 12165 -11245 12187 -11211
rect 12233 -11245 12259 -11211
rect 12301 -11245 12331 -11211
rect 12369 -11245 12403 -11211
rect 12437 -11245 12471 -11211
rect 12509 -11245 12539 -11211
rect 12581 -11245 12607 -11211
rect 12653 -11245 12675 -11211
rect 12725 -11245 12743 -11211
rect 12797 -11245 12811 -11211
rect 12869 -11245 12879 -11211
rect 12941 -11245 12947 -11211
rect 13013 -11245 13015 -11211
rect 13049 -11245 13051 -11211
rect 13117 -11245 13123 -11211
rect 13185 -11245 13195 -11211
rect 13253 -11245 13267 -11211
rect 13321 -11245 13339 -11211
rect 13389 -11245 13411 -11211
rect 13457 -11245 13483 -11211
rect 13525 -11245 13555 -11211
rect 13593 -11245 13627 -11211
rect 13661 -11245 13695 -11211
rect 13733 -11245 13763 -11211
rect 13805 -11245 13831 -11211
rect 13877 -11245 13899 -11211
rect 13949 -11245 13967 -11211
rect 14021 -11245 14035 -11211
rect 14093 -11245 14103 -11211
rect 14165 -11245 14171 -11211
rect 14237 -11245 14239 -11211
rect 14273 -11245 14275 -11211
rect 14341 -11245 14347 -11211
rect 14409 -11245 14419 -11211
rect 14477 -11245 14491 -11211
rect 14545 -11245 14563 -11211
rect 14613 -11245 14635 -11211
rect 14681 -11245 14707 -11211
rect 14749 -11245 14779 -11211
rect 14817 -11245 14851 -11211
rect 14885 -11245 14919 -11211
rect 14957 -11245 14987 -11211
rect 15029 -11245 15055 -11211
rect 15101 -11245 15123 -11211
rect 15173 -11245 15191 -11211
rect 15245 -11245 15259 -11211
rect 15317 -11245 15327 -11211
rect 15389 -11245 15395 -11211
rect 15461 -11245 15463 -11211
rect 15497 -11245 15499 -11211
rect 15565 -11245 15571 -11211
rect 15633 -11245 15643 -11211
rect 15701 -11245 15715 -11211
rect 15769 -11245 15787 -11211
rect 15837 -11245 15859 -11211
rect 15905 -11245 15931 -11211
rect 15973 -11245 16003 -11211
rect 16041 -11245 16075 -11211
rect 16109 -11245 16143 -11211
rect 16181 -11245 16211 -11211
rect 16253 -11245 16279 -11211
rect 16325 -11245 16347 -11211
rect 16397 -11245 16415 -11211
rect 16469 -11245 16483 -11211
rect 16541 -11245 16551 -11211
rect 16613 -11245 16619 -11211
rect 16685 -11245 16687 -11211
rect 16721 -11245 16723 -11211
rect 16789 -11245 16795 -11211
rect 16857 -11245 16867 -11211
rect 16925 -11245 16939 -11211
rect 16993 -11245 17011 -11211
rect 17061 -11245 17083 -11211
rect 17129 -11245 17155 -11211
rect 17197 -11245 17227 -11211
rect 17265 -11245 17299 -11211
rect 17333 -11245 17367 -11211
rect 17405 -11245 17435 -11211
rect 17477 -11245 17503 -11211
rect 17549 -11245 17571 -11211
rect 17621 -11245 17639 -11211
rect 17693 -11245 17707 -11211
rect 17765 -11245 17775 -11211
rect 17837 -11245 17843 -11211
rect 17909 -11245 17911 -11211
rect 17945 -11245 17947 -11211
rect 18013 -11245 18019 -11211
rect 18081 -11245 18091 -11211
rect 18149 -11245 18163 -11211
rect 18217 -11245 18235 -11211
rect 18285 -11245 18307 -11211
rect 18353 -11245 18379 -11211
rect 18421 -11245 18451 -11211
rect 18489 -11245 18523 -11211
rect 18557 -11245 18591 -11211
rect 18629 -11245 18659 -11211
rect 18701 -11245 18727 -11211
rect 18773 -11245 18795 -11211
rect 18845 -11245 18863 -11211
rect 18917 -11245 18931 -11211
rect 18989 -11245 18999 -11211
rect 19061 -11245 19067 -11211
rect 19133 -11245 19135 -11211
rect 19169 -11245 19171 -11211
rect 19237 -11245 19243 -11211
rect 19305 -11245 19315 -11211
rect 19373 -11245 19387 -11211
rect 19441 -11245 19459 -11211
rect 19509 -11245 19531 -11211
rect 19577 -11245 19603 -11211
rect 19645 -11245 19675 -11211
rect 19713 -11245 19747 -11211
rect 19781 -11245 19815 -11211
rect 19853 -11245 19883 -11211
rect 19925 -11245 19951 -11211
rect 19997 -11245 20019 -11211
rect 20069 -11245 20087 -11211
rect 20141 -11245 20155 -11211
rect 20213 -11245 20223 -11211
rect 20285 -11245 20291 -11211
rect 20357 -11245 20359 -11211
rect 20393 -11245 20395 -11211
rect 20461 -11245 20467 -11211
rect 20529 -11245 20539 -11211
rect 20597 -11245 20611 -11211
rect 20665 -11245 20683 -11211
rect 20733 -11245 20755 -11211
rect 20801 -11245 20827 -11211
rect 20869 -11245 20899 -11211
rect 20937 -11245 20971 -11211
rect 21005 -11245 21039 -11211
rect 21077 -11245 21107 -11211
rect 21149 -11245 21175 -11211
rect 21221 -11245 21243 -11211
rect 21293 -11245 21311 -11211
rect 21365 -11245 21379 -11211
rect 21437 -11245 21447 -11211
rect 21509 -11245 21515 -11211
rect 21581 -11245 21583 -11211
rect 21617 -11245 21619 -11211
rect 21685 -11245 21691 -11211
rect 21753 -11245 21763 -11211
rect 21821 -11245 21835 -11211
rect 21889 -11245 21907 -11211
rect 21957 -11245 21979 -11211
rect 22025 -11245 22051 -11211
rect 22093 -11245 22123 -11211
rect 22161 -11245 22195 -11211
rect 22229 -11245 22263 -11211
rect 22301 -11245 22331 -11211
rect 22373 -11245 22399 -11211
rect 22445 -11245 22467 -11211
rect 22517 -11245 22535 -11211
rect 22589 -11245 22603 -11211
rect 22661 -11245 22671 -11211
rect 22733 -11245 22739 -11211
rect 22805 -11245 22807 -11211
rect 22841 -11245 22843 -11211
rect 22909 -11245 22915 -11211
rect 22977 -11245 22987 -11211
rect 23045 -11245 23059 -11211
rect 23113 -11245 23131 -11211
rect 23181 -11245 23203 -11211
rect 23249 -11245 23275 -11211
rect 23317 -11245 23347 -11211
rect 23385 -11245 23419 -11211
rect 23453 -11245 23487 -11211
rect 23525 -11245 23555 -11211
rect 23597 -11245 23623 -11211
rect 23669 -11245 23691 -11211
rect 23741 -11245 23759 -11211
rect 23813 -11245 23827 -11211
rect 23885 -11245 23895 -11211
rect 23957 -11245 23963 -11211
rect 24029 -11245 24031 -11211
rect 24065 -11245 24067 -11211
rect 24133 -11245 24139 -11211
rect 24201 -11245 24211 -11211
rect 24269 -11245 24283 -11211
rect 24337 -11245 24355 -11211
rect 24405 -11245 24427 -11211
rect 24473 -11245 24499 -11211
rect 24541 -11245 24571 -11211
rect 24609 -11245 24643 -11211
rect 24677 -11245 24711 -11211
rect 24749 -11245 24787 -11211
rect 24821 -11245 24922 -11211
rect -12322 -11278 24922 -11245
rect -12322 -11363 -12222 -11278
rect -12322 -11397 -12289 -11363
rect -12255 -11397 -12222 -11363
rect -12322 -11431 -12222 -11397
rect -12322 -11465 -12289 -11431
rect -12255 -11465 -12222 -11431
rect -12322 -11499 -12222 -11465
rect -12322 -11533 -12289 -11499
rect -12255 -11533 -12222 -11499
rect -12322 -11567 -12222 -11533
rect -12322 -11601 -12289 -11567
rect -12255 -11601 -12222 -11567
rect -12322 -11635 -12222 -11601
rect -12322 -11669 -12289 -11635
rect -12255 -11669 -12222 -11635
rect -12322 -11703 -12222 -11669
rect -12322 -11737 -12289 -11703
rect -12255 -11737 -12222 -11703
rect -12322 -11771 -12222 -11737
rect -12322 -11805 -12289 -11771
rect -12255 -11805 -12222 -11771
rect -12322 -11839 -12222 -11805
rect -12322 -11873 -12289 -11839
rect -12255 -11873 -12222 -11839
rect -12322 -11907 -12222 -11873
rect -12322 -11941 -12289 -11907
rect -12255 -11941 -12222 -11907
rect -12322 -11975 -12222 -11941
rect -12322 -12009 -12289 -11975
rect -12255 -12009 -12222 -11975
rect -12322 -12043 -12222 -12009
rect -12322 -12077 -12289 -12043
rect -12255 -12077 -12222 -12043
rect -12322 -12091 -12222 -12077
rect -12322 -12145 -12289 -12091
rect -12255 -12145 -12222 -12091
rect -12322 -12163 -12222 -12145
rect -12322 -12213 -12289 -12163
rect -12255 -12213 -12222 -12163
rect -12322 -12235 -12222 -12213
rect -12322 -12281 -12289 -12235
rect -12255 -12281 -12222 -12235
rect -12322 -12307 -12222 -12281
rect -12322 -12349 -12289 -12307
rect -12255 -12349 -12222 -12307
rect -12322 -12379 -12222 -12349
rect -12322 -12417 -12289 -12379
rect -12255 -12417 -12222 -12379
rect -12322 -12451 -12222 -12417
rect 24822 -11363 24922 -11278
rect 24822 -11397 24855 -11363
rect 24889 -11397 24922 -11363
rect 24822 -11431 24922 -11397
rect 24822 -11465 24855 -11431
rect 24889 -11465 24922 -11431
rect 24822 -11499 24922 -11465
rect 24822 -11533 24855 -11499
rect 24889 -11533 24922 -11499
rect 24822 -11567 24922 -11533
rect 24822 -11601 24855 -11567
rect 24889 -11601 24922 -11567
rect 24822 -11635 24922 -11601
rect 24822 -11669 24855 -11635
rect 24889 -11669 24922 -11635
rect 24822 -11703 24922 -11669
rect 24822 -11737 24855 -11703
rect 24889 -11737 24922 -11703
rect 24822 -11771 24922 -11737
rect 24822 -11805 24855 -11771
rect 24889 -11805 24922 -11771
rect 24822 -11839 24922 -11805
rect 24822 -11873 24855 -11839
rect 24889 -11873 24922 -11839
rect 24822 -11907 24922 -11873
rect 24822 -11941 24855 -11907
rect 24889 -11941 24922 -11907
rect 24822 -11975 24922 -11941
rect 24822 -12009 24855 -11975
rect 24889 -12009 24922 -11975
rect 24822 -12043 24922 -12009
rect 24822 -12077 24855 -12043
rect 24889 -12077 24922 -12043
rect 24822 -12091 24922 -12077
rect 24822 -12145 24855 -12091
rect 24889 -12145 24922 -12091
rect 24822 -12163 24922 -12145
rect 24822 -12213 24855 -12163
rect 24889 -12213 24922 -12163
rect 24822 -12235 24922 -12213
rect 24822 -12281 24855 -12235
rect 24889 -12281 24922 -12235
rect 24822 -12307 24922 -12281
rect 24822 -12349 24855 -12307
rect 24889 -12349 24922 -12307
rect 24822 -12379 24922 -12349
rect 24822 -12417 24855 -12379
rect 24889 -12417 24922 -12379
rect -12322 -12485 -12289 -12451
rect -12255 -12485 -12222 -12451
rect -8952 -12474 -8913 -12440
rect -8879 -12474 -8855 -12440
rect -8811 -12474 -8783 -12440
rect -8743 -12474 -8711 -12440
rect -8675 -12474 -8641 -12440
rect -8605 -12474 -8573 -12440
rect -8533 -12474 -8505 -12440
rect -8461 -12474 -8437 -12440
rect -8403 -12474 -8364 -12440
rect -7934 -12474 -7895 -12440
rect -7861 -12474 -7837 -12440
rect -7793 -12474 -7765 -12440
rect -7725 -12474 -7693 -12440
rect -7657 -12474 -7623 -12440
rect -7587 -12474 -7555 -12440
rect -7515 -12474 -7487 -12440
rect -7443 -12474 -7419 -12440
rect -7385 -12474 -7346 -12440
rect -6916 -12474 -6877 -12440
rect -6843 -12474 -6819 -12440
rect -6775 -12474 -6747 -12440
rect -6707 -12474 -6675 -12440
rect -6639 -12474 -6605 -12440
rect -6569 -12474 -6537 -12440
rect -6497 -12474 -6469 -12440
rect -6425 -12474 -6401 -12440
rect -6367 -12474 -6328 -12440
rect -5898 -12474 -5859 -12440
rect -5825 -12474 -5801 -12440
rect -5757 -12474 -5729 -12440
rect -5689 -12474 -5657 -12440
rect -5621 -12474 -5587 -12440
rect -5551 -12474 -5519 -12440
rect -5479 -12474 -5451 -12440
rect -5407 -12474 -5383 -12440
rect -5349 -12474 -5310 -12440
rect -4880 -12474 -4841 -12440
rect -4807 -12474 -4783 -12440
rect -4739 -12474 -4711 -12440
rect -4671 -12474 -4639 -12440
rect -4603 -12474 -4569 -12440
rect -4533 -12474 -4501 -12440
rect -4461 -12474 -4433 -12440
rect -4389 -12474 -4365 -12440
rect -4331 -12474 -4292 -12440
rect -3862 -12474 -3823 -12440
rect -3789 -12474 -3765 -12440
rect -3721 -12474 -3693 -12440
rect -3653 -12474 -3621 -12440
rect -3585 -12474 -3551 -12440
rect -3515 -12474 -3483 -12440
rect -3443 -12474 -3415 -12440
rect -3371 -12474 -3347 -12440
rect -3313 -12474 -3274 -12440
rect -2844 -12474 -2805 -12440
rect -2771 -12474 -2747 -12440
rect -2703 -12474 -2675 -12440
rect -2635 -12474 -2603 -12440
rect -2567 -12474 -2533 -12440
rect -2497 -12474 -2465 -12440
rect -2425 -12474 -2397 -12440
rect -2353 -12474 -2329 -12440
rect -2295 -12474 -2256 -12440
rect -1826 -12474 -1787 -12440
rect -1753 -12474 -1729 -12440
rect -1685 -12474 -1657 -12440
rect -1617 -12474 -1585 -12440
rect -1549 -12474 -1515 -12440
rect -1479 -12474 -1447 -12440
rect -1407 -12474 -1379 -12440
rect -1335 -12474 -1311 -12440
rect -1277 -12474 -1238 -12440
rect -808 -12474 -769 -12440
rect -735 -12474 -711 -12440
rect -667 -12474 -639 -12440
rect -599 -12474 -567 -12440
rect -531 -12474 -497 -12440
rect -461 -12474 -429 -12440
rect -389 -12474 -361 -12440
rect -317 -12474 -293 -12440
rect -259 -12474 -220 -12440
rect 24822 -12451 24922 -12417
rect -12322 -12519 -12222 -12485
rect 24822 -12485 24855 -12451
rect 24889 -12485 24922 -12451
rect -12322 -12557 -12289 -12519
rect -12255 -12557 -12222 -12519
rect -12322 -12587 -12222 -12557
rect -12322 -12629 -12289 -12587
rect -12255 -12629 -12222 -12587
rect -12322 -12655 -12222 -12629
rect -12322 -12701 -12289 -12655
rect -12255 -12701 -12222 -12655
rect -12322 -12723 -12222 -12701
rect -12322 -12773 -12289 -12723
rect -12255 -12773 -12222 -12723
rect -12322 -12791 -12222 -12773
rect -12322 -12845 -12289 -12791
rect -12255 -12845 -12222 -12791
rect -12322 -12859 -12222 -12845
rect -12322 -12917 -12289 -12859
rect -12255 -12917 -12222 -12859
rect -12322 -12927 -12222 -12917
rect -12322 -12989 -12289 -12927
rect -12255 -12989 -12222 -12927
rect -12322 -12995 -12222 -12989
rect -12322 -13061 -12289 -12995
rect -12255 -13061 -12222 -12995
rect -12322 -13063 -12222 -13061
rect -12322 -13097 -12289 -13063
rect -12255 -13097 -12222 -13063
rect -12322 -13099 -12222 -13097
rect -12322 -13165 -12289 -13099
rect -12255 -13165 -12222 -13099
rect -9184 -12543 -9150 -12508
rect -9184 -12615 -9150 -12591
rect -9184 -12687 -9150 -12659
rect -9184 -12759 -9150 -12727
rect -9184 -12829 -9150 -12795
rect -9184 -12897 -9150 -12865
rect -9184 -12965 -9150 -12937
rect -9184 -13033 -9150 -13009
rect -9184 -13116 -9150 -13081
rect -8166 -12543 -8132 -12508
rect -8166 -12615 -8132 -12591
rect -8166 -12687 -8132 -12659
rect -8166 -12759 -8132 -12727
rect -8166 -12829 -8132 -12795
rect -8166 -12897 -8132 -12865
rect -8166 -12965 -8132 -12937
rect -8166 -13033 -8132 -13009
rect -8166 -13116 -8132 -13081
rect -7148 -12543 -7114 -12508
rect -7148 -12615 -7114 -12591
rect -7148 -12687 -7114 -12659
rect -7148 -12759 -7114 -12727
rect -7148 -12829 -7114 -12795
rect -7148 -12897 -7114 -12865
rect -7148 -12965 -7114 -12937
rect -7148 -13033 -7114 -13009
rect -7148 -13116 -7114 -13081
rect -6130 -12543 -6096 -12508
rect -6130 -12615 -6096 -12591
rect -6130 -12687 -6096 -12659
rect -6130 -12759 -6096 -12727
rect -6130 -12829 -6096 -12795
rect -6130 -12897 -6096 -12865
rect -6130 -12965 -6096 -12937
rect -6130 -13033 -6096 -13009
rect -6130 -13116 -6096 -13081
rect -5112 -12543 -5078 -12508
rect -5112 -12615 -5078 -12591
rect -5112 -12687 -5078 -12659
rect -5112 -12759 -5078 -12727
rect -5112 -12829 -5078 -12795
rect -5112 -12897 -5078 -12865
rect -5112 -12965 -5078 -12937
rect -5112 -13033 -5078 -13009
rect -5112 -13116 -5078 -13081
rect -4094 -12543 -4060 -12508
rect -4094 -12615 -4060 -12591
rect -4094 -12687 -4060 -12659
rect -4094 -12759 -4060 -12727
rect -4094 -12829 -4060 -12795
rect -4094 -12897 -4060 -12865
rect -4094 -12965 -4060 -12937
rect -4094 -13033 -4060 -13009
rect -4094 -13116 -4060 -13081
rect -3076 -12543 -3042 -12508
rect -3076 -12615 -3042 -12591
rect -3076 -12687 -3042 -12659
rect -3076 -12759 -3042 -12727
rect -3076 -12829 -3042 -12795
rect -3076 -12897 -3042 -12865
rect -3076 -12965 -3042 -12937
rect -3076 -13033 -3042 -13009
rect -3076 -13116 -3042 -13081
rect -2058 -12543 -2024 -12508
rect -2058 -12615 -2024 -12591
rect -2058 -12687 -2024 -12659
rect -2058 -12759 -2024 -12727
rect -2058 -12829 -2024 -12795
rect -2058 -12897 -2024 -12865
rect -2058 -12965 -2024 -12937
rect -2058 -13033 -2024 -13009
rect -2058 -13116 -2024 -13081
rect -1040 -12543 -1006 -12508
rect -1040 -12615 -1006 -12591
rect -1040 -12687 -1006 -12659
rect -1040 -12759 -1006 -12727
rect -1040 -12829 -1006 -12795
rect -1040 -12897 -1006 -12865
rect -1040 -12965 -1006 -12937
rect -1040 -13033 -1006 -13009
rect -1040 -13116 -1006 -13081
rect -22 -12543 12 -12508
rect -22 -12615 12 -12591
rect -22 -12687 12 -12659
rect -22 -12759 12 -12727
rect -22 -12829 12 -12795
rect -22 -12897 12 -12865
rect -22 -12965 12 -12937
rect -22 -13033 12 -13009
rect -22 -13116 12 -13081
rect 24822 -12519 24922 -12485
rect 24822 -12557 24855 -12519
rect 24889 -12557 24922 -12519
rect 24822 -12587 24922 -12557
rect 24822 -12629 24855 -12587
rect 24889 -12629 24922 -12587
rect 24822 -12655 24922 -12629
rect 24822 -12701 24855 -12655
rect 24889 -12701 24922 -12655
rect 24822 -12723 24922 -12701
rect 24822 -12773 24855 -12723
rect 24889 -12773 24922 -12723
rect 24822 -12791 24922 -12773
rect 24822 -12845 24855 -12791
rect 24889 -12845 24922 -12791
rect 24822 -12859 24922 -12845
rect 24822 -12917 24855 -12859
rect 24889 -12917 24922 -12859
rect 24822 -12927 24922 -12917
rect 24822 -12989 24855 -12927
rect 24889 -12989 24922 -12927
rect 24822 -12995 24922 -12989
rect 24822 -13061 24855 -12995
rect 24889 -13061 24922 -12995
rect 24822 -13063 24922 -13061
rect 24822 -13097 24855 -13063
rect 24889 -13097 24922 -13063
rect 24822 -13099 24922 -13097
rect -12322 -13171 -12222 -13165
rect -12322 -13233 -12289 -13171
rect -12255 -13233 -12222 -13171
rect -8952 -13184 -8913 -13150
rect -8879 -13184 -8855 -13150
rect -8811 -13184 -8783 -13150
rect -8743 -13184 -8711 -13150
rect -8675 -13184 -8641 -13150
rect -8605 -13184 -8573 -13150
rect -8533 -13184 -8505 -13150
rect -8461 -13184 -8437 -13150
rect -8403 -13184 -8364 -13150
rect -7934 -13184 -7895 -13150
rect -7861 -13184 -7837 -13150
rect -7793 -13184 -7765 -13150
rect -7725 -13184 -7693 -13150
rect -7657 -13184 -7623 -13150
rect -7587 -13184 -7555 -13150
rect -7515 -13184 -7487 -13150
rect -7443 -13184 -7419 -13150
rect -7385 -13184 -7346 -13150
rect -6916 -13184 -6877 -13150
rect -6843 -13184 -6819 -13150
rect -6775 -13184 -6747 -13150
rect -6707 -13184 -6675 -13150
rect -6639 -13184 -6605 -13150
rect -6569 -13184 -6537 -13150
rect -6497 -13184 -6469 -13150
rect -6425 -13184 -6401 -13150
rect -6367 -13184 -6328 -13150
rect -5898 -13184 -5859 -13150
rect -5825 -13184 -5801 -13150
rect -5757 -13184 -5729 -13150
rect -5689 -13184 -5657 -13150
rect -5621 -13184 -5587 -13150
rect -5551 -13184 -5519 -13150
rect -5479 -13184 -5451 -13150
rect -5407 -13184 -5383 -13150
rect -5349 -13184 -5310 -13150
rect -4880 -13184 -4841 -13150
rect -4807 -13184 -4783 -13150
rect -4739 -13184 -4711 -13150
rect -4671 -13184 -4639 -13150
rect -4603 -13184 -4569 -13150
rect -4533 -13184 -4501 -13150
rect -4461 -13184 -4433 -13150
rect -4389 -13184 -4365 -13150
rect -4331 -13184 -4292 -13150
rect -3862 -13184 -3823 -13150
rect -3789 -13184 -3765 -13150
rect -3721 -13184 -3693 -13150
rect -3653 -13184 -3621 -13150
rect -3585 -13184 -3551 -13150
rect -3515 -13184 -3483 -13150
rect -3443 -13184 -3415 -13150
rect -3371 -13184 -3347 -13150
rect -3313 -13184 -3274 -13150
rect -2844 -13184 -2805 -13150
rect -2771 -13184 -2747 -13150
rect -2703 -13184 -2675 -13150
rect -2635 -13184 -2603 -13150
rect -2567 -13184 -2533 -13150
rect -2497 -13184 -2465 -13150
rect -2425 -13184 -2397 -13150
rect -2353 -13184 -2329 -13150
rect -2295 -13184 -2256 -13150
rect -1826 -13184 -1787 -13150
rect -1753 -13184 -1729 -13150
rect -1685 -13184 -1657 -13150
rect -1617 -13184 -1585 -13150
rect -1549 -13184 -1515 -13150
rect -1479 -13184 -1447 -13150
rect -1407 -13184 -1379 -13150
rect -1335 -13184 -1311 -13150
rect -1277 -13184 -1238 -13150
rect -808 -13184 -769 -13150
rect -735 -13184 -711 -13150
rect -667 -13184 -639 -13150
rect -599 -13184 -567 -13150
rect -531 -13184 -497 -13150
rect -461 -13184 -429 -13150
rect -389 -13184 -361 -13150
rect -317 -13184 -293 -13150
rect -259 -13184 -220 -13150
rect 24822 -13165 24855 -13099
rect 24889 -13165 24922 -13099
rect 24822 -13171 24922 -13165
rect -12322 -13243 -12222 -13233
rect -12322 -13301 -12289 -13243
rect -12255 -13301 -12222 -13243
rect 24822 -13233 24855 -13171
rect 24889 -13233 24922 -13171
rect 24822 -13243 24922 -13233
rect -8952 -13292 -8913 -13258
rect -8879 -13292 -8855 -13258
rect -8811 -13292 -8783 -13258
rect -8743 -13292 -8711 -13258
rect -8675 -13292 -8641 -13258
rect -8605 -13292 -8573 -13258
rect -8533 -13292 -8505 -13258
rect -8461 -13292 -8437 -13258
rect -8403 -13292 -8364 -13258
rect -7934 -13292 -7895 -13258
rect -7861 -13292 -7837 -13258
rect -7793 -13292 -7765 -13258
rect -7725 -13292 -7693 -13258
rect -7657 -13292 -7623 -13258
rect -7587 -13292 -7555 -13258
rect -7515 -13292 -7487 -13258
rect -7443 -13292 -7419 -13258
rect -7385 -13292 -7346 -13258
rect -6916 -13292 -6877 -13258
rect -6843 -13292 -6819 -13258
rect -6775 -13292 -6747 -13258
rect -6707 -13292 -6675 -13258
rect -6639 -13292 -6605 -13258
rect -6569 -13292 -6537 -13258
rect -6497 -13292 -6469 -13258
rect -6425 -13292 -6401 -13258
rect -6367 -13292 -6328 -13258
rect -5898 -13292 -5859 -13258
rect -5825 -13292 -5801 -13258
rect -5757 -13292 -5729 -13258
rect -5689 -13292 -5657 -13258
rect -5621 -13292 -5587 -13258
rect -5551 -13292 -5519 -13258
rect -5479 -13292 -5451 -13258
rect -5407 -13292 -5383 -13258
rect -5349 -13292 -5310 -13258
rect -4880 -13292 -4841 -13258
rect -4807 -13292 -4783 -13258
rect -4739 -13292 -4711 -13258
rect -4671 -13292 -4639 -13258
rect -4603 -13292 -4569 -13258
rect -4533 -13292 -4501 -13258
rect -4461 -13292 -4433 -13258
rect -4389 -13292 -4365 -13258
rect -4331 -13292 -4292 -13258
rect -3862 -13292 -3823 -13258
rect -3789 -13292 -3765 -13258
rect -3721 -13292 -3693 -13258
rect -3653 -13292 -3621 -13258
rect -3585 -13292 -3551 -13258
rect -3515 -13292 -3483 -13258
rect -3443 -13292 -3415 -13258
rect -3371 -13292 -3347 -13258
rect -3313 -13292 -3274 -13258
rect -2844 -13292 -2805 -13258
rect -2771 -13292 -2747 -13258
rect -2703 -13292 -2675 -13258
rect -2635 -13292 -2603 -13258
rect -2567 -13292 -2533 -13258
rect -2497 -13292 -2465 -13258
rect -2425 -13292 -2397 -13258
rect -2353 -13292 -2329 -13258
rect -2295 -13292 -2256 -13258
rect -1826 -13292 -1787 -13258
rect -1753 -13292 -1729 -13258
rect -1685 -13292 -1657 -13258
rect -1617 -13292 -1585 -13258
rect -1549 -13292 -1515 -13258
rect -1479 -13292 -1447 -13258
rect -1407 -13292 -1379 -13258
rect -1335 -13292 -1311 -13258
rect -1277 -13292 -1238 -13258
rect -808 -13292 -769 -13258
rect -735 -13292 -711 -13258
rect -667 -13292 -639 -13258
rect -599 -13292 -567 -13258
rect -531 -13292 -497 -13258
rect -461 -13292 -429 -13258
rect -389 -13292 -361 -13258
rect -317 -13292 -293 -13258
rect -259 -13292 -220 -13258
rect -3592 -13294 -3532 -13292
rect -12322 -13315 -12222 -13301
rect -12322 -13369 -12289 -13315
rect -12255 -13369 -12222 -13315
rect 24822 -13301 24855 -13243
rect 24889 -13301 24922 -13243
rect 24822 -13315 24922 -13301
rect -12322 -13387 -12222 -13369
rect -12322 -13437 -12289 -13387
rect -12255 -13437 -12222 -13387
rect -12322 -13459 -12222 -13437
rect -12322 -13505 -12289 -13459
rect -12255 -13505 -12222 -13459
rect -12322 -13531 -12222 -13505
rect -12322 -13573 -12289 -13531
rect -12255 -13573 -12222 -13531
rect -12322 -13603 -12222 -13573
rect -12322 -13641 -12289 -13603
rect -12255 -13641 -12222 -13603
rect -12322 -13675 -12222 -13641
rect -12322 -13709 -12289 -13675
rect -12255 -13709 -12222 -13675
rect -12322 -13743 -12222 -13709
rect -12322 -13781 -12289 -13743
rect -12255 -13781 -12222 -13743
rect -12322 -13811 -12222 -13781
rect -12322 -13853 -12289 -13811
rect -12255 -13853 -12222 -13811
rect -12322 -13879 -12222 -13853
rect -12322 -13925 -12289 -13879
rect -12255 -13925 -12222 -13879
rect -12322 -13947 -12222 -13925
rect -9184 -13361 -9150 -13326
rect -9184 -13433 -9150 -13409
rect -9184 -13505 -9150 -13477
rect -9184 -13577 -9150 -13545
rect -9184 -13647 -9150 -13613
rect -9184 -13715 -9150 -13683
rect -9184 -13783 -9150 -13755
rect -9184 -13851 -9150 -13827
rect -9184 -13934 -9150 -13899
rect -8166 -13361 -8132 -13326
rect -8166 -13433 -8132 -13409
rect -8166 -13505 -8132 -13477
rect -8166 -13577 -8132 -13545
rect -8166 -13647 -8132 -13613
rect -8166 -13715 -8132 -13683
rect -8166 -13783 -8132 -13755
rect -8166 -13851 -8132 -13827
rect -8166 -13934 -8132 -13899
rect -7148 -13361 -7114 -13326
rect -7148 -13433 -7114 -13409
rect -7148 -13505 -7114 -13477
rect -7148 -13577 -7114 -13545
rect -7148 -13647 -7114 -13613
rect -7148 -13715 -7114 -13683
rect -7148 -13783 -7114 -13755
rect -7148 -13851 -7114 -13827
rect -7148 -13934 -7114 -13899
rect -6130 -13361 -6096 -13326
rect -6130 -13433 -6096 -13409
rect -6130 -13505 -6096 -13477
rect -6130 -13577 -6096 -13545
rect -6130 -13647 -6096 -13613
rect -6130 -13715 -6096 -13683
rect -6130 -13783 -6096 -13755
rect -6130 -13851 -6096 -13827
rect -6130 -13934 -6096 -13899
rect -5112 -13361 -5078 -13326
rect -5112 -13433 -5078 -13409
rect -5112 -13505 -5078 -13477
rect -5112 -13577 -5078 -13545
rect -5112 -13647 -5078 -13613
rect -5112 -13715 -5078 -13683
rect -5112 -13783 -5078 -13755
rect -5112 -13851 -5078 -13827
rect -5112 -13934 -5078 -13899
rect -4094 -13361 -4060 -13326
rect -4094 -13433 -4060 -13409
rect -4094 -13505 -4060 -13477
rect -4094 -13577 -4060 -13545
rect -4094 -13647 -4060 -13613
rect -4094 -13715 -4060 -13683
rect -4094 -13783 -4060 -13755
rect -4094 -13851 -4060 -13827
rect -4094 -13934 -4060 -13899
rect -3076 -13361 -3042 -13326
rect -3076 -13433 -3042 -13409
rect -3076 -13505 -3042 -13477
rect -3076 -13577 -3042 -13545
rect -3076 -13647 -3042 -13613
rect -3076 -13715 -3042 -13683
rect -3076 -13783 -3042 -13755
rect -3076 -13851 -3042 -13827
rect -3076 -13934 -3042 -13899
rect -2058 -13361 -2024 -13326
rect -2058 -13433 -2024 -13409
rect -2058 -13505 -2024 -13477
rect -2058 -13577 -2024 -13545
rect -2058 -13647 -2024 -13613
rect -2058 -13715 -2024 -13683
rect -2058 -13783 -2024 -13755
rect -2058 -13851 -2024 -13827
rect -2058 -13934 -2024 -13899
rect -1040 -13361 -1006 -13326
rect -1040 -13433 -1006 -13409
rect -1040 -13505 -1006 -13477
rect -1040 -13577 -1006 -13545
rect -1040 -13647 -1006 -13613
rect -1040 -13715 -1006 -13683
rect -1040 -13783 -1006 -13755
rect -1040 -13851 -1006 -13827
rect -1040 -13934 -1006 -13899
rect -22 -13361 12 -13326
rect -22 -13433 12 -13409
rect -22 -13505 12 -13477
rect -22 -13577 12 -13545
rect -22 -13647 12 -13613
rect -22 -13715 12 -13683
rect -22 -13783 12 -13755
rect -22 -13851 12 -13827
rect -22 -13934 12 -13899
rect 24822 -13369 24855 -13315
rect 24889 -13369 24922 -13315
rect 24822 -13387 24922 -13369
rect 24822 -13437 24855 -13387
rect 24889 -13437 24922 -13387
rect 24822 -13459 24922 -13437
rect 24822 -13505 24855 -13459
rect 24889 -13505 24922 -13459
rect 24822 -13531 24922 -13505
rect 24822 -13573 24855 -13531
rect 24889 -13573 24922 -13531
rect 24822 -13603 24922 -13573
rect 24822 -13641 24855 -13603
rect 24889 -13641 24922 -13603
rect 24822 -13675 24922 -13641
rect 24822 -13709 24855 -13675
rect 24889 -13709 24922 -13675
rect 24822 -13743 24922 -13709
rect 24822 -13781 24855 -13743
rect 24889 -13781 24922 -13743
rect 24822 -13811 24922 -13781
rect 24822 -13853 24855 -13811
rect 24889 -13853 24922 -13811
rect 24822 -13879 24922 -13853
rect 24822 -13925 24855 -13879
rect 24889 -13925 24922 -13879
rect -12322 -13997 -12289 -13947
rect -12255 -13997 -12222 -13947
rect 24822 -13947 24922 -13925
rect -7660 -13968 -7600 -13966
rect -6646 -13968 -6586 -13966
rect -2572 -13968 -2512 -13966
rect -1556 -13968 -1496 -13966
rect -12322 -14015 -12222 -13997
rect -8952 -14002 -8913 -13968
rect -8879 -14002 -8855 -13968
rect -8811 -14002 -8783 -13968
rect -8743 -14002 -8711 -13968
rect -8675 -14002 -8641 -13968
rect -8605 -14002 -8573 -13968
rect -8533 -14002 -8505 -13968
rect -8461 -14002 -8437 -13968
rect -8403 -14002 -8364 -13968
rect -7934 -14002 -7895 -13968
rect -7861 -14002 -7837 -13968
rect -7793 -14002 -7765 -13968
rect -7725 -14002 -7693 -13968
rect -7657 -14002 -7623 -13968
rect -7587 -14002 -7555 -13968
rect -7515 -14002 -7487 -13968
rect -7443 -14002 -7419 -13968
rect -7385 -14002 -7346 -13968
rect -6916 -14002 -6877 -13968
rect -6843 -14002 -6819 -13968
rect -6775 -14002 -6747 -13968
rect -6707 -14002 -6675 -13968
rect -6639 -14002 -6605 -13968
rect -6569 -14002 -6537 -13968
rect -6497 -14002 -6469 -13968
rect -6425 -14002 -6401 -13968
rect -6367 -14002 -6328 -13968
rect -5898 -14002 -5859 -13968
rect -5825 -14002 -5801 -13968
rect -5757 -14002 -5729 -13968
rect -5689 -14002 -5657 -13968
rect -5621 -14002 -5587 -13968
rect -5551 -14002 -5519 -13968
rect -5479 -14002 -5451 -13968
rect -5407 -14002 -5383 -13968
rect -5349 -14002 -5310 -13968
rect -4880 -14002 -4841 -13968
rect -4807 -14002 -4783 -13968
rect -4739 -14002 -4711 -13968
rect -4671 -14002 -4639 -13968
rect -4603 -14002 -4569 -13968
rect -4533 -14002 -4501 -13968
rect -4461 -14002 -4433 -13968
rect -4389 -14002 -4365 -13968
rect -4331 -14002 -4292 -13968
rect -3862 -14002 -3823 -13968
rect -3789 -14002 -3765 -13968
rect -3721 -14002 -3693 -13968
rect -3653 -14002 -3621 -13968
rect -3585 -14002 -3551 -13968
rect -3515 -14002 -3483 -13968
rect -3443 -14002 -3415 -13968
rect -3371 -14002 -3347 -13968
rect -3313 -14002 -3274 -13968
rect -2844 -14002 -2805 -13968
rect -2771 -14002 -2747 -13968
rect -2703 -14002 -2675 -13968
rect -2635 -14002 -2603 -13968
rect -2567 -14002 -2533 -13968
rect -2497 -14002 -2465 -13968
rect -2425 -14002 -2397 -13968
rect -2353 -14002 -2329 -13968
rect -2295 -14002 -2256 -13968
rect -1826 -14002 -1787 -13968
rect -1753 -14002 -1729 -13968
rect -1685 -14002 -1657 -13968
rect -1617 -14002 -1585 -13968
rect -1549 -14002 -1515 -13968
rect -1479 -14002 -1447 -13968
rect -1407 -14002 -1379 -13968
rect -1335 -14002 -1311 -13968
rect -1277 -14002 -1238 -13968
rect -808 -14002 -769 -13968
rect -735 -14002 -711 -13968
rect -667 -14002 -639 -13968
rect -599 -14002 -567 -13968
rect -531 -14002 -497 -13968
rect -461 -14002 -429 -13968
rect -389 -14002 -361 -13968
rect -317 -14002 -293 -13968
rect -259 -14002 -220 -13968
rect 24822 -13997 24855 -13947
rect 24889 -13997 24922 -13947
rect -12322 -14069 -12289 -14015
rect -12255 -14069 -12222 -14015
rect -12322 -14083 -12222 -14069
rect 24822 -14015 24922 -13997
rect 24822 -14069 24855 -14015
rect 24889 -14069 24922 -14015
rect -12322 -14141 -12289 -14083
rect -12255 -14141 -12222 -14083
rect -8952 -14110 -8913 -14076
rect -8879 -14110 -8855 -14076
rect -8811 -14110 -8783 -14076
rect -8743 -14110 -8711 -14076
rect -8675 -14110 -8641 -14076
rect -8605 -14110 -8573 -14076
rect -8533 -14110 -8505 -14076
rect -8461 -14110 -8437 -14076
rect -8403 -14110 -8364 -14076
rect -7934 -14110 -7895 -14076
rect -7861 -14110 -7837 -14076
rect -7793 -14110 -7765 -14076
rect -7725 -14110 -7693 -14076
rect -7657 -14110 -7623 -14076
rect -7587 -14110 -7555 -14076
rect -7515 -14110 -7487 -14076
rect -7443 -14110 -7419 -14076
rect -7385 -14110 -7346 -14076
rect -6916 -14110 -6877 -14076
rect -6843 -14110 -6819 -14076
rect -6775 -14110 -6747 -14076
rect -6707 -14110 -6675 -14076
rect -6639 -14110 -6605 -14076
rect -6569 -14110 -6537 -14076
rect -6497 -14110 -6469 -14076
rect -6425 -14110 -6401 -14076
rect -6367 -14110 -6328 -14076
rect -5898 -14110 -5859 -14076
rect -5825 -14110 -5801 -14076
rect -5757 -14110 -5729 -14076
rect -5689 -14110 -5657 -14076
rect -5621 -14110 -5587 -14076
rect -5551 -14110 -5519 -14076
rect -5479 -14110 -5451 -14076
rect -5407 -14110 -5383 -14076
rect -5349 -14110 -5310 -14076
rect -4880 -14110 -4841 -14076
rect -4807 -14110 -4783 -14076
rect -4739 -14110 -4711 -14076
rect -4671 -14110 -4639 -14076
rect -4603 -14110 -4569 -14076
rect -4533 -14110 -4501 -14076
rect -4461 -14110 -4433 -14076
rect -4389 -14110 -4365 -14076
rect -4331 -14110 -4292 -14076
rect -3862 -14110 -3823 -14076
rect -3789 -14110 -3765 -14076
rect -3721 -14110 -3693 -14076
rect -3653 -14110 -3621 -14076
rect -3585 -14110 -3551 -14076
rect -3515 -14110 -3483 -14076
rect -3443 -14110 -3415 -14076
rect -3371 -14110 -3347 -14076
rect -3313 -14110 -3274 -14076
rect -2844 -14110 -2805 -14076
rect -2771 -14110 -2747 -14076
rect -2703 -14110 -2675 -14076
rect -2635 -14110 -2603 -14076
rect -2567 -14110 -2533 -14076
rect -2497 -14110 -2465 -14076
rect -2425 -14110 -2397 -14076
rect -2353 -14110 -2329 -14076
rect -2295 -14110 -2256 -14076
rect -1826 -14110 -1787 -14076
rect -1753 -14110 -1729 -14076
rect -1685 -14110 -1657 -14076
rect -1617 -14110 -1585 -14076
rect -1549 -14110 -1515 -14076
rect -1479 -14110 -1447 -14076
rect -1407 -14110 -1379 -14076
rect -1335 -14110 -1311 -14076
rect -1277 -14110 -1238 -14076
rect -808 -14110 -769 -14076
rect -735 -14110 -711 -14076
rect -667 -14110 -639 -14076
rect -599 -14110 -567 -14076
rect -531 -14110 -497 -14076
rect -461 -14110 -429 -14076
rect -389 -14110 -361 -14076
rect -317 -14110 -293 -14076
rect -259 -14110 -220 -14076
rect 24822 -14083 24922 -14069
rect -12322 -14151 -12222 -14141
rect 24822 -14141 24855 -14083
rect 24889 -14141 24922 -14083
rect -12322 -14213 -12289 -14151
rect -12255 -14213 -12222 -14151
rect -12322 -14219 -12222 -14213
rect -12322 -14285 -12289 -14219
rect -12255 -14285 -12222 -14219
rect -12322 -14287 -12222 -14285
rect -12322 -14321 -12289 -14287
rect -12255 -14321 -12222 -14287
rect -12322 -14323 -12222 -14321
rect -12322 -14389 -12289 -14323
rect -12255 -14389 -12222 -14323
rect -12322 -14395 -12222 -14389
rect -12322 -14457 -12289 -14395
rect -12255 -14457 -12222 -14395
rect -12322 -14467 -12222 -14457
rect -12322 -14525 -12289 -14467
rect -12255 -14525 -12222 -14467
rect -12322 -14539 -12222 -14525
rect -12322 -14593 -12289 -14539
rect -12255 -14593 -12222 -14539
rect -12322 -14611 -12222 -14593
rect -12322 -14661 -12289 -14611
rect -12255 -14661 -12222 -14611
rect -12322 -14683 -12222 -14661
rect -12322 -14729 -12289 -14683
rect -12255 -14729 -12222 -14683
rect -12322 -14755 -12222 -14729
rect -9184 -14179 -9150 -14144
rect -9184 -14251 -9150 -14227
rect -9184 -14323 -9150 -14295
rect -9184 -14395 -9150 -14363
rect -9184 -14465 -9150 -14431
rect -9184 -14533 -9150 -14501
rect -9184 -14601 -9150 -14573
rect -9184 -14669 -9150 -14645
rect -9184 -14752 -9150 -14717
rect -8166 -14179 -8132 -14144
rect -8166 -14251 -8132 -14227
rect -8166 -14323 -8132 -14295
rect -8166 -14395 -8132 -14363
rect -8166 -14465 -8132 -14431
rect -8166 -14533 -8132 -14501
rect -8166 -14601 -8132 -14573
rect -8166 -14669 -8132 -14645
rect -8166 -14752 -8132 -14717
rect -7148 -14179 -7114 -14144
rect -7148 -14251 -7114 -14227
rect -7148 -14323 -7114 -14295
rect -7148 -14395 -7114 -14363
rect -7148 -14465 -7114 -14431
rect -7148 -14533 -7114 -14501
rect -7148 -14601 -7114 -14573
rect -7148 -14669 -7114 -14645
rect -7148 -14752 -7114 -14717
rect -6130 -14179 -6096 -14144
rect -6130 -14251 -6096 -14227
rect -6130 -14323 -6096 -14295
rect -6130 -14395 -6096 -14363
rect -6130 -14465 -6096 -14431
rect -6130 -14533 -6096 -14501
rect -6130 -14601 -6096 -14573
rect -6130 -14669 -6096 -14645
rect -6130 -14752 -6096 -14717
rect -5112 -14179 -5078 -14144
rect -5112 -14251 -5078 -14227
rect -5112 -14323 -5078 -14295
rect -5112 -14395 -5078 -14363
rect -5112 -14465 -5078 -14431
rect -5112 -14533 -5078 -14501
rect -5112 -14601 -5078 -14573
rect -5112 -14669 -5078 -14645
rect -5112 -14752 -5078 -14717
rect -4094 -14179 -4060 -14144
rect -4094 -14251 -4060 -14227
rect -4094 -14323 -4060 -14295
rect -4094 -14395 -4060 -14363
rect -4094 -14465 -4060 -14431
rect -4094 -14533 -4060 -14501
rect -4094 -14601 -4060 -14573
rect -4094 -14669 -4060 -14645
rect -4094 -14752 -4060 -14717
rect -3076 -14179 -3042 -14144
rect -3076 -14251 -3042 -14227
rect -3076 -14323 -3042 -14295
rect -3076 -14395 -3042 -14363
rect -3076 -14465 -3042 -14431
rect -3076 -14533 -3042 -14501
rect -3076 -14601 -3042 -14573
rect -3076 -14669 -3042 -14645
rect -3076 -14752 -3042 -14717
rect -2058 -14179 -2024 -14144
rect -2058 -14251 -2024 -14227
rect -2058 -14323 -2024 -14295
rect -2058 -14395 -2024 -14363
rect -2058 -14465 -2024 -14431
rect -2058 -14533 -2024 -14501
rect -2058 -14601 -2024 -14573
rect -2058 -14669 -2024 -14645
rect -2058 -14752 -2024 -14717
rect -1040 -14179 -1006 -14144
rect -1040 -14251 -1006 -14227
rect -1040 -14323 -1006 -14295
rect -1040 -14395 -1006 -14363
rect -1040 -14465 -1006 -14431
rect -1040 -14533 -1006 -14501
rect -1040 -14601 -1006 -14573
rect -1040 -14669 -1006 -14645
rect -1040 -14752 -1006 -14717
rect -22 -14179 12 -14144
rect 24822 -14151 24922 -14141
rect 2814 -14194 2853 -14160
rect 2887 -14194 2911 -14160
rect 2955 -14194 2983 -14160
rect 3023 -14194 3055 -14160
rect 3091 -14194 3125 -14160
rect 3161 -14194 3193 -14160
rect 3233 -14194 3261 -14160
rect 3305 -14194 3329 -14160
rect 3363 -14194 3402 -14160
rect 3832 -14194 3871 -14160
rect 3905 -14194 3929 -14160
rect 3973 -14194 4001 -14160
rect 4041 -14194 4073 -14160
rect 4109 -14194 4143 -14160
rect 4179 -14194 4211 -14160
rect 4251 -14194 4279 -14160
rect 4323 -14194 4347 -14160
rect 4381 -14194 4420 -14160
rect 4850 -14194 4889 -14160
rect 4923 -14194 4947 -14160
rect 4991 -14194 5019 -14160
rect 5059 -14194 5091 -14160
rect 5127 -14194 5161 -14160
rect 5197 -14194 5229 -14160
rect 5269 -14194 5297 -14160
rect 5341 -14194 5365 -14160
rect 5399 -14194 5438 -14160
rect 5868 -14194 5907 -14160
rect 5941 -14194 5965 -14160
rect 6009 -14194 6037 -14160
rect 6077 -14194 6109 -14160
rect 6145 -14194 6179 -14160
rect 6215 -14194 6247 -14160
rect 6287 -14194 6315 -14160
rect 6359 -14194 6383 -14160
rect 6417 -14194 6456 -14160
rect 6886 -14194 6925 -14160
rect 6959 -14194 6983 -14160
rect 7027 -14194 7055 -14160
rect 7095 -14194 7127 -14160
rect 7163 -14194 7197 -14160
rect 7233 -14194 7265 -14160
rect 7305 -14194 7333 -14160
rect 7377 -14194 7401 -14160
rect 7435 -14194 7474 -14160
rect 7904 -14194 7943 -14160
rect 7977 -14194 8001 -14160
rect 8045 -14194 8073 -14160
rect 8113 -14194 8145 -14160
rect 8181 -14194 8215 -14160
rect 8251 -14194 8283 -14160
rect 8323 -14194 8351 -14160
rect 8395 -14194 8419 -14160
rect 8453 -14194 8492 -14160
rect 8922 -14194 8961 -14160
rect 8995 -14194 9019 -14160
rect 9063 -14194 9091 -14160
rect 9131 -14194 9163 -14160
rect 9199 -14194 9233 -14160
rect 9269 -14194 9301 -14160
rect 9341 -14194 9369 -14160
rect 9413 -14194 9437 -14160
rect 9471 -14194 9510 -14160
rect 9940 -14194 9979 -14160
rect 10013 -14194 10037 -14160
rect 10081 -14194 10109 -14160
rect 10149 -14194 10181 -14160
rect 10217 -14194 10251 -14160
rect 10287 -14194 10319 -14160
rect 10359 -14194 10387 -14160
rect 10431 -14194 10455 -14160
rect 10489 -14194 10528 -14160
rect 10958 -14194 10997 -14160
rect 11031 -14194 11055 -14160
rect 11099 -14194 11127 -14160
rect 11167 -14194 11199 -14160
rect 11235 -14194 11269 -14160
rect 11305 -14194 11337 -14160
rect 11377 -14194 11405 -14160
rect 11449 -14194 11473 -14160
rect 11507 -14194 11546 -14160
rect 11976 -14194 12015 -14160
rect 12049 -14194 12073 -14160
rect 12117 -14194 12145 -14160
rect 12185 -14194 12217 -14160
rect 12253 -14194 12287 -14160
rect 12323 -14194 12355 -14160
rect 12395 -14194 12423 -14160
rect 12467 -14194 12491 -14160
rect 12525 -14194 12564 -14160
rect 12994 -14194 13033 -14160
rect 13067 -14194 13091 -14160
rect 13135 -14194 13163 -14160
rect 13203 -14194 13235 -14160
rect 13271 -14194 13305 -14160
rect 13341 -14194 13373 -14160
rect 13413 -14194 13441 -14160
rect 13485 -14194 13509 -14160
rect 13543 -14194 13582 -14160
rect 14012 -14194 14051 -14160
rect 14085 -14194 14109 -14160
rect 14153 -14194 14181 -14160
rect 14221 -14194 14253 -14160
rect 14289 -14194 14323 -14160
rect 14359 -14194 14391 -14160
rect 14431 -14194 14459 -14160
rect 14503 -14194 14527 -14160
rect 14561 -14194 14600 -14160
rect 15030 -14194 15069 -14160
rect 15103 -14194 15127 -14160
rect 15171 -14194 15199 -14160
rect 15239 -14194 15271 -14160
rect 15307 -14194 15341 -14160
rect 15377 -14194 15409 -14160
rect 15449 -14194 15477 -14160
rect 15521 -14194 15545 -14160
rect 15579 -14194 15618 -14160
rect 16048 -14194 16087 -14160
rect 16121 -14194 16145 -14160
rect 16189 -14194 16217 -14160
rect 16257 -14194 16289 -14160
rect 16325 -14194 16359 -14160
rect 16395 -14194 16427 -14160
rect 16467 -14194 16495 -14160
rect 16539 -14194 16563 -14160
rect 16597 -14194 16636 -14160
rect 17066 -14194 17105 -14160
rect 17139 -14194 17163 -14160
rect 17207 -14194 17235 -14160
rect 17275 -14194 17307 -14160
rect 17343 -14194 17377 -14160
rect 17413 -14194 17445 -14160
rect 17485 -14194 17513 -14160
rect 17557 -14194 17581 -14160
rect 17615 -14194 17654 -14160
rect 18084 -14194 18123 -14160
rect 18157 -14194 18181 -14160
rect 18225 -14194 18253 -14160
rect 18293 -14194 18325 -14160
rect 18361 -14194 18395 -14160
rect 18431 -14194 18463 -14160
rect 18503 -14194 18531 -14160
rect 18575 -14194 18599 -14160
rect 18633 -14194 18672 -14160
rect 19102 -14194 19141 -14160
rect 19175 -14194 19199 -14160
rect 19243 -14194 19271 -14160
rect 19311 -14194 19343 -14160
rect 19379 -14194 19413 -14160
rect 19449 -14194 19481 -14160
rect 19521 -14194 19549 -14160
rect 19593 -14194 19617 -14160
rect 19651 -14194 19690 -14160
rect 20120 -14194 20159 -14160
rect 20193 -14194 20217 -14160
rect 20261 -14194 20289 -14160
rect 20329 -14194 20361 -14160
rect 20397 -14194 20431 -14160
rect 20467 -14194 20499 -14160
rect 20539 -14194 20567 -14160
rect 20611 -14194 20635 -14160
rect 20669 -14194 20708 -14160
rect 21138 -14194 21177 -14160
rect 21211 -14194 21235 -14160
rect 21279 -14194 21307 -14160
rect 21347 -14194 21379 -14160
rect 21415 -14194 21449 -14160
rect 21485 -14194 21517 -14160
rect 21557 -14194 21585 -14160
rect 21629 -14194 21653 -14160
rect 21687 -14194 21726 -14160
rect 22156 -14194 22195 -14160
rect 22229 -14194 22253 -14160
rect 22297 -14194 22325 -14160
rect 22365 -14194 22397 -14160
rect 22433 -14194 22467 -14160
rect 22503 -14194 22535 -14160
rect 22575 -14194 22603 -14160
rect 22647 -14194 22671 -14160
rect 22705 -14194 22744 -14160
rect 12238 -14200 12298 -14194
rect -22 -14251 12 -14227
rect 24822 -14213 24855 -14151
rect 24889 -14213 24922 -14151
rect 24822 -14219 24922 -14213
rect -22 -14323 12 -14295
rect -22 -14395 12 -14363
rect -22 -14465 12 -14431
rect -22 -14533 12 -14501
rect -22 -14601 12 -14573
rect -22 -14669 12 -14645
rect -22 -14752 12 -14717
rect 2582 -14263 2616 -14228
rect 2582 -14335 2616 -14311
rect 2582 -14407 2616 -14379
rect 2582 -14479 2616 -14447
rect 2582 -14549 2616 -14515
rect 2582 -14617 2616 -14585
rect 2582 -14685 2616 -14657
rect -12322 -14797 -12289 -14755
rect -12255 -14797 -12222 -14755
rect 2582 -14753 2616 -14729
rect -7656 -14786 -7596 -14784
rect -6642 -14786 -6582 -14784
rect -2568 -14786 -2508 -14784
rect -1552 -14786 -1492 -14784
rect -12322 -14827 -12222 -14797
rect -8952 -14820 -8913 -14786
rect -8879 -14820 -8855 -14786
rect -8811 -14820 -8783 -14786
rect -8743 -14820 -8711 -14786
rect -8675 -14820 -8641 -14786
rect -8605 -14820 -8573 -14786
rect -8533 -14820 -8505 -14786
rect -8461 -14820 -8437 -14786
rect -8403 -14820 -8364 -14786
rect -7934 -14820 -7895 -14786
rect -7861 -14820 -7837 -14786
rect -7793 -14820 -7765 -14786
rect -7725 -14820 -7693 -14786
rect -7657 -14820 -7623 -14786
rect -7587 -14820 -7555 -14786
rect -7515 -14820 -7487 -14786
rect -7443 -14820 -7419 -14786
rect -7385 -14820 -7346 -14786
rect -6916 -14820 -6877 -14786
rect -6843 -14820 -6819 -14786
rect -6775 -14820 -6747 -14786
rect -6707 -14820 -6675 -14786
rect -6639 -14820 -6605 -14786
rect -6569 -14820 -6537 -14786
rect -6497 -14820 -6469 -14786
rect -6425 -14820 -6401 -14786
rect -6367 -14820 -6328 -14786
rect -5898 -14820 -5859 -14786
rect -5825 -14820 -5801 -14786
rect -5757 -14820 -5729 -14786
rect -5689 -14820 -5657 -14786
rect -5621 -14820 -5587 -14786
rect -5551 -14820 -5519 -14786
rect -5479 -14820 -5451 -14786
rect -5407 -14820 -5383 -14786
rect -5349 -14820 -5310 -14786
rect -4880 -14820 -4841 -14786
rect -4807 -14820 -4783 -14786
rect -4739 -14820 -4711 -14786
rect -4671 -14820 -4639 -14786
rect -4603 -14820 -4569 -14786
rect -4533 -14820 -4501 -14786
rect -4461 -14820 -4433 -14786
rect -4389 -14820 -4365 -14786
rect -4331 -14820 -4292 -14786
rect -3862 -14820 -3823 -14786
rect -3789 -14820 -3765 -14786
rect -3721 -14820 -3693 -14786
rect -3653 -14820 -3621 -14786
rect -3585 -14820 -3551 -14786
rect -3515 -14820 -3483 -14786
rect -3443 -14820 -3415 -14786
rect -3371 -14820 -3347 -14786
rect -3313 -14820 -3274 -14786
rect -2844 -14820 -2805 -14786
rect -2771 -14820 -2747 -14786
rect -2703 -14820 -2675 -14786
rect -2635 -14820 -2603 -14786
rect -2567 -14820 -2533 -14786
rect -2497 -14820 -2465 -14786
rect -2425 -14820 -2397 -14786
rect -2353 -14820 -2329 -14786
rect -2295 -14820 -2256 -14786
rect -1826 -14820 -1787 -14786
rect -1753 -14820 -1729 -14786
rect -1685 -14820 -1657 -14786
rect -1617 -14820 -1585 -14786
rect -1549 -14820 -1515 -14786
rect -1479 -14820 -1447 -14786
rect -1407 -14820 -1379 -14786
rect -1335 -14820 -1311 -14786
rect -1277 -14820 -1238 -14786
rect -808 -14820 -769 -14786
rect -735 -14820 -711 -14786
rect -667 -14820 -639 -14786
rect -599 -14820 -567 -14786
rect -531 -14820 -497 -14786
rect -461 -14820 -429 -14786
rect -389 -14820 -361 -14786
rect -317 -14820 -293 -14786
rect -259 -14820 -220 -14786
rect -12322 -14865 -12289 -14827
rect -12255 -14865 -12222 -14827
rect 2582 -14836 2616 -14801
rect 3600 -14263 3634 -14228
rect 3600 -14335 3634 -14311
rect 3600 -14407 3634 -14379
rect 3600 -14479 3634 -14447
rect 3600 -14549 3634 -14515
rect 3600 -14617 3634 -14585
rect 3600 -14685 3634 -14657
rect 3600 -14753 3634 -14729
rect 3600 -14836 3634 -14801
rect 4618 -14263 4652 -14228
rect 4618 -14335 4652 -14311
rect 4618 -14407 4652 -14379
rect 4618 -14479 4652 -14447
rect 4618 -14549 4652 -14515
rect 4618 -14617 4652 -14585
rect 4618 -14685 4652 -14657
rect 4618 -14753 4652 -14729
rect 4618 -14836 4652 -14801
rect 5636 -14263 5670 -14228
rect 5636 -14335 5670 -14311
rect 5636 -14407 5670 -14379
rect 5636 -14479 5670 -14447
rect 5636 -14549 5670 -14515
rect 5636 -14617 5670 -14585
rect 5636 -14685 5670 -14657
rect 5636 -14753 5670 -14729
rect 5636 -14836 5670 -14801
rect 6654 -14263 6688 -14228
rect 6654 -14335 6688 -14311
rect 6654 -14407 6688 -14379
rect 6654 -14479 6688 -14447
rect 6654 -14549 6688 -14515
rect 6654 -14617 6688 -14585
rect 6654 -14685 6688 -14657
rect 6654 -14753 6688 -14729
rect 6654 -14836 6688 -14801
rect 7672 -14263 7706 -14228
rect 7672 -14335 7706 -14311
rect 7672 -14407 7706 -14379
rect 7672 -14479 7706 -14447
rect 7672 -14549 7706 -14515
rect 7672 -14617 7706 -14585
rect 7672 -14685 7706 -14657
rect 7672 -14753 7706 -14729
rect 7672 -14836 7706 -14801
rect 8690 -14263 8724 -14228
rect 8690 -14335 8724 -14311
rect 8690 -14407 8724 -14379
rect 8690 -14479 8724 -14447
rect 8690 -14549 8724 -14515
rect 8690 -14617 8724 -14585
rect 8690 -14685 8724 -14657
rect 8690 -14753 8724 -14729
rect 8690 -14836 8724 -14801
rect 9708 -14263 9742 -14228
rect 9708 -14335 9742 -14311
rect 9708 -14407 9742 -14379
rect 9708 -14479 9742 -14447
rect 9708 -14549 9742 -14515
rect 9708 -14617 9742 -14585
rect 9708 -14685 9742 -14657
rect 9708 -14753 9742 -14729
rect 9708 -14836 9742 -14801
rect 10726 -14263 10760 -14228
rect 10726 -14335 10760 -14311
rect 10726 -14407 10760 -14379
rect 10726 -14479 10760 -14447
rect 10726 -14549 10760 -14515
rect 10726 -14617 10760 -14585
rect 10726 -14685 10760 -14657
rect 10726 -14753 10760 -14729
rect 10726 -14836 10760 -14801
rect 11744 -14263 11778 -14228
rect 11744 -14335 11778 -14311
rect 11744 -14407 11778 -14379
rect 11744 -14479 11778 -14447
rect 11744 -14549 11778 -14515
rect 11744 -14617 11778 -14585
rect 11744 -14685 11778 -14657
rect 11744 -14753 11778 -14729
rect 11744 -14836 11778 -14801
rect 12762 -14263 12796 -14228
rect 12762 -14335 12796 -14311
rect 12762 -14407 12796 -14379
rect 12762 -14479 12796 -14447
rect 12762 -14549 12796 -14515
rect 12762 -14617 12796 -14585
rect 12762 -14685 12796 -14657
rect 12762 -14753 12796 -14729
rect 12762 -14836 12796 -14801
rect 13780 -14263 13814 -14228
rect 13780 -14335 13814 -14311
rect 13780 -14407 13814 -14379
rect 13780 -14479 13814 -14447
rect 13780 -14549 13814 -14515
rect 13780 -14617 13814 -14585
rect 13780 -14685 13814 -14657
rect 13780 -14753 13814 -14729
rect 13780 -14836 13814 -14801
rect 14798 -14263 14832 -14228
rect 14798 -14335 14832 -14311
rect 14798 -14407 14832 -14379
rect 14798 -14479 14832 -14447
rect 14798 -14549 14832 -14515
rect 14798 -14617 14832 -14585
rect 14798 -14685 14832 -14657
rect 14798 -14753 14832 -14729
rect 14798 -14836 14832 -14801
rect 15816 -14263 15850 -14228
rect 15816 -14335 15850 -14311
rect 15816 -14407 15850 -14379
rect 15816 -14479 15850 -14447
rect 15816 -14549 15850 -14515
rect 15816 -14617 15850 -14585
rect 15816 -14685 15850 -14657
rect 15816 -14753 15850 -14729
rect 15816 -14836 15850 -14801
rect 16834 -14263 16868 -14228
rect 16834 -14335 16868 -14311
rect 16834 -14407 16868 -14379
rect 16834 -14479 16868 -14447
rect 16834 -14549 16868 -14515
rect 16834 -14617 16868 -14585
rect 16834 -14685 16868 -14657
rect 16834 -14753 16868 -14729
rect 16834 -14836 16868 -14801
rect 17852 -14263 17886 -14228
rect 17852 -14335 17886 -14311
rect 17852 -14407 17886 -14379
rect 17852 -14479 17886 -14447
rect 17852 -14549 17886 -14515
rect 17852 -14617 17886 -14585
rect 17852 -14685 17886 -14657
rect 17852 -14753 17886 -14729
rect 17852 -14836 17886 -14801
rect 18870 -14263 18904 -14228
rect 18870 -14335 18904 -14311
rect 18870 -14407 18904 -14379
rect 18870 -14479 18904 -14447
rect 18870 -14549 18904 -14515
rect 18870 -14617 18904 -14585
rect 18870 -14685 18904 -14657
rect 18870 -14753 18904 -14729
rect 18870 -14836 18904 -14801
rect 19888 -14263 19922 -14228
rect 19888 -14335 19922 -14311
rect 19888 -14407 19922 -14379
rect 19888 -14479 19922 -14447
rect 19888 -14549 19922 -14515
rect 19888 -14617 19922 -14585
rect 19888 -14685 19922 -14657
rect 19888 -14753 19922 -14729
rect 19888 -14836 19922 -14801
rect 20906 -14263 20940 -14228
rect 20906 -14335 20940 -14311
rect 20906 -14407 20940 -14379
rect 20906 -14479 20940 -14447
rect 20906 -14549 20940 -14515
rect 20906 -14617 20940 -14585
rect 20906 -14685 20940 -14657
rect 20906 -14753 20940 -14729
rect 20906 -14836 20940 -14801
rect 21924 -14263 21958 -14228
rect 21924 -14335 21958 -14311
rect 21924 -14407 21958 -14379
rect 21924 -14479 21958 -14447
rect 21924 -14549 21958 -14515
rect 21924 -14617 21958 -14585
rect 21924 -14685 21958 -14657
rect 21924 -14753 21958 -14729
rect 21924 -14836 21958 -14801
rect 22942 -14263 22976 -14228
rect 22942 -14335 22976 -14311
rect 22942 -14407 22976 -14379
rect 22942 -14479 22976 -14447
rect 22942 -14549 22976 -14515
rect 22942 -14617 22976 -14585
rect 22942 -14685 22976 -14657
rect 22942 -14753 22976 -14729
rect 22942 -14836 22976 -14801
rect 24822 -14285 24855 -14219
rect 24889 -14285 24922 -14219
rect 24822 -14287 24922 -14285
rect 24822 -14321 24855 -14287
rect 24889 -14321 24922 -14287
rect 24822 -14323 24922 -14321
rect 24822 -14389 24855 -14323
rect 24889 -14389 24922 -14323
rect 24822 -14395 24922 -14389
rect 24822 -14457 24855 -14395
rect 24889 -14457 24922 -14395
rect 24822 -14467 24922 -14457
rect 24822 -14525 24855 -14467
rect 24889 -14525 24922 -14467
rect 24822 -14539 24922 -14525
rect 24822 -14593 24855 -14539
rect 24889 -14593 24922 -14539
rect 24822 -14611 24922 -14593
rect 24822 -14661 24855 -14611
rect 24889 -14661 24922 -14611
rect 24822 -14683 24922 -14661
rect 24822 -14729 24855 -14683
rect 24889 -14729 24922 -14683
rect 24822 -14755 24922 -14729
rect 24822 -14797 24855 -14755
rect 24889 -14797 24922 -14755
rect 24822 -14827 24922 -14797
rect -12322 -14899 -12222 -14865
rect 8166 -14870 8226 -14864
rect 10202 -14870 10262 -14864
rect 11222 -14870 11282 -14864
rect 16294 -14870 16354 -14864
rect 24822 -14865 24855 -14827
rect 24889 -14865 24922 -14827
rect -12322 -14933 -12289 -14899
rect -12255 -14933 -12222 -14899
rect -8952 -14928 -8913 -14894
rect -8879 -14928 -8855 -14894
rect -8811 -14928 -8783 -14894
rect -8743 -14928 -8711 -14894
rect -8675 -14928 -8641 -14894
rect -8605 -14928 -8573 -14894
rect -8533 -14928 -8505 -14894
rect -8461 -14928 -8437 -14894
rect -8403 -14928 -8364 -14894
rect -7934 -14928 -7895 -14894
rect -7861 -14928 -7837 -14894
rect -7793 -14928 -7765 -14894
rect -7725 -14928 -7693 -14894
rect -7657 -14928 -7623 -14894
rect -7587 -14928 -7555 -14894
rect -7515 -14928 -7487 -14894
rect -7443 -14928 -7419 -14894
rect -7385 -14928 -7346 -14894
rect -6916 -14928 -6877 -14894
rect -6843 -14928 -6819 -14894
rect -6775 -14928 -6747 -14894
rect -6707 -14928 -6675 -14894
rect -6639 -14928 -6605 -14894
rect -6569 -14928 -6537 -14894
rect -6497 -14928 -6469 -14894
rect -6425 -14928 -6401 -14894
rect -6367 -14928 -6328 -14894
rect -5898 -14928 -5859 -14894
rect -5825 -14928 -5801 -14894
rect -5757 -14928 -5729 -14894
rect -5689 -14928 -5657 -14894
rect -5621 -14928 -5587 -14894
rect -5551 -14928 -5519 -14894
rect -5479 -14928 -5451 -14894
rect -5407 -14928 -5383 -14894
rect -5349 -14928 -5310 -14894
rect -4880 -14928 -4841 -14894
rect -4807 -14928 -4783 -14894
rect -4739 -14928 -4711 -14894
rect -4671 -14928 -4639 -14894
rect -4603 -14928 -4569 -14894
rect -4533 -14928 -4501 -14894
rect -4461 -14928 -4433 -14894
rect -4389 -14928 -4365 -14894
rect -4331 -14928 -4292 -14894
rect -3862 -14928 -3823 -14894
rect -3789 -14928 -3765 -14894
rect -3721 -14928 -3693 -14894
rect -3653 -14928 -3621 -14894
rect -3585 -14928 -3551 -14894
rect -3515 -14928 -3483 -14894
rect -3443 -14928 -3415 -14894
rect -3371 -14928 -3347 -14894
rect -3313 -14928 -3274 -14894
rect -2844 -14928 -2805 -14894
rect -2771 -14928 -2747 -14894
rect -2703 -14928 -2675 -14894
rect -2635 -14928 -2603 -14894
rect -2567 -14928 -2533 -14894
rect -2497 -14928 -2465 -14894
rect -2425 -14928 -2397 -14894
rect -2353 -14928 -2329 -14894
rect -2295 -14928 -2256 -14894
rect -1826 -14928 -1787 -14894
rect -1753 -14928 -1729 -14894
rect -1685 -14928 -1657 -14894
rect -1617 -14928 -1585 -14894
rect -1549 -14928 -1515 -14894
rect -1479 -14928 -1447 -14894
rect -1407 -14928 -1379 -14894
rect -1335 -14928 -1311 -14894
rect -1277 -14928 -1238 -14894
rect -808 -14928 -769 -14894
rect -735 -14928 -711 -14894
rect -667 -14928 -639 -14894
rect -599 -14928 -567 -14894
rect -531 -14928 -497 -14894
rect -461 -14928 -429 -14894
rect -389 -14928 -361 -14894
rect -317 -14928 -293 -14894
rect -259 -14928 -220 -14894
rect 2814 -14904 2853 -14870
rect 2887 -14904 2911 -14870
rect 2955 -14904 2983 -14870
rect 3023 -14904 3055 -14870
rect 3091 -14904 3125 -14870
rect 3161 -14904 3193 -14870
rect 3233 -14904 3261 -14870
rect 3305 -14904 3329 -14870
rect 3363 -14904 3402 -14870
rect 3832 -14904 3871 -14870
rect 3905 -14904 3929 -14870
rect 3973 -14904 4001 -14870
rect 4041 -14904 4073 -14870
rect 4109 -14904 4143 -14870
rect 4179 -14904 4211 -14870
rect 4251 -14904 4279 -14870
rect 4323 -14904 4347 -14870
rect 4381 -14904 4420 -14870
rect 4850 -14904 4889 -14870
rect 4923 -14904 4947 -14870
rect 4991 -14904 5019 -14870
rect 5059 -14904 5091 -14870
rect 5127 -14904 5161 -14870
rect 5197 -14904 5229 -14870
rect 5269 -14904 5297 -14870
rect 5341 -14904 5365 -14870
rect 5399 -14904 5438 -14870
rect 5868 -14904 5907 -14870
rect 5941 -14904 5965 -14870
rect 6009 -14904 6037 -14870
rect 6077 -14904 6109 -14870
rect 6145 -14904 6179 -14870
rect 6215 -14904 6247 -14870
rect 6287 -14904 6315 -14870
rect 6359 -14904 6383 -14870
rect 6417 -14904 6456 -14870
rect 6886 -14904 6925 -14870
rect 6959 -14904 6983 -14870
rect 7027 -14904 7055 -14870
rect 7095 -14904 7127 -14870
rect 7163 -14904 7197 -14870
rect 7233 -14904 7265 -14870
rect 7305 -14904 7333 -14870
rect 7377 -14904 7401 -14870
rect 7435 -14904 7474 -14870
rect 7904 -14904 7943 -14870
rect 7977 -14904 8001 -14870
rect 8045 -14904 8073 -14870
rect 8113 -14904 8145 -14870
rect 8181 -14904 8215 -14870
rect 8251 -14904 8283 -14870
rect 8323 -14904 8351 -14870
rect 8395 -14904 8419 -14870
rect 8453 -14904 8492 -14870
rect 8922 -14904 8961 -14870
rect 8995 -14904 9019 -14870
rect 9063 -14904 9091 -14870
rect 9131 -14904 9163 -14870
rect 9199 -14904 9233 -14870
rect 9269 -14904 9301 -14870
rect 9341 -14904 9369 -14870
rect 9413 -14904 9437 -14870
rect 9471 -14904 9510 -14870
rect 9940 -14904 9979 -14870
rect 10013 -14904 10037 -14870
rect 10081 -14904 10109 -14870
rect 10149 -14904 10181 -14870
rect 10217 -14904 10251 -14870
rect 10287 -14904 10319 -14870
rect 10359 -14904 10387 -14870
rect 10431 -14904 10455 -14870
rect 10489 -14904 10528 -14870
rect 10958 -14904 10997 -14870
rect 11031 -14904 11055 -14870
rect 11099 -14904 11127 -14870
rect 11167 -14904 11199 -14870
rect 11235 -14904 11269 -14870
rect 11305 -14904 11337 -14870
rect 11377 -14904 11405 -14870
rect 11449 -14904 11473 -14870
rect 11507 -14904 11546 -14870
rect 11976 -14904 12015 -14870
rect 12049 -14904 12073 -14870
rect 12117 -14904 12145 -14870
rect 12185 -14904 12217 -14870
rect 12253 -14904 12287 -14870
rect 12323 -14904 12355 -14870
rect 12395 -14904 12423 -14870
rect 12467 -14904 12491 -14870
rect 12525 -14904 12564 -14870
rect 12994 -14904 13033 -14870
rect 13067 -14904 13091 -14870
rect 13135 -14904 13163 -14870
rect 13203 -14904 13235 -14870
rect 13271 -14904 13305 -14870
rect 13341 -14904 13373 -14870
rect 13413 -14904 13441 -14870
rect 13485 -14904 13509 -14870
rect 13543 -14904 13582 -14870
rect 14012 -14904 14051 -14870
rect 14085 -14904 14109 -14870
rect 14153 -14904 14181 -14870
rect 14221 -14904 14253 -14870
rect 14289 -14904 14323 -14870
rect 14359 -14904 14391 -14870
rect 14431 -14904 14459 -14870
rect 14503 -14904 14527 -14870
rect 14561 -14904 14600 -14870
rect 15030 -14904 15069 -14870
rect 15103 -14904 15127 -14870
rect 15171 -14904 15199 -14870
rect 15239 -14904 15271 -14870
rect 15307 -14904 15341 -14870
rect 15377 -14904 15409 -14870
rect 15449 -14904 15477 -14870
rect 15521 -14904 15545 -14870
rect 15579 -14904 15618 -14870
rect 16048 -14904 16087 -14870
rect 16121 -14904 16145 -14870
rect 16189 -14904 16217 -14870
rect 16257 -14904 16289 -14870
rect 16325 -14904 16359 -14870
rect 16395 -14904 16427 -14870
rect 16467 -14904 16495 -14870
rect 16539 -14904 16563 -14870
rect 16597 -14904 16636 -14870
rect 17066 -14904 17105 -14870
rect 17139 -14904 17163 -14870
rect 17207 -14904 17235 -14870
rect 17275 -14904 17307 -14870
rect 17343 -14904 17377 -14870
rect 17413 -14904 17445 -14870
rect 17485 -14904 17513 -14870
rect 17557 -14904 17581 -14870
rect 17615 -14904 17654 -14870
rect 18084 -14904 18123 -14870
rect 18157 -14904 18181 -14870
rect 18225 -14904 18253 -14870
rect 18293 -14904 18325 -14870
rect 18361 -14904 18395 -14870
rect 18431 -14904 18463 -14870
rect 18503 -14904 18531 -14870
rect 18575 -14904 18599 -14870
rect 18633 -14904 18672 -14870
rect 19102 -14904 19141 -14870
rect 19175 -14904 19199 -14870
rect 19243 -14904 19271 -14870
rect 19311 -14904 19343 -14870
rect 19379 -14904 19413 -14870
rect 19449 -14904 19481 -14870
rect 19521 -14904 19549 -14870
rect 19593 -14904 19617 -14870
rect 19651 -14904 19690 -14870
rect 20120 -14904 20159 -14870
rect 20193 -14904 20217 -14870
rect 20261 -14904 20289 -14870
rect 20329 -14904 20361 -14870
rect 20397 -14904 20431 -14870
rect 20467 -14904 20499 -14870
rect 20539 -14904 20567 -14870
rect 20611 -14904 20635 -14870
rect 20669 -14904 20708 -14870
rect 21138 -14904 21177 -14870
rect 21211 -14904 21235 -14870
rect 21279 -14904 21307 -14870
rect 21347 -14904 21379 -14870
rect 21415 -14904 21449 -14870
rect 21485 -14904 21517 -14870
rect 21557 -14904 21585 -14870
rect 21629 -14904 21653 -14870
rect 21687 -14904 21726 -14870
rect 22156 -14904 22195 -14870
rect 22229 -14904 22253 -14870
rect 22297 -14904 22325 -14870
rect 22365 -14904 22397 -14870
rect 22433 -14904 22467 -14870
rect 22503 -14904 22535 -14870
rect 22575 -14904 22603 -14870
rect 22647 -14904 22671 -14870
rect 22705 -14904 22744 -14870
rect 24822 -14899 24922 -14865
rect -12322 -14967 -12222 -14933
rect 24822 -14933 24855 -14899
rect 24889 -14933 24922 -14899
rect -12322 -15005 -12289 -14967
rect -12255 -15005 -12222 -14967
rect -12322 -15035 -12222 -15005
rect -12322 -15077 -12289 -15035
rect -12255 -15077 -12222 -15035
rect -12322 -15103 -12222 -15077
rect -12322 -15149 -12289 -15103
rect -12255 -15149 -12222 -15103
rect -12322 -15171 -12222 -15149
rect -12322 -15221 -12289 -15171
rect -12255 -15221 -12222 -15171
rect -12322 -15239 -12222 -15221
rect -12322 -15293 -12289 -15239
rect -12255 -15293 -12222 -15239
rect -12322 -15307 -12222 -15293
rect -12322 -15365 -12289 -15307
rect -12255 -15365 -12222 -15307
rect -12322 -15375 -12222 -15365
rect -12322 -15437 -12289 -15375
rect -12255 -15437 -12222 -15375
rect -12322 -15443 -12222 -15437
rect -12322 -15509 -12289 -15443
rect -12255 -15509 -12222 -15443
rect -12322 -15511 -12222 -15509
rect -12322 -15545 -12289 -15511
rect -12255 -15545 -12222 -15511
rect -12322 -15547 -12222 -15545
rect -12322 -15613 -12289 -15547
rect -12255 -15613 -12222 -15547
rect -9184 -14997 -9150 -14962
rect -9184 -15069 -9150 -15045
rect -9184 -15141 -9150 -15113
rect -9184 -15213 -9150 -15181
rect -9184 -15283 -9150 -15249
rect -9184 -15351 -9150 -15319
rect -9184 -15419 -9150 -15391
rect -9184 -15487 -9150 -15463
rect -9184 -15570 -9150 -15535
rect -8166 -14997 -8132 -14962
rect -8166 -15069 -8132 -15045
rect -8166 -15141 -8132 -15113
rect -8166 -15213 -8132 -15181
rect -8166 -15283 -8132 -15249
rect -8166 -15351 -8132 -15319
rect -8166 -15419 -8132 -15391
rect -8166 -15487 -8132 -15463
rect -8166 -15570 -8132 -15535
rect -7148 -14997 -7114 -14962
rect -7148 -15069 -7114 -15045
rect -7148 -15141 -7114 -15113
rect -7148 -15213 -7114 -15181
rect -7148 -15283 -7114 -15249
rect -7148 -15351 -7114 -15319
rect -7148 -15419 -7114 -15391
rect -7148 -15487 -7114 -15463
rect -7148 -15570 -7114 -15535
rect -6130 -14997 -6096 -14962
rect -6130 -15069 -6096 -15045
rect -6130 -15141 -6096 -15113
rect -6130 -15213 -6096 -15181
rect -6130 -15283 -6096 -15249
rect -6130 -15351 -6096 -15319
rect -6130 -15419 -6096 -15391
rect -6130 -15487 -6096 -15463
rect -6130 -15570 -6096 -15535
rect -5112 -14997 -5078 -14962
rect -5112 -15069 -5078 -15045
rect -5112 -15141 -5078 -15113
rect -5112 -15213 -5078 -15181
rect -5112 -15283 -5078 -15249
rect -5112 -15351 -5078 -15319
rect -5112 -15419 -5078 -15391
rect -5112 -15487 -5078 -15463
rect -5112 -15570 -5078 -15535
rect -4094 -14997 -4060 -14962
rect -4094 -15069 -4060 -15045
rect -4094 -15141 -4060 -15113
rect -4094 -15213 -4060 -15181
rect -4094 -15283 -4060 -15249
rect -4094 -15351 -4060 -15319
rect -4094 -15419 -4060 -15391
rect -4094 -15487 -4060 -15463
rect -4094 -15570 -4060 -15535
rect -3076 -14997 -3042 -14962
rect -3076 -15069 -3042 -15045
rect -3076 -15141 -3042 -15113
rect -3076 -15213 -3042 -15181
rect -3076 -15283 -3042 -15249
rect -3076 -15351 -3042 -15319
rect -3076 -15419 -3042 -15391
rect -3076 -15487 -3042 -15463
rect -3076 -15570 -3042 -15535
rect -2058 -14997 -2024 -14962
rect -2058 -15069 -2024 -15045
rect -2058 -15141 -2024 -15113
rect -2058 -15213 -2024 -15181
rect -2058 -15283 -2024 -15249
rect -2058 -15351 -2024 -15319
rect -2058 -15419 -2024 -15391
rect -2058 -15487 -2024 -15463
rect -2058 -15570 -2024 -15535
rect -1040 -14997 -1006 -14962
rect -1040 -15069 -1006 -15045
rect -1040 -15141 -1006 -15113
rect -1040 -15213 -1006 -15181
rect -1040 -15283 -1006 -15249
rect -1040 -15351 -1006 -15319
rect -1040 -15419 -1006 -15391
rect -1040 -15487 -1006 -15463
rect -1040 -15570 -1006 -15535
rect -22 -14997 12 -14962
rect -22 -15069 12 -15045
rect -22 -15141 12 -15113
rect -22 -15213 12 -15181
rect -22 -15283 12 -15249
rect -22 -15351 12 -15319
rect -22 -15419 12 -15391
rect 24822 -14967 24922 -14933
rect 24822 -15005 24855 -14967
rect 24889 -15005 24922 -14967
rect 24822 -15035 24922 -15005
rect 24822 -15077 24855 -15035
rect 24889 -15077 24922 -15035
rect 24822 -15103 24922 -15077
rect 24822 -15149 24855 -15103
rect 24889 -15149 24922 -15103
rect 24822 -15171 24922 -15149
rect 24822 -15221 24855 -15171
rect 24889 -15221 24922 -15171
rect 24822 -15239 24922 -15221
rect 24822 -15293 24855 -15239
rect 24889 -15293 24922 -15239
rect 24822 -15307 24922 -15293
rect 24822 -15365 24855 -15307
rect 24889 -15365 24922 -15307
rect 24822 -15375 24922 -15365
rect 2814 -15426 2853 -15392
rect 2887 -15426 2911 -15392
rect 2955 -15426 2983 -15392
rect 3023 -15426 3055 -15392
rect 3091 -15426 3125 -15392
rect 3161 -15426 3193 -15392
rect 3233 -15426 3261 -15392
rect 3305 -15426 3329 -15392
rect 3363 -15426 3402 -15392
rect 3832 -15426 3871 -15392
rect 3905 -15426 3929 -15392
rect 3973 -15426 4001 -15392
rect 4041 -15426 4073 -15392
rect 4109 -15426 4143 -15392
rect 4179 -15426 4211 -15392
rect 4251 -15426 4279 -15392
rect 4323 -15426 4347 -15392
rect 4381 -15426 4420 -15392
rect 4850 -15426 4889 -15392
rect 4923 -15426 4947 -15392
rect 4991 -15426 5019 -15392
rect 5059 -15426 5091 -15392
rect 5127 -15426 5161 -15392
rect 5197 -15426 5229 -15392
rect 5269 -15426 5297 -15392
rect 5341 -15426 5365 -15392
rect 5399 -15426 5438 -15392
rect 5868 -15426 5907 -15392
rect 5941 -15426 5965 -15392
rect 6009 -15426 6037 -15392
rect 6077 -15426 6109 -15392
rect 6145 -15426 6179 -15392
rect 6215 -15426 6247 -15392
rect 6287 -15426 6315 -15392
rect 6359 -15426 6383 -15392
rect 6417 -15426 6456 -15392
rect 6886 -15426 6925 -15392
rect 6959 -15426 6983 -15392
rect 7027 -15426 7055 -15392
rect 7095 -15426 7127 -15392
rect 7163 -15426 7197 -15392
rect 7233 -15426 7265 -15392
rect 7305 -15426 7333 -15392
rect 7377 -15426 7401 -15392
rect 7435 -15426 7474 -15392
rect 7904 -15426 7943 -15392
rect 7977 -15426 8001 -15392
rect 8045 -15426 8073 -15392
rect 8113 -15426 8145 -15392
rect 8181 -15426 8215 -15392
rect 8251 -15426 8283 -15392
rect 8323 -15426 8351 -15392
rect 8395 -15426 8419 -15392
rect 8453 -15426 8492 -15392
rect 8922 -15426 8961 -15392
rect 8995 -15426 9019 -15392
rect 9063 -15426 9091 -15392
rect 9131 -15426 9163 -15392
rect 9199 -15426 9233 -15392
rect 9269 -15426 9301 -15392
rect 9341 -15426 9369 -15392
rect 9413 -15426 9437 -15392
rect 9471 -15426 9510 -15392
rect 9940 -15426 9979 -15392
rect 10013 -15426 10037 -15392
rect 10081 -15426 10109 -15392
rect 10149 -15426 10181 -15392
rect 10217 -15426 10251 -15392
rect 10287 -15426 10319 -15392
rect 10359 -15426 10387 -15392
rect 10431 -15426 10455 -15392
rect 10489 -15426 10528 -15392
rect 10958 -15426 10997 -15392
rect 11031 -15426 11055 -15392
rect 11099 -15426 11127 -15392
rect 11167 -15426 11199 -15392
rect 11235 -15426 11269 -15392
rect 11305 -15426 11337 -15392
rect 11377 -15426 11405 -15392
rect 11449 -15426 11473 -15392
rect 11507 -15426 11546 -15392
rect 11976 -15426 12015 -15392
rect 12049 -15426 12073 -15392
rect 12117 -15426 12145 -15392
rect 12185 -15426 12217 -15392
rect 12253 -15426 12287 -15392
rect 12323 -15426 12355 -15392
rect 12395 -15426 12423 -15392
rect 12467 -15426 12491 -15392
rect 12525 -15426 12564 -15392
rect 12994 -15426 13033 -15392
rect 13067 -15426 13091 -15392
rect 13135 -15426 13163 -15392
rect 13203 -15426 13235 -15392
rect 13271 -15426 13305 -15392
rect 13341 -15426 13373 -15392
rect 13413 -15426 13441 -15392
rect 13485 -15426 13509 -15392
rect 13543 -15426 13582 -15392
rect 14012 -15426 14051 -15392
rect 14085 -15426 14109 -15392
rect 14153 -15426 14181 -15392
rect 14221 -15426 14253 -15392
rect 14289 -15426 14323 -15392
rect 14359 -15426 14391 -15392
rect 14431 -15426 14459 -15392
rect 14503 -15426 14527 -15392
rect 14561 -15426 14600 -15392
rect 15030 -15426 15069 -15392
rect 15103 -15426 15127 -15392
rect 15171 -15426 15199 -15392
rect 15239 -15426 15271 -15392
rect 15307 -15426 15341 -15392
rect 15377 -15426 15409 -15392
rect 15449 -15426 15477 -15392
rect 15521 -15426 15545 -15392
rect 15579 -15426 15618 -15392
rect 16048 -15426 16087 -15392
rect 16121 -15426 16145 -15392
rect 16189 -15426 16217 -15392
rect 16257 -15426 16289 -15392
rect 16325 -15426 16359 -15392
rect 16395 -15426 16427 -15392
rect 16467 -15426 16495 -15392
rect 16539 -15426 16563 -15392
rect 16597 -15426 16636 -15392
rect 17066 -15426 17105 -15392
rect 17139 -15426 17163 -15392
rect 17207 -15426 17235 -15392
rect 17275 -15426 17307 -15392
rect 17343 -15426 17377 -15392
rect 17413 -15426 17445 -15392
rect 17485 -15426 17513 -15392
rect 17557 -15426 17581 -15392
rect 17615 -15426 17654 -15392
rect 18084 -15426 18123 -15392
rect 18157 -15426 18181 -15392
rect 18225 -15426 18253 -15392
rect 18293 -15426 18325 -15392
rect 18361 -15426 18395 -15392
rect 18431 -15426 18463 -15392
rect 18503 -15426 18531 -15392
rect 18575 -15426 18599 -15392
rect 18633 -15426 18672 -15392
rect 19102 -15426 19141 -15392
rect 19175 -15426 19199 -15392
rect 19243 -15426 19271 -15392
rect 19311 -15426 19343 -15392
rect 19379 -15426 19413 -15392
rect 19449 -15426 19481 -15392
rect 19521 -15426 19549 -15392
rect 19593 -15426 19617 -15392
rect 19651 -15426 19690 -15392
rect 20120 -15426 20159 -15392
rect 20193 -15426 20217 -15392
rect 20261 -15426 20289 -15392
rect 20329 -15426 20361 -15392
rect 20397 -15426 20431 -15392
rect 20467 -15426 20499 -15392
rect 20539 -15426 20567 -15392
rect 20611 -15426 20635 -15392
rect 20669 -15426 20708 -15392
rect 21138 -15426 21177 -15392
rect 21211 -15426 21235 -15392
rect 21279 -15426 21307 -15392
rect 21347 -15426 21379 -15392
rect 21415 -15426 21449 -15392
rect 21485 -15426 21517 -15392
rect 21557 -15426 21585 -15392
rect 21629 -15426 21653 -15392
rect 21687 -15426 21726 -15392
rect 22156 -15426 22195 -15392
rect 22229 -15426 22253 -15392
rect 22297 -15426 22325 -15392
rect 22365 -15426 22397 -15392
rect 22433 -15426 22467 -15392
rect 22503 -15426 22535 -15392
rect 22575 -15426 22603 -15392
rect 22647 -15426 22671 -15392
rect 22705 -15426 22744 -15392
rect 4100 -15430 4160 -15426
rect 5116 -15430 5176 -15426
rect 9192 -15434 9252 -15426
rect 13258 -15430 13318 -15426
rect 15292 -15430 15352 -15426
rect 21404 -15430 21464 -15426
rect 24822 -15437 24855 -15375
rect 24889 -15437 24922 -15375
rect 24822 -15443 24922 -15437
rect -22 -15487 12 -15463
rect -22 -15570 12 -15535
rect 2582 -15495 2616 -15460
rect 2582 -15567 2616 -15543
rect -12322 -15619 -12222 -15613
rect -12322 -15681 -12289 -15619
rect -12255 -15681 -12222 -15619
rect -8952 -15638 -8913 -15604
rect -8879 -15638 -8855 -15604
rect -8811 -15638 -8783 -15604
rect -8743 -15638 -8711 -15604
rect -8675 -15638 -8641 -15604
rect -8605 -15638 -8573 -15604
rect -8533 -15638 -8505 -15604
rect -8461 -15638 -8437 -15604
rect -8403 -15638 -8364 -15604
rect -7934 -15638 -7895 -15604
rect -7861 -15638 -7837 -15604
rect -7793 -15638 -7765 -15604
rect -7725 -15638 -7693 -15604
rect -7657 -15638 -7623 -15604
rect -7587 -15638 -7555 -15604
rect -7515 -15638 -7487 -15604
rect -7443 -15638 -7419 -15604
rect -7385 -15638 -7346 -15604
rect -6916 -15638 -6877 -15604
rect -6843 -15638 -6819 -15604
rect -6775 -15638 -6747 -15604
rect -6707 -15638 -6675 -15604
rect -6639 -15638 -6605 -15604
rect -6569 -15638 -6537 -15604
rect -6497 -15638 -6469 -15604
rect -6425 -15638 -6401 -15604
rect -6367 -15638 -6328 -15604
rect -5898 -15638 -5859 -15604
rect -5825 -15638 -5801 -15604
rect -5757 -15638 -5729 -15604
rect -5689 -15638 -5657 -15604
rect -5621 -15638 -5587 -15604
rect -5551 -15638 -5519 -15604
rect -5479 -15638 -5451 -15604
rect -5407 -15638 -5383 -15604
rect -5349 -15638 -5310 -15604
rect -4880 -15638 -4841 -15604
rect -4807 -15638 -4783 -15604
rect -4739 -15638 -4711 -15604
rect -4671 -15638 -4639 -15604
rect -4603 -15638 -4569 -15604
rect -4533 -15638 -4501 -15604
rect -4461 -15638 -4433 -15604
rect -4389 -15638 -4365 -15604
rect -4331 -15638 -4292 -15604
rect -3862 -15638 -3823 -15604
rect -3789 -15638 -3765 -15604
rect -3721 -15638 -3693 -15604
rect -3653 -15638 -3621 -15604
rect -3585 -15638 -3551 -15604
rect -3515 -15638 -3483 -15604
rect -3443 -15638 -3415 -15604
rect -3371 -15638 -3347 -15604
rect -3313 -15638 -3274 -15604
rect -2844 -15638 -2805 -15604
rect -2771 -15638 -2747 -15604
rect -2703 -15638 -2675 -15604
rect -2635 -15638 -2603 -15604
rect -2567 -15638 -2533 -15604
rect -2497 -15638 -2465 -15604
rect -2425 -15638 -2397 -15604
rect -2353 -15638 -2329 -15604
rect -2295 -15638 -2256 -15604
rect -1826 -15638 -1787 -15604
rect -1753 -15638 -1729 -15604
rect -1685 -15638 -1657 -15604
rect -1617 -15638 -1585 -15604
rect -1549 -15638 -1515 -15604
rect -1479 -15638 -1447 -15604
rect -1407 -15638 -1379 -15604
rect -1335 -15638 -1311 -15604
rect -1277 -15638 -1238 -15604
rect -808 -15638 -769 -15604
rect -735 -15638 -711 -15604
rect -667 -15638 -639 -15604
rect -599 -15638 -567 -15604
rect -531 -15638 -497 -15604
rect -461 -15638 -429 -15604
rect -389 -15638 -361 -15604
rect -317 -15638 -293 -15604
rect -259 -15638 -220 -15604
rect -12322 -15691 -12222 -15681
rect -12322 -15749 -12289 -15691
rect -12255 -15749 -12222 -15691
rect 2582 -15639 2616 -15611
rect 2582 -15711 2616 -15679
rect -8952 -15746 -8913 -15712
rect -8879 -15746 -8855 -15712
rect -8811 -15746 -8783 -15712
rect -8743 -15746 -8711 -15712
rect -8675 -15746 -8641 -15712
rect -8605 -15746 -8573 -15712
rect -8533 -15746 -8505 -15712
rect -8461 -15746 -8437 -15712
rect -8403 -15746 -8364 -15712
rect -7934 -15746 -7895 -15712
rect -7861 -15746 -7837 -15712
rect -7793 -15746 -7765 -15712
rect -7725 -15746 -7693 -15712
rect -7657 -15746 -7623 -15712
rect -7587 -15746 -7555 -15712
rect -7515 -15746 -7487 -15712
rect -7443 -15746 -7419 -15712
rect -7385 -15746 -7346 -15712
rect -6916 -15746 -6877 -15712
rect -6843 -15746 -6819 -15712
rect -6775 -15746 -6747 -15712
rect -6707 -15746 -6675 -15712
rect -6639 -15746 -6605 -15712
rect -6569 -15746 -6537 -15712
rect -6497 -15746 -6469 -15712
rect -6425 -15746 -6401 -15712
rect -6367 -15746 -6328 -15712
rect -5898 -15746 -5859 -15712
rect -5825 -15746 -5801 -15712
rect -5757 -15746 -5729 -15712
rect -5689 -15746 -5657 -15712
rect -5621 -15746 -5587 -15712
rect -5551 -15746 -5519 -15712
rect -5479 -15746 -5451 -15712
rect -5407 -15746 -5383 -15712
rect -5349 -15746 -5310 -15712
rect -4880 -15746 -4841 -15712
rect -4807 -15746 -4783 -15712
rect -4739 -15746 -4711 -15712
rect -4671 -15746 -4639 -15712
rect -4603 -15746 -4569 -15712
rect -4533 -15746 -4501 -15712
rect -4461 -15746 -4433 -15712
rect -4389 -15746 -4365 -15712
rect -4331 -15746 -4292 -15712
rect -3862 -15746 -3823 -15712
rect -3789 -15746 -3765 -15712
rect -3721 -15746 -3693 -15712
rect -3653 -15746 -3621 -15712
rect -3585 -15746 -3551 -15712
rect -3515 -15746 -3483 -15712
rect -3443 -15746 -3415 -15712
rect -3371 -15746 -3347 -15712
rect -3313 -15746 -3274 -15712
rect -2844 -15746 -2805 -15712
rect -2771 -15746 -2747 -15712
rect -2703 -15746 -2675 -15712
rect -2635 -15746 -2603 -15712
rect -2567 -15746 -2533 -15712
rect -2497 -15746 -2465 -15712
rect -2425 -15746 -2397 -15712
rect -2353 -15746 -2329 -15712
rect -2295 -15746 -2256 -15712
rect -1826 -15746 -1787 -15712
rect -1753 -15746 -1729 -15712
rect -1685 -15746 -1657 -15712
rect -1617 -15746 -1585 -15712
rect -1549 -15746 -1515 -15712
rect -1479 -15746 -1447 -15712
rect -1407 -15746 -1379 -15712
rect -1335 -15746 -1311 -15712
rect -1277 -15746 -1238 -15712
rect -808 -15746 -769 -15712
rect -735 -15746 -711 -15712
rect -667 -15746 -639 -15712
rect -599 -15746 -567 -15712
rect -531 -15746 -497 -15712
rect -461 -15746 -429 -15712
rect -389 -15746 -361 -15712
rect -317 -15746 -293 -15712
rect -259 -15746 -220 -15712
rect -3596 -15748 -3536 -15746
rect -12322 -15763 -12222 -15749
rect -12322 -15817 -12289 -15763
rect -12255 -15817 -12222 -15763
rect -12322 -15835 -12222 -15817
rect -12322 -15885 -12289 -15835
rect -12255 -15885 -12222 -15835
rect -12322 -15907 -12222 -15885
rect -12322 -15953 -12289 -15907
rect -12255 -15953 -12222 -15907
rect -12322 -15979 -12222 -15953
rect -12322 -16021 -12289 -15979
rect -12255 -16021 -12222 -15979
rect -12322 -16051 -12222 -16021
rect -12322 -16089 -12289 -16051
rect -12255 -16089 -12222 -16051
rect -12322 -16123 -12222 -16089
rect -12322 -16157 -12289 -16123
rect -12255 -16157 -12222 -16123
rect -12322 -16191 -12222 -16157
rect -12322 -16229 -12289 -16191
rect -12255 -16229 -12222 -16191
rect -12322 -16259 -12222 -16229
rect -12322 -16301 -12289 -16259
rect -12255 -16301 -12222 -16259
rect -12322 -16327 -12222 -16301
rect -12322 -16373 -12289 -16327
rect -12255 -16373 -12222 -16327
rect -12322 -16395 -12222 -16373
rect -9184 -15815 -9150 -15780
rect -9184 -15887 -9150 -15863
rect -9184 -15959 -9150 -15931
rect -9184 -16031 -9150 -15999
rect -9184 -16101 -9150 -16067
rect -9184 -16169 -9150 -16137
rect -9184 -16237 -9150 -16209
rect -9184 -16305 -9150 -16281
rect -9184 -16388 -9150 -16353
rect -8166 -15815 -8132 -15780
rect -8166 -15887 -8132 -15863
rect -8166 -15959 -8132 -15931
rect -8166 -16031 -8132 -15999
rect -8166 -16101 -8132 -16067
rect -8166 -16169 -8132 -16137
rect -8166 -16237 -8132 -16209
rect -8166 -16305 -8132 -16281
rect -8166 -16388 -8132 -16353
rect -7148 -15815 -7114 -15780
rect -7148 -15887 -7114 -15863
rect -7148 -15959 -7114 -15931
rect -7148 -16031 -7114 -15999
rect -7148 -16101 -7114 -16067
rect -7148 -16169 -7114 -16137
rect -7148 -16237 -7114 -16209
rect -7148 -16305 -7114 -16281
rect -7148 -16388 -7114 -16353
rect -6130 -15815 -6096 -15780
rect -6130 -15887 -6096 -15863
rect -6130 -15959 -6096 -15931
rect -6130 -16031 -6096 -15999
rect -6130 -16101 -6096 -16067
rect -6130 -16169 -6096 -16137
rect -6130 -16237 -6096 -16209
rect -6130 -16305 -6096 -16281
rect -6130 -16388 -6096 -16353
rect -5112 -15815 -5078 -15780
rect -5112 -15887 -5078 -15863
rect -5112 -15959 -5078 -15931
rect -5112 -16031 -5078 -15999
rect -5112 -16101 -5078 -16067
rect -5112 -16169 -5078 -16137
rect -5112 -16237 -5078 -16209
rect -5112 -16305 -5078 -16281
rect -5112 -16388 -5078 -16353
rect -4094 -15815 -4060 -15780
rect -4094 -15887 -4060 -15863
rect -4094 -15959 -4060 -15931
rect -4094 -16031 -4060 -15999
rect -4094 -16101 -4060 -16067
rect -4094 -16169 -4060 -16137
rect -4094 -16237 -4060 -16209
rect -4094 -16305 -4060 -16281
rect -4094 -16388 -4060 -16353
rect -3076 -15815 -3042 -15780
rect -3076 -15887 -3042 -15863
rect -3076 -15959 -3042 -15931
rect -3076 -16031 -3042 -15999
rect -3076 -16101 -3042 -16067
rect -3076 -16169 -3042 -16137
rect -3076 -16237 -3042 -16209
rect -3076 -16305 -3042 -16281
rect -3076 -16388 -3042 -16353
rect -2058 -15815 -2024 -15780
rect -2058 -15887 -2024 -15863
rect -2058 -15959 -2024 -15931
rect -2058 -16031 -2024 -15999
rect -2058 -16101 -2024 -16067
rect -2058 -16169 -2024 -16137
rect -2058 -16237 -2024 -16209
rect -2058 -16305 -2024 -16281
rect -2058 -16388 -2024 -16353
rect -1040 -15815 -1006 -15780
rect -1040 -15887 -1006 -15863
rect -1040 -15959 -1006 -15931
rect -1040 -16031 -1006 -15999
rect -1040 -16101 -1006 -16067
rect -1040 -16169 -1006 -16137
rect -1040 -16237 -1006 -16209
rect -1040 -16305 -1006 -16281
rect -1040 -16388 -1006 -16353
rect -22 -15815 12 -15780
rect -22 -15887 12 -15863
rect -22 -15959 12 -15931
rect -22 -16031 12 -15999
rect -22 -16101 12 -16067
rect 2582 -15781 2616 -15747
rect 2582 -15849 2616 -15817
rect 2582 -15917 2616 -15889
rect 2582 -15985 2616 -15961
rect 2582 -16068 2616 -16033
rect 3600 -15495 3634 -15460
rect 3600 -15567 3634 -15543
rect 3600 -15639 3634 -15611
rect 3600 -15711 3634 -15679
rect 3600 -15781 3634 -15747
rect 3600 -15849 3634 -15817
rect 3600 -15917 3634 -15889
rect 3600 -15985 3634 -15961
rect 3600 -16068 3634 -16033
rect 4618 -15495 4652 -15460
rect 4618 -15567 4652 -15543
rect 4618 -15639 4652 -15611
rect 4618 -15711 4652 -15679
rect 4618 -15781 4652 -15747
rect 4618 -15849 4652 -15817
rect 4618 -15917 4652 -15889
rect 4618 -15985 4652 -15961
rect 4618 -16068 4652 -16033
rect 5636 -15495 5670 -15460
rect 5636 -15567 5670 -15543
rect 5636 -15639 5670 -15611
rect 5636 -15711 5670 -15679
rect 5636 -15781 5670 -15747
rect 5636 -15849 5670 -15817
rect 5636 -15917 5670 -15889
rect 5636 -15985 5670 -15961
rect 5636 -16068 5670 -16033
rect 6654 -15495 6688 -15460
rect 6654 -15567 6688 -15543
rect 6654 -15639 6688 -15611
rect 6654 -15711 6688 -15679
rect 6654 -15781 6688 -15747
rect 6654 -15849 6688 -15817
rect 6654 -15917 6688 -15889
rect 6654 -15985 6688 -15961
rect 6654 -16068 6688 -16033
rect 7672 -15495 7706 -15460
rect 7672 -15567 7706 -15543
rect 7672 -15639 7706 -15611
rect 7672 -15711 7706 -15679
rect 7672 -15781 7706 -15747
rect 7672 -15849 7706 -15817
rect 7672 -15917 7706 -15889
rect 7672 -15985 7706 -15961
rect 7672 -16068 7706 -16033
rect 8690 -15495 8724 -15460
rect 8690 -15567 8724 -15543
rect 8690 -15639 8724 -15611
rect 8690 -15711 8724 -15679
rect 8690 -15781 8724 -15747
rect 8690 -15849 8724 -15817
rect 8690 -15917 8724 -15889
rect 8690 -15985 8724 -15961
rect 8690 -16068 8724 -16033
rect 9708 -15495 9742 -15460
rect 9708 -15567 9742 -15543
rect 9708 -15639 9742 -15611
rect 9708 -15711 9742 -15679
rect 9708 -15781 9742 -15747
rect 9708 -15849 9742 -15817
rect 9708 -15917 9742 -15889
rect 9708 -15985 9742 -15961
rect 9708 -16068 9742 -16033
rect 10726 -15495 10760 -15460
rect 10726 -15567 10760 -15543
rect 10726 -15639 10760 -15611
rect 10726 -15711 10760 -15679
rect 10726 -15781 10760 -15747
rect 10726 -15849 10760 -15817
rect 10726 -15917 10760 -15889
rect 10726 -15985 10760 -15961
rect 10726 -16068 10760 -16033
rect 11744 -15495 11778 -15460
rect 11744 -15567 11778 -15543
rect 11744 -15639 11778 -15611
rect 11744 -15711 11778 -15679
rect 11744 -15781 11778 -15747
rect 11744 -15849 11778 -15817
rect 11744 -15917 11778 -15889
rect 11744 -15985 11778 -15961
rect 11744 -16068 11778 -16033
rect 12762 -15495 12796 -15460
rect 12762 -15567 12796 -15543
rect 12762 -15639 12796 -15611
rect 12762 -15711 12796 -15679
rect 12762 -15781 12796 -15747
rect 12762 -15849 12796 -15817
rect 12762 -15917 12796 -15889
rect 12762 -15985 12796 -15961
rect 12762 -16068 12796 -16033
rect 13780 -15495 13814 -15460
rect 13780 -15567 13814 -15543
rect 13780 -15639 13814 -15611
rect 13780 -15711 13814 -15679
rect 13780 -15781 13814 -15747
rect 13780 -15849 13814 -15817
rect 13780 -15917 13814 -15889
rect 13780 -15985 13814 -15961
rect 13780 -16068 13814 -16033
rect 14798 -15495 14832 -15460
rect 14798 -15567 14832 -15543
rect 14798 -15639 14832 -15611
rect 14798 -15711 14832 -15679
rect 14798 -15781 14832 -15747
rect 14798 -15849 14832 -15817
rect 14798 -15917 14832 -15889
rect 14798 -15985 14832 -15961
rect 14798 -16068 14832 -16033
rect 15816 -15495 15850 -15460
rect 15816 -15567 15850 -15543
rect 15816 -15639 15850 -15611
rect 15816 -15711 15850 -15679
rect 15816 -15781 15850 -15747
rect 15816 -15849 15850 -15817
rect 15816 -15917 15850 -15889
rect 15816 -15985 15850 -15961
rect 15816 -16068 15850 -16033
rect 16834 -15495 16868 -15460
rect 16834 -15567 16868 -15543
rect 16834 -15639 16868 -15611
rect 16834 -15711 16868 -15679
rect 16834 -15781 16868 -15747
rect 16834 -15849 16868 -15817
rect 16834 -15917 16868 -15889
rect 16834 -15985 16868 -15961
rect 16834 -16068 16868 -16033
rect 17852 -15495 17886 -15460
rect 17852 -15567 17886 -15543
rect 17852 -15639 17886 -15611
rect 17852 -15711 17886 -15679
rect 17852 -15781 17886 -15747
rect 17852 -15849 17886 -15817
rect 17852 -15917 17886 -15889
rect 17852 -15985 17886 -15961
rect 17852 -16068 17886 -16033
rect 18870 -15495 18904 -15460
rect 18870 -15567 18904 -15543
rect 18870 -15639 18904 -15611
rect 18870 -15711 18904 -15679
rect 18870 -15781 18904 -15747
rect 18870 -15849 18904 -15817
rect 18870 -15917 18904 -15889
rect 18870 -15985 18904 -15961
rect 18870 -16068 18904 -16033
rect 19888 -15495 19922 -15460
rect 19888 -15567 19922 -15543
rect 19888 -15639 19922 -15611
rect 19888 -15711 19922 -15679
rect 19888 -15781 19922 -15747
rect 19888 -15849 19922 -15817
rect 19888 -15917 19922 -15889
rect 19888 -15985 19922 -15961
rect 19888 -16068 19922 -16033
rect 20906 -15495 20940 -15460
rect 20906 -15567 20940 -15543
rect 20906 -15639 20940 -15611
rect 20906 -15711 20940 -15679
rect 20906 -15781 20940 -15747
rect 20906 -15849 20940 -15817
rect 20906 -15917 20940 -15889
rect 20906 -15985 20940 -15961
rect 20906 -16068 20940 -16033
rect 21924 -15495 21958 -15460
rect 21924 -15567 21958 -15543
rect 21924 -15639 21958 -15611
rect 21924 -15711 21958 -15679
rect 21924 -15781 21958 -15747
rect 21924 -15849 21958 -15817
rect 21924 -15917 21958 -15889
rect 21924 -15985 21958 -15961
rect 21924 -16068 21958 -16033
rect 22942 -15495 22976 -15460
rect 22942 -15567 22976 -15543
rect 22942 -15639 22976 -15611
rect 22942 -15711 22976 -15679
rect 22942 -15781 22976 -15747
rect 22942 -15849 22976 -15817
rect 22942 -15917 22976 -15889
rect 22942 -15985 22976 -15961
rect 24822 -15509 24855 -15443
rect 24889 -15509 24922 -15443
rect 24822 -15511 24922 -15509
rect 24822 -15545 24855 -15511
rect 24889 -15545 24922 -15511
rect 24822 -15547 24922 -15545
rect 24822 -15613 24855 -15547
rect 24889 -15613 24922 -15547
rect 24822 -15619 24922 -15613
rect 24822 -15681 24855 -15619
rect 24889 -15681 24922 -15619
rect 24822 -15691 24922 -15681
rect 24822 -15749 24855 -15691
rect 24889 -15749 24922 -15691
rect 24822 -15763 24922 -15749
rect 24822 -15817 24855 -15763
rect 24889 -15817 24922 -15763
rect 24822 -15835 24922 -15817
rect 24822 -15885 24855 -15835
rect 24889 -15885 24922 -15835
rect 24822 -15907 24922 -15885
rect 24822 -15953 24855 -15907
rect 24889 -15953 24922 -15907
rect 24822 -15979 24922 -15953
rect 22976 -16033 22982 -16004
rect 22942 -16052 22982 -16033
rect 24822 -16021 24855 -15979
rect 24889 -16021 24922 -15979
rect 24822 -16051 24922 -16021
rect 22942 -16068 22976 -16052
rect 24822 -16089 24855 -16051
rect 24889 -16089 24922 -16051
rect 6126 -16102 6186 -16100
rect 2814 -16136 2853 -16102
rect 2887 -16136 2911 -16102
rect 2955 -16136 2983 -16102
rect 3023 -16136 3055 -16102
rect 3091 -16136 3125 -16102
rect 3161 -16136 3193 -16102
rect 3233 -16136 3261 -16102
rect 3305 -16136 3329 -16102
rect 3363 -16136 3402 -16102
rect 3832 -16136 3871 -16102
rect 3905 -16136 3929 -16102
rect 3973 -16136 4001 -16102
rect 4041 -16136 4073 -16102
rect 4109 -16136 4143 -16102
rect 4179 -16136 4211 -16102
rect 4251 -16136 4279 -16102
rect 4323 -16136 4347 -16102
rect 4381 -16136 4420 -16102
rect 4850 -16136 4889 -16102
rect 4923 -16136 4947 -16102
rect 4991 -16136 5019 -16102
rect 5059 -16136 5091 -16102
rect 5127 -16136 5161 -16102
rect 5197 -16136 5229 -16102
rect 5269 -16136 5297 -16102
rect 5341 -16136 5365 -16102
rect 5399 -16136 5438 -16102
rect 5868 -16136 5907 -16102
rect 5941 -16136 5965 -16102
rect 6009 -16136 6037 -16102
rect 6077 -16136 6109 -16102
rect 6145 -16136 6179 -16102
rect 6215 -16136 6247 -16102
rect 6287 -16136 6315 -16102
rect 6359 -16136 6383 -16102
rect 6417 -16136 6456 -16102
rect 6886 -16136 6925 -16102
rect 6959 -16136 6983 -16102
rect 7027 -16136 7055 -16102
rect 7095 -16136 7127 -16102
rect 7163 -16136 7197 -16102
rect 7233 -16136 7265 -16102
rect 7305 -16136 7333 -16102
rect 7377 -16136 7401 -16102
rect 7435 -16136 7474 -16102
rect 7904 -16136 7943 -16102
rect 7977 -16136 8001 -16102
rect 8045 -16136 8073 -16102
rect 8113 -16136 8145 -16102
rect 8181 -16136 8215 -16102
rect 8251 -16136 8283 -16102
rect 8323 -16136 8351 -16102
rect 8395 -16136 8419 -16102
rect 8453 -16136 8492 -16102
rect 8922 -16136 8961 -16102
rect 8995 -16136 9019 -16102
rect 9063 -16136 9091 -16102
rect 9131 -16136 9163 -16102
rect 9199 -16136 9233 -16102
rect 9269 -16136 9301 -16102
rect 9341 -16136 9369 -16102
rect 9413 -16136 9437 -16102
rect 9471 -16136 9510 -16102
rect 9940 -16136 9979 -16102
rect 10013 -16136 10037 -16102
rect 10081 -16136 10109 -16102
rect 10149 -16136 10181 -16102
rect 10217 -16136 10251 -16102
rect 10287 -16136 10319 -16102
rect 10359 -16136 10387 -16102
rect 10431 -16136 10455 -16102
rect 10489 -16136 10528 -16102
rect 10958 -16136 10997 -16102
rect 11031 -16136 11055 -16102
rect 11099 -16136 11127 -16102
rect 11167 -16136 11199 -16102
rect 11235 -16136 11269 -16102
rect 11305 -16136 11337 -16102
rect 11377 -16136 11405 -16102
rect 11449 -16136 11473 -16102
rect 11507 -16136 11546 -16102
rect 11976 -16136 12015 -16102
rect 12049 -16136 12073 -16102
rect 12117 -16136 12145 -16102
rect 12185 -16136 12217 -16102
rect 12253 -16136 12287 -16102
rect 12323 -16136 12355 -16102
rect 12395 -16136 12423 -16102
rect 12467 -16136 12491 -16102
rect 12525 -16136 12564 -16102
rect 12994 -16136 13033 -16102
rect 13067 -16136 13091 -16102
rect 13135 -16136 13163 -16102
rect 13203 -16136 13235 -16102
rect 13271 -16136 13305 -16102
rect 13341 -16136 13373 -16102
rect 13413 -16136 13441 -16102
rect 13485 -16136 13509 -16102
rect 13543 -16136 13582 -16102
rect 14012 -16136 14051 -16102
rect 14085 -16136 14109 -16102
rect 14153 -16136 14181 -16102
rect 14221 -16136 14253 -16102
rect 14289 -16136 14323 -16102
rect 14359 -16136 14391 -16102
rect 14431 -16136 14459 -16102
rect 14503 -16136 14527 -16102
rect 14561 -16136 14600 -16102
rect 15030 -16136 15069 -16102
rect 15103 -16136 15127 -16102
rect 15171 -16136 15199 -16102
rect 15239 -16136 15271 -16102
rect 15307 -16136 15341 -16102
rect 15377 -16136 15409 -16102
rect 15449 -16136 15477 -16102
rect 15521 -16136 15545 -16102
rect 15579 -16136 15618 -16102
rect 16048 -16136 16087 -16102
rect 16121 -16136 16145 -16102
rect 16189 -16136 16217 -16102
rect 16257 -16136 16289 -16102
rect 16325 -16136 16359 -16102
rect 16395 -16136 16427 -16102
rect 16467 -16136 16495 -16102
rect 16539 -16136 16563 -16102
rect 16597 -16136 16636 -16102
rect 17066 -16136 17105 -16102
rect 17139 -16136 17163 -16102
rect 17207 -16136 17235 -16102
rect 17275 -16136 17309 -16102
rect 17343 -16136 17377 -16102
rect 17413 -16136 17445 -16102
rect 17485 -16136 17513 -16102
rect 17557 -16136 17581 -16102
rect 17615 -16136 17654 -16102
rect 18084 -16136 18123 -16102
rect 18157 -16136 18181 -16102
rect 18225 -16136 18253 -16102
rect 18293 -16136 18327 -16102
rect 18361 -16136 18395 -16102
rect 18429 -16136 18463 -16102
rect 18503 -16136 18531 -16102
rect 18575 -16136 18599 -16102
rect 18633 -16136 18672 -16102
rect 19102 -16136 19141 -16102
rect 19175 -16136 19199 -16102
rect 19243 -16136 19271 -16102
rect 19311 -16136 19343 -16102
rect 19379 -16136 19413 -16102
rect 19449 -16136 19481 -16102
rect 19521 -16136 19549 -16102
rect 19593 -16136 19617 -16102
rect 19651 -16136 19690 -16102
rect 20120 -16136 20159 -16102
rect 20193 -16136 20217 -16102
rect 20261 -16136 20289 -16102
rect 20329 -16136 20361 -16102
rect 20397 -16136 20431 -16102
rect 20467 -16136 20499 -16102
rect 20539 -16136 20567 -16102
rect 20611 -16136 20635 -16102
rect 20669 -16136 20708 -16102
rect 21138 -16136 21177 -16102
rect 21211 -16136 21235 -16102
rect 21279 -16136 21307 -16102
rect 21347 -16136 21379 -16102
rect 21415 -16136 21449 -16102
rect 21485 -16136 21517 -16102
rect 21557 -16136 21585 -16102
rect 21629 -16136 21653 -16102
rect 21687 -16136 21726 -16102
rect 22156 -16136 22195 -16102
rect 22229 -16136 22253 -16102
rect 22297 -16136 22325 -16102
rect 22365 -16136 22397 -16102
rect 22433 -16136 22467 -16102
rect 22503 -16136 22535 -16102
rect 22575 -16136 22603 -16102
rect 22647 -16136 22671 -16102
rect 22705 -16136 22744 -16102
rect 24822 -16123 24922 -16089
rect -22 -16169 12 -16137
rect 8160 -16140 8220 -16136
rect 17318 -16150 17378 -16136
rect 18352 -16150 18412 -16136
rect -22 -16237 12 -16209
rect -22 -16305 12 -16281
rect -22 -16388 12 -16353
rect 24822 -16157 24855 -16123
rect 24889 -16157 24922 -16123
rect 24822 -16191 24922 -16157
rect 24822 -16229 24855 -16191
rect 24889 -16229 24922 -16191
rect 24822 -16259 24922 -16229
rect 24822 -16301 24855 -16259
rect 24889 -16301 24922 -16259
rect 24822 -16327 24922 -16301
rect 24822 -16373 24855 -16327
rect 24889 -16373 24922 -16327
rect -12322 -16445 -12289 -16395
rect -12255 -16445 -12222 -16395
rect 24822 -16395 24922 -16373
rect -7670 -16422 -7610 -16420
rect -6656 -16422 -6596 -16420
rect -2582 -16422 -2522 -16420
rect -1566 -16422 -1506 -16420
rect -12322 -16463 -12222 -16445
rect -8952 -16456 -8913 -16422
rect -8879 -16456 -8855 -16422
rect -8811 -16456 -8783 -16422
rect -8743 -16456 -8711 -16422
rect -8675 -16456 -8641 -16422
rect -8605 -16456 -8573 -16422
rect -8533 -16456 -8505 -16422
rect -8461 -16456 -8437 -16422
rect -8403 -16456 -8364 -16422
rect -7934 -16456 -7895 -16422
rect -7861 -16456 -7837 -16422
rect -7793 -16456 -7765 -16422
rect -7725 -16456 -7693 -16422
rect -7657 -16456 -7623 -16422
rect -7587 -16456 -7555 -16422
rect -7515 -16456 -7487 -16422
rect -7443 -16456 -7419 -16422
rect -7385 -16456 -7346 -16422
rect -6916 -16456 -6877 -16422
rect -6843 -16456 -6819 -16422
rect -6775 -16456 -6747 -16422
rect -6707 -16456 -6675 -16422
rect -6639 -16456 -6605 -16422
rect -6569 -16456 -6537 -16422
rect -6497 -16456 -6469 -16422
rect -6425 -16456 -6401 -16422
rect -6367 -16456 -6328 -16422
rect -5898 -16456 -5859 -16422
rect -5825 -16456 -5801 -16422
rect -5757 -16456 -5729 -16422
rect -5689 -16456 -5657 -16422
rect -5621 -16456 -5587 -16422
rect -5551 -16456 -5519 -16422
rect -5479 -16456 -5451 -16422
rect -5407 -16456 -5383 -16422
rect -5349 -16456 -5310 -16422
rect -4880 -16456 -4841 -16422
rect -4807 -16456 -4783 -16422
rect -4739 -16456 -4711 -16422
rect -4671 -16456 -4639 -16422
rect -4603 -16456 -4569 -16422
rect -4533 -16456 -4501 -16422
rect -4461 -16456 -4433 -16422
rect -4389 -16456 -4365 -16422
rect -4331 -16456 -4292 -16422
rect -3862 -16456 -3823 -16422
rect -3789 -16456 -3765 -16422
rect -3721 -16456 -3693 -16422
rect -3653 -16456 -3621 -16422
rect -3585 -16456 -3551 -16422
rect -3515 -16456 -3483 -16422
rect -3443 -16456 -3415 -16422
rect -3371 -16456 -3347 -16422
rect -3313 -16456 -3274 -16422
rect -2844 -16456 -2805 -16422
rect -2771 -16456 -2747 -16422
rect -2703 -16456 -2675 -16422
rect -2635 -16456 -2603 -16422
rect -2567 -16456 -2533 -16422
rect -2497 -16456 -2465 -16422
rect -2425 -16456 -2397 -16422
rect -2353 -16456 -2329 -16422
rect -2295 -16456 -2256 -16422
rect -1826 -16456 -1787 -16422
rect -1753 -16456 -1729 -16422
rect -1685 -16456 -1657 -16422
rect -1617 -16456 -1585 -16422
rect -1549 -16456 -1515 -16422
rect -1479 -16456 -1447 -16422
rect -1407 -16456 -1379 -16422
rect -1335 -16456 -1311 -16422
rect -1277 -16456 -1238 -16422
rect -808 -16456 -769 -16422
rect -735 -16456 -711 -16422
rect -667 -16456 -639 -16422
rect -599 -16456 -567 -16422
rect -531 -16456 -497 -16422
rect -461 -16456 -429 -16422
rect -389 -16456 -361 -16422
rect -317 -16456 -293 -16422
rect -259 -16456 -220 -16422
rect 24822 -16445 24855 -16395
rect 24889 -16445 24922 -16395
rect -12322 -16517 -12289 -16463
rect -12255 -16517 -12222 -16463
rect -12322 -16531 -12222 -16517
rect 24822 -16463 24922 -16445
rect 24822 -16517 24855 -16463
rect 24889 -16517 24922 -16463
rect -12322 -16589 -12289 -16531
rect -12255 -16589 -12222 -16531
rect -8952 -16564 -8913 -16530
rect -8879 -16564 -8855 -16530
rect -8811 -16564 -8783 -16530
rect -8743 -16564 -8711 -16530
rect -8675 -16564 -8641 -16530
rect -8605 -16564 -8573 -16530
rect -8533 -16564 -8505 -16530
rect -8461 -16564 -8437 -16530
rect -8403 -16564 -8364 -16530
rect -7934 -16564 -7895 -16530
rect -7861 -16564 -7837 -16530
rect -7793 -16564 -7765 -16530
rect -7725 -16564 -7693 -16530
rect -7657 -16564 -7623 -16530
rect -7587 -16564 -7555 -16530
rect -7515 -16564 -7487 -16530
rect -7443 -16564 -7419 -16530
rect -7385 -16564 -7346 -16530
rect -6916 -16564 -6877 -16530
rect -6843 -16564 -6819 -16530
rect -6775 -16564 -6747 -16530
rect -6707 -16564 -6675 -16530
rect -6639 -16564 -6605 -16530
rect -6569 -16564 -6537 -16530
rect -6497 -16564 -6469 -16530
rect -6425 -16564 -6401 -16530
rect -6367 -16564 -6328 -16530
rect -5898 -16564 -5859 -16530
rect -5825 -16564 -5801 -16530
rect -5757 -16564 -5729 -16530
rect -5689 -16564 -5657 -16530
rect -5621 -16564 -5587 -16530
rect -5551 -16564 -5519 -16530
rect -5479 -16564 -5451 -16530
rect -5407 -16564 -5383 -16530
rect -5349 -16564 -5310 -16530
rect -4880 -16564 -4841 -16530
rect -4807 -16564 -4783 -16530
rect -4739 -16564 -4711 -16530
rect -4671 -16564 -4639 -16530
rect -4603 -16564 -4569 -16530
rect -4533 -16564 -4501 -16530
rect -4461 -16564 -4433 -16530
rect -4389 -16564 -4365 -16530
rect -4331 -16564 -4292 -16530
rect -3862 -16564 -3823 -16530
rect -3789 -16564 -3765 -16530
rect -3721 -16564 -3693 -16530
rect -3653 -16564 -3621 -16530
rect -3585 -16564 -3551 -16530
rect -3515 -16564 -3483 -16530
rect -3443 -16564 -3415 -16530
rect -3371 -16564 -3347 -16530
rect -3313 -16564 -3274 -16530
rect -2844 -16564 -2805 -16530
rect -2771 -16564 -2747 -16530
rect -2703 -16564 -2675 -16530
rect -2635 -16564 -2603 -16530
rect -2567 -16564 -2533 -16530
rect -2497 -16564 -2465 -16530
rect -2425 -16564 -2397 -16530
rect -2353 -16564 -2329 -16530
rect -2295 -16564 -2256 -16530
rect -1826 -16564 -1787 -16530
rect -1753 -16564 -1729 -16530
rect -1685 -16564 -1657 -16530
rect -1617 -16564 -1585 -16530
rect -1549 -16564 -1515 -16530
rect -1479 -16564 -1447 -16530
rect -1407 -16564 -1379 -16530
rect -1335 -16564 -1311 -16530
rect -1277 -16564 -1238 -16530
rect -808 -16564 -769 -16530
rect -735 -16564 -711 -16530
rect -667 -16564 -639 -16530
rect -599 -16564 -567 -16530
rect -531 -16564 -497 -16530
rect -461 -16564 -429 -16530
rect -389 -16564 -361 -16530
rect -317 -16564 -293 -16530
rect -259 -16564 -220 -16530
rect 24822 -16531 24922 -16517
rect -12322 -16599 -12222 -16589
rect 24822 -16589 24855 -16531
rect 24889 -16589 24922 -16531
rect -12322 -16661 -12289 -16599
rect -12255 -16661 -12222 -16599
rect -12322 -16667 -12222 -16661
rect -12322 -16733 -12289 -16667
rect -12255 -16733 -12222 -16667
rect -12322 -16735 -12222 -16733
rect -12322 -16769 -12289 -16735
rect -12255 -16769 -12222 -16735
rect -12322 -16771 -12222 -16769
rect -12322 -16837 -12289 -16771
rect -12255 -16837 -12222 -16771
rect -12322 -16843 -12222 -16837
rect -12322 -16905 -12289 -16843
rect -12255 -16905 -12222 -16843
rect -12322 -16915 -12222 -16905
rect -12322 -16973 -12289 -16915
rect -12255 -16973 -12222 -16915
rect -12322 -16987 -12222 -16973
rect -12322 -17041 -12289 -16987
rect -12255 -17041 -12222 -16987
rect -12322 -17059 -12222 -17041
rect -12322 -17109 -12289 -17059
rect -12255 -17109 -12222 -17059
rect -12322 -17131 -12222 -17109
rect -12322 -17177 -12289 -17131
rect -12255 -17177 -12222 -17131
rect -12322 -17203 -12222 -17177
rect -12322 -17245 -12289 -17203
rect -12255 -17245 -12222 -17203
rect -9184 -16633 -9150 -16598
rect -9184 -16705 -9150 -16681
rect -9184 -16777 -9150 -16749
rect -9184 -16849 -9150 -16817
rect -9184 -16919 -9150 -16885
rect -9184 -16987 -9150 -16955
rect -9184 -17055 -9150 -17027
rect -9184 -17123 -9150 -17099
rect -9184 -17206 -9150 -17171
rect -8166 -16633 -8132 -16598
rect -8166 -16705 -8132 -16681
rect -8166 -16777 -8132 -16749
rect -8166 -16849 -8132 -16817
rect -8166 -16919 -8132 -16885
rect -8166 -16987 -8132 -16955
rect -8166 -17055 -8132 -17027
rect -8166 -17123 -8132 -17099
rect -8166 -17206 -8132 -17171
rect -7148 -16633 -7114 -16598
rect -7148 -16705 -7114 -16681
rect -7148 -16777 -7114 -16749
rect -7148 -16849 -7114 -16817
rect -7148 -16919 -7114 -16885
rect -7148 -16987 -7114 -16955
rect -7148 -17055 -7114 -17027
rect -7148 -17123 -7114 -17099
rect -7148 -17206 -7114 -17171
rect -6130 -16633 -6096 -16598
rect -6130 -16705 -6096 -16681
rect -6130 -16777 -6096 -16749
rect -6130 -16849 -6096 -16817
rect -6130 -16919 -6096 -16885
rect -6130 -16987 -6096 -16955
rect -6130 -17055 -6096 -17027
rect -6130 -17123 -6096 -17099
rect -6130 -17206 -6096 -17171
rect -5112 -16633 -5078 -16598
rect -5112 -16705 -5078 -16681
rect -5112 -16777 -5078 -16749
rect -5112 -16849 -5078 -16817
rect -5112 -16919 -5078 -16885
rect -5112 -16987 -5078 -16955
rect -5112 -17055 -5078 -17027
rect -5112 -17123 -5078 -17099
rect -5112 -17206 -5078 -17171
rect -4094 -16633 -4060 -16598
rect -4094 -16705 -4060 -16681
rect -4094 -16777 -4060 -16749
rect -4094 -16849 -4060 -16817
rect -4094 -16919 -4060 -16885
rect -4094 -16987 -4060 -16955
rect -4094 -17055 -4060 -17027
rect -4094 -17123 -4060 -17099
rect -4094 -17206 -4060 -17171
rect -3076 -16633 -3042 -16598
rect -3076 -16705 -3042 -16681
rect -3076 -16777 -3042 -16749
rect -3076 -16849 -3042 -16817
rect -3076 -16919 -3042 -16885
rect -3076 -16987 -3042 -16955
rect -3076 -17055 -3042 -17027
rect -3076 -17123 -3042 -17099
rect -3076 -17206 -3042 -17171
rect -2058 -16633 -2024 -16598
rect -2058 -16705 -2024 -16681
rect -2058 -16777 -2024 -16749
rect -2058 -16849 -2024 -16817
rect -2058 -16919 -2024 -16885
rect -2058 -16987 -2024 -16955
rect -2058 -17055 -2024 -17027
rect -2058 -17123 -2024 -17099
rect -2058 -17206 -2024 -17171
rect -1040 -16633 -1006 -16598
rect -1040 -16705 -1006 -16681
rect -1040 -16777 -1006 -16749
rect -1040 -16849 -1006 -16817
rect -1040 -16919 -1006 -16885
rect -1040 -16987 -1006 -16955
rect -1040 -17055 -1006 -17027
rect -1040 -17123 -1006 -17099
rect -1040 -17206 -1006 -17171
rect -22 -16633 12 -16598
rect 24822 -16599 24922 -16589
rect 2812 -16660 2851 -16626
rect 2885 -16660 2909 -16626
rect 2953 -16660 2981 -16626
rect 3021 -16660 3053 -16626
rect 3089 -16660 3123 -16626
rect 3159 -16660 3191 -16626
rect 3231 -16660 3259 -16626
rect 3303 -16660 3327 -16626
rect 3361 -16660 3400 -16626
rect 3830 -16660 3869 -16626
rect 3903 -16660 3927 -16626
rect 3971 -16660 3999 -16626
rect 4039 -16660 4071 -16626
rect 4107 -16660 4141 -16626
rect 4177 -16660 4209 -16626
rect 4249 -16660 4277 -16626
rect 4321 -16660 4345 -16626
rect 4379 -16660 4418 -16626
rect 4848 -16660 4887 -16626
rect 4921 -16660 4945 -16626
rect 4989 -16660 5017 -16626
rect 5057 -16660 5089 -16626
rect 5125 -16660 5159 -16626
rect 5195 -16660 5227 -16626
rect 5267 -16660 5295 -16626
rect 5339 -16660 5363 -16626
rect 5397 -16660 5436 -16626
rect 5866 -16660 5905 -16626
rect 5939 -16660 5963 -16626
rect 6007 -16660 6035 -16626
rect 6075 -16660 6107 -16626
rect 6143 -16660 6177 -16626
rect 6213 -16660 6245 -16626
rect 6285 -16660 6313 -16626
rect 6357 -16660 6381 -16626
rect 6415 -16660 6454 -16626
rect 6884 -16660 6923 -16626
rect 6957 -16660 6981 -16626
rect 7025 -16660 7053 -16626
rect 7093 -16660 7125 -16626
rect 7161 -16660 7195 -16626
rect 7231 -16660 7263 -16626
rect 7303 -16660 7331 -16626
rect 7375 -16660 7399 -16626
rect 7433 -16660 7472 -16626
rect 7902 -16660 7941 -16626
rect 7975 -16660 7999 -16626
rect 8043 -16660 8071 -16626
rect 8111 -16660 8143 -16626
rect 8179 -16660 8213 -16626
rect 8249 -16660 8281 -16626
rect 8321 -16660 8349 -16626
rect 8393 -16660 8417 -16626
rect 8451 -16660 8490 -16626
rect 8920 -16660 8959 -16626
rect 8993 -16660 9017 -16626
rect 9061 -16660 9089 -16626
rect 9129 -16660 9161 -16626
rect 9197 -16660 9231 -16626
rect 9267 -16660 9299 -16626
rect 9339 -16660 9367 -16626
rect 9411 -16660 9435 -16626
rect 9469 -16660 9508 -16626
rect 9938 -16660 9977 -16626
rect 10011 -16660 10035 -16626
rect 10079 -16660 10107 -16626
rect 10147 -16660 10179 -16626
rect 10215 -16660 10249 -16626
rect 10285 -16660 10317 -16626
rect 10357 -16660 10385 -16626
rect 10429 -16660 10453 -16626
rect 10487 -16660 10526 -16626
rect 10956 -16660 10995 -16626
rect 11029 -16660 11053 -16626
rect 11097 -16660 11125 -16626
rect 11165 -16660 11197 -16626
rect 11233 -16660 11267 -16626
rect 11303 -16660 11335 -16626
rect 11375 -16660 11403 -16626
rect 11447 -16660 11471 -16626
rect 11505 -16660 11544 -16626
rect 11974 -16660 12013 -16626
rect 12047 -16660 12071 -16626
rect 12115 -16660 12143 -16626
rect 12183 -16660 12215 -16626
rect 12251 -16660 12285 -16626
rect 12321 -16660 12353 -16626
rect 12393 -16660 12421 -16626
rect 12465 -16660 12489 -16626
rect 12523 -16660 12562 -16626
rect 12992 -16660 13031 -16626
rect 13065 -16660 13089 -16626
rect 13133 -16660 13161 -16626
rect 13201 -16660 13233 -16626
rect 13269 -16660 13303 -16626
rect 13339 -16660 13371 -16626
rect 13411 -16660 13439 -16626
rect 13483 -16660 13507 -16626
rect 13541 -16660 13580 -16626
rect 14010 -16660 14049 -16626
rect 14083 -16660 14107 -16626
rect 14151 -16660 14179 -16626
rect 14219 -16660 14251 -16626
rect 14287 -16660 14321 -16626
rect 14357 -16660 14389 -16626
rect 14429 -16660 14457 -16626
rect 14501 -16660 14525 -16626
rect 14559 -16660 14598 -16626
rect 15028 -16660 15067 -16626
rect 15101 -16660 15125 -16626
rect 15169 -16660 15197 -16626
rect 15237 -16660 15269 -16626
rect 15305 -16660 15339 -16626
rect 15375 -16660 15407 -16626
rect 15447 -16660 15475 -16626
rect 15519 -16660 15543 -16626
rect 15577 -16660 15616 -16626
rect 16046 -16660 16085 -16626
rect 16119 -16660 16143 -16626
rect 16187 -16660 16215 -16626
rect 16255 -16660 16287 -16626
rect 16323 -16660 16357 -16626
rect 16393 -16660 16425 -16626
rect 16465 -16660 16493 -16626
rect 16537 -16660 16561 -16626
rect 16595 -16660 16634 -16626
rect 17064 -16660 17103 -16626
rect 17137 -16660 17161 -16626
rect 17205 -16660 17233 -16626
rect 17273 -16660 17305 -16626
rect 17341 -16660 17375 -16626
rect 17411 -16660 17443 -16626
rect 17483 -16660 17511 -16626
rect 17555 -16660 17579 -16626
rect 17613 -16660 17652 -16626
rect 18082 -16660 18121 -16626
rect 18155 -16660 18179 -16626
rect 18223 -16660 18251 -16626
rect 18291 -16660 18323 -16626
rect 18359 -16660 18393 -16626
rect 18429 -16660 18461 -16626
rect 18501 -16660 18529 -16626
rect 18573 -16660 18597 -16626
rect 18631 -16660 18670 -16626
rect 19100 -16660 19139 -16626
rect 19173 -16660 19197 -16626
rect 19241 -16660 19269 -16626
rect 19309 -16660 19341 -16626
rect 19377 -16660 19411 -16626
rect 19447 -16660 19479 -16626
rect 19519 -16660 19547 -16626
rect 19591 -16660 19615 -16626
rect 19649 -16660 19688 -16626
rect 20118 -16660 20157 -16626
rect 20191 -16660 20215 -16626
rect 20259 -16660 20287 -16626
rect 20327 -16660 20359 -16626
rect 20395 -16660 20429 -16626
rect 20465 -16660 20497 -16626
rect 20537 -16660 20565 -16626
rect 20609 -16660 20633 -16626
rect 20667 -16660 20706 -16626
rect 21136 -16660 21175 -16626
rect 21209 -16660 21233 -16626
rect 21277 -16660 21305 -16626
rect 21345 -16660 21377 -16626
rect 21413 -16660 21447 -16626
rect 21483 -16660 21515 -16626
rect 21555 -16660 21583 -16626
rect 21627 -16660 21651 -16626
rect 21685 -16660 21724 -16626
rect 22154 -16660 22193 -16626
rect 22227 -16660 22251 -16626
rect 22295 -16660 22323 -16626
rect 22363 -16660 22395 -16626
rect 22431 -16660 22465 -16626
rect 22501 -16660 22533 -16626
rect 22573 -16660 22601 -16626
rect 22645 -16660 22669 -16626
rect 22703 -16660 22742 -16626
rect 5122 -16664 5182 -16660
rect 24822 -16661 24855 -16599
rect 24889 -16661 24922 -16599
rect -22 -16705 12 -16681
rect 24822 -16667 24922 -16661
rect -22 -16777 12 -16749
rect -22 -16849 12 -16817
rect -22 -16919 12 -16885
rect -22 -16987 12 -16955
rect -22 -17055 12 -17027
rect -22 -17123 12 -17099
rect -22 -17206 12 -17171
rect 2580 -16729 2614 -16694
rect 2580 -16801 2614 -16777
rect 2580 -16873 2614 -16845
rect 2580 -16945 2614 -16913
rect 2580 -17015 2614 -16981
rect 2580 -17083 2614 -17051
rect 2580 -17151 2614 -17123
rect 2580 -17219 2614 -17195
rect -7666 -17240 -7606 -17238
rect -6652 -17240 -6592 -17238
rect -2578 -17240 -2518 -17238
rect -1562 -17240 -1502 -17238
rect -12322 -17275 -12222 -17245
rect -8952 -17274 -8913 -17240
rect -8879 -17274 -8855 -17240
rect -8811 -17274 -8783 -17240
rect -8743 -17274 -8711 -17240
rect -8675 -17274 -8641 -17240
rect -8605 -17274 -8573 -17240
rect -8533 -17274 -8505 -17240
rect -8461 -17274 -8437 -17240
rect -8403 -17274 -8364 -17240
rect -7934 -17274 -7895 -17240
rect -7861 -17274 -7837 -17240
rect -7793 -17274 -7765 -17240
rect -7725 -17274 -7693 -17240
rect -7657 -17274 -7623 -17240
rect -7587 -17274 -7555 -17240
rect -7515 -17274 -7487 -17240
rect -7443 -17274 -7419 -17240
rect -7385 -17274 -7346 -17240
rect -6916 -17274 -6877 -17240
rect -6843 -17274 -6819 -17240
rect -6775 -17274 -6747 -17240
rect -6707 -17274 -6675 -17240
rect -6639 -17274 -6605 -17240
rect -6569 -17274 -6537 -17240
rect -6497 -17274 -6469 -17240
rect -6425 -17274 -6401 -17240
rect -6367 -17274 -6328 -17240
rect -5898 -17274 -5859 -17240
rect -5825 -17274 -5801 -17240
rect -5757 -17274 -5729 -17240
rect -5689 -17274 -5657 -17240
rect -5621 -17274 -5587 -17240
rect -5551 -17274 -5519 -17240
rect -5479 -17274 -5451 -17240
rect -5407 -17274 -5383 -17240
rect -5349 -17274 -5310 -17240
rect -4880 -17274 -4841 -17240
rect -4807 -17274 -4783 -17240
rect -4739 -17274 -4711 -17240
rect -4671 -17274 -4639 -17240
rect -4603 -17274 -4569 -17240
rect -4533 -17274 -4501 -17240
rect -4461 -17274 -4433 -17240
rect -4389 -17274 -4365 -17240
rect -4331 -17274 -4292 -17240
rect -3862 -17274 -3823 -17240
rect -3789 -17274 -3765 -17240
rect -3721 -17274 -3693 -17240
rect -3653 -17274 -3621 -17240
rect -3585 -17274 -3551 -17240
rect -3515 -17274 -3483 -17240
rect -3443 -17274 -3415 -17240
rect -3371 -17274 -3347 -17240
rect -3313 -17274 -3274 -17240
rect -2844 -17274 -2805 -17240
rect -2771 -17274 -2747 -17240
rect -2703 -17274 -2675 -17240
rect -2635 -17274 -2603 -17240
rect -2567 -17274 -2533 -17240
rect -2497 -17274 -2465 -17240
rect -2425 -17274 -2397 -17240
rect -2353 -17274 -2329 -17240
rect -2295 -17274 -2256 -17240
rect -1826 -17274 -1787 -17240
rect -1753 -17274 -1729 -17240
rect -1685 -17274 -1657 -17240
rect -1617 -17274 -1585 -17240
rect -1549 -17274 -1515 -17240
rect -1479 -17274 -1447 -17240
rect -1407 -17274 -1379 -17240
rect -1335 -17274 -1311 -17240
rect -1277 -17274 -1238 -17240
rect -808 -17274 -769 -17240
rect -735 -17274 -711 -17240
rect -667 -17274 -639 -17240
rect -599 -17274 -567 -17240
rect -531 -17274 -497 -17240
rect -461 -17274 -429 -17240
rect -389 -17274 -361 -17240
rect -317 -17274 -293 -17240
rect -259 -17274 -220 -17240
rect -12322 -17313 -12289 -17275
rect -12255 -17313 -12222 -17275
rect 2580 -17302 2614 -17267
rect 3598 -16729 3632 -16694
rect 3598 -16801 3632 -16777
rect 3598 -16873 3632 -16845
rect 3598 -16945 3632 -16913
rect 3598 -17015 3632 -16981
rect 3598 -17083 3632 -17051
rect 3598 -17151 3632 -17123
rect 3598 -17219 3632 -17195
rect 3598 -17302 3632 -17267
rect 4616 -16729 4650 -16694
rect 4616 -16801 4650 -16777
rect 4616 -16873 4650 -16845
rect 4616 -16945 4650 -16913
rect 4616 -17015 4650 -16981
rect 4616 -17083 4650 -17051
rect 4616 -17151 4650 -17123
rect 4616 -17219 4650 -17195
rect 4616 -17302 4650 -17267
rect 5634 -16729 5668 -16694
rect 5634 -16801 5668 -16777
rect 5634 -16873 5668 -16845
rect 5634 -16945 5668 -16913
rect 5634 -17015 5668 -16981
rect 5634 -17083 5668 -17051
rect 5634 -17151 5668 -17123
rect 5634 -17219 5668 -17195
rect 5634 -17302 5668 -17267
rect 6652 -16729 6686 -16694
rect 6652 -16801 6686 -16777
rect 6652 -16873 6686 -16845
rect 6652 -16945 6686 -16913
rect 6652 -17015 6686 -16981
rect 6652 -17083 6686 -17051
rect 6652 -17151 6686 -17123
rect 6652 -17219 6686 -17195
rect 6652 -17302 6686 -17267
rect 7670 -16729 7704 -16694
rect 7670 -16801 7704 -16777
rect 7670 -16873 7704 -16845
rect 7670 -16945 7704 -16913
rect 7670 -17015 7704 -16981
rect 7670 -17083 7704 -17051
rect 7670 -17151 7704 -17123
rect 7670 -17219 7704 -17195
rect 7670 -17302 7704 -17267
rect 8688 -16729 8722 -16694
rect 8688 -16801 8722 -16777
rect 8688 -16873 8722 -16845
rect 8688 -16945 8722 -16913
rect 8688 -17015 8722 -16981
rect 8688 -17083 8722 -17051
rect 8688 -17151 8722 -17123
rect 8688 -17219 8722 -17195
rect 8688 -17302 8722 -17267
rect 9706 -16729 9740 -16694
rect 9706 -16801 9740 -16777
rect 9706 -16873 9740 -16845
rect 9706 -16945 9740 -16913
rect 9706 -17015 9740 -16981
rect 9706 -17083 9740 -17051
rect 9706 -17151 9740 -17123
rect 9706 -17219 9740 -17195
rect 9706 -17302 9740 -17267
rect 10724 -16729 10758 -16694
rect 10724 -16801 10758 -16777
rect 10724 -16873 10758 -16845
rect 10724 -16945 10758 -16913
rect 10724 -17015 10758 -16981
rect 10724 -17083 10758 -17051
rect 10724 -17151 10758 -17123
rect 10724 -17219 10758 -17195
rect 10724 -17302 10758 -17267
rect 11742 -16729 11776 -16694
rect 11742 -16801 11776 -16777
rect 11742 -16873 11776 -16845
rect 11742 -16945 11776 -16913
rect 11742 -17015 11776 -16981
rect 11742 -17083 11776 -17051
rect 11742 -17151 11776 -17123
rect 11742 -17219 11776 -17195
rect 11742 -17302 11776 -17267
rect 12760 -16729 12794 -16694
rect 12760 -16801 12794 -16777
rect 12760 -16873 12794 -16845
rect 12760 -16945 12794 -16913
rect 12760 -17015 12794 -16981
rect 12760 -17083 12794 -17051
rect 12760 -17151 12794 -17123
rect 12760 -17219 12794 -17195
rect 12760 -17302 12794 -17267
rect 13778 -16729 13812 -16694
rect 13778 -16801 13812 -16777
rect 13778 -16873 13812 -16845
rect 13778 -16945 13812 -16913
rect 13778 -17015 13812 -16981
rect 13778 -17083 13812 -17051
rect 13778 -17151 13812 -17123
rect 13778 -17219 13812 -17195
rect 13778 -17302 13812 -17267
rect 14796 -16729 14830 -16694
rect 14796 -16801 14830 -16777
rect 14796 -16873 14830 -16845
rect 14796 -16945 14830 -16913
rect 14796 -17015 14830 -16981
rect 14796 -17083 14830 -17051
rect 14796 -17151 14830 -17123
rect 14796 -17219 14830 -17195
rect 14796 -17302 14830 -17267
rect 15814 -16729 15848 -16694
rect 15814 -16801 15848 -16777
rect 15814 -16873 15848 -16845
rect 15814 -16945 15848 -16913
rect 15814 -17015 15848 -16981
rect 15814 -17083 15848 -17051
rect 15814 -17151 15848 -17123
rect 15814 -17219 15848 -17195
rect 15814 -17302 15848 -17267
rect 16832 -16729 16866 -16694
rect 16832 -16801 16866 -16777
rect 16832 -16873 16866 -16845
rect 16832 -16945 16866 -16913
rect 16832 -17015 16866 -16981
rect 16832 -17083 16866 -17051
rect 16832 -17151 16866 -17123
rect 16832 -17219 16866 -17195
rect 16832 -17302 16866 -17267
rect 17850 -16729 17884 -16694
rect 17850 -16801 17884 -16777
rect 17850 -16873 17884 -16845
rect 17850 -16945 17884 -16913
rect 17850 -17015 17884 -16981
rect 17850 -17083 17884 -17051
rect 17850 -17151 17884 -17123
rect 17850 -17219 17884 -17195
rect 17850 -17302 17884 -17267
rect 18868 -16729 18902 -16694
rect 18868 -16801 18902 -16777
rect 18868 -16873 18902 -16845
rect 18868 -16945 18902 -16913
rect 18868 -17015 18902 -16981
rect 18868 -17083 18902 -17051
rect 18868 -17151 18902 -17123
rect 18868 -17219 18902 -17195
rect 18868 -17302 18902 -17267
rect 19886 -16729 19920 -16694
rect 19886 -16801 19920 -16777
rect 19886 -16873 19920 -16845
rect 19886 -16945 19920 -16913
rect 19886 -17015 19920 -16981
rect 19886 -17083 19920 -17051
rect 19886 -17151 19920 -17123
rect 19886 -17219 19920 -17195
rect 19886 -17302 19920 -17267
rect 20904 -16729 20938 -16694
rect 20904 -16801 20938 -16777
rect 20904 -16873 20938 -16845
rect 20904 -16945 20938 -16913
rect 20904 -17015 20938 -16981
rect 20904 -17083 20938 -17051
rect 20904 -17151 20938 -17123
rect 20904 -17219 20938 -17195
rect 20904 -17302 20938 -17267
rect 21922 -16729 21956 -16694
rect 21922 -16801 21956 -16777
rect 21922 -16873 21956 -16845
rect 21922 -16945 21956 -16913
rect 21922 -17015 21956 -16981
rect 21922 -17083 21956 -17051
rect 21922 -17151 21956 -17123
rect 21922 -17219 21956 -17195
rect 21922 -17302 21956 -17267
rect 22940 -16729 22974 -16694
rect 22940 -16801 22974 -16777
rect 22940 -16873 22974 -16845
rect 22940 -16945 22974 -16913
rect 22940 -17015 22974 -16981
rect 22940 -17083 22974 -17051
rect 22940 -17151 22974 -17123
rect 22940 -17219 22974 -17195
rect 22940 -17302 22974 -17267
rect 24822 -16733 24855 -16667
rect 24889 -16733 24922 -16667
rect 24822 -16735 24922 -16733
rect 24822 -16769 24855 -16735
rect 24889 -16769 24922 -16735
rect 24822 -16771 24922 -16769
rect 24822 -16837 24855 -16771
rect 24889 -16837 24922 -16771
rect 24822 -16843 24922 -16837
rect 24822 -16905 24855 -16843
rect 24889 -16905 24922 -16843
rect 24822 -16915 24922 -16905
rect 24822 -16973 24855 -16915
rect 24889 -16973 24922 -16915
rect 24822 -16987 24922 -16973
rect 24822 -17041 24855 -16987
rect 24889 -17041 24922 -16987
rect 24822 -17059 24922 -17041
rect 24822 -17109 24855 -17059
rect 24889 -17109 24922 -17059
rect 24822 -17131 24922 -17109
rect 24822 -17177 24855 -17131
rect 24889 -17177 24922 -17131
rect 24822 -17203 24922 -17177
rect 24822 -17245 24855 -17203
rect 24889 -17245 24922 -17203
rect 24822 -17275 24922 -17245
rect -12322 -17347 -12222 -17313
rect 24822 -17313 24855 -17275
rect 24889 -17313 24922 -17275
rect 10190 -17336 10250 -17332
rect 11218 -17336 11278 -17334
rect 13262 -17336 13322 -17332
rect -12322 -17381 -12289 -17347
rect -12255 -17381 -12222 -17347
rect -12322 -17415 -12222 -17381
rect -8952 -17382 -8913 -17348
rect -8879 -17382 -8855 -17348
rect -8811 -17382 -8783 -17348
rect -8743 -17382 -8711 -17348
rect -8675 -17382 -8641 -17348
rect -8605 -17382 -8573 -17348
rect -8533 -17382 -8505 -17348
rect -8461 -17382 -8437 -17348
rect -8403 -17382 -8364 -17348
rect -7934 -17382 -7895 -17348
rect -7861 -17382 -7837 -17348
rect -7793 -17382 -7765 -17348
rect -7725 -17382 -7693 -17348
rect -7657 -17382 -7623 -17348
rect -7587 -17382 -7555 -17348
rect -7515 -17382 -7487 -17348
rect -7443 -17382 -7419 -17348
rect -7385 -17382 -7346 -17348
rect -6916 -17382 -6877 -17348
rect -6843 -17382 -6819 -17348
rect -6775 -17382 -6747 -17348
rect -6707 -17382 -6675 -17348
rect -6639 -17382 -6605 -17348
rect -6569 -17382 -6537 -17348
rect -6497 -17382 -6469 -17348
rect -6425 -17382 -6401 -17348
rect -6367 -17382 -6328 -17348
rect -5898 -17382 -5859 -17348
rect -5825 -17382 -5801 -17348
rect -5757 -17382 -5729 -17348
rect -5689 -17382 -5657 -17348
rect -5621 -17382 -5587 -17348
rect -5551 -17382 -5519 -17348
rect -5479 -17382 -5451 -17348
rect -5407 -17382 -5383 -17348
rect -5349 -17382 -5310 -17348
rect -4880 -17382 -4841 -17348
rect -4807 -17382 -4783 -17348
rect -4739 -17382 -4711 -17348
rect -4671 -17382 -4639 -17348
rect -4603 -17382 -4569 -17348
rect -4533 -17382 -4501 -17348
rect -4461 -17382 -4433 -17348
rect -4389 -17382 -4365 -17348
rect -4331 -17382 -4292 -17348
rect -3862 -17382 -3823 -17348
rect -3789 -17382 -3765 -17348
rect -3721 -17382 -3693 -17348
rect -3653 -17382 -3621 -17348
rect -3585 -17382 -3551 -17348
rect -3515 -17382 -3483 -17348
rect -3443 -17382 -3415 -17348
rect -3371 -17382 -3347 -17348
rect -3313 -17382 -3274 -17348
rect -2844 -17382 -2805 -17348
rect -2771 -17382 -2747 -17348
rect -2703 -17382 -2675 -17348
rect -2635 -17382 -2603 -17348
rect -2567 -17382 -2533 -17348
rect -2497 -17382 -2465 -17348
rect -2425 -17382 -2397 -17348
rect -2353 -17382 -2329 -17348
rect -2295 -17382 -2256 -17348
rect -1826 -17382 -1787 -17348
rect -1753 -17382 -1729 -17348
rect -1685 -17382 -1657 -17348
rect -1617 -17382 -1585 -17348
rect -1549 -17382 -1515 -17348
rect -1479 -17382 -1447 -17348
rect -1407 -17382 -1379 -17348
rect -1335 -17382 -1311 -17348
rect -1277 -17382 -1238 -17348
rect -808 -17382 -769 -17348
rect -735 -17382 -711 -17348
rect -667 -17382 -639 -17348
rect -599 -17382 -567 -17348
rect -531 -17382 -497 -17348
rect -461 -17382 -429 -17348
rect -389 -17382 -361 -17348
rect -317 -17382 -293 -17348
rect -259 -17382 -220 -17348
rect 2812 -17370 2851 -17336
rect 2885 -17370 2909 -17336
rect 2953 -17370 2981 -17336
rect 3021 -17370 3053 -17336
rect 3089 -17370 3123 -17336
rect 3159 -17370 3191 -17336
rect 3231 -17370 3259 -17336
rect 3303 -17370 3327 -17336
rect 3361 -17370 3400 -17336
rect 3830 -17370 3869 -17336
rect 3903 -17370 3927 -17336
rect 3971 -17370 3999 -17336
rect 4039 -17370 4071 -17336
rect 4107 -17370 4141 -17336
rect 4177 -17370 4209 -17336
rect 4249 -17370 4277 -17336
rect 4321 -17370 4345 -17336
rect 4379 -17370 4418 -17336
rect 4848 -17370 4887 -17336
rect 4921 -17370 4945 -17336
rect 4989 -17370 5017 -17336
rect 5057 -17370 5089 -17336
rect 5125 -17370 5159 -17336
rect 5195 -17370 5227 -17336
rect 5267 -17370 5295 -17336
rect 5339 -17370 5363 -17336
rect 5397 -17370 5436 -17336
rect 5866 -17370 5905 -17336
rect 5939 -17370 5963 -17336
rect 6007 -17370 6035 -17336
rect 6075 -17370 6107 -17336
rect 6143 -17370 6177 -17336
rect 6213 -17370 6245 -17336
rect 6285 -17370 6313 -17336
rect 6357 -17370 6381 -17336
rect 6415 -17370 6454 -17336
rect 6884 -17370 6923 -17336
rect 6957 -17370 6981 -17336
rect 7025 -17370 7053 -17336
rect 7093 -17370 7125 -17336
rect 7161 -17370 7195 -17336
rect 7231 -17370 7263 -17336
rect 7303 -17370 7331 -17336
rect 7375 -17370 7399 -17336
rect 7433 -17370 7472 -17336
rect 7902 -17370 7941 -17336
rect 7975 -17370 7999 -17336
rect 8043 -17370 8071 -17336
rect 8111 -17370 8143 -17336
rect 8179 -17370 8213 -17336
rect 8249 -17370 8281 -17336
rect 8321 -17370 8349 -17336
rect 8393 -17370 8417 -17336
rect 8451 -17370 8490 -17336
rect 8920 -17370 8959 -17336
rect 8993 -17370 9017 -17336
rect 9061 -17370 9089 -17336
rect 9129 -17370 9161 -17336
rect 9197 -17370 9231 -17336
rect 9267 -17370 9299 -17336
rect 9339 -17370 9367 -17336
rect 9411 -17370 9435 -17336
rect 9469 -17370 9508 -17336
rect 9938 -17370 9977 -17336
rect 10011 -17370 10035 -17336
rect 10079 -17370 10107 -17336
rect 10147 -17370 10179 -17336
rect 10215 -17370 10249 -17336
rect 10285 -17370 10317 -17336
rect 10357 -17370 10385 -17336
rect 10429 -17370 10453 -17336
rect 10487 -17370 10526 -17336
rect 10956 -17370 10995 -17336
rect 11029 -17370 11053 -17336
rect 11097 -17370 11125 -17336
rect 11165 -17370 11197 -17336
rect 11233 -17370 11267 -17336
rect 11303 -17370 11335 -17336
rect 11375 -17370 11403 -17336
rect 11447 -17370 11471 -17336
rect 11505 -17370 11544 -17336
rect 11974 -17370 12013 -17336
rect 12047 -17370 12071 -17336
rect 12115 -17370 12143 -17336
rect 12183 -17370 12215 -17336
rect 12251 -17370 12285 -17336
rect 12321 -17370 12353 -17336
rect 12393 -17370 12421 -17336
rect 12465 -17370 12489 -17336
rect 12523 -17370 12562 -17336
rect 12992 -17370 13031 -17336
rect 13065 -17370 13089 -17336
rect 13133 -17370 13161 -17336
rect 13201 -17370 13233 -17336
rect 13269 -17370 13303 -17336
rect 13339 -17370 13371 -17336
rect 13411 -17370 13439 -17336
rect 13483 -17370 13507 -17336
rect 13541 -17370 13580 -17336
rect 14010 -17370 14049 -17336
rect 14083 -17370 14107 -17336
rect 14151 -17370 14179 -17336
rect 14219 -17370 14251 -17336
rect 14287 -17370 14321 -17336
rect 14357 -17370 14389 -17336
rect 14429 -17370 14457 -17336
rect 14501 -17370 14525 -17336
rect 14559 -17370 14598 -17336
rect 15028 -17370 15067 -17336
rect 15101 -17370 15125 -17336
rect 15169 -17370 15197 -17336
rect 15237 -17370 15269 -17336
rect 15305 -17370 15339 -17336
rect 15375 -17370 15407 -17336
rect 15447 -17370 15475 -17336
rect 15519 -17370 15543 -17336
rect 15577 -17370 15616 -17336
rect 16046 -17370 16085 -17336
rect 16119 -17370 16143 -17336
rect 16187 -17370 16215 -17336
rect 16255 -17370 16287 -17336
rect 16323 -17370 16357 -17336
rect 16393 -17370 16425 -17336
rect 16465 -17370 16493 -17336
rect 16537 -17370 16561 -17336
rect 16595 -17370 16634 -17336
rect 17064 -17370 17103 -17336
rect 17137 -17370 17161 -17336
rect 17205 -17370 17233 -17336
rect 17273 -17370 17305 -17336
rect 17341 -17370 17375 -17336
rect 17411 -17370 17443 -17336
rect 17483 -17370 17511 -17336
rect 17555 -17370 17579 -17336
rect 17613 -17370 17652 -17336
rect 18082 -17370 18121 -17336
rect 18155 -17370 18179 -17336
rect 18223 -17370 18251 -17336
rect 18291 -17370 18323 -17336
rect 18359 -17370 18393 -17336
rect 18429 -17370 18461 -17336
rect 18501 -17370 18529 -17336
rect 18573 -17370 18597 -17336
rect 18631 -17370 18670 -17336
rect 19100 -17370 19139 -17336
rect 19173 -17370 19197 -17336
rect 19241 -17370 19269 -17336
rect 19309 -17370 19341 -17336
rect 19377 -17370 19411 -17336
rect 19447 -17370 19479 -17336
rect 19519 -17370 19547 -17336
rect 19591 -17370 19615 -17336
rect 19649 -17370 19688 -17336
rect 20118 -17370 20157 -17336
rect 20191 -17370 20215 -17336
rect 20259 -17370 20287 -17336
rect 20327 -17370 20359 -17336
rect 20395 -17370 20429 -17336
rect 20465 -17370 20497 -17336
rect 20537 -17370 20565 -17336
rect 20609 -17370 20633 -17336
rect 20667 -17370 20706 -17336
rect 21136 -17370 21175 -17336
rect 21209 -17370 21233 -17336
rect 21277 -17370 21305 -17336
rect 21345 -17370 21377 -17336
rect 21413 -17370 21447 -17336
rect 21483 -17370 21515 -17336
rect 21555 -17370 21583 -17336
rect 21627 -17370 21651 -17336
rect 21685 -17370 21724 -17336
rect 22154 -17370 22193 -17336
rect 22227 -17370 22251 -17336
rect 22295 -17370 22323 -17336
rect 22363 -17370 22395 -17336
rect 22431 -17370 22465 -17336
rect 22501 -17370 22533 -17336
rect 22573 -17370 22601 -17336
rect 22645 -17370 22669 -17336
rect 22703 -17370 22742 -17336
rect 24822 -17347 24922 -17313
rect 24822 -17381 24855 -17347
rect 24889 -17381 24922 -17347
rect -12322 -17453 -12289 -17415
rect -12255 -17453 -12222 -17415
rect 24822 -17415 24922 -17381
rect -12322 -17483 -12222 -17453
rect -12322 -17525 -12289 -17483
rect -12255 -17525 -12222 -17483
rect -12322 -17551 -12222 -17525
rect -12322 -17597 -12289 -17551
rect -12255 -17597 -12222 -17551
rect -12322 -17619 -12222 -17597
rect -12322 -17669 -12289 -17619
rect -12255 -17669 -12222 -17619
rect -12322 -17687 -12222 -17669
rect -12322 -17741 -12289 -17687
rect -12255 -17741 -12222 -17687
rect -12322 -17755 -12222 -17741
rect -12322 -17813 -12289 -17755
rect -12255 -17813 -12222 -17755
rect -12322 -17823 -12222 -17813
rect -12322 -17885 -12289 -17823
rect -12255 -17885 -12222 -17823
rect -12322 -17891 -12222 -17885
rect -12322 -17957 -12289 -17891
rect -12255 -17957 -12222 -17891
rect -12322 -17959 -12222 -17957
rect -12322 -17993 -12289 -17959
rect -12255 -17993 -12222 -17959
rect -12322 -17995 -12222 -17993
rect -12322 -18061 -12289 -17995
rect -12255 -18061 -12222 -17995
rect -9184 -17451 -9150 -17416
rect -9184 -17523 -9150 -17499
rect -9184 -17595 -9150 -17567
rect -9184 -17667 -9150 -17635
rect -9184 -17737 -9150 -17703
rect -9184 -17805 -9150 -17773
rect -9184 -17873 -9150 -17845
rect -9184 -17941 -9150 -17917
rect -9184 -18024 -9150 -17989
rect -8166 -17451 -8132 -17416
rect -8166 -17523 -8132 -17499
rect -8166 -17595 -8132 -17567
rect -8166 -17667 -8132 -17635
rect -8166 -17737 -8132 -17703
rect -8166 -17805 -8132 -17773
rect -8166 -17873 -8132 -17845
rect -8166 -17941 -8132 -17917
rect -8166 -18024 -8132 -17989
rect -7148 -17451 -7114 -17416
rect -7148 -17523 -7114 -17499
rect -7148 -17595 -7114 -17567
rect -7148 -17667 -7114 -17635
rect -7148 -17737 -7114 -17703
rect -7148 -17805 -7114 -17773
rect -7148 -17873 -7114 -17845
rect -7148 -17941 -7114 -17917
rect -7148 -18024 -7114 -17989
rect -6130 -17451 -6096 -17416
rect -6130 -17523 -6096 -17499
rect -6130 -17595 -6096 -17567
rect -6130 -17667 -6096 -17635
rect -6130 -17737 -6096 -17703
rect -6130 -17805 -6096 -17773
rect -6130 -17873 -6096 -17845
rect -6130 -17941 -6096 -17917
rect -6130 -18024 -6096 -17989
rect -5112 -17451 -5078 -17416
rect -5112 -17523 -5078 -17499
rect -5112 -17595 -5078 -17567
rect -5112 -17667 -5078 -17635
rect -5112 -17737 -5078 -17703
rect -5112 -17805 -5078 -17773
rect -5112 -17873 -5078 -17845
rect -5112 -17941 -5078 -17917
rect -5112 -18024 -5078 -17989
rect -4094 -17451 -4060 -17416
rect -4094 -17523 -4060 -17499
rect -4094 -17595 -4060 -17567
rect -4094 -17667 -4060 -17635
rect -4094 -17737 -4060 -17703
rect -4094 -17805 -4060 -17773
rect -4094 -17873 -4060 -17845
rect -4094 -17941 -4060 -17917
rect -4094 -18024 -4060 -17989
rect -3076 -17451 -3042 -17416
rect -3076 -17523 -3042 -17499
rect -3076 -17595 -3042 -17567
rect -3076 -17667 -3042 -17635
rect -3076 -17737 -3042 -17703
rect -3076 -17805 -3042 -17773
rect -3076 -17873 -3042 -17845
rect -3076 -17941 -3042 -17917
rect -3076 -18024 -3042 -17989
rect -2058 -17451 -2024 -17416
rect -2058 -17523 -2024 -17499
rect -2058 -17595 -2024 -17567
rect -2058 -17667 -2024 -17635
rect -2058 -17737 -2024 -17703
rect -2058 -17805 -2024 -17773
rect -2058 -17873 -2024 -17845
rect -2058 -17941 -2024 -17917
rect -2058 -18024 -2024 -17989
rect -1040 -17451 -1006 -17416
rect -1040 -17523 -1006 -17499
rect -1040 -17595 -1006 -17567
rect -1040 -17667 -1006 -17635
rect -1040 -17737 -1006 -17703
rect -1040 -17805 -1006 -17773
rect -1040 -17873 -1006 -17845
rect -1040 -17941 -1006 -17917
rect -1040 -18024 -1006 -17989
rect -22 -17451 12 -17416
rect -22 -17523 12 -17499
rect -22 -17595 12 -17567
rect -22 -17667 12 -17635
rect -22 -17737 12 -17703
rect -22 -17805 12 -17773
rect -22 -17873 12 -17845
rect 24822 -17453 24855 -17415
rect 24889 -17453 24922 -17415
rect 24822 -17483 24922 -17453
rect 24822 -17525 24855 -17483
rect 24889 -17525 24922 -17483
rect 24822 -17551 24922 -17525
rect 24822 -17597 24855 -17551
rect 24889 -17597 24922 -17551
rect 24822 -17619 24922 -17597
rect 24822 -17669 24855 -17619
rect 24889 -17669 24922 -17619
rect 24822 -17687 24922 -17669
rect 24822 -17741 24855 -17687
rect 24889 -17741 24922 -17687
rect 24822 -17755 24922 -17741
rect 24822 -17813 24855 -17755
rect 24889 -17813 24922 -17755
rect 24822 -17823 24922 -17813
rect 2812 -17894 2851 -17860
rect 2885 -17894 2909 -17860
rect 2953 -17894 2981 -17860
rect 3021 -17894 3053 -17860
rect 3089 -17894 3123 -17860
rect 3159 -17894 3191 -17860
rect 3231 -17894 3259 -17860
rect 3303 -17894 3327 -17860
rect 3361 -17894 3400 -17860
rect 3830 -17894 3869 -17860
rect 3903 -17894 3927 -17860
rect 3971 -17894 3999 -17860
rect 4039 -17894 4071 -17860
rect 4107 -17894 4141 -17860
rect 4177 -17894 4209 -17860
rect 4249 -17894 4277 -17860
rect 4321 -17894 4345 -17860
rect 4379 -17894 4418 -17860
rect 4848 -17894 4887 -17860
rect 4921 -17894 4945 -17860
rect 4989 -17894 5017 -17860
rect 5057 -17894 5089 -17860
rect 5125 -17894 5159 -17860
rect 5195 -17894 5227 -17860
rect 5267 -17894 5295 -17860
rect 5339 -17894 5363 -17860
rect 5397 -17894 5436 -17860
rect 5866 -17894 5905 -17860
rect 5939 -17894 5963 -17860
rect 6007 -17894 6035 -17860
rect 6075 -17894 6107 -17860
rect 6143 -17894 6177 -17860
rect 6213 -17894 6245 -17860
rect 6285 -17894 6313 -17860
rect 6357 -17894 6381 -17860
rect 6415 -17894 6454 -17860
rect 6884 -17894 6923 -17860
rect 6957 -17894 6981 -17860
rect 7025 -17894 7053 -17860
rect 7093 -17894 7125 -17860
rect 7161 -17894 7195 -17860
rect 7231 -17894 7263 -17860
rect 7303 -17894 7331 -17860
rect 7375 -17894 7399 -17860
rect 7433 -17894 7472 -17860
rect 7902 -17894 7941 -17860
rect 7975 -17894 7999 -17860
rect 8043 -17894 8071 -17860
rect 8111 -17894 8143 -17860
rect 8179 -17894 8213 -17860
rect 8249 -17894 8281 -17860
rect 8321 -17894 8349 -17860
rect 8393 -17894 8417 -17860
rect 8451 -17894 8490 -17860
rect 8920 -17894 8959 -17860
rect 8993 -17894 9017 -17860
rect 9061 -17894 9089 -17860
rect 9129 -17894 9161 -17860
rect 9197 -17894 9231 -17860
rect 9267 -17894 9299 -17860
rect 9339 -17894 9367 -17860
rect 9411 -17894 9435 -17860
rect 9469 -17894 9508 -17860
rect 9938 -17894 9977 -17860
rect 10011 -17894 10035 -17860
rect 10079 -17894 10107 -17860
rect 10147 -17894 10179 -17860
rect 10215 -17894 10249 -17860
rect 10285 -17894 10317 -17860
rect 10357 -17894 10385 -17860
rect 10429 -17894 10453 -17860
rect 10487 -17894 10526 -17860
rect 10956 -17894 10995 -17860
rect 11029 -17894 11053 -17860
rect 11097 -17894 11125 -17860
rect 11165 -17894 11197 -17860
rect 11233 -17894 11267 -17860
rect 11303 -17894 11335 -17860
rect 11375 -17894 11403 -17860
rect 11447 -17894 11471 -17860
rect 11505 -17894 11544 -17860
rect 11974 -17894 12013 -17860
rect 12047 -17894 12071 -17860
rect 12115 -17894 12143 -17860
rect 12183 -17894 12215 -17860
rect 12251 -17894 12285 -17860
rect 12321 -17894 12353 -17860
rect 12393 -17894 12421 -17860
rect 12465 -17894 12489 -17860
rect 12523 -17894 12562 -17860
rect 12992 -17894 13031 -17860
rect 13065 -17894 13089 -17860
rect 13133 -17894 13161 -17860
rect 13201 -17894 13233 -17860
rect 13269 -17894 13303 -17860
rect 13339 -17894 13371 -17860
rect 13411 -17894 13439 -17860
rect 13483 -17894 13507 -17860
rect 13541 -17894 13580 -17860
rect 14010 -17894 14049 -17860
rect 14083 -17894 14107 -17860
rect 14151 -17894 14179 -17860
rect 14219 -17894 14251 -17860
rect 14287 -17894 14321 -17860
rect 14357 -17894 14389 -17860
rect 14429 -17894 14457 -17860
rect 14501 -17894 14525 -17860
rect 14559 -17894 14598 -17860
rect 15028 -17894 15067 -17860
rect 15101 -17894 15125 -17860
rect 15169 -17894 15197 -17860
rect 15237 -17894 15269 -17860
rect 15305 -17894 15339 -17860
rect 15375 -17894 15407 -17860
rect 15447 -17894 15475 -17860
rect 15519 -17894 15543 -17860
rect 15577 -17894 15616 -17860
rect 16046 -17894 16085 -17860
rect 16119 -17894 16143 -17860
rect 16187 -17894 16215 -17860
rect 16255 -17894 16287 -17860
rect 16323 -17894 16357 -17860
rect 16393 -17894 16425 -17860
rect 16465 -17894 16493 -17860
rect 16537 -17894 16561 -17860
rect 16595 -17894 16634 -17860
rect 17064 -17894 17103 -17860
rect 17137 -17894 17161 -17860
rect 17205 -17894 17233 -17860
rect 17273 -17894 17305 -17860
rect 17341 -17894 17375 -17860
rect 17411 -17894 17443 -17860
rect 17483 -17894 17511 -17860
rect 17555 -17894 17579 -17860
rect 17613 -17894 17652 -17860
rect 18082 -17894 18121 -17860
rect 18155 -17894 18179 -17860
rect 18223 -17894 18251 -17860
rect 18291 -17894 18323 -17860
rect 18359 -17894 18393 -17860
rect 18429 -17894 18461 -17860
rect 18501 -17894 18529 -17860
rect 18573 -17894 18597 -17860
rect 18631 -17894 18670 -17860
rect 19100 -17894 19139 -17860
rect 19173 -17894 19197 -17860
rect 19241 -17894 19269 -17860
rect 19309 -17894 19341 -17860
rect 19377 -17894 19411 -17860
rect 19447 -17894 19479 -17860
rect 19519 -17894 19547 -17860
rect 19591 -17894 19615 -17860
rect 19649 -17894 19688 -17860
rect 20118 -17894 20157 -17860
rect 20191 -17894 20215 -17860
rect 20259 -17894 20287 -17860
rect 20327 -17894 20359 -17860
rect 20395 -17894 20429 -17860
rect 20465 -17894 20497 -17860
rect 20537 -17894 20565 -17860
rect 20609 -17894 20633 -17860
rect 20667 -17894 20706 -17860
rect 21136 -17894 21175 -17860
rect 21209 -17894 21233 -17860
rect 21277 -17894 21305 -17860
rect 21345 -17894 21377 -17860
rect 21413 -17894 21447 -17860
rect 21483 -17894 21515 -17860
rect 21555 -17894 21583 -17860
rect 21627 -17894 21651 -17860
rect 21685 -17894 21724 -17860
rect 22154 -17894 22193 -17860
rect 22227 -17894 22251 -17860
rect 22295 -17894 22323 -17860
rect 22363 -17894 22395 -17860
rect 22431 -17894 22465 -17860
rect 22501 -17894 22533 -17860
rect 22573 -17894 22601 -17860
rect 22645 -17894 22669 -17860
rect 22703 -17894 22742 -17860
rect 24822 -17885 24855 -17823
rect 24889 -17885 24922 -17823
rect 24822 -17891 24922 -17885
rect -22 -17941 12 -17917
rect -22 -18024 12 -17989
rect 2580 -17963 2614 -17928
rect 2580 -18035 2614 -18011
rect -8692 -18058 -8632 -18056
rect -7666 -18058 -7606 -18054
rect -6652 -18058 -6592 -18054
rect -5632 -18058 -5572 -18056
rect -4610 -18058 -4550 -18056
rect -2578 -18058 -2518 -18054
rect -1562 -18058 -1502 -18054
rect -542 -18058 -482 -18056
rect -12322 -18067 -12222 -18061
rect -12322 -18129 -12289 -18067
rect -12255 -18129 -12222 -18067
rect -8952 -18092 -8913 -18058
rect -8879 -18092 -8855 -18058
rect -8811 -18092 -8783 -18058
rect -8743 -18092 -8711 -18058
rect -8675 -18092 -8641 -18058
rect -8605 -18092 -8573 -18058
rect -8533 -18092 -8505 -18058
rect -8461 -18092 -8437 -18058
rect -8403 -18092 -8364 -18058
rect -7934 -18092 -7895 -18058
rect -7861 -18092 -7837 -18058
rect -7793 -18092 -7765 -18058
rect -7725 -18092 -7693 -18058
rect -7657 -18092 -7623 -18058
rect -7587 -18092 -7555 -18058
rect -7515 -18092 -7487 -18058
rect -7443 -18092 -7419 -18058
rect -7385 -18092 -7346 -18058
rect -6916 -18092 -6877 -18058
rect -6843 -18092 -6819 -18058
rect -6775 -18092 -6747 -18058
rect -6707 -18092 -6675 -18058
rect -6639 -18092 -6605 -18058
rect -6569 -18092 -6537 -18058
rect -6497 -18092 -6469 -18058
rect -6425 -18092 -6401 -18058
rect -6367 -18092 -6328 -18058
rect -5898 -18092 -5859 -18058
rect -5825 -18092 -5801 -18058
rect -5757 -18092 -5729 -18058
rect -5689 -18092 -5657 -18058
rect -5621 -18092 -5587 -18058
rect -5551 -18092 -5519 -18058
rect -5479 -18092 -5451 -18058
rect -5407 -18092 -5383 -18058
rect -5349 -18092 -5310 -18058
rect -4880 -18092 -4841 -18058
rect -4807 -18092 -4783 -18058
rect -4739 -18092 -4711 -18058
rect -4671 -18092 -4639 -18058
rect -4603 -18092 -4569 -18058
rect -4533 -18092 -4501 -18058
rect -4461 -18092 -4433 -18058
rect -4389 -18092 -4365 -18058
rect -4331 -18092 -4292 -18058
rect -3862 -18092 -3823 -18058
rect -3789 -18092 -3765 -18058
rect -3721 -18092 -3693 -18058
rect -3653 -18092 -3621 -18058
rect -3585 -18092 -3551 -18058
rect -3515 -18092 -3483 -18058
rect -3443 -18092 -3415 -18058
rect -3371 -18092 -3347 -18058
rect -3313 -18092 -3274 -18058
rect -2844 -18092 -2805 -18058
rect -2771 -18092 -2747 -18058
rect -2703 -18092 -2675 -18058
rect -2635 -18092 -2603 -18058
rect -2567 -18092 -2533 -18058
rect -2497 -18092 -2465 -18058
rect -2425 -18092 -2397 -18058
rect -2353 -18092 -2329 -18058
rect -2295 -18092 -2256 -18058
rect -1826 -18092 -1787 -18058
rect -1753 -18092 -1729 -18058
rect -1685 -18092 -1657 -18058
rect -1617 -18092 -1585 -18058
rect -1549 -18092 -1515 -18058
rect -1479 -18092 -1447 -18058
rect -1407 -18092 -1379 -18058
rect -1335 -18092 -1311 -18058
rect -1277 -18092 -1238 -18058
rect -808 -18092 -769 -18058
rect -735 -18092 -711 -18058
rect -667 -18092 -639 -18058
rect -599 -18092 -567 -18058
rect -531 -18092 -497 -18058
rect -461 -18092 -429 -18058
rect -389 -18092 -361 -18058
rect -317 -18092 -293 -18058
rect -259 -18092 -220 -18058
rect -12322 -18139 -12222 -18129
rect -12322 -18197 -12289 -18139
rect -12255 -18197 -12222 -18139
rect 2580 -18107 2614 -18079
rect -12322 -18211 -12222 -18197
rect -8952 -18200 -8913 -18166
rect -8879 -18200 -8855 -18166
rect -8811 -18200 -8783 -18166
rect -8743 -18200 -8711 -18166
rect -8675 -18200 -8641 -18166
rect -8605 -18200 -8573 -18166
rect -8533 -18200 -8505 -18166
rect -8461 -18200 -8437 -18166
rect -8403 -18200 -8364 -18166
rect -7934 -18200 -7895 -18166
rect -7861 -18200 -7837 -18166
rect -7793 -18200 -7765 -18166
rect -7725 -18200 -7693 -18166
rect -7657 -18200 -7623 -18166
rect -7587 -18200 -7555 -18166
rect -7515 -18200 -7487 -18166
rect -7443 -18200 -7419 -18166
rect -7385 -18200 -7346 -18166
rect -6916 -18200 -6877 -18166
rect -6843 -18200 -6819 -18166
rect -6775 -18200 -6747 -18166
rect -6707 -18200 -6675 -18166
rect -6639 -18200 -6605 -18166
rect -6569 -18200 -6537 -18166
rect -6497 -18200 -6469 -18166
rect -6425 -18200 -6401 -18166
rect -6367 -18200 -6328 -18166
rect -5898 -18200 -5859 -18166
rect -5825 -18200 -5801 -18166
rect -5757 -18200 -5729 -18166
rect -5689 -18200 -5657 -18166
rect -5621 -18200 -5587 -18166
rect -5551 -18200 -5519 -18166
rect -5479 -18200 -5451 -18166
rect -5407 -18200 -5383 -18166
rect -5349 -18200 -5310 -18166
rect -4880 -18200 -4841 -18166
rect -4807 -18200 -4783 -18166
rect -4739 -18200 -4711 -18166
rect -4671 -18200 -4639 -18166
rect -4603 -18200 -4569 -18166
rect -4533 -18200 -4501 -18166
rect -4461 -18200 -4433 -18166
rect -4389 -18200 -4365 -18166
rect -4331 -18200 -4292 -18166
rect -3862 -18200 -3823 -18166
rect -3789 -18200 -3765 -18166
rect -3721 -18200 -3693 -18166
rect -3653 -18200 -3621 -18166
rect -3585 -18200 -3551 -18166
rect -3515 -18200 -3483 -18166
rect -3443 -18200 -3415 -18166
rect -3371 -18200 -3347 -18166
rect -3313 -18200 -3274 -18166
rect -2844 -18200 -2805 -18166
rect -2771 -18200 -2747 -18166
rect -2703 -18200 -2675 -18166
rect -2635 -18200 -2603 -18166
rect -2567 -18200 -2533 -18166
rect -2497 -18200 -2465 -18166
rect -2425 -18200 -2397 -18166
rect -2353 -18200 -2329 -18166
rect -2295 -18200 -2256 -18166
rect -1826 -18200 -1787 -18166
rect -1753 -18200 -1729 -18166
rect -1685 -18200 -1657 -18166
rect -1617 -18200 -1585 -18166
rect -1549 -18200 -1515 -18166
rect -1479 -18200 -1447 -18166
rect -1407 -18200 -1379 -18166
rect -1335 -18200 -1311 -18166
rect -1277 -18200 -1238 -18166
rect -808 -18200 -769 -18166
rect -735 -18200 -711 -18166
rect -667 -18200 -639 -18166
rect -599 -18200 -567 -18166
rect -531 -18200 -497 -18166
rect -461 -18200 -429 -18166
rect -389 -18200 -361 -18166
rect -317 -18200 -293 -18166
rect -259 -18200 -220 -18166
rect 2580 -18179 2614 -18147
rect -12322 -18265 -12289 -18211
rect -12255 -18265 -12222 -18211
rect -12322 -18283 -12222 -18265
rect -12322 -18333 -12289 -18283
rect -12255 -18333 -12222 -18283
rect -12322 -18355 -12222 -18333
rect -12322 -18401 -12289 -18355
rect -12255 -18401 -12222 -18355
rect -12322 -18427 -12222 -18401
rect -12322 -18469 -12289 -18427
rect -12255 -18469 -12222 -18427
rect -12322 -18499 -12222 -18469
rect -12322 -18537 -12289 -18499
rect -12255 -18537 -12222 -18499
rect -12322 -18571 -12222 -18537
rect -12322 -18605 -12289 -18571
rect -12255 -18605 -12222 -18571
rect -12322 -18639 -12222 -18605
rect -12322 -18677 -12289 -18639
rect -12255 -18677 -12222 -18639
rect -12322 -18707 -12222 -18677
rect -12322 -18749 -12289 -18707
rect -12255 -18749 -12222 -18707
rect -12322 -18775 -12222 -18749
rect -12322 -18821 -12289 -18775
rect -12255 -18821 -12222 -18775
rect -12322 -18843 -12222 -18821
rect -9184 -18269 -9150 -18234
rect -9184 -18341 -9150 -18317
rect -9184 -18413 -9150 -18385
rect -9184 -18485 -9150 -18453
rect -9184 -18555 -9150 -18521
rect -9184 -18623 -9150 -18591
rect -9184 -18691 -9150 -18663
rect -9184 -18759 -9150 -18735
rect -9184 -18842 -9150 -18807
rect -8166 -18269 -8132 -18234
rect -8166 -18341 -8132 -18317
rect -8166 -18413 -8132 -18385
rect -8166 -18485 -8132 -18453
rect -8166 -18555 -8132 -18521
rect -8166 -18623 -8132 -18591
rect -8166 -18691 -8132 -18663
rect -8166 -18759 -8132 -18735
rect -8166 -18842 -8132 -18807
rect -7148 -18269 -7114 -18234
rect -7148 -18341 -7114 -18317
rect -7148 -18413 -7114 -18385
rect -7148 -18485 -7114 -18453
rect -7148 -18555 -7114 -18521
rect -7148 -18623 -7114 -18591
rect -7148 -18691 -7114 -18663
rect -7148 -18759 -7114 -18735
rect -7148 -18842 -7114 -18807
rect -6130 -18269 -6096 -18234
rect -6130 -18341 -6096 -18317
rect -6130 -18413 -6096 -18385
rect -6130 -18485 -6096 -18453
rect -6130 -18555 -6096 -18521
rect -6130 -18623 -6096 -18591
rect -6130 -18691 -6096 -18663
rect -6130 -18759 -6096 -18735
rect -6130 -18842 -6096 -18807
rect -5112 -18269 -5078 -18234
rect -5112 -18341 -5078 -18317
rect -5112 -18413 -5078 -18385
rect -5112 -18485 -5078 -18453
rect -5112 -18555 -5078 -18521
rect -5112 -18623 -5078 -18591
rect -5112 -18691 -5078 -18663
rect -5112 -18759 -5078 -18735
rect -5112 -18842 -5078 -18807
rect -4094 -18269 -4060 -18234
rect -4094 -18341 -4060 -18317
rect -4094 -18413 -4060 -18385
rect -4094 -18485 -4060 -18453
rect -4094 -18555 -4060 -18521
rect -4094 -18623 -4060 -18591
rect -4094 -18691 -4060 -18663
rect -4094 -18759 -4060 -18735
rect -4094 -18842 -4060 -18807
rect -3076 -18269 -3042 -18234
rect -3076 -18341 -3042 -18317
rect -3076 -18413 -3042 -18385
rect -3076 -18485 -3042 -18453
rect -3076 -18555 -3042 -18521
rect -3076 -18623 -3042 -18591
rect -3076 -18691 -3042 -18663
rect -3076 -18759 -3042 -18735
rect -3076 -18842 -3042 -18807
rect -2058 -18269 -2024 -18234
rect -2058 -18341 -2024 -18317
rect -2058 -18413 -2024 -18385
rect -2058 -18485 -2024 -18453
rect -2058 -18555 -2024 -18521
rect -2058 -18623 -2024 -18591
rect -2058 -18691 -2024 -18663
rect -2058 -18759 -2024 -18735
rect -2058 -18842 -2024 -18807
rect -1040 -18269 -1006 -18234
rect -1040 -18341 -1006 -18317
rect -1040 -18413 -1006 -18385
rect -1040 -18485 -1006 -18453
rect -1040 -18555 -1006 -18521
rect -1040 -18623 -1006 -18591
rect -1040 -18691 -1006 -18663
rect -1040 -18759 -1006 -18735
rect -1040 -18842 -1006 -18807
rect -22 -18269 12 -18234
rect -22 -18341 12 -18317
rect -22 -18413 12 -18385
rect -22 -18485 12 -18453
rect -22 -18555 12 -18521
rect 2580 -18249 2614 -18215
rect 2580 -18317 2614 -18285
rect 2580 -18385 2614 -18357
rect 2580 -18453 2614 -18429
rect 2580 -18536 2614 -18501
rect 3598 -17963 3632 -17928
rect 3598 -18035 3632 -18011
rect 3598 -18107 3632 -18079
rect 3598 -18179 3632 -18147
rect 3598 -18249 3632 -18215
rect 3598 -18317 3632 -18285
rect 3598 -18385 3632 -18357
rect 3598 -18453 3632 -18429
rect 3598 -18536 3632 -18501
rect 4616 -17963 4650 -17928
rect 4616 -18035 4650 -18011
rect 4616 -18107 4650 -18079
rect 4616 -18179 4650 -18147
rect 4616 -18249 4650 -18215
rect 4616 -18317 4650 -18285
rect 4616 -18385 4650 -18357
rect 4616 -18453 4650 -18429
rect 4616 -18536 4650 -18501
rect 5634 -17963 5668 -17928
rect 5634 -18035 5668 -18011
rect 5634 -18107 5668 -18079
rect 5634 -18179 5668 -18147
rect 5634 -18249 5668 -18215
rect 5634 -18317 5668 -18285
rect 5634 -18385 5668 -18357
rect 5634 -18453 5668 -18429
rect 5634 -18536 5668 -18501
rect 6652 -17963 6686 -17928
rect 6652 -18035 6686 -18011
rect 6652 -18107 6686 -18079
rect 6652 -18179 6686 -18147
rect 6652 -18249 6686 -18215
rect 6652 -18317 6686 -18285
rect 6652 -18385 6686 -18357
rect 6652 -18453 6686 -18429
rect 6652 -18536 6686 -18501
rect 7670 -17963 7704 -17928
rect 7670 -18035 7704 -18011
rect 7670 -18107 7704 -18079
rect 7670 -18179 7704 -18147
rect 7670 -18249 7704 -18215
rect 7670 -18317 7704 -18285
rect 7670 -18385 7704 -18357
rect 7670 -18453 7704 -18429
rect 7670 -18536 7704 -18501
rect 8688 -17963 8722 -17928
rect 8688 -18035 8722 -18011
rect 8688 -18107 8722 -18079
rect 8688 -18179 8722 -18147
rect 8688 -18249 8722 -18215
rect 8688 -18317 8722 -18285
rect 8688 -18385 8722 -18357
rect 8688 -18453 8722 -18429
rect 8688 -18536 8722 -18501
rect 9706 -17963 9740 -17928
rect 9706 -18035 9740 -18011
rect 9706 -18107 9740 -18079
rect 9706 -18179 9740 -18147
rect 9706 -18249 9740 -18215
rect 9706 -18317 9740 -18285
rect 9706 -18385 9740 -18357
rect 9706 -18453 9740 -18429
rect 9706 -18536 9740 -18501
rect 10724 -17963 10758 -17928
rect 10724 -18035 10758 -18011
rect 10724 -18107 10758 -18079
rect 10724 -18179 10758 -18147
rect 10724 -18249 10758 -18215
rect 10724 -18317 10758 -18285
rect 10724 -18385 10758 -18357
rect 10724 -18453 10758 -18429
rect 10724 -18536 10758 -18501
rect 11742 -17963 11776 -17928
rect 11742 -18035 11776 -18011
rect 11742 -18107 11776 -18079
rect 11742 -18179 11776 -18147
rect 11742 -18249 11776 -18215
rect 11742 -18317 11776 -18285
rect 11742 -18385 11776 -18357
rect 11742 -18453 11776 -18429
rect 11742 -18536 11776 -18501
rect 12760 -17963 12794 -17928
rect 12760 -18035 12794 -18011
rect 12760 -18107 12794 -18079
rect 12760 -18179 12794 -18147
rect 12760 -18249 12794 -18215
rect 12760 -18317 12794 -18285
rect 12760 -18385 12794 -18357
rect 12760 -18453 12794 -18429
rect 12760 -18536 12794 -18501
rect 13778 -17963 13812 -17928
rect 13778 -18035 13812 -18011
rect 13778 -18107 13812 -18079
rect 13778 -18179 13812 -18147
rect 13778 -18249 13812 -18215
rect 13778 -18317 13812 -18285
rect 13778 -18385 13812 -18357
rect 13778 -18453 13812 -18429
rect 13778 -18536 13812 -18501
rect 14796 -17963 14830 -17928
rect 14796 -18035 14830 -18011
rect 14796 -18107 14830 -18079
rect 14796 -18179 14830 -18147
rect 14796 -18249 14830 -18215
rect 14796 -18317 14830 -18285
rect 14796 -18385 14830 -18357
rect 14796 -18453 14830 -18429
rect 14796 -18536 14830 -18501
rect 15814 -17963 15848 -17928
rect 15814 -18035 15848 -18011
rect 15814 -18107 15848 -18079
rect 15814 -18179 15848 -18147
rect 15814 -18249 15848 -18215
rect 15814 -18317 15848 -18285
rect 15814 -18385 15848 -18357
rect 15814 -18453 15848 -18429
rect 15814 -18536 15848 -18501
rect 16832 -17963 16866 -17928
rect 16832 -18035 16866 -18011
rect 16832 -18107 16866 -18079
rect 16832 -18179 16866 -18147
rect 16832 -18249 16866 -18215
rect 16832 -18317 16866 -18285
rect 16832 -18385 16866 -18357
rect 16832 -18453 16866 -18429
rect 16832 -18536 16866 -18501
rect 17850 -17963 17884 -17928
rect 17850 -18035 17884 -18011
rect 17850 -18107 17884 -18079
rect 17850 -18179 17884 -18147
rect 17850 -18249 17884 -18215
rect 17850 -18317 17884 -18285
rect 17850 -18385 17884 -18357
rect 17850 -18453 17884 -18429
rect 17850 -18536 17884 -18501
rect 18868 -17963 18902 -17928
rect 18868 -18035 18902 -18011
rect 18868 -18107 18902 -18079
rect 18868 -18179 18902 -18147
rect 18868 -18249 18902 -18215
rect 18868 -18317 18902 -18285
rect 18868 -18385 18902 -18357
rect 18868 -18453 18902 -18429
rect 18868 -18536 18902 -18501
rect 19886 -17963 19920 -17928
rect 19886 -18035 19920 -18011
rect 19886 -18107 19920 -18079
rect 19886 -18179 19920 -18147
rect 19886 -18249 19920 -18215
rect 19886 -18317 19920 -18285
rect 19886 -18385 19920 -18357
rect 19886 -18453 19920 -18429
rect 19886 -18536 19920 -18501
rect 20904 -17963 20938 -17928
rect 20904 -18035 20938 -18011
rect 20904 -18107 20938 -18079
rect 20904 -18179 20938 -18147
rect 20904 -18249 20938 -18215
rect 20904 -18317 20938 -18285
rect 20904 -18385 20938 -18357
rect 20904 -18453 20938 -18429
rect 20904 -18536 20938 -18501
rect 21922 -17963 21956 -17928
rect 21922 -18035 21956 -18011
rect 21922 -18107 21956 -18079
rect 21922 -18179 21956 -18147
rect 21922 -18249 21956 -18215
rect 21922 -18317 21956 -18285
rect 21922 -18385 21956 -18357
rect 21922 -18453 21956 -18429
rect 21922 -18536 21956 -18501
rect 22940 -17963 22974 -17928
rect 22940 -18035 22974 -18011
rect 22940 -18107 22974 -18079
rect 22940 -18179 22974 -18147
rect 22940 -18249 22974 -18215
rect 22940 -18317 22974 -18285
rect 22940 -18385 22974 -18357
rect 22940 -18453 22974 -18429
rect 22940 -18536 22974 -18501
rect 24822 -17957 24855 -17891
rect 24889 -17957 24922 -17891
rect 24822 -17959 24922 -17957
rect 24822 -17993 24855 -17959
rect 24889 -17993 24922 -17959
rect 24822 -17995 24922 -17993
rect 24822 -18061 24855 -17995
rect 24889 -18061 24922 -17995
rect 24822 -18067 24922 -18061
rect 24822 -18129 24855 -18067
rect 24889 -18129 24922 -18067
rect 24822 -18139 24922 -18129
rect 24822 -18197 24855 -18139
rect 24889 -18197 24922 -18139
rect 24822 -18211 24922 -18197
rect 24822 -18265 24855 -18211
rect 24889 -18265 24922 -18211
rect 24822 -18283 24922 -18265
rect 24822 -18333 24855 -18283
rect 24889 -18333 24922 -18283
rect 24822 -18355 24922 -18333
rect 24822 -18401 24855 -18355
rect 24889 -18401 24922 -18355
rect 24822 -18427 24922 -18401
rect 24822 -18469 24855 -18427
rect 24889 -18469 24922 -18427
rect 24822 -18499 24922 -18469
rect 24822 -18537 24855 -18499
rect 24889 -18537 24922 -18499
rect -22 -18623 12 -18591
rect 2812 -18604 2851 -18570
rect 2885 -18604 2909 -18570
rect 2953 -18604 2981 -18570
rect 3021 -18604 3053 -18570
rect 3089 -18604 3123 -18570
rect 3159 -18604 3191 -18570
rect 3231 -18604 3259 -18570
rect 3303 -18604 3327 -18570
rect 3361 -18604 3400 -18570
rect 3830 -18604 3869 -18570
rect 3903 -18604 3927 -18570
rect 3971 -18604 3999 -18570
rect 4039 -18604 4071 -18570
rect 4107 -18604 4141 -18570
rect 4177 -18604 4209 -18570
rect 4249 -18604 4277 -18570
rect 4321 -18604 4345 -18570
rect 4379 -18604 4418 -18570
rect 4848 -18604 4887 -18570
rect 4921 -18604 4945 -18570
rect 4989 -18604 5017 -18570
rect 5057 -18604 5089 -18570
rect 5125 -18604 5159 -18570
rect 5195 -18604 5227 -18570
rect 5267 -18604 5295 -18570
rect 5339 -18604 5363 -18570
rect 5397 -18604 5436 -18570
rect 5866 -18604 5905 -18570
rect 5939 -18604 5963 -18570
rect 6007 -18604 6035 -18570
rect 6075 -18604 6107 -18570
rect 6143 -18604 6177 -18570
rect 6213 -18604 6245 -18570
rect 6285 -18604 6313 -18570
rect 6357 -18604 6381 -18570
rect 6415 -18604 6454 -18570
rect 6884 -18604 6923 -18570
rect 6957 -18604 6981 -18570
rect 7025 -18604 7053 -18570
rect 7093 -18604 7125 -18570
rect 7161 -18604 7195 -18570
rect 7231 -18604 7263 -18570
rect 7303 -18604 7331 -18570
rect 7375 -18604 7399 -18570
rect 7433 -18604 7472 -18570
rect 7902 -18604 7941 -18570
rect 7975 -18604 7999 -18570
rect 8043 -18604 8071 -18570
rect 8111 -18604 8143 -18570
rect 8179 -18604 8213 -18570
rect 8249 -18604 8281 -18570
rect 8321 -18604 8349 -18570
rect 8393 -18604 8417 -18570
rect 8451 -18604 8490 -18570
rect 8920 -18604 8959 -18570
rect 8993 -18604 9017 -18570
rect 9061 -18604 9089 -18570
rect 9129 -18604 9161 -18570
rect 9197 -18604 9231 -18570
rect 9267 -18604 9299 -18570
rect 9339 -18604 9367 -18570
rect 9411 -18604 9435 -18570
rect 9469 -18604 9508 -18570
rect 9938 -18604 9977 -18570
rect 10011 -18604 10035 -18570
rect 10079 -18604 10107 -18570
rect 10147 -18604 10179 -18570
rect 10215 -18604 10249 -18570
rect 10285 -18604 10317 -18570
rect 10357 -18604 10385 -18570
rect 10429 -18604 10453 -18570
rect 10487 -18604 10526 -18570
rect 10956 -18604 10995 -18570
rect 11029 -18604 11053 -18570
rect 11097 -18604 11125 -18570
rect 11165 -18604 11197 -18570
rect 11233 -18604 11267 -18570
rect 11303 -18604 11335 -18570
rect 11375 -18604 11403 -18570
rect 11447 -18604 11471 -18570
rect 11505 -18604 11544 -18570
rect 11974 -18604 12013 -18570
rect 12047 -18604 12071 -18570
rect 12115 -18604 12143 -18570
rect 12183 -18604 12215 -18570
rect 12251 -18604 12285 -18570
rect 12321 -18604 12353 -18570
rect 12393 -18604 12421 -18570
rect 12465 -18604 12489 -18570
rect 12523 -18604 12562 -18570
rect 12992 -18604 13031 -18570
rect 13065 -18604 13089 -18570
rect 13133 -18604 13161 -18570
rect 13201 -18604 13233 -18570
rect 13269 -18604 13303 -18570
rect 13339 -18604 13371 -18570
rect 13411 -18604 13439 -18570
rect 13483 -18604 13507 -18570
rect 13541 -18604 13580 -18570
rect 14010 -18604 14049 -18570
rect 14083 -18604 14107 -18570
rect 14151 -18604 14179 -18570
rect 14219 -18604 14251 -18570
rect 14287 -18604 14321 -18570
rect 14357 -18604 14389 -18570
rect 14429 -18604 14457 -18570
rect 14501 -18604 14525 -18570
rect 14559 -18604 14598 -18570
rect 15028 -18604 15067 -18570
rect 15101 -18604 15125 -18570
rect 15169 -18604 15197 -18570
rect 15237 -18604 15269 -18570
rect 15305 -18604 15339 -18570
rect 15375 -18604 15407 -18570
rect 15447 -18604 15475 -18570
rect 15519 -18604 15543 -18570
rect 15577 -18604 15616 -18570
rect 16046 -18604 16085 -18570
rect 16119 -18604 16143 -18570
rect 16187 -18604 16215 -18570
rect 16255 -18604 16287 -18570
rect 16323 -18604 16357 -18570
rect 16393 -18604 16425 -18570
rect 16465 -18604 16493 -18570
rect 16537 -18604 16561 -18570
rect 16595 -18604 16634 -18570
rect 17064 -18604 17103 -18570
rect 17137 -18604 17161 -18570
rect 17205 -18604 17233 -18570
rect 17273 -18604 17305 -18570
rect 17341 -18604 17375 -18570
rect 17411 -18604 17443 -18570
rect 17483 -18604 17511 -18570
rect 17555 -18604 17579 -18570
rect 17613 -18604 17652 -18570
rect 18082 -18604 18121 -18570
rect 18155 -18604 18179 -18570
rect 18223 -18604 18251 -18570
rect 18291 -18604 18323 -18570
rect 18359 -18604 18393 -18570
rect 18429 -18604 18461 -18570
rect 18501 -18604 18529 -18570
rect 18573 -18604 18597 -18570
rect 18631 -18604 18670 -18570
rect 19100 -18604 19139 -18570
rect 19173 -18604 19197 -18570
rect 19241 -18604 19269 -18570
rect 19309 -18604 19341 -18570
rect 19377 -18604 19411 -18570
rect 19447 -18604 19479 -18570
rect 19519 -18604 19547 -18570
rect 19591 -18604 19615 -18570
rect 19649 -18604 19688 -18570
rect 20118 -18604 20157 -18570
rect 20191 -18604 20215 -18570
rect 20259 -18604 20287 -18570
rect 20327 -18604 20359 -18570
rect 20395 -18604 20429 -18570
rect 20465 -18604 20497 -18570
rect 20537 -18604 20565 -18570
rect 20609 -18604 20633 -18570
rect 20667 -18604 20706 -18570
rect 21136 -18604 21175 -18570
rect 21209 -18604 21233 -18570
rect 21277 -18604 21305 -18570
rect 21345 -18604 21377 -18570
rect 21413 -18604 21447 -18570
rect 21483 -18604 21515 -18570
rect 21555 -18604 21583 -18570
rect 21627 -18604 21651 -18570
rect 21685 -18604 21724 -18570
rect 22154 -18604 22193 -18570
rect 22227 -18604 22251 -18570
rect 22295 -18604 22323 -18570
rect 22363 -18604 22395 -18570
rect 22431 -18604 22465 -18570
rect 22501 -18604 22533 -18570
rect 22573 -18604 22601 -18570
rect 22645 -18604 22669 -18570
rect 22703 -18604 22742 -18570
rect 24822 -18571 24922 -18537
rect -22 -18691 12 -18663
rect -22 -18759 12 -18735
rect -22 -18842 12 -18807
rect 24822 -18605 24855 -18571
rect 24889 -18605 24922 -18571
rect 24822 -18639 24922 -18605
rect 24822 -18677 24855 -18639
rect 24889 -18677 24922 -18639
rect 24822 -18707 24922 -18677
rect 24822 -18749 24855 -18707
rect 24889 -18749 24922 -18707
rect 24822 -18775 24922 -18749
rect 24822 -18821 24855 -18775
rect 24889 -18821 24922 -18775
rect -12322 -18893 -12289 -18843
rect -12255 -18893 -12222 -18843
rect 24822 -18843 24922 -18821
rect -12322 -18911 -12222 -18893
rect -8952 -18910 -8913 -18876
rect -8879 -18910 -8855 -18876
rect -8811 -18910 -8783 -18876
rect -8743 -18910 -8711 -18876
rect -8675 -18910 -8641 -18876
rect -8605 -18910 -8573 -18876
rect -8533 -18910 -8505 -18876
rect -8461 -18910 -8437 -18876
rect -8403 -18910 -8364 -18876
rect -7934 -18910 -7895 -18876
rect -7861 -18910 -7837 -18876
rect -7793 -18910 -7765 -18876
rect -7725 -18910 -7693 -18876
rect -7657 -18910 -7623 -18876
rect -7587 -18910 -7555 -18876
rect -7515 -18910 -7487 -18876
rect -7443 -18910 -7419 -18876
rect -7385 -18910 -7346 -18876
rect -6916 -18910 -6877 -18876
rect -6843 -18910 -6819 -18876
rect -6775 -18910 -6747 -18876
rect -6707 -18910 -6675 -18876
rect -6639 -18910 -6605 -18876
rect -6569 -18910 -6537 -18876
rect -6497 -18910 -6469 -18876
rect -6425 -18910 -6401 -18876
rect -6367 -18910 -6328 -18876
rect -5898 -18910 -5859 -18876
rect -5825 -18910 -5801 -18876
rect -5757 -18910 -5729 -18876
rect -5689 -18910 -5657 -18876
rect -5621 -18910 -5587 -18876
rect -5551 -18910 -5519 -18876
rect -5479 -18910 -5451 -18876
rect -5407 -18910 -5383 -18876
rect -5349 -18910 -5310 -18876
rect -4880 -18910 -4841 -18876
rect -4807 -18910 -4783 -18876
rect -4739 -18910 -4711 -18876
rect -4671 -18910 -4639 -18876
rect -4603 -18910 -4569 -18876
rect -4533 -18910 -4501 -18876
rect -4461 -18910 -4433 -18876
rect -4389 -18910 -4365 -18876
rect -4331 -18910 -4292 -18876
rect -3862 -18910 -3823 -18876
rect -3789 -18910 -3765 -18876
rect -3721 -18910 -3693 -18876
rect -3653 -18910 -3621 -18876
rect -3585 -18910 -3551 -18876
rect -3515 -18910 -3483 -18876
rect -3443 -18910 -3415 -18876
rect -3371 -18910 -3347 -18876
rect -3313 -18910 -3274 -18876
rect -2844 -18910 -2805 -18876
rect -2771 -18910 -2747 -18876
rect -2703 -18910 -2675 -18876
rect -2635 -18910 -2603 -18876
rect -2567 -18910 -2533 -18876
rect -2497 -18910 -2465 -18876
rect -2425 -18910 -2397 -18876
rect -2353 -18910 -2329 -18876
rect -2295 -18910 -2256 -18876
rect -1826 -18910 -1787 -18876
rect -1753 -18910 -1729 -18876
rect -1685 -18910 -1657 -18876
rect -1617 -18910 -1585 -18876
rect -1549 -18910 -1515 -18876
rect -1479 -18910 -1447 -18876
rect -1407 -18910 -1379 -18876
rect -1335 -18910 -1311 -18876
rect -1277 -18910 -1238 -18876
rect -808 -18910 -769 -18876
rect -735 -18910 -711 -18876
rect -667 -18910 -639 -18876
rect -599 -18910 -567 -18876
rect -531 -18910 -497 -18876
rect -461 -18910 -429 -18876
rect -389 -18910 -361 -18876
rect -317 -18910 -293 -18876
rect -259 -18910 -220 -18876
rect 24822 -18893 24855 -18843
rect 24889 -18893 24922 -18843
rect -12322 -18965 -12289 -18911
rect -12255 -18965 -12222 -18911
rect -12322 -18979 -12222 -18965
rect -12322 -19037 -12289 -18979
rect -12255 -19037 -12222 -18979
rect -12322 -19047 -12222 -19037
rect -12322 -19109 -12289 -19047
rect -12255 -19109 -12222 -19047
rect 24822 -18911 24922 -18893
rect 24822 -18965 24855 -18911
rect 24889 -18965 24922 -18911
rect 24822 -18979 24922 -18965
rect 24822 -19037 24855 -18979
rect 24889 -19037 24922 -18979
rect 24822 -19047 24922 -19037
rect -12322 -19115 -12222 -19109
rect -12322 -19181 -12289 -19115
rect -12255 -19181 -12222 -19115
rect 2812 -19126 2851 -19092
rect 2885 -19126 2909 -19092
rect 2953 -19126 2981 -19092
rect 3021 -19126 3053 -19092
rect 3089 -19126 3123 -19092
rect 3159 -19126 3191 -19092
rect 3231 -19126 3259 -19092
rect 3303 -19126 3327 -19092
rect 3361 -19126 3400 -19092
rect 3830 -19126 3869 -19092
rect 3903 -19126 3927 -19092
rect 3971 -19126 3999 -19092
rect 4039 -19126 4071 -19092
rect 4107 -19126 4141 -19092
rect 4177 -19126 4209 -19092
rect 4249 -19126 4277 -19092
rect 4321 -19126 4345 -19092
rect 4379 -19126 4418 -19092
rect 4848 -19126 4887 -19092
rect 4921 -19126 4945 -19092
rect 4989 -19126 5017 -19092
rect 5057 -19126 5089 -19092
rect 5125 -19126 5159 -19092
rect 5195 -19126 5227 -19092
rect 5267 -19126 5295 -19092
rect 5339 -19126 5363 -19092
rect 5397 -19126 5436 -19092
rect 5866 -19126 5905 -19092
rect 5939 -19126 5963 -19092
rect 6007 -19126 6035 -19092
rect 6075 -19126 6107 -19092
rect 6143 -19126 6177 -19092
rect 6213 -19126 6245 -19092
rect 6285 -19126 6313 -19092
rect 6357 -19126 6381 -19092
rect 6415 -19126 6454 -19092
rect 6884 -19126 6923 -19092
rect 6957 -19126 6981 -19092
rect 7025 -19126 7053 -19092
rect 7093 -19126 7125 -19092
rect 7161 -19126 7195 -19092
rect 7231 -19126 7263 -19092
rect 7303 -19126 7331 -19092
rect 7375 -19126 7399 -19092
rect 7433 -19126 7472 -19092
rect 7902 -19126 7941 -19092
rect 7975 -19126 7999 -19092
rect 8043 -19126 8071 -19092
rect 8111 -19126 8143 -19092
rect 8179 -19126 8213 -19092
rect 8249 -19126 8281 -19092
rect 8321 -19126 8349 -19092
rect 8393 -19126 8417 -19092
rect 8451 -19126 8490 -19092
rect 8920 -19126 8959 -19092
rect 8993 -19126 9017 -19092
rect 9061 -19126 9089 -19092
rect 9129 -19126 9161 -19092
rect 9197 -19126 9231 -19092
rect 9267 -19126 9299 -19092
rect 9339 -19126 9367 -19092
rect 9411 -19126 9435 -19092
rect 9469 -19126 9508 -19092
rect 9938 -19126 9977 -19092
rect 10011 -19126 10035 -19092
rect 10079 -19126 10107 -19092
rect 10147 -19126 10179 -19092
rect 10215 -19126 10249 -19092
rect 10285 -19126 10317 -19092
rect 10357 -19126 10385 -19092
rect 10429 -19126 10453 -19092
rect 10487 -19126 10526 -19092
rect 10956 -19126 10995 -19092
rect 11029 -19126 11053 -19092
rect 11097 -19126 11125 -19092
rect 11165 -19126 11197 -19092
rect 11233 -19126 11267 -19092
rect 11303 -19126 11335 -19092
rect 11375 -19126 11403 -19092
rect 11447 -19126 11471 -19092
rect 11505 -19126 11544 -19092
rect 11974 -19126 12013 -19092
rect 12047 -19126 12071 -19092
rect 12115 -19126 12143 -19092
rect 12183 -19126 12215 -19092
rect 12251 -19126 12285 -19092
rect 12321 -19126 12353 -19092
rect 12393 -19126 12421 -19092
rect 12465 -19126 12489 -19092
rect 12523 -19126 12562 -19092
rect 12992 -19126 13031 -19092
rect 13065 -19126 13089 -19092
rect 13133 -19126 13161 -19092
rect 13201 -19126 13233 -19092
rect 13269 -19126 13303 -19092
rect 13339 -19126 13371 -19092
rect 13411 -19126 13439 -19092
rect 13483 -19126 13507 -19092
rect 13541 -19126 13580 -19092
rect 14010 -19126 14049 -19092
rect 14083 -19126 14107 -19092
rect 14151 -19126 14179 -19092
rect 14219 -19126 14251 -19092
rect 14287 -19126 14321 -19092
rect 14357 -19126 14389 -19092
rect 14429 -19126 14457 -19092
rect 14501 -19126 14525 -19092
rect 14559 -19126 14598 -19092
rect 15028 -19126 15067 -19092
rect 15101 -19126 15125 -19092
rect 15169 -19126 15197 -19092
rect 15237 -19126 15269 -19092
rect 15305 -19126 15339 -19092
rect 15375 -19126 15407 -19092
rect 15447 -19126 15475 -19092
rect 15519 -19126 15543 -19092
rect 15577 -19126 15616 -19092
rect 16046 -19126 16085 -19092
rect 16119 -19126 16143 -19092
rect 16187 -19126 16215 -19092
rect 16255 -19126 16287 -19092
rect 16323 -19126 16357 -19092
rect 16393 -19126 16425 -19092
rect 16465 -19126 16493 -19092
rect 16537 -19126 16561 -19092
rect 16595 -19126 16634 -19092
rect 17064 -19126 17103 -19092
rect 17137 -19126 17161 -19092
rect 17205 -19126 17233 -19092
rect 17273 -19126 17305 -19092
rect 17341 -19126 17375 -19092
rect 17411 -19126 17443 -19092
rect 17483 -19126 17511 -19092
rect 17555 -19126 17579 -19092
rect 17613 -19126 17652 -19092
rect 18082 -19126 18121 -19092
rect 18155 -19126 18179 -19092
rect 18223 -19126 18251 -19092
rect 18291 -19126 18323 -19092
rect 18359 -19126 18393 -19092
rect 18429 -19126 18461 -19092
rect 18501 -19126 18529 -19092
rect 18573 -19126 18597 -19092
rect 18631 -19126 18670 -19092
rect 19100 -19126 19139 -19092
rect 19173 -19126 19197 -19092
rect 19241 -19126 19269 -19092
rect 19309 -19126 19341 -19092
rect 19377 -19126 19411 -19092
rect 19447 -19126 19479 -19092
rect 19519 -19126 19547 -19092
rect 19591 -19126 19615 -19092
rect 19649 -19126 19688 -19092
rect 20118 -19126 20157 -19092
rect 20191 -19126 20215 -19092
rect 20259 -19126 20287 -19092
rect 20327 -19126 20359 -19092
rect 20395 -19126 20429 -19092
rect 20465 -19126 20497 -19092
rect 20537 -19126 20565 -19092
rect 20609 -19126 20633 -19092
rect 20667 -19126 20706 -19092
rect 21136 -19126 21175 -19092
rect 21209 -19126 21233 -19092
rect 21277 -19126 21305 -19092
rect 21345 -19126 21377 -19092
rect 21413 -19126 21447 -19092
rect 21483 -19126 21515 -19092
rect 21555 -19126 21583 -19092
rect 21627 -19126 21651 -19092
rect 21685 -19126 21724 -19092
rect 22154 -19126 22193 -19092
rect 22227 -19126 22251 -19092
rect 22295 -19126 22323 -19092
rect 22363 -19126 22395 -19092
rect 22431 -19126 22465 -19092
rect 22501 -19126 22533 -19092
rect 22573 -19126 22601 -19092
rect 22645 -19126 22669 -19092
rect 22703 -19126 22742 -19092
rect 24822 -19109 24855 -19047
rect 24889 -19109 24922 -19047
rect 24822 -19115 24922 -19109
rect -12322 -19183 -12222 -19181
rect -12322 -19217 -12289 -19183
rect -12255 -19217 -12222 -19183
rect -12322 -19219 -12222 -19217
rect -12322 -19285 -12289 -19219
rect -12255 -19285 -12222 -19219
rect -12322 -19291 -12222 -19285
rect -12322 -19353 -12289 -19291
rect -12255 -19353 -12222 -19291
rect -12322 -19363 -12222 -19353
rect -12322 -19421 -12289 -19363
rect -12255 -19421 -12222 -19363
rect -12322 -19435 -12222 -19421
rect -12322 -19489 -12289 -19435
rect -12255 -19489 -12222 -19435
rect -12322 -19507 -12222 -19489
rect -12322 -19557 -12289 -19507
rect -12255 -19557 -12222 -19507
rect -12322 -19579 -12222 -19557
rect -12322 -19625 -12289 -19579
rect -12255 -19625 -12222 -19579
rect -12322 -19651 -12222 -19625
rect -12322 -19693 -12289 -19651
rect -12255 -19693 -12222 -19651
rect -12322 -19723 -12222 -19693
rect -12322 -19761 -12289 -19723
rect -12255 -19761 -12222 -19723
rect -12322 -19795 -12222 -19761
rect 2580 -19195 2614 -19160
rect 2580 -19267 2614 -19243
rect 2580 -19339 2614 -19311
rect 2580 -19411 2614 -19379
rect 2580 -19481 2614 -19447
rect 2580 -19549 2614 -19517
rect 2580 -19617 2614 -19589
rect 2580 -19685 2614 -19661
rect 2580 -19768 2614 -19733
rect 3598 -19195 3632 -19160
rect 3598 -19267 3632 -19243
rect 3598 -19339 3632 -19311
rect 3598 -19411 3632 -19379
rect 3598 -19481 3632 -19447
rect 3598 -19549 3632 -19517
rect 3598 -19617 3632 -19589
rect 3598 -19685 3632 -19661
rect 3598 -19768 3632 -19733
rect 4616 -19195 4650 -19160
rect 4616 -19267 4650 -19243
rect 4616 -19339 4650 -19311
rect 4616 -19411 4650 -19379
rect 4616 -19481 4650 -19447
rect 4616 -19549 4650 -19517
rect 4616 -19617 4650 -19589
rect 4616 -19685 4650 -19661
rect 4616 -19768 4650 -19733
rect 5634 -19195 5668 -19160
rect 5634 -19267 5668 -19243
rect 5634 -19339 5668 -19311
rect 5634 -19411 5668 -19379
rect 5634 -19481 5668 -19447
rect 5634 -19549 5668 -19517
rect 5634 -19617 5668 -19589
rect 5634 -19685 5668 -19661
rect 5634 -19768 5668 -19733
rect 6652 -19195 6686 -19160
rect 6652 -19267 6686 -19243
rect 6652 -19339 6686 -19311
rect 6652 -19411 6686 -19379
rect 6652 -19481 6686 -19447
rect 6652 -19549 6686 -19517
rect 6652 -19617 6686 -19589
rect 6652 -19685 6686 -19661
rect 6652 -19768 6686 -19733
rect 7670 -19195 7704 -19160
rect 7670 -19267 7704 -19243
rect 7670 -19339 7704 -19311
rect 7670 -19411 7704 -19379
rect 7670 -19481 7704 -19447
rect 7670 -19549 7704 -19517
rect 7670 -19617 7704 -19589
rect 7670 -19685 7704 -19661
rect 7670 -19768 7704 -19733
rect 8688 -19195 8722 -19160
rect 8688 -19267 8722 -19243
rect 8688 -19339 8722 -19311
rect 8688 -19411 8722 -19379
rect 8688 -19481 8722 -19447
rect 8688 -19549 8722 -19517
rect 8688 -19617 8722 -19589
rect 8688 -19685 8722 -19661
rect 8688 -19768 8722 -19733
rect 9706 -19195 9740 -19160
rect 9706 -19267 9740 -19243
rect 9706 -19339 9740 -19311
rect 9706 -19411 9740 -19379
rect 9706 -19481 9740 -19447
rect 9706 -19549 9740 -19517
rect 9706 -19617 9740 -19589
rect 9706 -19685 9740 -19661
rect 9706 -19768 9740 -19733
rect 10724 -19195 10758 -19160
rect 10724 -19267 10758 -19243
rect 10724 -19339 10758 -19311
rect 10724 -19411 10758 -19379
rect 10724 -19481 10758 -19447
rect 10724 -19549 10758 -19517
rect 10724 -19617 10758 -19589
rect 10724 -19685 10758 -19661
rect 10724 -19768 10758 -19733
rect 11742 -19195 11776 -19160
rect 11742 -19267 11776 -19243
rect 11742 -19339 11776 -19311
rect 11742 -19411 11776 -19379
rect 11742 -19481 11776 -19447
rect 11742 -19549 11776 -19517
rect 11742 -19617 11776 -19589
rect 11742 -19685 11776 -19661
rect 11742 -19768 11776 -19733
rect 12760 -19195 12794 -19160
rect 12760 -19267 12794 -19243
rect 12760 -19339 12794 -19311
rect 12760 -19411 12794 -19379
rect 12760 -19481 12794 -19447
rect 12760 -19549 12794 -19517
rect 12760 -19617 12794 -19589
rect 12760 -19685 12794 -19661
rect 12760 -19768 12794 -19733
rect 13778 -19195 13812 -19160
rect 13778 -19267 13812 -19243
rect 13778 -19339 13812 -19311
rect 13778 -19411 13812 -19379
rect 13778 -19481 13812 -19447
rect 13778 -19549 13812 -19517
rect 13778 -19617 13812 -19589
rect 13778 -19685 13812 -19661
rect 13778 -19768 13812 -19733
rect 14796 -19195 14830 -19160
rect 14796 -19267 14830 -19243
rect 14796 -19339 14830 -19311
rect 14796 -19411 14830 -19379
rect 14796 -19481 14830 -19447
rect 14796 -19549 14830 -19517
rect 14796 -19617 14830 -19589
rect 14796 -19685 14830 -19661
rect 14796 -19768 14830 -19733
rect 15814 -19195 15848 -19160
rect 15814 -19267 15848 -19243
rect 15814 -19339 15848 -19311
rect 15814 -19411 15848 -19379
rect 15814 -19481 15848 -19447
rect 15814 -19549 15848 -19517
rect 15814 -19617 15848 -19589
rect 15814 -19685 15848 -19661
rect 15814 -19768 15848 -19733
rect 16832 -19195 16866 -19160
rect 16832 -19267 16866 -19243
rect 16832 -19339 16866 -19311
rect 16832 -19411 16866 -19379
rect 16832 -19481 16866 -19447
rect 16832 -19549 16866 -19517
rect 16832 -19617 16866 -19589
rect 16832 -19685 16866 -19661
rect 16832 -19768 16866 -19733
rect 17850 -19195 17884 -19160
rect 17850 -19267 17884 -19243
rect 17850 -19339 17884 -19311
rect 17850 -19411 17884 -19379
rect 17850 -19481 17884 -19447
rect 17850 -19549 17884 -19517
rect 17850 -19617 17884 -19589
rect 17850 -19685 17884 -19661
rect 17850 -19768 17884 -19733
rect 18868 -19195 18902 -19160
rect 18868 -19267 18902 -19243
rect 18868 -19339 18902 -19311
rect 18868 -19411 18902 -19379
rect 18868 -19481 18902 -19447
rect 18868 -19549 18902 -19517
rect 18868 -19617 18902 -19589
rect 18868 -19685 18902 -19661
rect 18868 -19768 18902 -19733
rect 19886 -19195 19920 -19160
rect 19886 -19267 19920 -19243
rect 19886 -19339 19920 -19311
rect 19886 -19411 19920 -19379
rect 19886 -19481 19920 -19447
rect 19886 -19549 19920 -19517
rect 19886 -19617 19920 -19589
rect 19886 -19685 19920 -19661
rect 19886 -19768 19920 -19733
rect 20904 -19195 20938 -19160
rect 20904 -19267 20938 -19243
rect 20904 -19339 20938 -19311
rect 20904 -19411 20938 -19379
rect 20904 -19481 20938 -19447
rect 20904 -19549 20938 -19517
rect 20904 -19617 20938 -19589
rect 20904 -19685 20938 -19661
rect 20904 -19768 20938 -19733
rect 21922 -19195 21956 -19160
rect 21922 -19267 21956 -19243
rect 21922 -19339 21956 -19311
rect 21922 -19411 21956 -19379
rect 21922 -19481 21956 -19447
rect 21922 -19549 21956 -19517
rect 21922 -19617 21956 -19589
rect 21922 -19685 21956 -19661
rect 21922 -19768 21956 -19733
rect 22940 -19195 22974 -19160
rect 22940 -19267 22974 -19243
rect 22940 -19339 22974 -19311
rect 22940 -19411 22974 -19379
rect 22940 -19481 22974 -19447
rect 22940 -19549 22974 -19517
rect 22940 -19617 22974 -19589
rect 22940 -19685 22974 -19661
rect 22940 -19768 22974 -19733
rect 24822 -19181 24855 -19115
rect 24889 -19181 24922 -19115
rect 24822 -19183 24922 -19181
rect 24822 -19217 24855 -19183
rect 24889 -19217 24922 -19183
rect 24822 -19219 24922 -19217
rect 24822 -19285 24855 -19219
rect 24889 -19285 24922 -19219
rect 24822 -19291 24922 -19285
rect 24822 -19353 24855 -19291
rect 24889 -19353 24922 -19291
rect 24822 -19363 24922 -19353
rect 24822 -19421 24855 -19363
rect 24889 -19421 24922 -19363
rect 24822 -19435 24922 -19421
rect 24822 -19489 24855 -19435
rect 24889 -19489 24922 -19435
rect 24822 -19507 24922 -19489
rect 24822 -19557 24855 -19507
rect 24889 -19557 24922 -19507
rect 24822 -19579 24922 -19557
rect 24822 -19625 24855 -19579
rect 24889 -19625 24922 -19579
rect 24822 -19651 24922 -19625
rect 24822 -19693 24855 -19651
rect 24889 -19693 24922 -19651
rect 24822 -19723 24922 -19693
rect 24822 -19761 24855 -19723
rect 24889 -19761 24922 -19723
rect -12322 -19829 -12289 -19795
rect -12255 -19829 -12222 -19795
rect 24822 -19795 24922 -19761
rect 11230 -19802 11290 -19800
rect 13274 -19802 13334 -19798
rect 21408 -19802 21468 -19800
rect -12322 -19863 -12222 -19829
rect 2812 -19836 2851 -19802
rect 2885 -19836 2909 -19802
rect 2953 -19836 2981 -19802
rect 3021 -19836 3053 -19802
rect 3089 -19836 3123 -19802
rect 3159 -19836 3191 -19802
rect 3231 -19836 3259 -19802
rect 3303 -19836 3327 -19802
rect 3361 -19836 3400 -19802
rect 3830 -19836 3869 -19802
rect 3903 -19836 3927 -19802
rect 3971 -19836 3999 -19802
rect 4039 -19836 4071 -19802
rect 4107 -19836 4141 -19802
rect 4177 -19836 4209 -19802
rect 4249 -19836 4277 -19802
rect 4321 -19836 4345 -19802
rect 4379 -19836 4418 -19802
rect 4848 -19836 4887 -19802
rect 4921 -19836 4945 -19802
rect 4989 -19836 5017 -19802
rect 5057 -19836 5089 -19802
rect 5125 -19836 5159 -19802
rect 5195 -19836 5227 -19802
rect 5267 -19836 5295 -19802
rect 5339 -19836 5363 -19802
rect 5397 -19836 5436 -19802
rect 5866 -19836 5905 -19802
rect 5939 -19836 5963 -19802
rect 6007 -19836 6035 -19802
rect 6075 -19836 6107 -19802
rect 6143 -19836 6177 -19802
rect 6213 -19836 6245 -19802
rect 6285 -19836 6313 -19802
rect 6357 -19836 6381 -19802
rect 6415 -19836 6454 -19802
rect 6884 -19836 6923 -19802
rect 6957 -19836 6981 -19802
rect 7025 -19836 7053 -19802
rect 7093 -19836 7125 -19802
rect 7161 -19836 7195 -19802
rect 7231 -19836 7263 -19802
rect 7303 -19836 7331 -19802
rect 7375 -19836 7399 -19802
rect 7433 -19836 7472 -19802
rect 7902 -19836 7941 -19802
rect 7975 -19836 7999 -19802
rect 8043 -19836 8071 -19802
rect 8111 -19836 8143 -19802
rect 8179 -19836 8213 -19802
rect 8249 -19836 8281 -19802
rect 8321 -19836 8349 -19802
rect 8393 -19836 8417 -19802
rect 8451 -19836 8490 -19802
rect 8920 -19836 8959 -19802
rect 8993 -19836 9017 -19802
rect 9061 -19836 9089 -19802
rect 9129 -19836 9161 -19802
rect 9197 -19836 9231 -19802
rect 9267 -19836 9299 -19802
rect 9339 -19836 9367 -19802
rect 9411 -19836 9435 -19802
rect 9469 -19836 9508 -19802
rect 9938 -19836 9977 -19802
rect 10011 -19836 10035 -19802
rect 10079 -19836 10107 -19802
rect 10147 -19836 10179 -19802
rect 10215 -19836 10249 -19802
rect 10285 -19836 10317 -19802
rect 10357 -19836 10385 -19802
rect 10429 -19836 10453 -19802
rect 10487 -19836 10526 -19802
rect 10956 -19836 10995 -19802
rect 11029 -19836 11053 -19802
rect 11097 -19836 11125 -19802
rect 11165 -19836 11197 -19802
rect 11233 -19836 11267 -19802
rect 11303 -19836 11335 -19802
rect 11375 -19836 11403 -19802
rect 11447 -19836 11471 -19802
rect 11505 -19836 11544 -19802
rect 11974 -19836 12013 -19802
rect 12047 -19836 12071 -19802
rect 12115 -19836 12143 -19802
rect 12183 -19836 12215 -19802
rect 12251 -19836 12285 -19802
rect 12321 -19836 12353 -19802
rect 12393 -19836 12421 -19802
rect 12465 -19836 12489 -19802
rect 12523 -19836 12562 -19802
rect 12992 -19836 13031 -19802
rect 13065 -19836 13089 -19802
rect 13133 -19836 13161 -19802
rect 13201 -19836 13233 -19802
rect 13269 -19836 13303 -19802
rect 13339 -19836 13371 -19802
rect 13411 -19836 13439 -19802
rect 13483 -19836 13507 -19802
rect 13541 -19836 13580 -19802
rect 14010 -19836 14049 -19802
rect 14083 -19836 14107 -19802
rect 14151 -19836 14179 -19802
rect 14219 -19836 14251 -19802
rect 14287 -19836 14321 -19802
rect 14357 -19836 14389 -19802
rect 14429 -19836 14457 -19802
rect 14501 -19836 14525 -19802
rect 14559 -19836 14598 -19802
rect 15028 -19836 15067 -19802
rect 15101 -19836 15125 -19802
rect 15169 -19836 15197 -19802
rect 15237 -19836 15269 -19802
rect 15305 -19836 15339 -19802
rect 15375 -19836 15407 -19802
rect 15447 -19836 15475 -19802
rect 15519 -19836 15543 -19802
rect 15577 -19836 15616 -19802
rect 16046 -19836 16085 -19802
rect 16119 -19836 16143 -19802
rect 16187 -19836 16215 -19802
rect 16255 -19836 16287 -19802
rect 16323 -19836 16357 -19802
rect 16393 -19836 16425 -19802
rect 16465 -19836 16493 -19802
rect 16537 -19836 16561 -19802
rect 16595 -19836 16634 -19802
rect 17064 -19836 17103 -19802
rect 17137 -19836 17161 -19802
rect 17205 -19836 17233 -19802
rect 17273 -19836 17305 -19802
rect 17341 -19836 17375 -19802
rect 17411 -19836 17443 -19802
rect 17483 -19836 17511 -19802
rect 17555 -19836 17579 -19802
rect 17613 -19836 17652 -19802
rect 18082 -19836 18121 -19802
rect 18155 -19836 18179 -19802
rect 18223 -19836 18251 -19802
rect 18291 -19836 18323 -19802
rect 18359 -19836 18393 -19802
rect 18429 -19836 18461 -19802
rect 18501 -19836 18529 -19802
rect 18573 -19836 18597 -19802
rect 18631 -19836 18670 -19802
rect 19100 -19836 19139 -19802
rect 19173 -19836 19197 -19802
rect 19241 -19836 19269 -19802
rect 19309 -19836 19341 -19802
rect 19377 -19836 19411 -19802
rect 19447 -19836 19479 -19802
rect 19519 -19836 19547 -19802
rect 19591 -19836 19615 -19802
rect 19649 -19836 19688 -19802
rect 20118 -19836 20157 -19802
rect 20191 -19836 20215 -19802
rect 20259 -19836 20287 -19802
rect 20327 -19836 20359 -19802
rect 20395 -19836 20429 -19802
rect 20465 -19836 20497 -19802
rect 20537 -19836 20565 -19802
rect 20609 -19836 20633 -19802
rect 20667 -19836 20706 -19802
rect 21136 -19836 21175 -19802
rect 21209 -19836 21233 -19802
rect 21277 -19836 21305 -19802
rect 21345 -19836 21377 -19802
rect 21413 -19836 21447 -19802
rect 21483 -19836 21515 -19802
rect 21555 -19836 21583 -19802
rect 21627 -19836 21651 -19802
rect 21685 -19836 21724 -19802
rect 22154 -19836 22193 -19802
rect 22227 -19836 22251 -19802
rect 22295 -19836 22323 -19802
rect 22363 -19836 22395 -19802
rect 22431 -19836 22465 -19802
rect 22501 -19836 22533 -19802
rect 22573 -19836 22601 -19802
rect 22645 -19836 22669 -19802
rect 22703 -19836 22742 -19802
rect 24822 -19829 24855 -19795
rect 24889 -19829 24922 -19795
rect -12322 -19901 -12289 -19863
rect -12255 -19901 -12222 -19863
rect -12322 -19931 -12222 -19901
rect -12322 -19973 -12289 -19931
rect -12255 -19973 -12222 -19931
rect -12322 -19999 -12222 -19973
rect -12322 -20045 -12289 -19999
rect -12255 -20045 -12222 -19999
rect -12322 -20067 -12222 -20045
rect -12322 -20117 -12289 -20067
rect -12255 -20117 -12222 -20067
rect -12322 -20135 -12222 -20117
rect -12322 -20189 -12289 -20135
rect -12255 -20189 -12222 -20135
rect -12322 -20203 -12222 -20189
rect -12322 -20261 -12289 -20203
rect -12255 -20261 -12222 -20203
rect -12322 -20271 -12222 -20261
rect -12322 -20333 -12289 -20271
rect -12255 -20333 -12222 -20271
rect 24822 -19863 24922 -19829
rect 24822 -19901 24855 -19863
rect 24889 -19901 24922 -19863
rect 24822 -19931 24922 -19901
rect 24822 -19973 24855 -19931
rect 24889 -19973 24922 -19931
rect 24822 -19999 24922 -19973
rect 24822 -20045 24855 -19999
rect 24889 -20045 24922 -19999
rect 24822 -20067 24922 -20045
rect 24822 -20117 24855 -20067
rect 24889 -20117 24922 -20067
rect 24822 -20135 24922 -20117
rect 24822 -20189 24855 -20135
rect 24889 -20189 24922 -20135
rect 24822 -20203 24922 -20189
rect 24822 -20261 24855 -20203
rect 24889 -20261 24922 -20203
rect 24822 -20271 24922 -20261
rect -12322 -20339 -12222 -20333
rect -12322 -20405 -12289 -20339
rect -12255 -20405 -12222 -20339
rect 2812 -20360 2851 -20326
rect 2885 -20360 2909 -20326
rect 2953 -20360 2981 -20326
rect 3021 -20360 3053 -20326
rect 3089 -20360 3123 -20326
rect 3159 -20360 3191 -20326
rect 3231 -20360 3259 -20326
rect 3303 -20360 3327 -20326
rect 3361 -20360 3400 -20326
rect 3830 -20360 3869 -20326
rect 3903 -20360 3927 -20326
rect 3971 -20360 3999 -20326
rect 4039 -20360 4071 -20326
rect 4107 -20360 4141 -20326
rect 4177 -20360 4209 -20326
rect 4249 -20360 4277 -20326
rect 4321 -20360 4345 -20326
rect 4379 -20360 4418 -20326
rect 4848 -20360 4887 -20326
rect 4921 -20360 4945 -20326
rect 4989 -20360 5017 -20326
rect 5057 -20360 5089 -20326
rect 5125 -20360 5159 -20326
rect 5195 -20360 5227 -20326
rect 5267 -20360 5295 -20326
rect 5339 -20360 5363 -20326
rect 5397 -20360 5436 -20326
rect 5866 -20360 5905 -20326
rect 5939 -20360 5963 -20326
rect 6007 -20360 6035 -20326
rect 6075 -20360 6107 -20326
rect 6143 -20360 6177 -20326
rect 6213 -20360 6245 -20326
rect 6285 -20360 6313 -20326
rect 6357 -20360 6381 -20326
rect 6415 -20360 6454 -20326
rect 6884 -20360 6923 -20326
rect 6957 -20360 6981 -20326
rect 7025 -20360 7053 -20326
rect 7093 -20360 7125 -20326
rect 7161 -20360 7195 -20326
rect 7231 -20360 7263 -20326
rect 7303 -20360 7331 -20326
rect 7375 -20360 7399 -20326
rect 7433 -20360 7472 -20326
rect 7902 -20360 7941 -20326
rect 7975 -20360 7999 -20326
rect 8043 -20360 8071 -20326
rect 8111 -20360 8143 -20326
rect 8179 -20360 8213 -20326
rect 8249 -20360 8281 -20326
rect 8321 -20360 8349 -20326
rect 8393 -20360 8417 -20326
rect 8451 -20360 8490 -20326
rect 8920 -20360 8959 -20326
rect 8993 -20360 9017 -20326
rect 9061 -20360 9089 -20326
rect 9129 -20360 9161 -20326
rect 9197 -20360 9231 -20326
rect 9267 -20360 9299 -20326
rect 9339 -20360 9367 -20326
rect 9411 -20360 9435 -20326
rect 9469 -20360 9508 -20326
rect 9938 -20360 9977 -20326
rect 10011 -20360 10035 -20326
rect 10079 -20360 10107 -20326
rect 10147 -20360 10179 -20326
rect 10215 -20360 10249 -20326
rect 10285 -20360 10317 -20326
rect 10357 -20360 10385 -20326
rect 10429 -20360 10453 -20326
rect 10487 -20360 10526 -20326
rect 10956 -20360 10995 -20326
rect 11029 -20360 11053 -20326
rect 11097 -20360 11125 -20326
rect 11165 -20360 11197 -20326
rect 11233 -20360 11267 -20326
rect 11303 -20360 11335 -20326
rect 11375 -20360 11403 -20326
rect 11447 -20360 11471 -20326
rect 11505 -20360 11544 -20326
rect 11974 -20360 12013 -20326
rect 12047 -20360 12071 -20326
rect 12115 -20360 12143 -20326
rect 12183 -20360 12215 -20326
rect 12251 -20360 12285 -20326
rect 12321 -20360 12353 -20326
rect 12393 -20360 12421 -20326
rect 12465 -20360 12489 -20326
rect 12523 -20360 12562 -20326
rect 12992 -20360 13031 -20326
rect 13065 -20360 13089 -20326
rect 13133 -20360 13161 -20326
rect 13201 -20360 13233 -20326
rect 13269 -20360 13303 -20326
rect 13339 -20360 13371 -20326
rect 13411 -20360 13439 -20326
rect 13483 -20360 13507 -20326
rect 13541 -20360 13580 -20326
rect 14010 -20360 14049 -20326
rect 14083 -20360 14107 -20326
rect 14151 -20360 14179 -20326
rect 14219 -20360 14251 -20326
rect 14287 -20360 14321 -20326
rect 14357 -20360 14389 -20326
rect 14429 -20360 14457 -20326
rect 14501 -20360 14525 -20326
rect 14559 -20360 14598 -20326
rect 15028 -20360 15067 -20326
rect 15101 -20360 15125 -20326
rect 15169 -20360 15197 -20326
rect 15237 -20360 15269 -20326
rect 15305 -20360 15339 -20326
rect 15375 -20360 15407 -20326
rect 15447 -20360 15475 -20326
rect 15519 -20360 15543 -20326
rect 15577 -20360 15616 -20326
rect 16046 -20360 16085 -20326
rect 16119 -20360 16143 -20326
rect 16187 -20360 16215 -20326
rect 16255 -20360 16287 -20326
rect 16323 -20360 16357 -20326
rect 16393 -20360 16425 -20326
rect 16465 -20360 16493 -20326
rect 16537 -20360 16561 -20326
rect 16595 -20360 16634 -20326
rect 17064 -20360 17103 -20326
rect 17137 -20360 17161 -20326
rect 17205 -20360 17233 -20326
rect 17273 -20360 17305 -20326
rect 17341 -20360 17375 -20326
rect 17411 -20360 17443 -20326
rect 17483 -20360 17511 -20326
rect 17555 -20360 17579 -20326
rect 17613 -20360 17652 -20326
rect 18082 -20360 18121 -20326
rect 18155 -20360 18179 -20326
rect 18223 -20360 18251 -20326
rect 18291 -20360 18323 -20326
rect 18359 -20360 18393 -20326
rect 18429 -20360 18461 -20326
rect 18501 -20360 18529 -20326
rect 18573 -20360 18597 -20326
rect 18631 -20360 18670 -20326
rect 19100 -20360 19139 -20326
rect 19173 -20360 19197 -20326
rect 19241 -20360 19269 -20326
rect 19309 -20360 19341 -20326
rect 19377 -20360 19411 -20326
rect 19447 -20360 19479 -20326
rect 19519 -20360 19547 -20326
rect 19591 -20360 19615 -20326
rect 19649 -20360 19688 -20326
rect 20118 -20360 20157 -20326
rect 20191 -20360 20215 -20326
rect 20259 -20360 20287 -20326
rect 20327 -20360 20359 -20326
rect 20395 -20360 20429 -20326
rect 20465 -20360 20497 -20326
rect 20537 -20360 20565 -20326
rect 20609 -20360 20633 -20326
rect 20667 -20360 20706 -20326
rect 21136 -20360 21175 -20326
rect 21209 -20360 21233 -20326
rect 21277 -20360 21305 -20326
rect 21345 -20360 21377 -20326
rect 21413 -20360 21447 -20326
rect 21483 -20360 21515 -20326
rect 21555 -20360 21583 -20326
rect 21627 -20360 21651 -20326
rect 21685 -20360 21724 -20326
rect 22154 -20360 22193 -20326
rect 22227 -20360 22251 -20326
rect 22295 -20360 22323 -20326
rect 22363 -20360 22395 -20326
rect 22431 -20360 22465 -20326
rect 22501 -20360 22533 -20326
rect 22573 -20360 22601 -20326
rect 22645 -20360 22669 -20326
rect 22703 -20360 22742 -20326
rect 24822 -20333 24855 -20271
rect 24889 -20333 24922 -20271
rect 24822 -20339 24922 -20333
rect -12322 -20407 -12222 -20405
rect -12322 -20441 -12289 -20407
rect -12255 -20441 -12222 -20407
rect -12322 -20443 -12222 -20441
rect -12322 -20509 -12289 -20443
rect -12255 -20509 -12222 -20443
rect -12322 -20515 -12222 -20509
rect -12322 -20577 -12289 -20515
rect -12255 -20577 -12222 -20515
rect -12322 -20587 -12222 -20577
rect -12322 -20645 -12289 -20587
rect -12255 -20645 -12222 -20587
rect -12322 -20659 -12222 -20645
rect -12322 -20713 -12289 -20659
rect -12255 -20713 -12222 -20659
rect -12322 -20731 -12222 -20713
rect -12322 -20781 -12289 -20731
rect -12255 -20781 -12222 -20731
rect -12322 -20803 -12222 -20781
rect -12322 -20849 -12289 -20803
rect -12255 -20849 -12222 -20803
rect -12322 -20875 -12222 -20849
rect -12322 -20917 -12289 -20875
rect -12255 -20917 -12222 -20875
rect -12322 -20947 -12222 -20917
rect -12322 -20985 -12289 -20947
rect -12255 -20985 -12222 -20947
rect -12322 -21019 -12222 -20985
rect 2580 -20429 2614 -20394
rect 2580 -20501 2614 -20477
rect 2580 -20573 2614 -20545
rect 2580 -20645 2614 -20613
rect 2580 -20715 2614 -20681
rect 2580 -20783 2614 -20751
rect 2580 -20851 2614 -20823
rect 2580 -20919 2614 -20895
rect 2580 -21002 2614 -20967
rect 3598 -20429 3632 -20394
rect 3598 -20501 3632 -20477
rect 3598 -20573 3632 -20545
rect 3598 -20645 3632 -20613
rect 3598 -20715 3632 -20681
rect 3598 -20783 3632 -20751
rect 3598 -20851 3632 -20823
rect 3598 -20919 3632 -20895
rect 3598 -21002 3632 -20967
rect 4616 -20429 4650 -20394
rect 4616 -20501 4650 -20477
rect 4616 -20573 4650 -20545
rect 4616 -20645 4650 -20613
rect 4616 -20715 4650 -20681
rect 4616 -20783 4650 -20751
rect 4616 -20851 4650 -20823
rect 4616 -20919 4650 -20895
rect 4616 -21002 4650 -20967
rect 5634 -20429 5668 -20394
rect 5634 -20501 5668 -20477
rect 5634 -20573 5668 -20545
rect 5634 -20645 5668 -20613
rect 5634 -20715 5668 -20681
rect 5634 -20783 5668 -20751
rect 5634 -20851 5668 -20823
rect 5634 -20919 5668 -20895
rect 5634 -21002 5668 -20967
rect 6652 -20429 6686 -20394
rect 6652 -20501 6686 -20477
rect 6652 -20573 6686 -20545
rect 6652 -20645 6686 -20613
rect 6652 -20715 6686 -20681
rect 6652 -20783 6686 -20751
rect 6652 -20851 6686 -20823
rect 6652 -20919 6686 -20895
rect 6652 -21002 6686 -20967
rect 7670 -20429 7704 -20394
rect 7670 -20501 7704 -20477
rect 7670 -20573 7704 -20545
rect 7670 -20645 7704 -20613
rect 7670 -20715 7704 -20681
rect 7670 -20783 7704 -20751
rect 7670 -20851 7704 -20823
rect 7670 -20919 7704 -20895
rect 7670 -21002 7704 -20967
rect 8688 -20429 8722 -20394
rect 8688 -20501 8722 -20477
rect 8688 -20573 8722 -20545
rect 8688 -20645 8722 -20613
rect 8688 -20715 8722 -20681
rect 8688 -20783 8722 -20751
rect 8688 -20851 8722 -20823
rect 8688 -20919 8722 -20895
rect 8688 -21002 8722 -20967
rect 9706 -20429 9740 -20394
rect 9706 -20501 9740 -20477
rect 9706 -20573 9740 -20545
rect 9706 -20645 9740 -20613
rect 9706 -20715 9740 -20681
rect 9706 -20783 9740 -20751
rect 9706 -20851 9740 -20823
rect 9706 -20919 9740 -20895
rect 9706 -21002 9740 -20967
rect 10724 -20429 10758 -20394
rect 10724 -20501 10758 -20477
rect 10724 -20573 10758 -20545
rect 10724 -20645 10758 -20613
rect 10724 -20715 10758 -20681
rect 10724 -20783 10758 -20751
rect 10724 -20851 10758 -20823
rect 10724 -20919 10758 -20895
rect 10724 -21002 10758 -20967
rect 11742 -20429 11776 -20394
rect 11742 -20501 11776 -20477
rect 11742 -20573 11776 -20545
rect 11742 -20645 11776 -20613
rect 11742 -20715 11776 -20681
rect 11742 -20783 11776 -20751
rect 11742 -20851 11776 -20823
rect 11742 -20919 11776 -20895
rect 11742 -21002 11776 -20967
rect 12760 -20429 12794 -20394
rect 12760 -20501 12794 -20477
rect 12760 -20573 12794 -20545
rect 12760 -20645 12794 -20613
rect 12760 -20715 12794 -20681
rect 12760 -20783 12794 -20751
rect 12760 -20851 12794 -20823
rect 12760 -20919 12794 -20895
rect 12760 -21002 12794 -20967
rect 13778 -20429 13812 -20394
rect 13778 -20501 13812 -20477
rect 13778 -20573 13812 -20545
rect 13778 -20645 13812 -20613
rect 13778 -20715 13812 -20681
rect 13778 -20783 13812 -20751
rect 13778 -20851 13812 -20823
rect 13778 -20919 13812 -20895
rect 13778 -21002 13812 -20967
rect 14796 -20429 14830 -20394
rect 14796 -20501 14830 -20477
rect 14796 -20573 14830 -20545
rect 14796 -20645 14830 -20613
rect 14796 -20715 14830 -20681
rect 14796 -20783 14830 -20751
rect 14796 -20851 14830 -20823
rect 14796 -20919 14830 -20895
rect 14796 -21002 14830 -20967
rect 15814 -20429 15848 -20394
rect 15814 -20501 15848 -20477
rect 15814 -20573 15848 -20545
rect 15814 -20645 15848 -20613
rect 15814 -20715 15848 -20681
rect 15814 -20783 15848 -20751
rect 15814 -20851 15848 -20823
rect 15814 -20919 15848 -20895
rect 15814 -21002 15848 -20967
rect 16832 -20429 16866 -20394
rect 16832 -20501 16866 -20477
rect 16832 -20573 16866 -20545
rect 16832 -20645 16866 -20613
rect 16832 -20715 16866 -20681
rect 16832 -20783 16866 -20751
rect 16832 -20851 16866 -20823
rect 16832 -20919 16866 -20895
rect 16832 -21002 16866 -20967
rect 17850 -20429 17884 -20394
rect 17850 -20501 17884 -20477
rect 17850 -20573 17884 -20545
rect 17850 -20645 17884 -20613
rect 17850 -20715 17884 -20681
rect 17850 -20783 17884 -20751
rect 17850 -20851 17884 -20823
rect 17850 -20919 17884 -20895
rect 17850 -21002 17884 -20967
rect 18868 -20429 18902 -20394
rect 18868 -20501 18902 -20477
rect 18868 -20573 18902 -20545
rect 18868 -20645 18902 -20613
rect 18868 -20715 18902 -20681
rect 18868 -20783 18902 -20751
rect 18868 -20851 18902 -20823
rect 18868 -20919 18902 -20895
rect 18868 -21002 18902 -20967
rect 19886 -20429 19920 -20394
rect 19886 -20501 19920 -20477
rect 19886 -20573 19920 -20545
rect 19886 -20645 19920 -20613
rect 19886 -20715 19920 -20681
rect 19886 -20783 19920 -20751
rect 19886 -20851 19920 -20823
rect 19886 -20919 19920 -20895
rect 19886 -21002 19920 -20967
rect 20904 -20429 20938 -20394
rect 20904 -20501 20938 -20477
rect 20904 -20573 20938 -20545
rect 20904 -20645 20938 -20613
rect 20904 -20715 20938 -20681
rect 20904 -20783 20938 -20751
rect 20904 -20851 20938 -20823
rect 20904 -20919 20938 -20895
rect 20904 -21002 20938 -20967
rect 21922 -20429 21956 -20394
rect 21922 -20501 21956 -20477
rect 21922 -20573 21956 -20545
rect 21922 -20645 21956 -20613
rect 21922 -20715 21956 -20681
rect 21922 -20783 21956 -20751
rect 21922 -20851 21956 -20823
rect 21922 -20919 21956 -20895
rect 21922 -21002 21956 -20967
rect 22940 -20429 22974 -20394
rect 22940 -20501 22974 -20477
rect 22940 -20573 22974 -20545
rect 22940 -20645 22974 -20613
rect 22940 -20715 22974 -20681
rect 22940 -20783 22974 -20751
rect 22940 -20851 22974 -20823
rect 22940 -20919 22974 -20895
rect 22940 -21002 22974 -20967
rect 24822 -20405 24855 -20339
rect 24889 -20405 24922 -20339
rect 24822 -20407 24922 -20405
rect 24822 -20441 24855 -20407
rect 24889 -20441 24922 -20407
rect 24822 -20443 24922 -20441
rect 24822 -20509 24855 -20443
rect 24889 -20509 24922 -20443
rect 24822 -20515 24922 -20509
rect 24822 -20577 24855 -20515
rect 24889 -20577 24922 -20515
rect 24822 -20587 24922 -20577
rect 24822 -20645 24855 -20587
rect 24889 -20645 24922 -20587
rect 24822 -20659 24922 -20645
rect 24822 -20713 24855 -20659
rect 24889 -20713 24922 -20659
rect 24822 -20731 24922 -20713
rect 24822 -20781 24855 -20731
rect 24889 -20781 24922 -20731
rect 24822 -20803 24922 -20781
rect 24822 -20849 24855 -20803
rect 24889 -20849 24922 -20803
rect 24822 -20875 24922 -20849
rect 24822 -20917 24855 -20875
rect 24889 -20917 24922 -20875
rect 24822 -20947 24922 -20917
rect 24822 -20985 24855 -20947
rect 24889 -20985 24922 -20947
rect -12322 -21053 -12289 -21019
rect -12255 -21053 -12222 -21019
rect 24822 -21019 24922 -20985
rect 5106 -21036 5166 -21032
rect -12322 -21087 -12222 -21053
rect 2812 -21070 2851 -21036
rect 2885 -21070 2909 -21036
rect 2953 -21070 2981 -21036
rect 3021 -21070 3053 -21036
rect 3089 -21070 3123 -21036
rect 3159 -21070 3191 -21036
rect 3231 -21070 3259 -21036
rect 3303 -21070 3327 -21036
rect 3361 -21070 3400 -21036
rect 3830 -21070 3869 -21036
rect 3903 -21070 3927 -21036
rect 3971 -21070 3999 -21036
rect 4039 -21070 4071 -21036
rect 4107 -21070 4141 -21036
rect 4177 -21070 4209 -21036
rect 4249 -21070 4277 -21036
rect 4321 -21070 4345 -21036
rect 4379 -21070 4418 -21036
rect 4848 -21070 4887 -21036
rect 4921 -21070 4945 -21036
rect 4989 -21070 5017 -21036
rect 5057 -21070 5089 -21036
rect 5125 -21070 5159 -21036
rect 5195 -21070 5227 -21036
rect 5267 -21070 5295 -21036
rect 5339 -21070 5363 -21036
rect 5397 -21070 5436 -21036
rect 5866 -21070 5905 -21036
rect 5939 -21070 5963 -21036
rect 6007 -21070 6035 -21036
rect 6075 -21070 6107 -21036
rect 6143 -21070 6177 -21036
rect 6213 -21070 6245 -21036
rect 6285 -21070 6313 -21036
rect 6357 -21070 6381 -21036
rect 6415 -21070 6454 -21036
rect 6884 -21070 6923 -21036
rect 6957 -21070 6981 -21036
rect 7025 -21070 7053 -21036
rect 7093 -21070 7125 -21036
rect 7161 -21070 7195 -21036
rect 7231 -21070 7263 -21036
rect 7303 -21070 7331 -21036
rect 7375 -21070 7399 -21036
rect 7433 -21070 7472 -21036
rect 7902 -21070 7941 -21036
rect 7975 -21070 7999 -21036
rect 8043 -21070 8071 -21036
rect 8111 -21070 8143 -21036
rect 8179 -21070 8213 -21036
rect 8249 -21070 8281 -21036
rect 8321 -21070 8349 -21036
rect 8393 -21070 8417 -21036
rect 8451 -21070 8490 -21036
rect 8920 -21070 8959 -21036
rect 8993 -21070 9017 -21036
rect 9061 -21070 9089 -21036
rect 9129 -21070 9161 -21036
rect 9197 -21070 9231 -21036
rect 9267 -21070 9299 -21036
rect 9339 -21070 9367 -21036
rect 9411 -21070 9435 -21036
rect 9469 -21070 9508 -21036
rect 9938 -21070 9977 -21036
rect 10011 -21070 10035 -21036
rect 10079 -21070 10107 -21036
rect 10147 -21070 10179 -21036
rect 10215 -21070 10249 -21036
rect 10285 -21070 10317 -21036
rect 10357 -21070 10385 -21036
rect 10429 -21070 10453 -21036
rect 10487 -21070 10526 -21036
rect 10956 -21070 10995 -21036
rect 11029 -21070 11053 -21036
rect 11097 -21070 11125 -21036
rect 11165 -21070 11197 -21036
rect 11233 -21070 11267 -21036
rect 11303 -21070 11335 -21036
rect 11375 -21070 11403 -21036
rect 11447 -21070 11471 -21036
rect 11505 -21070 11544 -21036
rect 11974 -21070 12013 -21036
rect 12047 -21070 12071 -21036
rect 12115 -21070 12143 -21036
rect 12183 -21070 12215 -21036
rect 12251 -21070 12285 -21036
rect 12321 -21070 12353 -21036
rect 12393 -21070 12421 -21036
rect 12465 -21070 12489 -21036
rect 12523 -21070 12562 -21036
rect 12992 -21070 13031 -21036
rect 13065 -21070 13089 -21036
rect 13133 -21070 13161 -21036
rect 13201 -21070 13233 -21036
rect 13269 -21070 13303 -21036
rect 13339 -21070 13371 -21036
rect 13411 -21070 13439 -21036
rect 13483 -21070 13507 -21036
rect 13541 -21070 13580 -21036
rect 14010 -21070 14049 -21036
rect 14083 -21070 14107 -21036
rect 14151 -21070 14179 -21036
rect 14219 -21070 14251 -21036
rect 14287 -21070 14321 -21036
rect 14357 -21070 14389 -21036
rect 14429 -21070 14457 -21036
rect 14501 -21070 14525 -21036
rect 14559 -21070 14598 -21036
rect 15028 -21070 15067 -21036
rect 15101 -21070 15125 -21036
rect 15169 -21070 15197 -21036
rect 15237 -21070 15269 -21036
rect 15305 -21070 15339 -21036
rect 15375 -21070 15407 -21036
rect 15447 -21070 15475 -21036
rect 15519 -21070 15543 -21036
rect 15577 -21070 15616 -21036
rect 16046 -21070 16085 -21036
rect 16119 -21070 16143 -21036
rect 16187 -21070 16215 -21036
rect 16255 -21070 16287 -21036
rect 16323 -21070 16357 -21036
rect 16393 -21070 16425 -21036
rect 16465 -21070 16493 -21036
rect 16537 -21070 16561 -21036
rect 16595 -21070 16634 -21036
rect 17064 -21070 17103 -21036
rect 17137 -21070 17161 -21036
rect 17205 -21070 17233 -21036
rect 17273 -21070 17305 -21036
rect 17341 -21070 17375 -21036
rect 17411 -21070 17443 -21036
rect 17483 -21070 17511 -21036
rect 17555 -21070 17579 -21036
rect 17613 -21070 17652 -21036
rect 18082 -21070 18121 -21036
rect 18155 -21070 18179 -21036
rect 18223 -21070 18251 -21036
rect 18291 -21070 18323 -21036
rect 18359 -21070 18393 -21036
rect 18429 -21070 18461 -21036
rect 18501 -21070 18529 -21036
rect 18573 -21070 18597 -21036
rect 18631 -21070 18670 -21036
rect 19100 -21070 19139 -21036
rect 19173 -21070 19197 -21036
rect 19241 -21070 19269 -21036
rect 19309 -21070 19341 -21036
rect 19377 -21070 19411 -21036
rect 19447 -21070 19479 -21036
rect 19519 -21070 19547 -21036
rect 19591 -21070 19615 -21036
rect 19649 -21070 19688 -21036
rect 20118 -21070 20157 -21036
rect 20191 -21070 20215 -21036
rect 20259 -21070 20287 -21036
rect 20327 -21070 20359 -21036
rect 20395 -21070 20429 -21036
rect 20465 -21070 20497 -21036
rect 20537 -21070 20565 -21036
rect 20609 -21070 20633 -21036
rect 20667 -21070 20706 -21036
rect 21136 -21070 21175 -21036
rect 21209 -21070 21233 -21036
rect 21277 -21070 21305 -21036
rect 21345 -21070 21377 -21036
rect 21413 -21070 21447 -21036
rect 21483 -21070 21515 -21036
rect 21555 -21070 21583 -21036
rect 21627 -21070 21651 -21036
rect 21685 -21070 21724 -21036
rect 22154 -21070 22193 -21036
rect 22227 -21070 22251 -21036
rect 22295 -21070 22323 -21036
rect 22363 -21070 22395 -21036
rect 22431 -21070 22465 -21036
rect 22501 -21070 22533 -21036
rect 22573 -21070 22601 -21036
rect 22645 -21070 22669 -21036
rect 22703 -21070 22742 -21036
rect 24822 -21053 24855 -21019
rect 24889 -21053 24922 -21019
rect -12322 -21125 -12289 -21087
rect -12255 -21125 -12222 -21087
rect -12322 -21155 -12222 -21125
rect -12322 -21197 -12289 -21155
rect -12255 -21197 -12222 -21155
rect -12322 -21223 -12222 -21197
rect -12322 -21269 -12289 -21223
rect -12255 -21269 -12222 -21223
rect -12322 -21291 -12222 -21269
rect -12322 -21341 -12289 -21291
rect -12255 -21341 -12222 -21291
rect -12322 -21359 -12222 -21341
rect -12322 -21413 -12289 -21359
rect -12255 -21413 -12222 -21359
rect -12322 -21427 -12222 -21413
rect -12322 -21485 -12289 -21427
rect -12255 -21485 -12222 -21427
rect -12322 -21495 -12222 -21485
rect -12322 -21557 -12289 -21495
rect -12255 -21557 -12222 -21495
rect -12322 -21563 -12222 -21557
rect 24822 -21087 24922 -21053
rect 24822 -21125 24855 -21087
rect 24889 -21125 24922 -21087
rect 24822 -21155 24922 -21125
rect 24822 -21197 24855 -21155
rect 24889 -21197 24922 -21155
rect 24822 -21223 24922 -21197
rect 24822 -21269 24855 -21223
rect 24889 -21269 24922 -21223
rect 24822 -21291 24922 -21269
rect 24822 -21341 24855 -21291
rect 24889 -21341 24922 -21291
rect 24822 -21359 24922 -21341
rect 24822 -21413 24855 -21359
rect 24889 -21413 24922 -21359
rect 24822 -21427 24922 -21413
rect 24822 -21485 24855 -21427
rect 24889 -21485 24922 -21427
rect 24822 -21495 24922 -21485
rect 24822 -21557 24855 -21495
rect 24889 -21557 24922 -21495
rect -12322 -21629 -12289 -21563
rect -12255 -21629 -12222 -21563
rect 2812 -21594 2851 -21560
rect 2885 -21594 2909 -21560
rect 2953 -21594 2981 -21560
rect 3021 -21594 3053 -21560
rect 3089 -21594 3123 -21560
rect 3159 -21594 3191 -21560
rect 3231 -21594 3259 -21560
rect 3303 -21594 3327 -21560
rect 3361 -21594 3400 -21560
rect 3830 -21594 3869 -21560
rect 3903 -21594 3927 -21560
rect 3971 -21594 3999 -21560
rect 4039 -21594 4071 -21560
rect 4107 -21594 4141 -21560
rect 4177 -21594 4209 -21560
rect 4249 -21594 4277 -21560
rect 4321 -21594 4345 -21560
rect 4379 -21594 4418 -21560
rect 4848 -21594 4887 -21560
rect 4921 -21594 4945 -21560
rect 4989 -21594 5017 -21560
rect 5057 -21594 5089 -21560
rect 5125 -21594 5159 -21560
rect 5195 -21594 5227 -21560
rect 5267 -21594 5295 -21560
rect 5339 -21594 5363 -21560
rect 5397 -21594 5436 -21560
rect 5866 -21594 5905 -21560
rect 5939 -21594 5963 -21560
rect 6007 -21594 6035 -21560
rect 6075 -21594 6107 -21560
rect 6143 -21594 6177 -21560
rect 6213 -21594 6245 -21560
rect 6285 -21594 6313 -21560
rect 6357 -21594 6381 -21560
rect 6415 -21594 6454 -21560
rect 6884 -21594 6923 -21560
rect 6957 -21594 6981 -21560
rect 7025 -21594 7053 -21560
rect 7093 -21594 7125 -21560
rect 7161 -21594 7195 -21560
rect 7231 -21594 7263 -21560
rect 7303 -21594 7331 -21560
rect 7375 -21594 7399 -21560
rect 7433 -21594 7472 -21560
rect 7902 -21594 7941 -21560
rect 7975 -21594 7999 -21560
rect 8043 -21594 8071 -21560
rect 8111 -21594 8143 -21560
rect 8179 -21594 8213 -21560
rect 8249 -21594 8281 -21560
rect 8321 -21594 8349 -21560
rect 8393 -21594 8417 -21560
rect 8451 -21594 8490 -21560
rect 8920 -21594 8959 -21560
rect 8993 -21594 9017 -21560
rect 9061 -21594 9089 -21560
rect 9129 -21594 9161 -21560
rect 9197 -21594 9231 -21560
rect 9267 -21594 9299 -21560
rect 9339 -21594 9367 -21560
rect 9411 -21594 9435 -21560
rect 9469 -21594 9508 -21560
rect 9938 -21594 9977 -21560
rect 10011 -21594 10035 -21560
rect 10079 -21594 10107 -21560
rect 10147 -21594 10179 -21560
rect 10215 -21594 10249 -21560
rect 10285 -21594 10317 -21560
rect 10357 -21594 10385 -21560
rect 10429 -21594 10453 -21560
rect 10487 -21594 10526 -21560
rect 10956 -21594 10995 -21560
rect 11029 -21594 11053 -21560
rect 11097 -21594 11125 -21560
rect 11165 -21594 11197 -21560
rect 11233 -21594 11267 -21560
rect 11303 -21594 11335 -21560
rect 11375 -21594 11403 -21560
rect 11447 -21594 11471 -21560
rect 11505 -21594 11544 -21560
rect 11974 -21594 12013 -21560
rect 12047 -21594 12071 -21560
rect 12115 -21594 12143 -21560
rect 12183 -21594 12215 -21560
rect 12251 -21594 12285 -21560
rect 12321 -21594 12353 -21560
rect 12393 -21594 12421 -21560
rect 12465 -21594 12489 -21560
rect 12523 -21594 12562 -21560
rect 12992 -21594 13031 -21560
rect 13065 -21594 13089 -21560
rect 13133 -21594 13161 -21560
rect 13201 -21594 13233 -21560
rect 13269 -21594 13303 -21560
rect 13339 -21594 13371 -21560
rect 13411 -21594 13439 -21560
rect 13483 -21594 13507 -21560
rect 13541 -21594 13580 -21560
rect 14010 -21594 14049 -21560
rect 14083 -21594 14107 -21560
rect 14151 -21594 14179 -21560
rect 14219 -21594 14251 -21560
rect 14287 -21594 14321 -21560
rect 14357 -21594 14389 -21560
rect 14429 -21594 14457 -21560
rect 14501 -21594 14525 -21560
rect 14559 -21594 14598 -21560
rect 15028 -21594 15067 -21560
rect 15101 -21594 15125 -21560
rect 15169 -21594 15197 -21560
rect 15237 -21594 15269 -21560
rect 15305 -21594 15339 -21560
rect 15375 -21594 15407 -21560
rect 15447 -21594 15475 -21560
rect 15519 -21594 15543 -21560
rect 15577 -21594 15616 -21560
rect 16046 -21594 16085 -21560
rect 16119 -21594 16143 -21560
rect 16187 -21594 16215 -21560
rect 16255 -21594 16287 -21560
rect 16323 -21594 16357 -21560
rect 16393 -21594 16425 -21560
rect 16465 -21594 16493 -21560
rect 16537 -21594 16561 -21560
rect 16595 -21594 16634 -21560
rect 17064 -21594 17103 -21560
rect 17137 -21594 17161 -21560
rect 17205 -21594 17233 -21560
rect 17273 -21594 17305 -21560
rect 17341 -21594 17375 -21560
rect 17411 -21594 17443 -21560
rect 17483 -21594 17511 -21560
rect 17555 -21594 17579 -21560
rect 17613 -21594 17652 -21560
rect 18082 -21594 18121 -21560
rect 18155 -21594 18179 -21560
rect 18223 -21594 18251 -21560
rect 18291 -21594 18323 -21560
rect 18359 -21594 18393 -21560
rect 18429 -21594 18461 -21560
rect 18501 -21594 18529 -21560
rect 18573 -21594 18597 -21560
rect 18631 -21594 18670 -21560
rect 19100 -21594 19139 -21560
rect 19173 -21594 19197 -21560
rect 19241 -21594 19269 -21560
rect 19309 -21594 19341 -21560
rect 19377 -21594 19411 -21560
rect 19447 -21594 19479 -21560
rect 19519 -21594 19547 -21560
rect 19591 -21594 19615 -21560
rect 19649 -21594 19688 -21560
rect 20118 -21594 20157 -21560
rect 20191 -21594 20215 -21560
rect 20259 -21594 20287 -21560
rect 20327 -21594 20359 -21560
rect 20395 -21594 20429 -21560
rect 20465 -21594 20497 -21560
rect 20537 -21594 20565 -21560
rect 20609 -21594 20633 -21560
rect 20667 -21594 20706 -21560
rect 21136 -21594 21175 -21560
rect 21209 -21594 21233 -21560
rect 21277 -21594 21305 -21560
rect 21345 -21594 21377 -21560
rect 21413 -21594 21447 -21560
rect 21483 -21594 21515 -21560
rect 21555 -21594 21583 -21560
rect 21627 -21594 21651 -21560
rect 21685 -21594 21724 -21560
rect 22154 -21594 22193 -21560
rect 22227 -21594 22251 -21560
rect 22295 -21594 22323 -21560
rect 22363 -21594 22395 -21560
rect 22431 -21594 22465 -21560
rect 22501 -21594 22533 -21560
rect 22573 -21594 22601 -21560
rect 22645 -21594 22669 -21560
rect 22703 -21594 22742 -21560
rect 24822 -21563 24922 -21557
rect -12322 -21631 -12222 -21629
rect -12322 -21665 -12289 -21631
rect -12255 -21665 -12222 -21631
rect -12322 -21667 -12222 -21665
rect -12322 -21733 -12289 -21667
rect -12255 -21733 -12222 -21667
rect -12322 -21739 -12222 -21733
rect -12322 -21801 -12289 -21739
rect -12255 -21801 -12222 -21739
rect -12322 -21811 -12222 -21801
rect -12322 -21869 -12289 -21811
rect -12255 -21869 -12222 -21811
rect -12322 -21883 -12222 -21869
rect -12322 -21937 -12289 -21883
rect -12255 -21937 -12222 -21883
rect -12322 -21955 -12222 -21937
rect -12322 -22005 -12289 -21955
rect -12255 -22005 -12222 -21955
rect -12322 -22027 -12222 -22005
rect -12322 -22073 -12289 -22027
rect -12255 -22073 -12222 -22027
rect -12322 -22099 -12222 -22073
rect -12322 -22141 -12289 -22099
rect -12255 -22141 -12222 -22099
rect -12322 -22171 -12222 -22141
rect -12322 -22209 -12289 -22171
rect -12255 -22209 -12222 -22171
rect -12322 -22243 -12222 -22209
rect 2580 -21663 2614 -21628
rect 2580 -21735 2614 -21711
rect 2580 -21807 2614 -21779
rect 2580 -21879 2614 -21847
rect 2580 -21949 2614 -21915
rect 2580 -22017 2614 -21985
rect 2580 -22085 2614 -22057
rect 2580 -22153 2614 -22129
rect 2580 -22236 2614 -22201
rect 3598 -21663 3632 -21628
rect 3598 -21735 3632 -21711
rect 3598 -21807 3632 -21779
rect 3598 -21879 3632 -21847
rect 3598 -21949 3632 -21915
rect 3598 -22017 3632 -21985
rect 3598 -22085 3632 -22057
rect 3598 -22153 3632 -22129
rect 3598 -22236 3632 -22201
rect 4616 -21663 4650 -21628
rect 4616 -21735 4650 -21711
rect 4616 -21807 4650 -21779
rect 4616 -21879 4650 -21847
rect 4616 -21949 4650 -21915
rect 4616 -22017 4650 -21985
rect 4616 -22085 4650 -22057
rect 4616 -22153 4650 -22129
rect 4616 -22236 4650 -22201
rect 5634 -21663 5668 -21628
rect 5634 -21735 5668 -21711
rect 5634 -21807 5668 -21779
rect 5634 -21879 5668 -21847
rect 5634 -21949 5668 -21915
rect 5634 -22017 5668 -21985
rect 5634 -22085 5668 -22057
rect 5634 -22153 5668 -22129
rect 5634 -22236 5668 -22201
rect 6652 -21663 6686 -21628
rect 6652 -21735 6686 -21711
rect 6652 -21807 6686 -21779
rect 6652 -21879 6686 -21847
rect 6652 -21949 6686 -21915
rect 6652 -22017 6686 -21985
rect 6652 -22085 6686 -22057
rect 6652 -22153 6686 -22129
rect 6652 -22236 6686 -22201
rect 7670 -21663 7704 -21628
rect 7670 -21735 7704 -21711
rect 7670 -21807 7704 -21779
rect 7670 -21879 7704 -21847
rect 7670 -21949 7704 -21915
rect 7670 -22017 7704 -21985
rect 7670 -22085 7704 -22057
rect 7670 -22153 7704 -22129
rect 7670 -22236 7704 -22201
rect 8688 -21663 8722 -21628
rect 8688 -21735 8722 -21711
rect 8688 -21807 8722 -21779
rect 8688 -21879 8722 -21847
rect 8688 -21949 8722 -21915
rect 8688 -22017 8722 -21985
rect 8688 -22085 8722 -22057
rect 8688 -22153 8722 -22129
rect 8688 -22236 8722 -22201
rect 9706 -21663 9740 -21628
rect 9706 -21735 9740 -21711
rect 9706 -21807 9740 -21779
rect 9706 -21879 9740 -21847
rect 9706 -21949 9740 -21915
rect 9706 -22017 9740 -21985
rect 9706 -22085 9740 -22057
rect 9706 -22153 9740 -22129
rect 9706 -22236 9740 -22201
rect 10724 -21663 10758 -21628
rect 10724 -21735 10758 -21711
rect 10724 -21807 10758 -21779
rect 10724 -21879 10758 -21847
rect 10724 -21949 10758 -21915
rect 10724 -22017 10758 -21985
rect 10724 -22085 10758 -22057
rect 10724 -22153 10758 -22129
rect 10724 -22236 10758 -22201
rect 11742 -21663 11776 -21628
rect 11742 -21735 11776 -21711
rect 11742 -21807 11776 -21779
rect 11742 -21879 11776 -21847
rect 11742 -21949 11776 -21915
rect 11742 -22017 11776 -21985
rect 11742 -22085 11776 -22057
rect 11742 -22153 11776 -22129
rect 11742 -22236 11776 -22201
rect 12760 -21663 12794 -21628
rect 12760 -21735 12794 -21711
rect 12760 -21807 12794 -21779
rect 12760 -21879 12794 -21847
rect 12760 -21949 12794 -21915
rect 12760 -22017 12794 -21985
rect 12760 -22085 12794 -22057
rect 12760 -22153 12794 -22129
rect 12760 -22236 12794 -22201
rect 13778 -21663 13812 -21628
rect 13778 -21735 13812 -21711
rect 13778 -21807 13812 -21779
rect 13778 -21879 13812 -21847
rect 13778 -21949 13812 -21915
rect 13778 -22017 13812 -21985
rect 13778 -22085 13812 -22057
rect 13778 -22153 13812 -22129
rect 13778 -22236 13812 -22201
rect 14796 -21663 14830 -21628
rect 14796 -21735 14830 -21711
rect 14796 -21807 14830 -21779
rect 14796 -21879 14830 -21847
rect 14796 -21949 14830 -21915
rect 14796 -22017 14830 -21985
rect 14796 -22085 14830 -22057
rect 14796 -22153 14830 -22129
rect 14796 -22236 14830 -22201
rect 15814 -21663 15848 -21628
rect 15814 -21735 15848 -21711
rect 15814 -21807 15848 -21779
rect 15814 -21879 15848 -21847
rect 15814 -21949 15848 -21915
rect 15814 -22017 15848 -21985
rect 15814 -22085 15848 -22057
rect 15814 -22153 15848 -22129
rect 15814 -22236 15848 -22201
rect 16832 -21663 16866 -21628
rect 16832 -21735 16866 -21711
rect 16832 -21807 16866 -21779
rect 16832 -21879 16866 -21847
rect 16832 -21949 16866 -21915
rect 16832 -22017 16866 -21985
rect 16832 -22085 16866 -22057
rect 16832 -22153 16866 -22129
rect 16832 -22236 16866 -22201
rect 17850 -21663 17884 -21628
rect 17850 -21735 17884 -21711
rect 17850 -21807 17884 -21779
rect 17850 -21879 17884 -21847
rect 17850 -21949 17884 -21915
rect 17850 -22017 17884 -21985
rect 17850 -22085 17884 -22057
rect 17850 -22153 17884 -22129
rect 17850 -22236 17884 -22201
rect 18868 -21663 18902 -21628
rect 18868 -21735 18902 -21711
rect 18868 -21807 18902 -21779
rect 18868 -21879 18902 -21847
rect 18868 -21949 18902 -21915
rect 18868 -22017 18902 -21985
rect 18868 -22085 18902 -22057
rect 18868 -22153 18902 -22129
rect 18868 -22236 18902 -22201
rect 19886 -21663 19920 -21628
rect 19886 -21735 19920 -21711
rect 19886 -21807 19920 -21779
rect 19886 -21879 19920 -21847
rect 19886 -21949 19920 -21915
rect 19886 -22017 19920 -21985
rect 19886 -22085 19920 -22057
rect 19886 -22153 19920 -22129
rect 19886 -22236 19920 -22201
rect 20904 -21663 20938 -21628
rect 20904 -21735 20938 -21711
rect 20904 -21807 20938 -21779
rect 20904 -21879 20938 -21847
rect 20904 -21949 20938 -21915
rect 20904 -22017 20938 -21985
rect 20904 -22085 20938 -22057
rect 20904 -22153 20938 -22129
rect 20904 -22236 20938 -22201
rect 21922 -21663 21956 -21628
rect 21922 -21735 21956 -21711
rect 21922 -21807 21956 -21779
rect 21922 -21879 21956 -21847
rect 21922 -21949 21956 -21915
rect 21922 -22017 21956 -21985
rect 21922 -22085 21956 -22057
rect 21922 -22153 21956 -22129
rect 21922 -22236 21956 -22201
rect 22940 -21663 22974 -21628
rect 22940 -21735 22974 -21711
rect 22940 -21807 22974 -21779
rect 22940 -21879 22974 -21847
rect 22940 -21949 22974 -21915
rect 22940 -22017 22974 -21985
rect 22940 -22085 22974 -22057
rect 22940 -22153 22974 -22129
rect 22940 -22236 22974 -22201
rect 24822 -21629 24855 -21563
rect 24889 -21629 24922 -21563
rect 24822 -21631 24922 -21629
rect 24822 -21665 24855 -21631
rect 24889 -21665 24922 -21631
rect 24822 -21667 24922 -21665
rect 24822 -21733 24855 -21667
rect 24889 -21733 24922 -21667
rect 24822 -21739 24922 -21733
rect 24822 -21801 24855 -21739
rect 24889 -21801 24922 -21739
rect 24822 -21811 24922 -21801
rect 24822 -21869 24855 -21811
rect 24889 -21869 24922 -21811
rect 24822 -21883 24922 -21869
rect 24822 -21937 24855 -21883
rect 24889 -21937 24922 -21883
rect 24822 -21955 24922 -21937
rect 24822 -22005 24855 -21955
rect 24889 -22005 24922 -21955
rect 24822 -22027 24922 -22005
rect 24822 -22073 24855 -22027
rect 24889 -22073 24922 -22027
rect 24822 -22099 24922 -22073
rect 24822 -22141 24855 -22099
rect 24889 -22141 24922 -22099
rect 24822 -22171 24922 -22141
rect 24822 -22209 24855 -22171
rect 24889 -22209 24922 -22171
rect -12322 -22277 -12289 -22243
rect -12255 -22277 -12222 -22243
rect 24822 -22243 24922 -22209
rect 11230 -22270 11290 -22268
rect 13274 -22270 13334 -22266
rect 16312 -22270 16372 -22266
rect -12322 -22311 -12222 -22277
rect 2812 -22304 2851 -22270
rect 2885 -22304 2909 -22270
rect 2953 -22304 2981 -22270
rect 3021 -22304 3053 -22270
rect 3089 -22304 3123 -22270
rect 3159 -22304 3191 -22270
rect 3231 -22304 3259 -22270
rect 3303 -22304 3327 -22270
rect 3361 -22304 3400 -22270
rect 3830 -22304 3869 -22270
rect 3903 -22304 3927 -22270
rect 3971 -22304 3999 -22270
rect 4039 -22304 4071 -22270
rect 4107 -22304 4141 -22270
rect 4177 -22304 4209 -22270
rect 4249 -22304 4277 -22270
rect 4321 -22304 4345 -22270
rect 4379 -22304 4418 -22270
rect 4848 -22304 4887 -22270
rect 4921 -22304 4945 -22270
rect 4989 -22304 5017 -22270
rect 5057 -22304 5089 -22270
rect 5125 -22304 5159 -22270
rect 5195 -22304 5227 -22270
rect 5267 -22304 5295 -22270
rect 5339 -22304 5363 -22270
rect 5397 -22304 5436 -22270
rect 5866 -22304 5905 -22270
rect 5939 -22304 5963 -22270
rect 6007 -22304 6035 -22270
rect 6075 -22304 6107 -22270
rect 6143 -22304 6177 -22270
rect 6213 -22304 6245 -22270
rect 6285 -22304 6313 -22270
rect 6357 -22304 6381 -22270
rect 6415 -22304 6454 -22270
rect 6884 -22304 6923 -22270
rect 6957 -22304 6981 -22270
rect 7025 -22304 7053 -22270
rect 7093 -22304 7125 -22270
rect 7161 -22304 7195 -22270
rect 7231 -22304 7263 -22270
rect 7303 -22304 7331 -22270
rect 7375 -22304 7399 -22270
rect 7433 -22304 7472 -22270
rect 7902 -22304 7941 -22270
rect 7975 -22304 7999 -22270
rect 8043 -22304 8071 -22270
rect 8111 -22304 8143 -22270
rect 8179 -22304 8213 -22270
rect 8249 -22304 8281 -22270
rect 8321 -22304 8349 -22270
rect 8393 -22304 8417 -22270
rect 8451 -22304 8490 -22270
rect 8920 -22304 8959 -22270
rect 8993 -22304 9017 -22270
rect 9061 -22304 9089 -22270
rect 9129 -22304 9161 -22270
rect 9197 -22304 9231 -22270
rect 9267 -22304 9299 -22270
rect 9339 -22304 9367 -22270
rect 9411 -22304 9435 -22270
rect 9469 -22304 9508 -22270
rect 9938 -22304 9977 -22270
rect 10011 -22304 10035 -22270
rect 10079 -22304 10107 -22270
rect 10147 -22304 10179 -22270
rect 10215 -22304 10249 -22270
rect 10285 -22304 10317 -22270
rect 10357 -22304 10385 -22270
rect 10429 -22304 10453 -22270
rect 10487 -22304 10526 -22270
rect 10956 -22304 10995 -22270
rect 11029 -22304 11053 -22270
rect 11097 -22304 11125 -22270
rect 11165 -22304 11197 -22270
rect 11233 -22304 11267 -22270
rect 11303 -22304 11335 -22270
rect 11375 -22304 11403 -22270
rect 11447 -22304 11471 -22270
rect 11505 -22304 11544 -22270
rect 11974 -22304 12013 -22270
rect 12047 -22304 12071 -22270
rect 12115 -22304 12143 -22270
rect 12183 -22304 12215 -22270
rect 12251 -22304 12285 -22270
rect 12321 -22304 12353 -22270
rect 12393 -22304 12421 -22270
rect 12465 -22304 12489 -22270
rect 12523 -22304 12562 -22270
rect 12992 -22304 13031 -22270
rect 13065 -22304 13089 -22270
rect 13133 -22304 13161 -22270
rect 13201 -22304 13233 -22270
rect 13269 -22304 13303 -22270
rect 13339 -22304 13371 -22270
rect 13411 -22304 13439 -22270
rect 13483 -22304 13507 -22270
rect 13541 -22304 13580 -22270
rect 14010 -22304 14049 -22270
rect 14083 -22304 14107 -22270
rect 14151 -22304 14179 -22270
rect 14219 -22304 14251 -22270
rect 14287 -22304 14321 -22270
rect 14357 -22304 14389 -22270
rect 14429 -22304 14457 -22270
rect 14501 -22304 14525 -22270
rect 14559 -22304 14598 -22270
rect 15028 -22304 15067 -22270
rect 15101 -22304 15125 -22270
rect 15169 -22304 15197 -22270
rect 15237 -22304 15269 -22270
rect 15305 -22304 15339 -22270
rect 15375 -22304 15407 -22270
rect 15447 -22304 15475 -22270
rect 15519 -22304 15543 -22270
rect 15577 -22304 15616 -22270
rect 16046 -22304 16085 -22270
rect 16119 -22304 16143 -22270
rect 16187 -22304 16215 -22270
rect 16255 -22304 16287 -22270
rect 16323 -22304 16357 -22270
rect 16393 -22304 16425 -22270
rect 16465 -22304 16493 -22270
rect 16537 -22304 16561 -22270
rect 16595 -22304 16634 -22270
rect 17064 -22304 17103 -22270
rect 17137 -22304 17161 -22270
rect 17205 -22304 17233 -22270
rect 17273 -22304 17305 -22270
rect 17341 -22304 17375 -22270
rect 17411 -22304 17443 -22270
rect 17483 -22304 17511 -22270
rect 17555 -22304 17579 -22270
rect 17613 -22304 17652 -22270
rect 18082 -22304 18121 -22270
rect 18155 -22304 18179 -22270
rect 18223 -22304 18251 -22270
rect 18291 -22304 18323 -22270
rect 18359 -22304 18393 -22270
rect 18429 -22304 18461 -22270
rect 18501 -22304 18529 -22270
rect 18573 -22304 18597 -22270
rect 18631 -22304 18670 -22270
rect 19100 -22304 19139 -22270
rect 19173 -22304 19197 -22270
rect 19241 -22304 19269 -22270
rect 19309 -22304 19341 -22270
rect 19377 -22304 19411 -22270
rect 19447 -22304 19479 -22270
rect 19519 -22304 19547 -22270
rect 19591 -22304 19615 -22270
rect 19649 -22304 19688 -22270
rect 20118 -22304 20157 -22270
rect 20191 -22304 20215 -22270
rect 20259 -22304 20287 -22270
rect 20327 -22304 20359 -22270
rect 20395 -22304 20429 -22270
rect 20465 -22304 20497 -22270
rect 20537 -22304 20565 -22270
rect 20609 -22304 20633 -22270
rect 20667 -22304 20706 -22270
rect 21136 -22304 21175 -22270
rect 21209 -22304 21233 -22270
rect 21277 -22304 21305 -22270
rect 21345 -22304 21377 -22270
rect 21413 -22304 21447 -22270
rect 21483 -22304 21515 -22270
rect 21555 -22304 21583 -22270
rect 21627 -22304 21651 -22270
rect 21685 -22304 21724 -22270
rect 22154 -22304 22193 -22270
rect 22227 -22304 22251 -22270
rect 22295 -22304 22323 -22270
rect 22363 -22304 22395 -22270
rect 22431 -22304 22465 -22270
rect 22501 -22304 22533 -22270
rect 22573 -22304 22601 -22270
rect 22645 -22304 22669 -22270
rect 22703 -22304 22742 -22270
rect 24822 -22277 24855 -22243
rect 24889 -22277 24922 -22243
rect -12322 -22349 -12289 -22311
rect -12255 -22349 -12222 -22311
rect -12322 -22379 -12222 -22349
rect -12322 -22421 -12289 -22379
rect -12255 -22421 -12222 -22379
rect -12322 -22447 -12222 -22421
rect -12322 -22493 -12289 -22447
rect -12255 -22493 -12222 -22447
rect -12322 -22515 -12222 -22493
rect -12322 -22565 -12289 -22515
rect -12255 -22565 -12222 -22515
rect -12322 -22583 -12222 -22565
rect -12322 -22637 -12289 -22583
rect -12255 -22637 -12222 -22583
rect -12322 -22651 -12222 -22637
rect -12322 -22709 -12289 -22651
rect -12255 -22709 -12222 -22651
rect -12322 -22719 -12222 -22709
rect -12322 -22781 -12289 -22719
rect -12255 -22781 -12222 -22719
rect -12322 -22787 -12222 -22781
rect -12322 -22853 -12289 -22787
rect -12255 -22853 -12222 -22787
rect 24822 -22311 24922 -22277
rect 24822 -22349 24855 -22311
rect 24889 -22349 24922 -22311
rect 24822 -22379 24922 -22349
rect 24822 -22421 24855 -22379
rect 24889 -22421 24922 -22379
rect 24822 -22447 24922 -22421
rect 24822 -22493 24855 -22447
rect 24889 -22493 24922 -22447
rect 24822 -22515 24922 -22493
rect 24822 -22565 24855 -22515
rect 24889 -22565 24922 -22515
rect 24822 -22583 24922 -22565
rect 24822 -22637 24855 -22583
rect 24889 -22637 24922 -22583
rect 24822 -22651 24922 -22637
rect 24822 -22709 24855 -22651
rect 24889 -22709 24922 -22651
rect 24822 -22719 24922 -22709
rect 24822 -22781 24855 -22719
rect 24889 -22781 24922 -22719
rect 24822 -22787 24922 -22781
rect 2812 -22826 2851 -22792
rect 2885 -22826 2909 -22792
rect 2953 -22826 2981 -22792
rect 3021 -22826 3053 -22792
rect 3089 -22826 3123 -22792
rect 3159 -22826 3191 -22792
rect 3231 -22826 3259 -22792
rect 3303 -22826 3327 -22792
rect 3361 -22826 3400 -22792
rect 3830 -22826 3869 -22792
rect 3903 -22826 3927 -22792
rect 3971 -22826 3999 -22792
rect 4039 -22826 4071 -22792
rect 4107 -22826 4141 -22792
rect 4177 -22826 4209 -22792
rect 4249 -22826 4277 -22792
rect 4321 -22826 4345 -22792
rect 4379 -22826 4418 -22792
rect 4848 -22826 4887 -22792
rect 4921 -22826 4945 -22792
rect 4989 -22826 5017 -22792
rect 5057 -22826 5089 -22792
rect 5125 -22826 5159 -22792
rect 5195 -22826 5227 -22792
rect 5267 -22826 5295 -22792
rect 5339 -22826 5363 -22792
rect 5397 -22826 5436 -22792
rect 5866 -22826 5905 -22792
rect 5939 -22826 5963 -22792
rect 6007 -22826 6035 -22792
rect 6075 -22826 6107 -22792
rect 6143 -22826 6177 -22792
rect 6213 -22826 6245 -22792
rect 6285 -22826 6313 -22792
rect 6357 -22826 6381 -22792
rect 6415 -22826 6454 -22792
rect 6884 -22826 6923 -22792
rect 6957 -22826 6981 -22792
rect 7025 -22826 7053 -22792
rect 7093 -22826 7125 -22792
rect 7161 -22826 7195 -22792
rect 7231 -22826 7263 -22792
rect 7303 -22826 7331 -22792
rect 7375 -22826 7399 -22792
rect 7433 -22826 7472 -22792
rect 7902 -22826 7941 -22792
rect 7975 -22826 7999 -22792
rect 8043 -22826 8071 -22792
rect 8111 -22826 8143 -22792
rect 8179 -22826 8213 -22792
rect 8249 -22826 8281 -22792
rect 8321 -22826 8349 -22792
rect 8393 -22826 8417 -22792
rect 8451 -22826 8490 -22792
rect 8920 -22826 8959 -22792
rect 8993 -22826 9017 -22792
rect 9061 -22826 9089 -22792
rect 9129 -22826 9161 -22792
rect 9197 -22826 9231 -22792
rect 9267 -22826 9299 -22792
rect 9339 -22826 9367 -22792
rect 9411 -22826 9435 -22792
rect 9469 -22826 9508 -22792
rect 9938 -22826 9977 -22792
rect 10011 -22826 10035 -22792
rect 10079 -22826 10107 -22792
rect 10147 -22826 10179 -22792
rect 10215 -22826 10249 -22792
rect 10285 -22826 10317 -22792
rect 10357 -22826 10385 -22792
rect 10429 -22826 10453 -22792
rect 10487 -22826 10526 -22792
rect 10956 -22826 10995 -22792
rect 11029 -22826 11053 -22792
rect 11097 -22826 11125 -22792
rect 11165 -22826 11197 -22792
rect 11233 -22826 11267 -22792
rect 11303 -22826 11335 -22792
rect 11375 -22826 11403 -22792
rect 11447 -22826 11471 -22792
rect 11505 -22826 11544 -22792
rect 11974 -22826 12013 -22792
rect 12047 -22826 12071 -22792
rect 12115 -22826 12143 -22792
rect 12183 -22826 12215 -22792
rect 12251 -22826 12285 -22792
rect 12321 -22826 12353 -22792
rect 12393 -22826 12421 -22792
rect 12465 -22826 12489 -22792
rect 12523 -22826 12562 -22792
rect 12992 -22826 13031 -22792
rect 13065 -22826 13089 -22792
rect 13133 -22826 13161 -22792
rect 13201 -22826 13233 -22792
rect 13269 -22826 13303 -22792
rect 13339 -22826 13371 -22792
rect 13411 -22826 13439 -22792
rect 13483 -22826 13507 -22792
rect 13541 -22826 13580 -22792
rect 14010 -22826 14049 -22792
rect 14083 -22826 14107 -22792
rect 14151 -22826 14179 -22792
rect 14219 -22826 14251 -22792
rect 14287 -22826 14321 -22792
rect 14357 -22826 14389 -22792
rect 14429 -22826 14457 -22792
rect 14501 -22826 14525 -22792
rect 14559 -22826 14598 -22792
rect 15028 -22826 15067 -22792
rect 15101 -22826 15125 -22792
rect 15169 -22826 15197 -22792
rect 15237 -22826 15269 -22792
rect 15305 -22826 15339 -22792
rect 15375 -22826 15407 -22792
rect 15447 -22826 15475 -22792
rect 15519 -22826 15543 -22792
rect 15577 -22826 15616 -22792
rect 16046 -22826 16085 -22792
rect 16119 -22826 16143 -22792
rect 16187 -22826 16215 -22792
rect 16255 -22826 16287 -22792
rect 16323 -22826 16357 -22792
rect 16393 -22826 16425 -22792
rect 16465 -22826 16493 -22792
rect 16537 -22826 16561 -22792
rect 16595 -22826 16634 -22792
rect 17064 -22826 17103 -22792
rect 17137 -22826 17161 -22792
rect 17205 -22826 17233 -22792
rect 17273 -22826 17305 -22792
rect 17341 -22826 17375 -22792
rect 17411 -22826 17443 -22792
rect 17483 -22826 17511 -22792
rect 17555 -22826 17579 -22792
rect 17613 -22826 17652 -22792
rect 18082 -22826 18121 -22792
rect 18155 -22826 18179 -22792
rect 18223 -22826 18251 -22792
rect 18291 -22826 18323 -22792
rect 18359 -22826 18393 -22792
rect 18429 -22826 18461 -22792
rect 18501 -22826 18529 -22792
rect 18573 -22826 18597 -22792
rect 18631 -22826 18670 -22792
rect 19100 -22826 19139 -22792
rect 19173 -22826 19197 -22792
rect 19241 -22826 19269 -22792
rect 19309 -22826 19341 -22792
rect 19377 -22826 19411 -22792
rect 19447 -22826 19479 -22792
rect 19519 -22826 19547 -22792
rect 19591 -22826 19615 -22792
rect 19649 -22826 19688 -22792
rect 20118 -22826 20157 -22792
rect 20191 -22826 20215 -22792
rect 20259 -22826 20287 -22792
rect 20327 -22826 20359 -22792
rect 20395 -22826 20429 -22792
rect 20465 -22826 20497 -22792
rect 20537 -22826 20565 -22792
rect 20609 -22826 20633 -22792
rect 20667 -22826 20706 -22792
rect 21136 -22826 21175 -22792
rect 21209 -22826 21233 -22792
rect 21277 -22826 21305 -22792
rect 21345 -22826 21377 -22792
rect 21413 -22826 21447 -22792
rect 21483 -22826 21515 -22792
rect 21555 -22826 21583 -22792
rect 21627 -22826 21651 -22792
rect 21685 -22826 21724 -22792
rect 22154 -22826 22193 -22792
rect 22227 -22826 22251 -22792
rect 22295 -22826 22323 -22792
rect 22363 -22826 22395 -22792
rect 22431 -22826 22465 -22792
rect 22501 -22826 22533 -22792
rect 22573 -22826 22601 -22792
rect 22645 -22826 22669 -22792
rect 22703 -22826 22742 -22792
rect 6134 -22828 6194 -22826
rect -12322 -22855 -12222 -22853
rect -12322 -22889 -12289 -22855
rect -12255 -22889 -12222 -22855
rect 24822 -22853 24855 -22787
rect 24889 -22853 24922 -22787
rect 24822 -22855 24922 -22853
rect -12322 -22891 -12222 -22889
rect -12322 -22957 -12289 -22891
rect -12255 -22957 -12222 -22891
rect -12322 -22963 -12222 -22957
rect -12322 -23025 -12289 -22963
rect -12255 -23025 -12222 -22963
rect -12322 -23035 -12222 -23025
rect -12322 -23093 -12289 -23035
rect -12255 -23093 -12222 -23035
rect -12322 -23107 -12222 -23093
rect -12322 -23161 -12289 -23107
rect -12255 -23161 -12222 -23107
rect -12322 -23179 -12222 -23161
rect -12322 -23229 -12289 -23179
rect -12255 -23229 -12222 -23179
rect -12322 -23251 -12222 -23229
rect -12322 -23297 -12289 -23251
rect -12255 -23297 -12222 -23251
rect -12322 -23323 -12222 -23297
rect -12322 -23365 -12289 -23323
rect -12255 -23365 -12222 -23323
rect -12322 -23395 -12222 -23365
rect -12322 -23433 -12289 -23395
rect -12255 -23433 -12222 -23395
rect -12322 -23467 -12222 -23433
rect -12322 -23501 -12289 -23467
rect -12255 -23501 -12222 -23467
rect 2580 -22895 2614 -22860
rect 2580 -22967 2614 -22943
rect 2580 -23039 2614 -23011
rect 2580 -23111 2614 -23079
rect 2580 -23181 2614 -23147
rect 2580 -23249 2614 -23217
rect 2580 -23317 2614 -23289
rect 2580 -23385 2614 -23361
rect 2580 -23468 2614 -23433
rect 3598 -22895 3632 -22860
rect 3598 -22967 3632 -22943
rect 3598 -23039 3632 -23011
rect 3598 -23111 3632 -23079
rect 3598 -23181 3632 -23147
rect 3598 -23249 3632 -23217
rect 3598 -23317 3632 -23289
rect 3598 -23385 3632 -23361
rect 3598 -23468 3632 -23433
rect 4616 -22895 4650 -22860
rect 4616 -22967 4650 -22943
rect 4616 -23039 4650 -23011
rect 4616 -23111 4650 -23079
rect 4616 -23181 4650 -23147
rect 4616 -23249 4650 -23217
rect 4616 -23317 4650 -23289
rect 4616 -23385 4650 -23361
rect 4616 -23468 4650 -23433
rect 5634 -22895 5668 -22860
rect 5634 -22967 5668 -22943
rect 5634 -23039 5668 -23011
rect 5634 -23111 5668 -23079
rect 5634 -23181 5668 -23147
rect 5634 -23249 5668 -23217
rect 5634 -23317 5668 -23289
rect 5634 -23385 5668 -23361
rect 5634 -23468 5668 -23433
rect 6652 -22895 6686 -22860
rect 6652 -22967 6686 -22943
rect 6652 -23039 6686 -23011
rect 6652 -23111 6686 -23079
rect 6652 -23181 6686 -23147
rect 6652 -23249 6686 -23217
rect 6652 -23317 6686 -23289
rect 6652 -23385 6686 -23361
rect 6652 -23468 6686 -23433
rect 7670 -22895 7704 -22860
rect 7670 -22967 7704 -22943
rect 7670 -23039 7704 -23011
rect 7670 -23111 7704 -23079
rect 7670 -23181 7704 -23147
rect 7670 -23249 7704 -23217
rect 7670 -23317 7704 -23289
rect 7670 -23385 7704 -23361
rect 7670 -23468 7704 -23433
rect 8688 -22895 8722 -22860
rect 8688 -22967 8722 -22943
rect 8688 -23039 8722 -23011
rect 8688 -23111 8722 -23079
rect 8688 -23181 8722 -23147
rect 8688 -23249 8722 -23217
rect 8688 -23317 8722 -23289
rect 8688 -23385 8722 -23361
rect 8688 -23468 8722 -23433
rect 9706 -22895 9740 -22860
rect 9706 -22967 9740 -22943
rect 9706 -23039 9740 -23011
rect 9706 -23111 9740 -23079
rect 9706 -23181 9740 -23147
rect 9706 -23249 9740 -23217
rect 9706 -23317 9740 -23289
rect 9706 -23385 9740 -23361
rect 9706 -23468 9740 -23433
rect 10724 -22895 10758 -22860
rect 10724 -22967 10758 -22943
rect 10724 -23039 10758 -23011
rect 10724 -23111 10758 -23079
rect 10724 -23181 10758 -23147
rect 10724 -23249 10758 -23217
rect 10724 -23317 10758 -23289
rect 10724 -23385 10758 -23361
rect 10724 -23468 10758 -23433
rect 11742 -22895 11776 -22860
rect 11742 -22967 11776 -22943
rect 11742 -23039 11776 -23011
rect 11742 -23111 11776 -23079
rect 11742 -23181 11776 -23147
rect 11742 -23249 11776 -23217
rect 11742 -23317 11776 -23289
rect 11742 -23385 11776 -23361
rect 11742 -23468 11776 -23433
rect 12760 -22895 12794 -22860
rect 12760 -22967 12794 -22943
rect 12760 -23039 12794 -23011
rect 12760 -23111 12794 -23079
rect 12760 -23181 12794 -23147
rect 12760 -23249 12794 -23217
rect 12760 -23317 12794 -23289
rect 12760 -23385 12794 -23361
rect 12760 -23468 12794 -23433
rect 13778 -22895 13812 -22860
rect 13778 -22967 13812 -22943
rect 13778 -23039 13812 -23011
rect 13778 -23111 13812 -23079
rect 13778 -23181 13812 -23147
rect 13778 -23249 13812 -23217
rect 13778 -23317 13812 -23289
rect 13778 -23385 13812 -23361
rect 13778 -23468 13812 -23433
rect 14796 -22895 14830 -22860
rect 14796 -22967 14830 -22943
rect 14796 -23039 14830 -23011
rect 14796 -23111 14830 -23079
rect 14796 -23181 14830 -23147
rect 14796 -23249 14830 -23217
rect 14796 -23317 14830 -23289
rect 14796 -23385 14830 -23361
rect 14796 -23468 14830 -23433
rect 15814 -22895 15848 -22860
rect 15814 -22967 15848 -22943
rect 15814 -23039 15848 -23011
rect 15814 -23111 15848 -23079
rect 15814 -23181 15848 -23147
rect 15814 -23249 15848 -23217
rect 15814 -23317 15848 -23289
rect 15814 -23385 15848 -23361
rect 15814 -23468 15848 -23433
rect 16832 -22895 16866 -22860
rect 16832 -22967 16866 -22943
rect 16832 -23039 16866 -23011
rect 16832 -23111 16866 -23079
rect 16832 -23181 16866 -23147
rect 16832 -23249 16866 -23217
rect 16832 -23317 16866 -23289
rect 16832 -23385 16866 -23361
rect 16832 -23468 16866 -23433
rect 17850 -22895 17884 -22860
rect 17850 -22967 17884 -22943
rect 17850 -23039 17884 -23011
rect 17850 -23111 17884 -23079
rect 17850 -23181 17884 -23147
rect 17850 -23249 17884 -23217
rect 17850 -23317 17884 -23289
rect 17850 -23385 17884 -23361
rect 17850 -23468 17884 -23433
rect 18868 -22895 18902 -22860
rect 18868 -22967 18902 -22943
rect 18868 -23039 18902 -23011
rect 18868 -23111 18902 -23079
rect 18868 -23181 18902 -23147
rect 18868 -23249 18902 -23217
rect 18868 -23317 18902 -23289
rect 18868 -23385 18902 -23361
rect 18868 -23468 18902 -23433
rect 19886 -22895 19920 -22860
rect 19886 -22967 19920 -22943
rect 19886 -23039 19920 -23011
rect 19886 -23111 19920 -23079
rect 19886 -23181 19920 -23147
rect 19886 -23249 19920 -23217
rect 19886 -23317 19920 -23289
rect 19886 -23385 19920 -23361
rect 19886 -23468 19920 -23433
rect 20904 -22895 20938 -22860
rect 20904 -22967 20938 -22943
rect 20904 -23039 20938 -23011
rect 20904 -23111 20938 -23079
rect 20904 -23181 20938 -23147
rect 20904 -23249 20938 -23217
rect 20904 -23317 20938 -23289
rect 20904 -23385 20938 -23361
rect 20904 -23468 20938 -23433
rect 21922 -22895 21956 -22860
rect 21922 -22967 21956 -22943
rect 21922 -23039 21956 -23011
rect 21922 -23111 21956 -23079
rect 21922 -23181 21956 -23147
rect 21922 -23249 21956 -23217
rect 21922 -23317 21956 -23289
rect 21922 -23385 21956 -23361
rect 21922 -23452 21956 -23433
rect 22940 -22895 22974 -22860
rect 22940 -22967 22974 -22943
rect 22940 -23039 22974 -23011
rect 22940 -23111 22974 -23079
rect 22940 -23181 22974 -23147
rect 22940 -23249 22974 -23217
rect 22940 -23317 22974 -23289
rect 22940 -23385 22974 -23361
rect 22940 -23468 22974 -23433
rect 24822 -22889 24855 -22855
rect 24889 -22889 24922 -22855
rect 24822 -22891 24922 -22889
rect 24822 -22957 24855 -22891
rect 24889 -22957 24922 -22891
rect 24822 -22963 24922 -22957
rect 24822 -23025 24855 -22963
rect 24889 -23025 24922 -22963
rect 24822 -23035 24922 -23025
rect 24822 -23093 24855 -23035
rect 24889 -23093 24922 -23035
rect 24822 -23107 24922 -23093
rect 24822 -23161 24855 -23107
rect 24889 -23161 24922 -23107
rect 24822 -23179 24922 -23161
rect 24822 -23229 24855 -23179
rect 24889 -23229 24922 -23179
rect 24822 -23251 24922 -23229
rect 24822 -23297 24855 -23251
rect 24889 -23297 24922 -23251
rect 24822 -23323 24922 -23297
rect 24822 -23365 24855 -23323
rect 24889 -23365 24922 -23323
rect 24822 -23395 24922 -23365
rect 24822 -23433 24855 -23395
rect 24889 -23433 24922 -23395
rect 24822 -23467 24922 -23433
rect -12322 -23535 -12222 -23501
rect 10206 -23502 10266 -23492
rect 24822 -23501 24855 -23467
rect 24889 -23501 24922 -23467
rect -12322 -23573 -12289 -23535
rect -12255 -23573 -12222 -23535
rect 2812 -23536 2851 -23502
rect 2885 -23536 2909 -23502
rect 2953 -23536 2981 -23502
rect 3021 -23536 3053 -23502
rect 3089 -23536 3123 -23502
rect 3159 -23536 3191 -23502
rect 3231 -23536 3259 -23502
rect 3303 -23536 3327 -23502
rect 3361 -23536 3400 -23502
rect 3830 -23536 3869 -23502
rect 3903 -23536 3927 -23502
rect 3971 -23536 3999 -23502
rect 4039 -23536 4071 -23502
rect 4107 -23536 4141 -23502
rect 4177 -23536 4209 -23502
rect 4249 -23536 4277 -23502
rect 4321 -23536 4345 -23502
rect 4379 -23536 4418 -23502
rect 4848 -23536 4887 -23502
rect 4921 -23536 4945 -23502
rect 4989 -23536 5017 -23502
rect 5057 -23536 5089 -23502
rect 5125 -23536 5159 -23502
rect 5195 -23536 5227 -23502
rect 5267 -23536 5295 -23502
rect 5339 -23536 5363 -23502
rect 5397 -23536 5436 -23502
rect 5866 -23536 5905 -23502
rect 5939 -23536 5963 -23502
rect 6007 -23536 6035 -23502
rect 6075 -23536 6107 -23502
rect 6143 -23536 6177 -23502
rect 6213 -23536 6245 -23502
rect 6285 -23536 6313 -23502
rect 6357 -23536 6381 -23502
rect 6415 -23536 6454 -23502
rect 6884 -23536 6923 -23502
rect 6957 -23536 6981 -23502
rect 7025 -23536 7053 -23502
rect 7093 -23536 7125 -23502
rect 7161 -23536 7195 -23502
rect 7231 -23536 7263 -23502
rect 7303 -23536 7331 -23502
rect 7375 -23536 7399 -23502
rect 7433 -23536 7472 -23502
rect 7902 -23536 7941 -23502
rect 7975 -23536 7999 -23502
rect 8043 -23536 8071 -23502
rect 8111 -23536 8143 -23502
rect 8179 -23536 8213 -23502
rect 8249 -23536 8281 -23502
rect 8321 -23536 8349 -23502
rect 8393 -23536 8417 -23502
rect 8451 -23536 8490 -23502
rect 8920 -23536 8959 -23502
rect 8993 -23536 9017 -23502
rect 9061 -23536 9089 -23502
rect 9129 -23536 9161 -23502
rect 9197 -23536 9231 -23502
rect 9267 -23536 9299 -23502
rect 9339 -23536 9367 -23502
rect 9411 -23536 9435 -23502
rect 9469 -23536 9508 -23502
rect 9938 -23536 9977 -23502
rect 10011 -23536 10035 -23502
rect 10079 -23536 10107 -23502
rect 10147 -23536 10179 -23502
rect 10215 -23536 10249 -23502
rect 10285 -23536 10317 -23502
rect 10357 -23536 10385 -23502
rect 10429 -23536 10453 -23502
rect 10487 -23536 10526 -23502
rect 10956 -23536 10995 -23502
rect 11029 -23536 11053 -23502
rect 11097 -23536 11125 -23502
rect 11165 -23536 11197 -23502
rect 11233 -23536 11267 -23502
rect 11303 -23536 11335 -23502
rect 11375 -23536 11403 -23502
rect 11447 -23536 11471 -23502
rect 11505 -23536 11544 -23502
rect 11974 -23536 12013 -23502
rect 12047 -23536 12071 -23502
rect 12115 -23536 12143 -23502
rect 12183 -23536 12215 -23502
rect 12251 -23536 12285 -23502
rect 12321 -23536 12353 -23502
rect 12393 -23536 12421 -23502
rect 12465 -23536 12489 -23502
rect 12523 -23536 12562 -23502
rect 12992 -23536 13031 -23502
rect 13065 -23536 13089 -23502
rect 13133 -23536 13161 -23502
rect 13201 -23536 13233 -23502
rect 13269 -23536 13303 -23502
rect 13339 -23536 13371 -23502
rect 13411 -23536 13439 -23502
rect 13483 -23536 13507 -23502
rect 13541 -23536 13580 -23502
rect 14010 -23536 14049 -23502
rect 14083 -23536 14107 -23502
rect 14151 -23536 14179 -23502
rect 14219 -23536 14251 -23502
rect 14287 -23536 14321 -23502
rect 14357 -23536 14389 -23502
rect 14429 -23536 14457 -23502
rect 14501 -23536 14525 -23502
rect 14559 -23536 14598 -23502
rect 15028 -23536 15067 -23502
rect 15101 -23536 15125 -23502
rect 15169 -23536 15197 -23502
rect 15237 -23536 15269 -23502
rect 15305 -23536 15339 -23502
rect 15375 -23536 15407 -23502
rect 15447 -23536 15475 -23502
rect 15519 -23536 15543 -23502
rect 15577 -23536 15616 -23502
rect 16046 -23536 16085 -23502
rect 16119 -23536 16143 -23502
rect 16187 -23536 16215 -23502
rect 16255 -23536 16287 -23502
rect 16323 -23536 16357 -23502
rect 16393 -23536 16425 -23502
rect 16465 -23536 16493 -23502
rect 16537 -23536 16561 -23502
rect 16595 -23536 16634 -23502
rect 17064 -23536 17103 -23502
rect 17137 -23536 17161 -23502
rect 17205 -23536 17233 -23502
rect 17273 -23536 17305 -23502
rect 17341 -23536 17375 -23502
rect 17411 -23536 17443 -23502
rect 17483 -23536 17511 -23502
rect 17555 -23536 17579 -23502
rect 17613 -23536 17652 -23502
rect 18082 -23536 18121 -23502
rect 18155 -23536 18179 -23502
rect 18223 -23536 18251 -23502
rect 18291 -23536 18323 -23502
rect 18359 -23536 18393 -23502
rect 18429 -23536 18461 -23502
rect 18501 -23536 18529 -23502
rect 18573 -23536 18597 -23502
rect 18631 -23536 18670 -23502
rect 19100 -23536 19139 -23502
rect 19173 -23536 19197 -23502
rect 19241 -23536 19269 -23502
rect 19309 -23536 19341 -23502
rect 19377 -23536 19411 -23502
rect 19447 -23536 19479 -23502
rect 19519 -23536 19547 -23502
rect 19591 -23536 19615 -23502
rect 19649 -23536 19688 -23502
rect 20118 -23536 20157 -23502
rect 20191 -23536 20215 -23502
rect 20259 -23536 20287 -23502
rect 20327 -23536 20359 -23502
rect 20395 -23536 20429 -23502
rect 20465 -23536 20497 -23502
rect 20537 -23536 20565 -23502
rect 20609 -23536 20633 -23502
rect 20667 -23536 20706 -23502
rect 21136 -23536 21175 -23502
rect 21209 -23536 21233 -23502
rect 21277 -23536 21305 -23502
rect 21345 -23536 21377 -23502
rect 21413 -23536 21447 -23502
rect 21483 -23536 21515 -23502
rect 21555 -23536 21583 -23502
rect 21627 -23536 21651 -23502
rect 21685 -23536 21724 -23502
rect 22154 -23536 22193 -23502
rect 22227 -23536 22251 -23502
rect 22295 -23536 22323 -23502
rect 22363 -23536 22395 -23502
rect 22431 -23536 22465 -23502
rect 22501 -23536 22533 -23502
rect 22573 -23536 22601 -23502
rect 22645 -23536 22669 -23502
rect 22703 -23536 22742 -23502
rect 24822 -23535 24922 -23501
rect -12322 -23603 -12222 -23573
rect -12322 -23645 -12289 -23603
rect -12255 -23645 -12222 -23603
rect -12322 -23671 -12222 -23645
rect -12322 -23717 -12289 -23671
rect -12255 -23717 -12222 -23671
rect -12322 -23739 -12222 -23717
rect -12322 -23789 -12289 -23739
rect -12255 -23789 -12222 -23739
rect -12322 -23807 -12222 -23789
rect -12322 -23861 -12289 -23807
rect -12255 -23861 -12222 -23807
rect -12322 -23875 -12222 -23861
rect -12322 -23933 -12289 -23875
rect -12255 -23933 -12222 -23875
rect -12322 -23943 -12222 -23933
rect -12322 -24005 -12289 -23943
rect -12255 -24005 -12222 -23943
rect -12322 -24011 -12222 -24005
rect -12322 -24077 -12289 -24011
rect -12255 -24077 -12222 -24011
rect 24822 -23573 24855 -23535
rect 24889 -23573 24922 -23535
rect 24822 -23603 24922 -23573
rect 24822 -23645 24855 -23603
rect 24889 -23645 24922 -23603
rect 24822 -23671 24922 -23645
rect 24822 -23717 24855 -23671
rect 24889 -23717 24922 -23671
rect 24822 -23739 24922 -23717
rect 24822 -23789 24855 -23739
rect 24889 -23789 24922 -23739
rect 24822 -23807 24922 -23789
rect 24822 -23861 24855 -23807
rect 24889 -23861 24922 -23807
rect 24822 -23875 24922 -23861
rect 24822 -23933 24855 -23875
rect 24889 -23933 24922 -23875
rect 24822 -23943 24922 -23933
rect 24822 -24005 24855 -23943
rect 24889 -24005 24922 -23943
rect 24822 -24011 24922 -24005
rect 2812 -24060 2851 -24026
rect 2885 -24060 2909 -24026
rect 2953 -24060 2981 -24026
rect 3021 -24060 3053 -24026
rect 3089 -24060 3123 -24026
rect 3159 -24060 3191 -24026
rect 3231 -24060 3259 -24026
rect 3303 -24060 3327 -24026
rect 3361 -24060 3400 -24026
rect 3830 -24060 3869 -24026
rect 3903 -24060 3927 -24026
rect 3971 -24060 3999 -24026
rect 4039 -24060 4071 -24026
rect 4107 -24060 4141 -24026
rect 4177 -24060 4209 -24026
rect 4249 -24060 4277 -24026
rect 4321 -24060 4345 -24026
rect 4379 -24060 4418 -24026
rect 4848 -24060 4887 -24026
rect 4921 -24060 4945 -24026
rect 4989 -24060 5017 -24026
rect 5057 -24060 5089 -24026
rect 5125 -24060 5159 -24026
rect 5195 -24060 5227 -24026
rect 5267 -24060 5295 -24026
rect 5339 -24060 5363 -24026
rect 5397 -24060 5436 -24026
rect 5866 -24060 5905 -24026
rect 5939 -24060 5963 -24026
rect 6007 -24060 6035 -24026
rect 6075 -24060 6107 -24026
rect 6143 -24060 6177 -24026
rect 6213 -24060 6245 -24026
rect 6285 -24060 6313 -24026
rect 6357 -24060 6381 -24026
rect 6415 -24060 6454 -24026
rect 6884 -24060 6923 -24026
rect 6957 -24060 6981 -24026
rect 7025 -24060 7053 -24026
rect 7093 -24060 7125 -24026
rect 7161 -24060 7195 -24026
rect 7231 -24060 7263 -24026
rect 7303 -24060 7331 -24026
rect 7375 -24060 7399 -24026
rect 7433 -24060 7472 -24026
rect 7902 -24060 7941 -24026
rect 7975 -24060 7999 -24026
rect 8043 -24060 8071 -24026
rect 8111 -24060 8143 -24026
rect 8179 -24060 8213 -24026
rect 8249 -24060 8281 -24026
rect 8321 -24060 8349 -24026
rect 8393 -24060 8417 -24026
rect 8451 -24060 8490 -24026
rect 8920 -24060 8959 -24026
rect 8993 -24060 9017 -24026
rect 9061 -24060 9089 -24026
rect 9129 -24060 9161 -24026
rect 9197 -24060 9231 -24026
rect 9267 -24060 9299 -24026
rect 9339 -24060 9367 -24026
rect 9411 -24060 9435 -24026
rect 9469 -24060 9508 -24026
rect 9938 -24060 9977 -24026
rect 10011 -24060 10035 -24026
rect 10079 -24060 10107 -24026
rect 10147 -24060 10179 -24026
rect 10215 -24060 10249 -24026
rect 10285 -24060 10317 -24026
rect 10357 -24060 10385 -24026
rect 10429 -24060 10453 -24026
rect 10487 -24060 10526 -24026
rect 10956 -24060 10995 -24026
rect 11029 -24060 11053 -24026
rect 11097 -24060 11125 -24026
rect 11165 -24060 11197 -24026
rect 11233 -24060 11267 -24026
rect 11303 -24060 11335 -24026
rect 11375 -24060 11403 -24026
rect 11447 -24060 11471 -24026
rect 11505 -24060 11544 -24026
rect 11974 -24060 12013 -24026
rect 12047 -24060 12071 -24026
rect 12115 -24060 12143 -24026
rect 12183 -24060 12215 -24026
rect 12251 -24060 12285 -24026
rect 12321 -24060 12353 -24026
rect 12393 -24060 12421 -24026
rect 12465 -24060 12489 -24026
rect 12523 -24060 12562 -24026
rect 12992 -24060 13031 -24026
rect 13065 -24060 13089 -24026
rect 13133 -24060 13161 -24026
rect 13201 -24060 13233 -24026
rect 13269 -24060 13303 -24026
rect 13339 -24060 13371 -24026
rect 13411 -24060 13439 -24026
rect 13483 -24060 13507 -24026
rect 13541 -24060 13580 -24026
rect 14010 -24060 14049 -24026
rect 14083 -24060 14107 -24026
rect 14151 -24060 14179 -24026
rect 14219 -24060 14251 -24026
rect 14287 -24060 14321 -24026
rect 14357 -24060 14389 -24026
rect 14429 -24060 14457 -24026
rect 14501 -24060 14525 -24026
rect 14559 -24060 14598 -24026
rect 15028 -24060 15067 -24026
rect 15101 -24060 15125 -24026
rect 15169 -24060 15197 -24026
rect 15237 -24060 15269 -24026
rect 15305 -24060 15339 -24026
rect 15375 -24060 15407 -24026
rect 15447 -24060 15475 -24026
rect 15519 -24060 15543 -24026
rect 15577 -24060 15616 -24026
rect 16046 -24060 16085 -24026
rect 16119 -24060 16143 -24026
rect 16187 -24060 16215 -24026
rect 16255 -24060 16287 -24026
rect 16323 -24060 16357 -24026
rect 16393 -24060 16425 -24026
rect 16465 -24060 16493 -24026
rect 16537 -24060 16561 -24026
rect 16595 -24060 16634 -24026
rect 17064 -24060 17103 -24026
rect 17137 -24060 17161 -24026
rect 17205 -24060 17233 -24026
rect 17273 -24060 17305 -24026
rect 17341 -24060 17375 -24026
rect 17411 -24060 17443 -24026
rect 17483 -24060 17511 -24026
rect 17555 -24060 17579 -24026
rect 17613 -24060 17652 -24026
rect 18082 -24060 18121 -24026
rect 18155 -24060 18179 -24026
rect 18223 -24060 18251 -24026
rect 18291 -24060 18323 -24026
rect 18359 -24060 18393 -24026
rect 18429 -24060 18461 -24026
rect 18501 -24060 18529 -24026
rect 18573 -24060 18597 -24026
rect 18631 -24060 18670 -24026
rect 19100 -24060 19139 -24026
rect 19173 -24060 19197 -24026
rect 19241 -24060 19269 -24026
rect 19309 -24060 19341 -24026
rect 19377 -24060 19411 -24026
rect 19447 -24060 19479 -24026
rect 19519 -24060 19547 -24026
rect 19591 -24060 19615 -24026
rect 19649 -24060 19688 -24026
rect 20118 -24060 20157 -24026
rect 20191 -24060 20215 -24026
rect 20259 -24060 20287 -24026
rect 20327 -24060 20359 -24026
rect 20395 -24060 20429 -24026
rect 20465 -24060 20497 -24026
rect 20537 -24060 20565 -24026
rect 20609 -24060 20633 -24026
rect 20667 -24060 20706 -24026
rect 21136 -24060 21175 -24026
rect 21209 -24060 21233 -24026
rect 21277 -24060 21305 -24026
rect 21345 -24060 21377 -24026
rect 21413 -24060 21447 -24026
rect 21483 -24060 21515 -24026
rect 21555 -24060 21583 -24026
rect 21627 -24060 21651 -24026
rect 21685 -24060 21724 -24026
rect 22154 -24060 22193 -24026
rect 22227 -24060 22251 -24026
rect 22295 -24060 22323 -24026
rect 22363 -24060 22395 -24026
rect 22431 -24060 22465 -24026
rect 22501 -24060 22533 -24026
rect 22573 -24060 22601 -24026
rect 22645 -24060 22669 -24026
rect 22703 -24060 22742 -24026
rect 6120 -24062 6180 -24060
rect -12322 -24079 -12222 -24077
rect -12322 -24113 -12289 -24079
rect -12255 -24113 -12222 -24079
rect 24822 -24077 24855 -24011
rect 24889 -24077 24922 -24011
rect 24822 -24079 24922 -24077
rect -12322 -24115 -12222 -24113
rect -12322 -24181 -12289 -24115
rect -12255 -24181 -12222 -24115
rect -12322 -24187 -12222 -24181
rect -12322 -24249 -12289 -24187
rect -12255 -24249 -12222 -24187
rect -12322 -24259 -12222 -24249
rect -12322 -24317 -12289 -24259
rect -12255 -24317 -12222 -24259
rect -12322 -24331 -12222 -24317
rect -12322 -24385 -12289 -24331
rect -12255 -24385 -12222 -24331
rect -12322 -24403 -12222 -24385
rect -12322 -24453 -12289 -24403
rect -12255 -24453 -12222 -24403
rect -12322 -24475 -12222 -24453
rect -12322 -24521 -12289 -24475
rect -12255 -24521 -12222 -24475
rect -12322 -24547 -12222 -24521
rect -12322 -24589 -12289 -24547
rect -12255 -24589 -12222 -24547
rect -12322 -24619 -12222 -24589
rect -12322 -24657 -12289 -24619
rect -12255 -24657 -12222 -24619
rect -12322 -24691 -12222 -24657
rect -12322 -24725 -12289 -24691
rect -12255 -24725 -12222 -24691
rect 2580 -24129 2614 -24094
rect 2580 -24201 2614 -24177
rect 2580 -24273 2614 -24245
rect 2580 -24345 2614 -24313
rect 2580 -24415 2614 -24381
rect 2580 -24483 2614 -24451
rect 2580 -24551 2614 -24523
rect 2580 -24619 2614 -24595
rect 2580 -24702 2614 -24667
rect 3598 -24129 3632 -24094
rect 3598 -24201 3632 -24177
rect 3598 -24273 3632 -24245
rect 3598 -24345 3632 -24313
rect 3598 -24415 3632 -24381
rect 3598 -24483 3632 -24451
rect 3598 -24551 3632 -24523
rect 3598 -24619 3632 -24595
rect 3598 -24702 3632 -24667
rect 4616 -24129 4650 -24094
rect 4616 -24201 4650 -24177
rect 4616 -24273 4650 -24245
rect 4616 -24345 4650 -24313
rect 4616 -24415 4650 -24381
rect 4616 -24483 4650 -24451
rect 4616 -24551 4650 -24523
rect 4616 -24619 4650 -24595
rect 4616 -24702 4650 -24667
rect 5634 -24129 5668 -24094
rect 5634 -24201 5668 -24177
rect 5634 -24273 5668 -24245
rect 5634 -24345 5668 -24313
rect 5634 -24415 5668 -24381
rect 5634 -24483 5668 -24451
rect 5634 -24551 5668 -24523
rect 5634 -24619 5668 -24595
rect 5634 -24702 5668 -24667
rect 6652 -24129 6686 -24094
rect 6652 -24201 6686 -24177
rect 6652 -24273 6686 -24245
rect 6652 -24345 6686 -24313
rect 6652 -24415 6686 -24381
rect 6652 -24483 6686 -24451
rect 6652 -24551 6686 -24523
rect 6652 -24619 6686 -24595
rect 6652 -24702 6686 -24667
rect 7670 -24129 7704 -24094
rect 7670 -24201 7704 -24177
rect 7670 -24273 7704 -24245
rect 7670 -24345 7704 -24313
rect 7670 -24415 7704 -24381
rect 7670 -24483 7704 -24451
rect 7670 -24551 7704 -24523
rect 7670 -24619 7704 -24595
rect 7670 -24702 7704 -24667
rect 8688 -24129 8722 -24094
rect 8688 -24201 8722 -24177
rect 8688 -24273 8722 -24245
rect 8688 -24345 8722 -24313
rect 8688 -24415 8722 -24381
rect 8688 -24483 8722 -24451
rect 8688 -24551 8722 -24523
rect 8688 -24619 8722 -24595
rect 8688 -24702 8722 -24667
rect 9706 -24129 9740 -24094
rect 9706 -24201 9740 -24177
rect 9706 -24273 9740 -24245
rect 9706 -24345 9740 -24313
rect 9706 -24415 9740 -24381
rect 9706 -24483 9740 -24451
rect 9706 -24551 9740 -24523
rect 9706 -24619 9740 -24595
rect 9706 -24702 9740 -24667
rect 10724 -24129 10758 -24094
rect 10724 -24201 10758 -24177
rect 10724 -24273 10758 -24245
rect 10724 -24345 10758 -24313
rect 10724 -24415 10758 -24381
rect 10724 -24483 10758 -24451
rect 10724 -24551 10758 -24523
rect 10724 -24619 10758 -24595
rect 10724 -24702 10758 -24667
rect 11742 -24129 11776 -24094
rect 11742 -24201 11776 -24177
rect 11742 -24273 11776 -24245
rect 11742 -24345 11776 -24313
rect 11742 -24415 11776 -24381
rect 11742 -24483 11776 -24451
rect 11742 -24551 11776 -24523
rect 11742 -24619 11776 -24595
rect 11742 -24702 11776 -24667
rect 12760 -24129 12794 -24094
rect 12760 -24201 12794 -24177
rect 12760 -24273 12794 -24245
rect 12760 -24345 12794 -24313
rect 12760 -24415 12794 -24381
rect 12760 -24483 12794 -24451
rect 12760 -24551 12794 -24523
rect 12760 -24619 12794 -24595
rect 12760 -24702 12794 -24667
rect 13778 -24129 13812 -24094
rect 13778 -24201 13812 -24177
rect 13778 -24273 13812 -24245
rect 13778 -24345 13812 -24313
rect 13778 -24415 13812 -24381
rect 13778 -24483 13812 -24451
rect 13778 -24551 13812 -24523
rect 13778 -24619 13812 -24595
rect 13778 -24702 13812 -24667
rect 14796 -24129 14830 -24094
rect 14796 -24201 14830 -24177
rect 14796 -24273 14830 -24245
rect 14796 -24345 14830 -24313
rect 14796 -24415 14830 -24381
rect 14796 -24483 14830 -24451
rect 14796 -24551 14830 -24523
rect 14796 -24619 14830 -24595
rect 14796 -24702 14830 -24667
rect 15814 -24129 15848 -24094
rect 15814 -24201 15848 -24177
rect 15814 -24273 15848 -24245
rect 15814 -24345 15848 -24313
rect 15814 -24415 15848 -24381
rect 15814 -24483 15848 -24451
rect 15814 -24551 15848 -24523
rect 15814 -24619 15848 -24595
rect 15814 -24702 15848 -24667
rect 16832 -24129 16866 -24094
rect 16832 -24201 16866 -24177
rect 16832 -24273 16866 -24245
rect 16832 -24345 16866 -24313
rect 16832 -24415 16866 -24381
rect 16832 -24483 16866 -24451
rect 16832 -24551 16866 -24523
rect 16832 -24619 16866 -24595
rect 16832 -24702 16866 -24667
rect 17850 -24129 17884 -24094
rect 17850 -24201 17884 -24177
rect 17850 -24273 17884 -24245
rect 17850 -24345 17884 -24313
rect 17850 -24415 17884 -24381
rect 17850 -24483 17884 -24451
rect 17850 -24551 17884 -24523
rect 17850 -24619 17884 -24595
rect 17850 -24702 17884 -24667
rect 18868 -24129 18902 -24094
rect 18868 -24201 18902 -24177
rect 18868 -24273 18902 -24245
rect 18868 -24345 18902 -24313
rect 18868 -24415 18902 -24381
rect 18868 -24483 18902 -24451
rect 18868 -24551 18902 -24523
rect 18868 -24619 18902 -24595
rect 18868 -24702 18902 -24667
rect 19886 -24129 19920 -24094
rect 19886 -24201 19920 -24177
rect 19886 -24273 19920 -24245
rect 19886 -24345 19920 -24313
rect 19886 -24415 19920 -24381
rect 19886 -24483 19920 -24451
rect 19886 -24551 19920 -24523
rect 19886 -24619 19920 -24595
rect 19886 -24702 19920 -24667
rect 20904 -24129 20938 -24094
rect 20904 -24201 20938 -24177
rect 20904 -24273 20938 -24245
rect 20904 -24345 20938 -24313
rect 20904 -24415 20938 -24381
rect 20904 -24483 20938 -24451
rect 20904 -24551 20938 -24523
rect 20904 -24619 20938 -24595
rect 20904 -24702 20938 -24667
rect 21922 -24129 21956 -24094
rect 21922 -24201 21956 -24177
rect 21922 -24273 21956 -24245
rect 21922 -24345 21956 -24313
rect 21922 -24415 21956 -24381
rect 21922 -24483 21956 -24451
rect 21922 -24551 21956 -24523
rect 21922 -24619 21956 -24595
rect 21922 -24702 21956 -24667
rect 22940 -24129 22974 -24094
rect 22940 -24201 22974 -24177
rect 22940 -24273 22974 -24245
rect 22940 -24345 22974 -24313
rect 22940 -24415 22974 -24381
rect 22940 -24483 22974 -24451
rect 22940 -24551 22974 -24523
rect 22940 -24619 22974 -24595
rect 22940 -24702 22974 -24667
rect 24822 -24113 24855 -24079
rect 24889 -24113 24922 -24079
rect 24822 -24115 24922 -24113
rect 24822 -24181 24855 -24115
rect 24889 -24181 24922 -24115
rect 24822 -24187 24922 -24181
rect 24822 -24249 24855 -24187
rect 24889 -24249 24922 -24187
rect 24822 -24259 24922 -24249
rect 24822 -24317 24855 -24259
rect 24889 -24317 24922 -24259
rect 24822 -24331 24922 -24317
rect 24822 -24385 24855 -24331
rect 24889 -24385 24922 -24331
rect 24822 -24403 24922 -24385
rect 24822 -24453 24855 -24403
rect 24889 -24453 24922 -24403
rect 24822 -24475 24922 -24453
rect 24822 -24521 24855 -24475
rect 24889 -24521 24922 -24475
rect 24822 -24547 24922 -24521
rect 24822 -24589 24855 -24547
rect 24889 -24589 24922 -24547
rect 24822 -24619 24922 -24589
rect 24822 -24657 24855 -24619
rect 24889 -24657 24922 -24619
rect 24822 -24691 24922 -24657
rect -12322 -24759 -12222 -24725
rect 24822 -24725 24855 -24691
rect 24889 -24725 24922 -24691
rect 4088 -24736 4148 -24734
rect 10200 -24736 10260 -24734
rect 12234 -24736 12294 -24734
rect 16300 -24736 16360 -24730
rect 20376 -24736 20436 -24734
rect 21392 -24736 21452 -24734
rect -12322 -24797 -12289 -24759
rect -12255 -24797 -12222 -24759
rect 2812 -24770 2851 -24736
rect 2885 -24770 2909 -24736
rect 2953 -24770 2981 -24736
rect 3021 -24770 3053 -24736
rect 3089 -24770 3123 -24736
rect 3159 -24770 3191 -24736
rect 3231 -24770 3259 -24736
rect 3303 -24770 3327 -24736
rect 3361 -24770 3400 -24736
rect 3830 -24770 3869 -24736
rect 3903 -24770 3927 -24736
rect 3971 -24770 3999 -24736
rect 4039 -24770 4071 -24736
rect 4107 -24770 4141 -24736
rect 4177 -24770 4209 -24736
rect 4249 -24770 4277 -24736
rect 4321 -24770 4345 -24736
rect 4379 -24770 4418 -24736
rect 4848 -24770 4887 -24736
rect 4921 -24770 4945 -24736
rect 4989 -24770 5017 -24736
rect 5057 -24770 5089 -24736
rect 5125 -24770 5159 -24736
rect 5195 -24770 5227 -24736
rect 5267 -24770 5295 -24736
rect 5339 -24770 5363 -24736
rect 5397 -24770 5436 -24736
rect 5866 -24770 5905 -24736
rect 5939 -24770 5963 -24736
rect 6007 -24770 6035 -24736
rect 6075 -24770 6107 -24736
rect 6143 -24770 6177 -24736
rect 6213 -24770 6245 -24736
rect 6285 -24770 6313 -24736
rect 6357 -24770 6381 -24736
rect 6415 -24770 6454 -24736
rect 6884 -24770 6923 -24736
rect 6957 -24770 6981 -24736
rect 7025 -24770 7053 -24736
rect 7093 -24770 7125 -24736
rect 7161 -24770 7195 -24736
rect 7231 -24770 7263 -24736
rect 7303 -24770 7331 -24736
rect 7375 -24770 7399 -24736
rect 7433 -24770 7472 -24736
rect 7902 -24770 7941 -24736
rect 7975 -24770 7999 -24736
rect 8043 -24770 8071 -24736
rect 8111 -24770 8143 -24736
rect 8179 -24770 8213 -24736
rect 8249 -24770 8281 -24736
rect 8321 -24770 8349 -24736
rect 8393 -24770 8417 -24736
rect 8451 -24770 8490 -24736
rect 8920 -24770 8959 -24736
rect 8993 -24770 9017 -24736
rect 9061 -24770 9089 -24736
rect 9129 -24770 9161 -24736
rect 9197 -24770 9231 -24736
rect 9267 -24770 9299 -24736
rect 9339 -24770 9367 -24736
rect 9411 -24770 9435 -24736
rect 9469 -24770 9508 -24736
rect 9938 -24770 9977 -24736
rect 10011 -24770 10035 -24736
rect 10079 -24770 10107 -24736
rect 10147 -24770 10179 -24736
rect 10215 -24770 10249 -24736
rect 10285 -24770 10317 -24736
rect 10357 -24770 10385 -24736
rect 10429 -24770 10453 -24736
rect 10487 -24770 10526 -24736
rect 10956 -24770 10995 -24736
rect 11029 -24770 11053 -24736
rect 11097 -24770 11125 -24736
rect 11165 -24770 11197 -24736
rect 11233 -24770 11267 -24736
rect 11303 -24770 11335 -24736
rect 11375 -24770 11403 -24736
rect 11447 -24770 11471 -24736
rect 11505 -24770 11544 -24736
rect 11974 -24770 12013 -24736
rect 12047 -24770 12071 -24736
rect 12115 -24770 12143 -24736
rect 12183 -24770 12215 -24736
rect 12251 -24770 12285 -24736
rect 12321 -24770 12353 -24736
rect 12393 -24770 12421 -24736
rect 12465 -24770 12489 -24736
rect 12523 -24770 12562 -24736
rect 12992 -24770 13031 -24736
rect 13065 -24770 13089 -24736
rect 13133 -24770 13161 -24736
rect 13201 -24770 13233 -24736
rect 13269 -24770 13303 -24736
rect 13339 -24770 13371 -24736
rect 13411 -24770 13439 -24736
rect 13483 -24770 13507 -24736
rect 13541 -24770 13580 -24736
rect 14010 -24770 14049 -24736
rect 14083 -24770 14107 -24736
rect 14151 -24770 14179 -24736
rect 14219 -24770 14251 -24736
rect 14287 -24770 14321 -24736
rect 14357 -24770 14389 -24736
rect 14429 -24770 14457 -24736
rect 14501 -24770 14525 -24736
rect 14559 -24770 14598 -24736
rect 15028 -24770 15067 -24736
rect 15101 -24770 15125 -24736
rect 15169 -24770 15197 -24736
rect 15237 -24770 15269 -24736
rect 15305 -24770 15339 -24736
rect 15375 -24770 15407 -24736
rect 15447 -24770 15475 -24736
rect 15519 -24770 15543 -24736
rect 15577 -24770 15616 -24736
rect 16046 -24770 16085 -24736
rect 16119 -24770 16143 -24736
rect 16187 -24770 16215 -24736
rect 16255 -24770 16287 -24736
rect 16323 -24770 16357 -24736
rect 16393 -24770 16425 -24736
rect 16465 -24770 16493 -24736
rect 16537 -24770 16561 -24736
rect 16595 -24770 16634 -24736
rect 17064 -24770 17103 -24736
rect 17137 -24770 17161 -24736
rect 17205 -24770 17233 -24736
rect 17273 -24770 17305 -24736
rect 17341 -24770 17375 -24736
rect 17411 -24770 17443 -24736
rect 17483 -24770 17511 -24736
rect 17555 -24770 17579 -24736
rect 17613 -24770 17652 -24736
rect 18082 -24770 18121 -24736
rect 18155 -24770 18179 -24736
rect 18223 -24770 18251 -24736
rect 18291 -24770 18323 -24736
rect 18359 -24770 18393 -24736
rect 18429 -24770 18461 -24736
rect 18501 -24770 18529 -24736
rect 18573 -24770 18597 -24736
rect 18631 -24770 18670 -24736
rect 19100 -24770 19139 -24736
rect 19173 -24770 19197 -24736
rect 19241 -24770 19269 -24736
rect 19309 -24770 19341 -24736
rect 19377 -24770 19411 -24736
rect 19447 -24770 19479 -24736
rect 19519 -24770 19547 -24736
rect 19591 -24770 19615 -24736
rect 19649 -24770 19688 -24736
rect 20118 -24770 20157 -24736
rect 20191 -24770 20215 -24736
rect 20259 -24770 20287 -24736
rect 20327 -24770 20359 -24736
rect 20395 -24770 20429 -24736
rect 20465 -24770 20497 -24736
rect 20537 -24770 20565 -24736
rect 20609 -24770 20633 -24736
rect 20667 -24770 20706 -24736
rect 21136 -24770 21175 -24736
rect 21209 -24770 21233 -24736
rect 21277 -24770 21305 -24736
rect 21345 -24770 21377 -24736
rect 21413 -24770 21447 -24736
rect 21483 -24770 21515 -24736
rect 21555 -24770 21583 -24736
rect 21627 -24770 21651 -24736
rect 21685 -24770 21724 -24736
rect 22154 -24770 22193 -24736
rect 22227 -24770 22251 -24736
rect 22295 -24770 22323 -24736
rect 22363 -24770 22395 -24736
rect 22431 -24770 22465 -24736
rect 22501 -24770 22533 -24736
rect 22573 -24770 22601 -24736
rect 22645 -24770 22669 -24736
rect 22703 -24770 22742 -24736
rect 24822 -24759 24922 -24725
rect -12322 -24827 -12222 -24797
rect -12322 -24869 -12289 -24827
rect -12255 -24869 -12222 -24827
rect -12322 -24895 -12222 -24869
rect -12322 -24941 -12289 -24895
rect -12255 -24941 -12222 -24895
rect -12322 -24963 -12222 -24941
rect -12322 -25013 -12289 -24963
rect -12255 -25013 -12222 -24963
rect -12322 -25031 -12222 -25013
rect -12322 -25085 -12289 -25031
rect -12255 -25085 -12222 -25031
rect -12322 -25099 -12222 -25085
rect -12322 -25157 -12289 -25099
rect -12255 -25157 -12222 -25099
rect -12322 -25167 -12222 -25157
rect -12322 -25229 -12289 -25167
rect -12255 -25229 -12222 -25167
rect -12322 -25235 -12222 -25229
rect -12322 -25301 -12289 -25235
rect -12255 -25301 -12222 -25235
rect -12322 -25303 -12222 -25301
rect -12322 -25337 -12289 -25303
rect -12255 -25337 -12222 -25303
rect -12322 -25339 -12222 -25337
rect -12322 -25405 -12289 -25339
rect -12255 -25405 -12222 -25339
rect -12322 -25411 -12222 -25405
rect -12322 -25473 -12289 -25411
rect -12255 -25473 -12222 -25411
rect -12322 -25483 -12222 -25473
rect -12322 -25541 -12289 -25483
rect -12255 -25541 -12222 -25483
rect -12322 -25555 -12222 -25541
rect -12322 -25609 -12289 -25555
rect -12255 -25609 -12222 -25555
rect -12322 -25627 -12222 -25609
rect -12322 -25677 -12289 -25627
rect -12255 -25677 -12222 -25627
rect -12322 -25699 -12222 -25677
rect -12322 -25745 -12289 -25699
rect -12255 -25745 -12222 -25699
rect -12322 -25771 -12222 -25745
rect -12322 -25813 -12289 -25771
rect -12255 -25813 -12222 -25771
rect -12322 -25843 -12222 -25813
rect -12322 -25881 -12289 -25843
rect -12255 -25881 -12222 -25843
rect -12322 -25915 -12222 -25881
rect -12322 -25949 -12289 -25915
rect -12255 -25949 -12222 -25915
rect -12322 -25983 -12222 -25949
rect -12322 -26021 -12289 -25983
rect -12255 -26021 -12222 -25983
rect -12322 -26051 -12222 -26021
rect -12322 -26093 -12289 -26051
rect -12255 -26093 -12222 -26051
rect -12322 -26119 -12222 -26093
rect -12322 -26165 -12289 -26119
rect -12255 -26165 -12222 -26119
rect -12322 -26187 -12222 -26165
rect -12322 -26237 -12289 -26187
rect -12255 -26237 -12222 -26187
rect -12322 -26255 -12222 -26237
rect -12322 -26309 -12289 -26255
rect -12255 -26309 -12222 -26255
rect -12322 -26323 -12222 -26309
rect -12322 -26357 -12289 -26323
rect -12255 -26357 -12222 -26323
rect -12322 -26391 -12222 -26357
rect -12322 -26425 -12289 -26391
rect -12255 -26425 -12222 -26391
rect -12322 -26459 -12222 -26425
rect -12322 -26493 -12289 -26459
rect -12255 -26493 -12222 -26459
rect -12322 -26527 -12222 -26493
rect -12322 -26561 -12289 -26527
rect -12255 -26561 -12222 -26527
rect -12322 -26595 -12222 -26561
rect -12322 -26629 -12289 -26595
rect -12255 -26629 -12222 -26595
rect -12322 -26663 -12222 -26629
rect -12322 -26697 -12289 -26663
rect -12255 -26697 -12222 -26663
rect -12322 -26731 -12222 -26697
rect -12322 -26765 -12289 -26731
rect -12255 -26765 -12222 -26731
rect -12322 -26799 -12222 -26765
rect -12322 -26833 -12289 -26799
rect -12255 -26833 -12222 -26799
rect -12322 -26867 -12222 -26833
rect -12322 -26901 -12289 -26867
rect -12255 -26901 -12222 -26867
rect -12322 -26935 -12222 -26901
rect -12322 -26969 -12289 -26935
rect -12255 -26969 -12222 -26935
rect -12322 -27003 -12222 -26969
rect -12322 -27037 -12289 -27003
rect -12255 -27037 -12222 -27003
rect -12322 -27122 -12222 -27037
rect 24822 -24797 24855 -24759
rect 24889 -24797 24922 -24759
rect 24822 -24827 24922 -24797
rect 24822 -24869 24855 -24827
rect 24889 -24869 24922 -24827
rect 24822 -24895 24922 -24869
rect 24822 -24941 24855 -24895
rect 24889 -24941 24922 -24895
rect 24822 -24963 24922 -24941
rect 24822 -25013 24855 -24963
rect 24889 -25013 24922 -24963
rect 24822 -25031 24922 -25013
rect 24822 -25085 24855 -25031
rect 24889 -25085 24922 -25031
rect 24822 -25099 24922 -25085
rect 24822 -25157 24855 -25099
rect 24889 -25157 24922 -25099
rect 24822 -25167 24922 -25157
rect 24822 -25229 24855 -25167
rect 24889 -25229 24922 -25167
rect 24822 -25235 24922 -25229
rect 24822 -25301 24855 -25235
rect 24889 -25301 24922 -25235
rect 24822 -25303 24922 -25301
rect 24822 -25337 24855 -25303
rect 24889 -25337 24922 -25303
rect 24822 -25339 24922 -25337
rect 24822 -25405 24855 -25339
rect 24889 -25405 24922 -25339
rect 24822 -25411 24922 -25405
rect 24822 -25473 24855 -25411
rect 24889 -25473 24922 -25411
rect 24822 -25483 24922 -25473
rect 24822 -25541 24855 -25483
rect 24889 -25541 24922 -25483
rect 24822 -25555 24922 -25541
rect 24822 -25609 24855 -25555
rect 24889 -25609 24922 -25555
rect 24822 -25627 24922 -25609
rect 24822 -25677 24855 -25627
rect 24889 -25677 24922 -25627
rect 24822 -25699 24922 -25677
rect 24822 -25745 24855 -25699
rect 24889 -25745 24922 -25699
rect 24822 -25771 24922 -25745
rect 24822 -25813 24855 -25771
rect 24889 -25813 24922 -25771
rect 24822 -25843 24922 -25813
rect 24822 -25881 24855 -25843
rect 24889 -25881 24922 -25843
rect 24822 -25915 24922 -25881
rect 24822 -25949 24855 -25915
rect 24889 -25949 24922 -25915
rect 24822 -25983 24922 -25949
rect 24822 -26021 24855 -25983
rect 24889 -26021 24922 -25983
rect 24822 -26051 24922 -26021
rect 24822 -26093 24855 -26051
rect 24889 -26093 24922 -26051
rect 24822 -26119 24922 -26093
rect 24822 -26165 24855 -26119
rect 24889 -26165 24922 -26119
rect 24822 -26187 24922 -26165
rect 24822 -26237 24855 -26187
rect 24889 -26237 24922 -26187
rect 24822 -26255 24922 -26237
rect 24822 -26309 24855 -26255
rect 24889 -26309 24922 -26255
rect 24822 -26323 24922 -26309
rect 24822 -26357 24855 -26323
rect 24889 -26357 24922 -26323
rect 24822 -26391 24922 -26357
rect 24822 -26425 24855 -26391
rect 24889 -26425 24922 -26391
rect 24822 -26459 24922 -26425
rect 24822 -26493 24855 -26459
rect 24889 -26493 24922 -26459
rect 24822 -26527 24922 -26493
rect 24822 -26561 24855 -26527
rect 24889 -26561 24922 -26527
rect 24822 -26595 24922 -26561
rect 24822 -26629 24855 -26595
rect 24889 -26629 24922 -26595
rect 24822 -26663 24922 -26629
rect 24822 -26697 24855 -26663
rect 24889 -26697 24922 -26663
rect 24822 -26731 24922 -26697
rect 24822 -26765 24855 -26731
rect 24889 -26765 24922 -26731
rect 24822 -26799 24922 -26765
rect 24822 -26833 24855 -26799
rect 24889 -26833 24922 -26799
rect 24822 -26867 24922 -26833
rect 24822 -26901 24855 -26867
rect 24889 -26901 24922 -26867
rect 24822 -26935 24922 -26901
rect 24822 -26969 24855 -26935
rect 24889 -26969 24922 -26935
rect 24822 -27003 24922 -26969
rect 24822 -27037 24855 -27003
rect 24889 -27037 24922 -27003
rect 24822 -27122 24922 -27037
rect -12322 -27155 24922 -27122
rect -12322 -27189 -12221 -27155
rect -12187 -27189 -12149 -27155
rect -12111 -27189 -12077 -27155
rect -12043 -27189 -12009 -27155
rect -11971 -27189 -11941 -27155
rect -11899 -27189 -11873 -27155
rect -11827 -27189 -11805 -27155
rect -11755 -27189 -11737 -27155
rect -11683 -27189 -11669 -27155
rect -11611 -27189 -11601 -27155
rect -11539 -27189 -11533 -27155
rect -11467 -27189 -11465 -27155
rect -11431 -27189 -11429 -27155
rect -11363 -27189 -11357 -27155
rect -11295 -27189 -11285 -27155
rect -11227 -27189 -11213 -27155
rect -11159 -27189 -11141 -27155
rect -11091 -27189 -11069 -27155
rect -11023 -27189 -10997 -27155
rect -10955 -27189 -10925 -27155
rect -10887 -27189 -10853 -27155
rect -10819 -27189 -10785 -27155
rect -10747 -27189 -10717 -27155
rect -10675 -27189 -10649 -27155
rect -10603 -27189 -10581 -27155
rect -10531 -27189 -10513 -27155
rect -10459 -27189 -10445 -27155
rect -10387 -27189 -10377 -27155
rect -10315 -27189 -10309 -27155
rect -10243 -27189 -10241 -27155
rect -10207 -27189 -10205 -27155
rect -10139 -27189 -10133 -27155
rect -10071 -27189 -10061 -27155
rect -10003 -27189 -9989 -27155
rect -9935 -27189 -9917 -27155
rect -9867 -27189 -9845 -27155
rect -9799 -27189 -9773 -27155
rect -9731 -27189 -9701 -27155
rect -9663 -27189 -9629 -27155
rect -9595 -27189 -9561 -27155
rect -9523 -27189 -9493 -27155
rect -9451 -27189 -9425 -27155
rect -9379 -27189 -9357 -27155
rect -9307 -27189 -9289 -27155
rect -9235 -27189 -9221 -27155
rect -9163 -27189 -9153 -27155
rect -9091 -27189 -9085 -27155
rect -9019 -27189 -9017 -27155
rect -8983 -27189 -8981 -27155
rect -8915 -27189 -8909 -27155
rect -8847 -27189 -8837 -27155
rect -8779 -27189 -8765 -27155
rect -8711 -27189 -8693 -27155
rect -8643 -27189 -8621 -27155
rect -8575 -27189 -8549 -27155
rect -8507 -27189 -8477 -27155
rect -8439 -27189 -8405 -27155
rect -8371 -27189 -8337 -27155
rect -8299 -27189 -8269 -27155
rect -8227 -27189 -8201 -27155
rect -8155 -27189 -8133 -27155
rect -8083 -27189 -8065 -27155
rect -8011 -27189 -7997 -27155
rect -7939 -27189 -7929 -27155
rect -7867 -27189 -7861 -27155
rect -7795 -27189 -7793 -27155
rect -7759 -27189 -7757 -27155
rect -7691 -27189 -7685 -27155
rect -7623 -27189 -7613 -27155
rect -7555 -27189 -7541 -27155
rect -7487 -27189 -7469 -27155
rect -7419 -27189 -7397 -27155
rect -7351 -27189 -7325 -27155
rect -7283 -27189 -7253 -27155
rect -7215 -27189 -7181 -27155
rect -7147 -27189 -7113 -27155
rect -7075 -27189 -7045 -27155
rect -7003 -27189 -6977 -27155
rect -6931 -27189 -6909 -27155
rect -6859 -27189 -6841 -27155
rect -6787 -27189 -6773 -27155
rect -6715 -27189 -6705 -27155
rect -6643 -27189 -6637 -27155
rect -6571 -27189 -6569 -27155
rect -6535 -27189 -6533 -27155
rect -6467 -27189 -6461 -27155
rect -6399 -27189 -6389 -27155
rect -6331 -27189 -6317 -27155
rect -6263 -27189 -6245 -27155
rect -6195 -27189 -6173 -27155
rect -6127 -27189 -6101 -27155
rect -6059 -27189 -6029 -27155
rect -5991 -27189 -5957 -27155
rect -5923 -27189 -5889 -27155
rect -5851 -27189 -5821 -27155
rect -5779 -27189 -5753 -27155
rect -5707 -27189 -5685 -27155
rect -5635 -27189 -5617 -27155
rect -5563 -27189 -5549 -27155
rect -5491 -27189 -5481 -27155
rect -5419 -27189 -5413 -27155
rect -5347 -27189 -5345 -27155
rect -5311 -27189 -5309 -27155
rect -5243 -27189 -5237 -27155
rect -5175 -27189 -5165 -27155
rect -5107 -27189 -5093 -27155
rect -5039 -27189 -5021 -27155
rect -4971 -27189 -4949 -27155
rect -4903 -27189 -4877 -27155
rect -4835 -27189 -4805 -27155
rect -4767 -27189 -4733 -27155
rect -4699 -27189 -4665 -27155
rect -4627 -27189 -4597 -27155
rect -4555 -27189 -4529 -27155
rect -4483 -27189 -4461 -27155
rect -4411 -27189 -4393 -27155
rect -4339 -27189 -4325 -27155
rect -4267 -27189 -4257 -27155
rect -4195 -27189 -4189 -27155
rect -4123 -27189 -4121 -27155
rect -4087 -27189 -4085 -27155
rect -4019 -27189 -4013 -27155
rect -3951 -27189 -3941 -27155
rect -3883 -27189 -3869 -27155
rect -3815 -27189 -3797 -27155
rect -3747 -27189 -3725 -27155
rect -3679 -27189 -3653 -27155
rect -3611 -27189 -3581 -27155
rect -3543 -27189 -3509 -27155
rect -3475 -27189 -3441 -27155
rect -3403 -27189 -3373 -27155
rect -3331 -27189 -3305 -27155
rect -3259 -27189 -3237 -27155
rect -3187 -27189 -3169 -27155
rect -3115 -27189 -3101 -27155
rect -3043 -27189 -3033 -27155
rect -2971 -27189 -2965 -27155
rect -2899 -27189 -2897 -27155
rect -2863 -27189 -2861 -27155
rect -2795 -27189 -2789 -27155
rect -2727 -27189 -2717 -27155
rect -2659 -27189 -2645 -27155
rect -2591 -27189 -2573 -27155
rect -2523 -27189 -2501 -27155
rect -2455 -27189 -2429 -27155
rect -2387 -27189 -2357 -27155
rect -2319 -27189 -2285 -27155
rect -2251 -27189 -2217 -27155
rect -2179 -27189 -2149 -27155
rect -2107 -27189 -2081 -27155
rect -2035 -27189 -2013 -27155
rect -1963 -27189 -1945 -27155
rect -1891 -27189 -1877 -27155
rect -1819 -27189 -1809 -27155
rect -1747 -27189 -1741 -27155
rect -1675 -27189 -1673 -27155
rect -1639 -27189 -1637 -27155
rect -1571 -27189 -1565 -27155
rect -1503 -27189 -1493 -27155
rect -1435 -27189 -1421 -27155
rect -1367 -27189 -1349 -27155
rect -1299 -27189 -1277 -27155
rect -1231 -27189 -1205 -27155
rect -1163 -27189 -1133 -27155
rect -1095 -27189 -1061 -27155
rect -1027 -27189 -993 -27155
rect -955 -27189 -925 -27155
rect -883 -27189 -857 -27155
rect -811 -27189 -789 -27155
rect -739 -27189 -721 -27155
rect -667 -27189 -653 -27155
rect -595 -27189 -585 -27155
rect -523 -27189 -517 -27155
rect -451 -27189 -449 -27155
rect -415 -27189 -413 -27155
rect -347 -27189 -341 -27155
rect -279 -27189 -269 -27155
rect -211 -27189 -197 -27155
rect -143 -27189 -125 -27155
rect -75 -27189 -53 -27155
rect -7 -27189 19 -27155
rect 61 -27189 91 -27155
rect 129 -27189 163 -27155
rect 197 -27189 231 -27155
rect 269 -27189 299 -27155
rect 341 -27189 367 -27155
rect 413 -27189 435 -27155
rect 485 -27189 503 -27155
rect 557 -27189 571 -27155
rect 629 -27189 639 -27155
rect 701 -27189 707 -27155
rect 773 -27189 775 -27155
rect 809 -27189 811 -27155
rect 877 -27189 883 -27155
rect 945 -27189 955 -27155
rect 1013 -27189 1027 -27155
rect 1081 -27189 1099 -27155
rect 1149 -27189 1171 -27155
rect 1217 -27189 1243 -27155
rect 1285 -27189 1315 -27155
rect 1353 -27189 1387 -27155
rect 1421 -27189 1455 -27155
rect 1493 -27189 1523 -27155
rect 1565 -27189 1591 -27155
rect 1637 -27189 1659 -27155
rect 1709 -27189 1727 -27155
rect 1781 -27189 1795 -27155
rect 1853 -27189 1863 -27155
rect 1925 -27189 1931 -27155
rect 1997 -27189 1999 -27155
rect 2033 -27189 2035 -27155
rect 2101 -27189 2107 -27155
rect 2169 -27189 2179 -27155
rect 2237 -27189 2251 -27155
rect 2305 -27189 2323 -27155
rect 2373 -27189 2395 -27155
rect 2441 -27189 2467 -27155
rect 2509 -27189 2539 -27155
rect 2577 -27189 2611 -27155
rect 2645 -27189 2679 -27155
rect 2717 -27189 2747 -27155
rect 2789 -27189 2815 -27155
rect 2861 -27189 2883 -27155
rect 2933 -27189 2951 -27155
rect 3005 -27189 3019 -27155
rect 3077 -27189 3087 -27155
rect 3149 -27189 3155 -27155
rect 3221 -27189 3223 -27155
rect 3257 -27189 3259 -27155
rect 3325 -27189 3331 -27155
rect 3393 -27189 3403 -27155
rect 3461 -27189 3475 -27155
rect 3529 -27189 3547 -27155
rect 3597 -27189 3619 -27155
rect 3665 -27189 3691 -27155
rect 3733 -27189 3763 -27155
rect 3801 -27189 3835 -27155
rect 3869 -27189 3903 -27155
rect 3941 -27189 3971 -27155
rect 4013 -27189 4039 -27155
rect 4085 -27189 4107 -27155
rect 4157 -27189 4175 -27155
rect 4229 -27189 4243 -27155
rect 4301 -27189 4311 -27155
rect 4373 -27189 4379 -27155
rect 4445 -27189 4447 -27155
rect 4481 -27189 4483 -27155
rect 4549 -27189 4555 -27155
rect 4617 -27189 4627 -27155
rect 4685 -27189 4699 -27155
rect 4753 -27189 4771 -27155
rect 4821 -27189 4843 -27155
rect 4889 -27189 4915 -27155
rect 4957 -27189 4987 -27155
rect 5025 -27189 5059 -27155
rect 5093 -27189 5127 -27155
rect 5165 -27189 5195 -27155
rect 5237 -27189 5263 -27155
rect 5309 -27189 5331 -27155
rect 5381 -27189 5399 -27155
rect 5453 -27189 5467 -27155
rect 5525 -27189 5535 -27155
rect 5597 -27189 5603 -27155
rect 5669 -27189 5671 -27155
rect 5705 -27189 5707 -27155
rect 5773 -27189 5779 -27155
rect 5841 -27189 5851 -27155
rect 5909 -27189 5923 -27155
rect 5977 -27189 5995 -27155
rect 6045 -27189 6067 -27155
rect 6113 -27189 6139 -27155
rect 6181 -27189 6211 -27155
rect 6249 -27189 6283 -27155
rect 6317 -27189 6351 -27155
rect 6389 -27189 6419 -27155
rect 6461 -27189 6487 -27155
rect 6533 -27189 6555 -27155
rect 6605 -27189 6623 -27155
rect 6677 -27189 6691 -27155
rect 6749 -27189 6759 -27155
rect 6821 -27189 6827 -27155
rect 6893 -27189 6895 -27155
rect 6929 -27189 6931 -27155
rect 6997 -27189 7003 -27155
rect 7065 -27189 7075 -27155
rect 7133 -27189 7147 -27155
rect 7201 -27189 7219 -27155
rect 7269 -27189 7291 -27155
rect 7337 -27189 7363 -27155
rect 7405 -27189 7435 -27155
rect 7473 -27189 7507 -27155
rect 7541 -27189 7575 -27155
rect 7613 -27189 7643 -27155
rect 7685 -27189 7711 -27155
rect 7757 -27189 7779 -27155
rect 7829 -27189 7847 -27155
rect 7901 -27189 7915 -27155
rect 7973 -27189 7983 -27155
rect 8045 -27189 8051 -27155
rect 8117 -27189 8119 -27155
rect 8153 -27189 8155 -27155
rect 8221 -27189 8227 -27155
rect 8289 -27189 8299 -27155
rect 8357 -27189 8371 -27155
rect 8425 -27189 8443 -27155
rect 8493 -27189 8515 -27155
rect 8561 -27189 8587 -27155
rect 8629 -27189 8659 -27155
rect 8697 -27189 8731 -27155
rect 8765 -27189 8799 -27155
rect 8837 -27189 8867 -27155
rect 8909 -27189 8935 -27155
rect 8981 -27189 9003 -27155
rect 9053 -27189 9071 -27155
rect 9125 -27189 9139 -27155
rect 9197 -27189 9207 -27155
rect 9269 -27189 9275 -27155
rect 9341 -27189 9343 -27155
rect 9377 -27189 9379 -27155
rect 9445 -27189 9451 -27155
rect 9513 -27189 9523 -27155
rect 9581 -27189 9595 -27155
rect 9649 -27189 9667 -27155
rect 9717 -27189 9739 -27155
rect 9785 -27189 9811 -27155
rect 9853 -27189 9883 -27155
rect 9921 -27189 9955 -27155
rect 9989 -27189 10023 -27155
rect 10061 -27189 10091 -27155
rect 10133 -27189 10159 -27155
rect 10205 -27189 10227 -27155
rect 10277 -27189 10295 -27155
rect 10349 -27189 10363 -27155
rect 10421 -27189 10431 -27155
rect 10493 -27189 10499 -27155
rect 10565 -27189 10567 -27155
rect 10601 -27189 10603 -27155
rect 10669 -27189 10675 -27155
rect 10737 -27189 10747 -27155
rect 10805 -27189 10819 -27155
rect 10873 -27189 10891 -27155
rect 10941 -27189 10963 -27155
rect 11009 -27189 11035 -27155
rect 11077 -27189 11107 -27155
rect 11145 -27189 11179 -27155
rect 11213 -27189 11247 -27155
rect 11285 -27189 11315 -27155
rect 11357 -27189 11383 -27155
rect 11429 -27189 11451 -27155
rect 11501 -27189 11519 -27155
rect 11573 -27189 11587 -27155
rect 11645 -27189 11655 -27155
rect 11717 -27189 11723 -27155
rect 11789 -27189 11791 -27155
rect 11825 -27189 11827 -27155
rect 11893 -27189 11899 -27155
rect 11961 -27189 11971 -27155
rect 12029 -27189 12043 -27155
rect 12097 -27189 12115 -27155
rect 12165 -27189 12187 -27155
rect 12233 -27189 12259 -27155
rect 12301 -27189 12331 -27155
rect 12369 -27189 12403 -27155
rect 12437 -27189 12471 -27155
rect 12509 -27189 12539 -27155
rect 12581 -27189 12607 -27155
rect 12653 -27189 12675 -27155
rect 12725 -27189 12743 -27155
rect 12797 -27189 12811 -27155
rect 12869 -27189 12879 -27155
rect 12941 -27189 12947 -27155
rect 13013 -27189 13015 -27155
rect 13049 -27189 13051 -27155
rect 13117 -27189 13123 -27155
rect 13185 -27189 13195 -27155
rect 13253 -27189 13267 -27155
rect 13321 -27189 13339 -27155
rect 13389 -27189 13411 -27155
rect 13457 -27189 13483 -27155
rect 13525 -27189 13555 -27155
rect 13593 -27189 13627 -27155
rect 13661 -27189 13695 -27155
rect 13733 -27189 13763 -27155
rect 13805 -27189 13831 -27155
rect 13877 -27189 13899 -27155
rect 13949 -27189 13967 -27155
rect 14021 -27189 14035 -27155
rect 14093 -27189 14103 -27155
rect 14165 -27189 14171 -27155
rect 14237 -27189 14239 -27155
rect 14273 -27189 14275 -27155
rect 14341 -27189 14347 -27155
rect 14409 -27189 14419 -27155
rect 14477 -27189 14491 -27155
rect 14545 -27189 14563 -27155
rect 14613 -27189 14635 -27155
rect 14681 -27189 14707 -27155
rect 14749 -27189 14779 -27155
rect 14817 -27189 14851 -27155
rect 14885 -27189 14919 -27155
rect 14957 -27189 14987 -27155
rect 15029 -27189 15055 -27155
rect 15101 -27189 15123 -27155
rect 15173 -27189 15191 -27155
rect 15245 -27189 15259 -27155
rect 15317 -27189 15327 -27155
rect 15389 -27189 15395 -27155
rect 15461 -27189 15463 -27155
rect 15497 -27189 15499 -27155
rect 15565 -27189 15571 -27155
rect 15633 -27189 15643 -27155
rect 15701 -27189 15715 -27155
rect 15769 -27189 15787 -27155
rect 15837 -27189 15859 -27155
rect 15905 -27189 15931 -27155
rect 15973 -27189 16003 -27155
rect 16041 -27189 16075 -27155
rect 16109 -27189 16143 -27155
rect 16181 -27189 16211 -27155
rect 16253 -27189 16279 -27155
rect 16325 -27189 16347 -27155
rect 16397 -27189 16415 -27155
rect 16469 -27189 16483 -27155
rect 16541 -27189 16551 -27155
rect 16613 -27189 16619 -27155
rect 16685 -27189 16687 -27155
rect 16721 -27189 16723 -27155
rect 16789 -27189 16795 -27155
rect 16857 -27189 16867 -27155
rect 16925 -27189 16939 -27155
rect 16993 -27189 17011 -27155
rect 17061 -27189 17083 -27155
rect 17129 -27189 17155 -27155
rect 17197 -27189 17227 -27155
rect 17265 -27189 17299 -27155
rect 17333 -27189 17367 -27155
rect 17405 -27189 17435 -27155
rect 17477 -27189 17503 -27155
rect 17549 -27189 17571 -27155
rect 17621 -27189 17639 -27155
rect 17693 -27189 17707 -27155
rect 17765 -27189 17775 -27155
rect 17837 -27189 17843 -27155
rect 17909 -27189 17911 -27155
rect 17945 -27189 17947 -27155
rect 18013 -27189 18019 -27155
rect 18081 -27189 18091 -27155
rect 18149 -27189 18163 -27155
rect 18217 -27189 18235 -27155
rect 18285 -27189 18307 -27155
rect 18353 -27189 18379 -27155
rect 18421 -27189 18451 -27155
rect 18489 -27189 18523 -27155
rect 18557 -27189 18591 -27155
rect 18629 -27189 18659 -27155
rect 18701 -27189 18727 -27155
rect 18773 -27189 18795 -27155
rect 18845 -27189 18863 -27155
rect 18917 -27189 18931 -27155
rect 18989 -27189 18999 -27155
rect 19061 -27189 19067 -27155
rect 19133 -27189 19135 -27155
rect 19169 -27189 19171 -27155
rect 19237 -27189 19243 -27155
rect 19305 -27189 19315 -27155
rect 19373 -27189 19387 -27155
rect 19441 -27189 19459 -27155
rect 19509 -27189 19531 -27155
rect 19577 -27189 19603 -27155
rect 19645 -27189 19675 -27155
rect 19713 -27189 19747 -27155
rect 19781 -27189 19815 -27155
rect 19853 -27189 19883 -27155
rect 19925 -27189 19951 -27155
rect 19997 -27189 20019 -27155
rect 20069 -27189 20087 -27155
rect 20141 -27189 20155 -27155
rect 20213 -27189 20223 -27155
rect 20285 -27189 20291 -27155
rect 20357 -27189 20359 -27155
rect 20393 -27189 20395 -27155
rect 20461 -27189 20467 -27155
rect 20529 -27189 20539 -27155
rect 20597 -27189 20611 -27155
rect 20665 -27189 20683 -27155
rect 20733 -27189 20755 -27155
rect 20801 -27189 20827 -27155
rect 20869 -27189 20899 -27155
rect 20937 -27189 20971 -27155
rect 21005 -27189 21039 -27155
rect 21077 -27189 21107 -27155
rect 21149 -27189 21175 -27155
rect 21221 -27189 21243 -27155
rect 21293 -27189 21311 -27155
rect 21365 -27189 21379 -27155
rect 21437 -27189 21447 -27155
rect 21509 -27189 21515 -27155
rect 21581 -27189 21583 -27155
rect 21617 -27189 21619 -27155
rect 21685 -27189 21691 -27155
rect 21753 -27189 21763 -27155
rect 21821 -27189 21835 -27155
rect 21889 -27189 21907 -27155
rect 21957 -27189 21979 -27155
rect 22025 -27189 22051 -27155
rect 22093 -27189 22123 -27155
rect 22161 -27189 22195 -27155
rect 22229 -27189 22263 -27155
rect 22301 -27189 22331 -27155
rect 22373 -27189 22399 -27155
rect 22445 -27189 22467 -27155
rect 22517 -27189 22535 -27155
rect 22589 -27189 22603 -27155
rect 22661 -27189 22671 -27155
rect 22733 -27189 22739 -27155
rect 22805 -27189 22807 -27155
rect 22841 -27189 22843 -27155
rect 22909 -27189 22915 -27155
rect 22977 -27189 22987 -27155
rect 23045 -27189 23059 -27155
rect 23113 -27189 23131 -27155
rect 23181 -27189 23203 -27155
rect 23249 -27189 23275 -27155
rect 23317 -27189 23347 -27155
rect 23385 -27189 23419 -27155
rect 23453 -27189 23487 -27155
rect 23525 -27189 23555 -27155
rect 23597 -27189 23623 -27155
rect 23669 -27189 23691 -27155
rect 23741 -27189 23759 -27155
rect 23813 -27189 23827 -27155
rect 23885 -27189 23895 -27155
rect 23957 -27189 23963 -27155
rect 24029 -27189 24031 -27155
rect 24065 -27189 24067 -27155
rect 24133 -27189 24139 -27155
rect 24201 -27189 24211 -27155
rect 24269 -27189 24283 -27155
rect 24337 -27189 24355 -27155
rect 24405 -27189 24427 -27155
rect 24473 -27189 24499 -27155
rect 24541 -27189 24571 -27155
rect 24609 -27189 24643 -27155
rect 24677 -27189 24711 -27155
rect 24749 -27189 24787 -27155
rect 24821 -27189 24922 -27155
rect -12322 -27222 24922 -27189
<< viali >>
rect 487 4255 521 4289
rect 559 4255 581 4289
rect 581 4255 593 4289
rect 631 4255 649 4289
rect 649 4255 665 4289
rect 703 4255 717 4289
rect 717 4255 737 4289
rect 775 4255 785 4289
rect 785 4255 809 4289
rect 847 4255 853 4289
rect 853 4255 881 4289
rect 919 4255 921 4289
rect 921 4255 953 4289
rect 991 4255 1023 4289
rect 1023 4255 1025 4289
rect 1063 4255 1091 4289
rect 1091 4255 1097 4289
rect 1135 4255 1159 4289
rect 1159 4255 1169 4289
rect 1207 4255 1227 4289
rect 1227 4255 1241 4289
rect 1279 4255 1295 4289
rect 1295 4255 1313 4289
rect 1351 4255 1363 4289
rect 1363 4255 1385 4289
rect 1423 4255 1431 4289
rect 1431 4255 1457 4289
rect 1495 4255 1499 4289
rect 1499 4255 1529 4289
rect 1567 4255 1601 4289
rect 1639 4255 1669 4289
rect 1669 4255 1673 4289
rect 1711 4255 1737 4289
rect 1737 4255 1745 4289
rect 1783 4255 1805 4289
rect 1805 4255 1817 4289
rect 1855 4255 1873 4289
rect 1873 4255 1889 4289
rect 1927 4255 1941 4289
rect 1941 4255 1961 4289
rect 1999 4255 2009 4289
rect 2009 4255 2033 4289
rect 2071 4255 2077 4289
rect 2077 4255 2105 4289
rect 2143 4255 2145 4289
rect 2145 4255 2177 4289
rect 2215 4255 2247 4289
rect 2247 4255 2249 4289
rect 2287 4255 2315 4289
rect 2315 4255 2321 4289
rect 2359 4255 2383 4289
rect 2383 4255 2393 4289
rect 2431 4255 2451 4289
rect 2451 4255 2465 4289
rect 2503 4255 2519 4289
rect 2519 4255 2537 4289
rect 2575 4255 2587 4289
rect 2587 4255 2609 4289
rect 2647 4255 2655 4289
rect 2655 4255 2681 4289
rect 2719 4255 2723 4289
rect 2723 4255 2753 4289
rect 2791 4255 2825 4289
rect 2863 4255 2893 4289
rect 2893 4255 2897 4289
rect 2935 4255 2961 4289
rect 2961 4255 2969 4289
rect 3007 4255 3029 4289
rect 3029 4255 3041 4289
rect 3079 4255 3097 4289
rect 3097 4255 3113 4289
rect 3151 4255 3165 4289
rect 3165 4255 3185 4289
rect 3223 4255 3233 4289
rect 3233 4255 3257 4289
rect 3295 4255 3301 4289
rect 3301 4255 3329 4289
rect 3367 4255 3369 4289
rect 3369 4255 3401 4289
rect 3439 4255 3471 4289
rect 3471 4255 3473 4289
rect 3511 4255 3539 4289
rect 3539 4255 3545 4289
rect 3583 4255 3607 4289
rect 3607 4255 3617 4289
rect 3655 4255 3675 4289
rect 3675 4255 3689 4289
rect 3727 4255 3743 4289
rect 3743 4255 3761 4289
rect 3799 4255 3811 4289
rect 3811 4255 3833 4289
rect 3871 4255 3879 4289
rect 3879 4255 3905 4289
rect 3943 4255 3947 4289
rect 3947 4255 3977 4289
rect 4015 4255 4049 4289
rect 4087 4255 4117 4289
rect 4117 4255 4121 4289
rect 4159 4255 4185 4289
rect 4185 4255 4193 4289
rect 4231 4255 4253 4289
rect 4253 4255 4265 4289
rect 4303 4255 4321 4289
rect 4321 4255 4337 4289
rect 4375 4255 4389 4289
rect 4389 4255 4409 4289
rect 4447 4255 4457 4289
rect 4457 4255 4481 4289
rect 4519 4255 4525 4289
rect 4525 4255 4553 4289
rect 4591 4255 4593 4289
rect 4593 4255 4625 4289
rect 4663 4255 4695 4289
rect 4695 4255 4697 4289
rect 4735 4255 4763 4289
rect 4763 4255 4769 4289
rect 4807 4255 4831 4289
rect 4831 4255 4841 4289
rect 4879 4255 4899 4289
rect 4899 4255 4913 4289
rect 4951 4255 4967 4289
rect 4967 4255 4985 4289
rect 5023 4255 5035 4289
rect 5035 4255 5057 4289
rect 5095 4255 5103 4289
rect 5103 4255 5129 4289
rect 5167 4255 5171 4289
rect 5171 4255 5201 4289
rect 5239 4255 5273 4289
rect 5311 4255 5341 4289
rect 5341 4255 5345 4289
rect 5383 4255 5409 4289
rect 5409 4255 5417 4289
rect 5455 4255 5477 4289
rect 5477 4255 5489 4289
rect 5527 4255 5545 4289
rect 5545 4255 5561 4289
rect 5599 4255 5613 4289
rect 5613 4255 5633 4289
rect 5671 4255 5681 4289
rect 5681 4255 5705 4289
rect 5743 4255 5749 4289
rect 5749 4255 5777 4289
rect 5815 4255 5817 4289
rect 5817 4255 5849 4289
rect 5887 4255 5919 4289
rect 5919 4255 5921 4289
rect 5959 4255 5987 4289
rect 5987 4255 5993 4289
rect 6031 4255 6055 4289
rect 6055 4255 6065 4289
rect 6103 4255 6123 4289
rect 6123 4255 6137 4289
rect 6175 4255 6191 4289
rect 6191 4255 6209 4289
rect 6247 4255 6259 4289
rect 6259 4255 6281 4289
rect 6319 4255 6327 4289
rect 6327 4255 6353 4289
rect 6391 4255 6395 4289
rect 6395 4255 6425 4289
rect 6463 4255 6497 4289
rect 6535 4255 6565 4289
rect 6565 4255 6569 4289
rect 6607 4255 6633 4289
rect 6633 4255 6641 4289
rect 6679 4255 6701 4289
rect 6701 4255 6713 4289
rect 6751 4255 6769 4289
rect 6769 4255 6785 4289
rect 6823 4255 6837 4289
rect 6837 4255 6857 4289
rect 6895 4255 6905 4289
rect 6905 4255 6929 4289
rect 6967 4255 6973 4289
rect 6973 4255 7001 4289
rect 7039 4255 7041 4289
rect 7041 4255 7073 4289
rect 7111 4255 7143 4289
rect 7143 4255 7145 4289
rect 7183 4255 7211 4289
rect 7211 4255 7217 4289
rect 7255 4255 7279 4289
rect 7279 4255 7289 4289
rect 7327 4255 7347 4289
rect 7347 4255 7361 4289
rect 7399 4255 7415 4289
rect 7415 4255 7433 4289
rect 7471 4255 7483 4289
rect 7483 4255 7505 4289
rect 7543 4255 7551 4289
rect 7551 4255 7577 4289
rect 7615 4255 7619 4289
rect 7619 4255 7649 4289
rect 7687 4255 7721 4289
rect 7759 4255 7789 4289
rect 7789 4255 7793 4289
rect 7831 4255 7857 4289
rect 7857 4255 7865 4289
rect 7903 4255 7925 4289
rect 7925 4255 7937 4289
rect 7975 4255 7993 4289
rect 7993 4255 8009 4289
rect 8047 4255 8061 4289
rect 8061 4255 8081 4289
rect 8119 4255 8129 4289
rect 8129 4255 8153 4289
rect 8191 4255 8197 4289
rect 8197 4255 8225 4289
rect 8263 4255 8265 4289
rect 8265 4255 8297 4289
rect 8335 4255 8367 4289
rect 8367 4255 8369 4289
rect 8407 4255 8435 4289
rect 8435 4255 8441 4289
rect 8479 4255 8503 4289
rect 8503 4255 8513 4289
rect 8551 4255 8571 4289
rect 8571 4255 8585 4289
rect 8623 4255 8639 4289
rect 8639 4255 8657 4289
rect 8695 4255 8707 4289
rect 8707 4255 8729 4289
rect 8767 4255 8775 4289
rect 8775 4255 8801 4289
rect 8839 4255 8843 4289
rect 8843 4255 8873 4289
rect 8911 4255 8945 4289
rect 8983 4255 9013 4289
rect 9013 4255 9017 4289
rect 9055 4255 9081 4289
rect 9081 4255 9089 4289
rect 9127 4255 9149 4289
rect 9149 4255 9161 4289
rect 9199 4255 9217 4289
rect 9217 4255 9233 4289
rect 9271 4255 9285 4289
rect 9285 4255 9305 4289
rect 9343 4255 9353 4289
rect 9353 4255 9377 4289
rect 9415 4255 9421 4289
rect 9421 4255 9449 4289
rect 9487 4255 9489 4289
rect 9489 4255 9521 4289
rect 9559 4255 9591 4289
rect 9591 4255 9593 4289
rect 9631 4255 9659 4289
rect 9659 4255 9665 4289
rect 9703 4255 9727 4289
rect 9727 4255 9737 4289
rect 9775 4255 9795 4289
rect 9795 4255 9809 4289
rect 9847 4255 9863 4289
rect 9863 4255 9881 4289
rect 9919 4255 9931 4289
rect 9931 4255 9953 4289
rect 9991 4255 9999 4289
rect 9999 4255 10025 4289
rect 10063 4255 10067 4289
rect 10067 4255 10097 4289
rect 10135 4255 10169 4289
rect 10207 4255 10237 4289
rect 10237 4255 10241 4289
rect 10279 4255 10305 4289
rect 10305 4255 10313 4289
rect 10351 4255 10373 4289
rect 10373 4255 10385 4289
rect 10423 4255 10441 4289
rect 10441 4255 10457 4289
rect 10495 4255 10509 4289
rect 10509 4255 10529 4289
rect 10567 4255 10577 4289
rect 10577 4255 10601 4289
rect 10639 4255 10645 4289
rect 10645 4255 10673 4289
rect 10711 4255 10713 4289
rect 10713 4255 10745 4289
rect 10783 4255 10815 4289
rect 10815 4255 10817 4289
rect 10855 4255 10883 4289
rect 10883 4255 10889 4289
rect 10927 4255 10951 4289
rect 10951 4255 10961 4289
rect 10999 4255 11019 4289
rect 11019 4255 11033 4289
rect 11071 4255 11087 4289
rect 11087 4255 11105 4289
rect 11143 4255 11155 4289
rect 11155 4255 11177 4289
rect 11215 4255 11223 4289
rect 11223 4255 11249 4289
rect 11287 4255 11291 4289
rect 11291 4255 11321 4289
rect 11359 4255 11393 4289
rect 11431 4255 11461 4289
rect 11461 4255 11465 4289
rect 11503 4255 11529 4289
rect 11529 4255 11537 4289
rect 11575 4255 11597 4289
rect 11597 4255 11609 4289
rect 11647 4255 11665 4289
rect 11665 4255 11681 4289
rect 11719 4255 11733 4289
rect 11733 4255 11753 4289
rect 11791 4255 11801 4289
rect 11801 4255 11825 4289
rect 11863 4255 11869 4289
rect 11869 4255 11897 4289
rect 11935 4255 11937 4289
rect 11937 4255 11969 4289
rect 12007 4255 12039 4289
rect 12039 4255 12041 4289
rect 12079 4255 12107 4289
rect 12107 4255 12113 4289
rect 12151 4255 12175 4289
rect 12175 4255 12185 4289
rect 12223 4255 12243 4289
rect 12243 4255 12257 4289
rect 12295 4255 12311 4289
rect 12311 4255 12329 4289
rect 12367 4255 12379 4289
rect 12379 4255 12401 4289
rect 12439 4255 12447 4289
rect 12447 4255 12473 4289
rect 12511 4255 12515 4289
rect 12515 4255 12545 4289
rect 12583 4255 12617 4289
rect 12655 4255 12685 4289
rect 12685 4255 12689 4289
rect 12727 4255 12753 4289
rect 12753 4255 12761 4289
rect 12799 4255 12821 4289
rect 12821 4255 12833 4289
rect 12871 4255 12889 4289
rect 12889 4255 12905 4289
rect 12943 4255 12957 4289
rect 12957 4255 12977 4289
rect 13015 4255 13025 4289
rect 13025 4255 13049 4289
rect 13087 4255 13093 4289
rect 13093 4255 13121 4289
rect 13159 4255 13161 4289
rect 13161 4255 13193 4289
rect 13231 4255 13263 4289
rect 13263 4255 13265 4289
rect 13303 4255 13331 4289
rect 13331 4255 13337 4289
rect 13375 4255 13399 4289
rect 13399 4255 13409 4289
rect 13447 4255 13467 4289
rect 13467 4255 13481 4289
rect 13519 4255 13535 4289
rect 13535 4255 13553 4289
rect 13591 4255 13603 4289
rect 13603 4255 13625 4289
rect 13663 4255 13671 4289
rect 13671 4255 13697 4289
rect 13735 4255 13739 4289
rect 13739 4255 13769 4289
rect 13807 4255 13841 4289
rect 13879 4255 13909 4289
rect 13909 4255 13913 4289
rect 13951 4255 13977 4289
rect 13977 4255 13985 4289
rect 14023 4255 14045 4289
rect 14045 4255 14057 4289
rect 14095 4255 14113 4289
rect 14113 4255 14129 4289
rect 14167 4255 14181 4289
rect 14181 4255 14201 4289
rect 14239 4255 14249 4289
rect 14249 4255 14273 4289
rect 14311 4255 14317 4289
rect 14317 4255 14345 4289
rect 14383 4255 14385 4289
rect 14385 4255 14417 4289
rect 14455 4255 14487 4289
rect 14487 4255 14489 4289
rect 14527 4255 14555 4289
rect 14555 4255 14561 4289
rect 14599 4255 14623 4289
rect 14623 4255 14633 4289
rect 14671 4255 14691 4289
rect 14691 4255 14705 4289
rect 14743 4255 14759 4289
rect 14759 4255 14777 4289
rect 14815 4255 14827 4289
rect 14827 4255 14849 4289
rect 14887 4255 14895 4289
rect 14895 4255 14921 4289
rect 14959 4255 14963 4289
rect 14963 4255 14993 4289
rect 15031 4255 15065 4289
rect 15103 4255 15133 4289
rect 15133 4255 15137 4289
rect 15175 4255 15201 4289
rect 15201 4255 15209 4289
rect 15247 4255 15269 4289
rect 15269 4255 15281 4289
rect 15319 4255 15337 4289
rect 15337 4255 15353 4289
rect 15391 4255 15405 4289
rect 15405 4255 15425 4289
rect 15463 4255 15473 4289
rect 15473 4255 15497 4289
rect 15535 4255 15541 4289
rect 15541 4255 15569 4289
rect 15607 4255 15609 4289
rect 15609 4255 15641 4289
rect 15679 4255 15711 4289
rect 15711 4255 15713 4289
rect 15751 4255 15779 4289
rect 15779 4255 15785 4289
rect 15823 4255 15847 4289
rect 15847 4255 15857 4289
rect 15895 4255 15915 4289
rect 15915 4255 15929 4289
rect 15967 4255 15983 4289
rect 15983 4255 16001 4289
rect 16039 4255 16051 4289
rect 16051 4255 16073 4289
rect 16111 4255 16119 4289
rect 16119 4255 16145 4289
rect 16183 4255 16187 4289
rect 16187 4255 16217 4289
rect 16255 4255 16289 4289
rect 16327 4255 16357 4289
rect 16357 4255 16361 4289
rect 16399 4255 16425 4289
rect 16425 4255 16433 4289
rect 16471 4255 16493 4289
rect 16493 4255 16505 4289
rect 16543 4255 16561 4289
rect 16561 4255 16577 4289
rect 16615 4255 16629 4289
rect 16629 4255 16649 4289
rect 16687 4255 16697 4289
rect 16697 4255 16721 4289
rect 16759 4255 16765 4289
rect 16765 4255 16793 4289
rect 16831 4255 16833 4289
rect 16833 4255 16865 4289
rect 16903 4255 16935 4289
rect 16935 4255 16937 4289
rect 16975 4255 17003 4289
rect 17003 4255 17009 4289
rect 17047 4255 17071 4289
rect 17071 4255 17081 4289
rect 17119 4255 17139 4289
rect 17139 4255 17153 4289
rect 17191 4255 17207 4289
rect 17207 4255 17225 4289
rect 17263 4255 17275 4289
rect 17275 4255 17297 4289
rect 17335 4255 17343 4289
rect 17343 4255 17369 4289
rect 17407 4255 17411 4289
rect 17411 4255 17441 4289
rect 17479 4255 17513 4289
rect 17551 4255 17581 4289
rect 17581 4255 17585 4289
rect 17623 4255 17649 4289
rect 17649 4255 17657 4289
rect 17695 4255 17717 4289
rect 17717 4255 17729 4289
rect 17767 4255 17785 4289
rect 17785 4255 17801 4289
rect 17839 4255 17853 4289
rect 17853 4255 17873 4289
rect 17911 4255 17921 4289
rect 17921 4255 17945 4289
rect 17983 4255 17989 4289
rect 17989 4255 18017 4289
rect 18055 4255 18057 4289
rect 18057 4255 18089 4289
rect 18127 4255 18159 4289
rect 18159 4255 18161 4289
rect 18199 4255 18227 4289
rect 18227 4255 18233 4289
rect 18271 4255 18295 4289
rect 18295 4255 18305 4289
rect 18343 4255 18363 4289
rect 18363 4255 18377 4289
rect 18415 4255 18431 4289
rect 18431 4255 18449 4289
rect 18487 4255 18499 4289
rect 18499 4255 18521 4289
rect 18559 4255 18567 4289
rect 18567 4255 18593 4289
rect 18631 4255 18635 4289
rect 18635 4255 18665 4289
rect 18703 4255 18737 4289
rect 18775 4255 18805 4289
rect 18805 4255 18809 4289
rect 18847 4255 18873 4289
rect 18873 4255 18881 4289
rect 18919 4255 18941 4289
rect 18941 4255 18953 4289
rect 18991 4255 19009 4289
rect 19009 4255 19025 4289
rect 19063 4255 19077 4289
rect 19077 4255 19097 4289
rect 19135 4255 19145 4289
rect 19145 4255 19169 4289
rect 19207 4255 19213 4289
rect 19213 4255 19241 4289
rect 19279 4255 19281 4289
rect 19281 4255 19313 4289
rect 19351 4255 19383 4289
rect 19383 4255 19385 4289
rect 19423 4255 19451 4289
rect 19451 4255 19457 4289
rect 19495 4255 19519 4289
rect 19519 4255 19529 4289
rect 19567 4255 19587 4289
rect 19587 4255 19601 4289
rect 19639 4255 19655 4289
rect 19655 4255 19673 4289
rect 19711 4255 19723 4289
rect 19723 4255 19745 4289
rect 19783 4255 19791 4289
rect 19791 4255 19817 4289
rect 19855 4255 19859 4289
rect 19859 4255 19889 4289
rect 19927 4255 19961 4289
rect 19999 4255 20029 4289
rect 20029 4255 20033 4289
rect 20071 4255 20097 4289
rect 20097 4255 20105 4289
rect 20143 4255 20165 4289
rect 20165 4255 20177 4289
rect 20215 4255 20233 4289
rect 20233 4255 20249 4289
rect 20287 4255 20301 4289
rect 20301 4255 20321 4289
rect 20359 4255 20369 4289
rect 20369 4255 20393 4289
rect 20431 4255 20437 4289
rect 20437 4255 20465 4289
rect 20503 4255 20505 4289
rect 20505 4255 20537 4289
rect 20575 4255 20607 4289
rect 20607 4255 20609 4289
rect 20647 4255 20675 4289
rect 20675 4255 20681 4289
rect 20719 4255 20743 4289
rect 20743 4255 20753 4289
rect 20791 4255 20811 4289
rect 20811 4255 20825 4289
rect 20863 4255 20879 4289
rect 20879 4255 20897 4289
rect 20935 4255 20947 4289
rect 20947 4255 20969 4289
rect 21007 4255 21015 4289
rect 21015 4255 21041 4289
rect 21079 4255 21083 4289
rect 21083 4255 21113 4289
rect 21151 4255 21185 4289
rect 21223 4255 21253 4289
rect 21253 4255 21257 4289
rect 21295 4255 21321 4289
rect 21321 4255 21329 4289
rect 21367 4255 21389 4289
rect 21389 4255 21401 4289
rect 21439 4255 21457 4289
rect 21457 4255 21473 4289
rect 21511 4255 21525 4289
rect 21525 4255 21545 4289
rect 21583 4255 21593 4289
rect 21593 4255 21617 4289
rect 21655 4255 21661 4289
rect 21661 4255 21689 4289
rect 21727 4255 21729 4289
rect 21729 4255 21761 4289
rect 21799 4255 21831 4289
rect 21831 4255 21833 4289
rect 21871 4255 21899 4289
rect 21899 4255 21905 4289
rect 21943 4255 21967 4289
rect 21967 4255 21977 4289
rect 22015 4255 22035 4289
rect 22035 4255 22049 4289
rect 22087 4255 22103 4289
rect 22103 4255 22121 4289
rect 22159 4255 22171 4289
rect 22171 4255 22193 4289
rect 22231 4255 22239 4289
rect 22239 4255 22265 4289
rect 22303 4255 22307 4289
rect 22307 4255 22337 4289
rect 22375 4255 22409 4289
rect 22447 4255 22477 4289
rect 22477 4255 22481 4289
rect 22519 4255 22545 4289
rect 22545 4255 22553 4289
rect 22591 4255 22613 4289
rect 22613 4255 22625 4289
rect 22663 4255 22681 4289
rect 22681 4255 22697 4289
rect 22735 4255 22749 4289
rect 22749 4255 22769 4289
rect 22807 4255 22817 4289
rect 22817 4255 22841 4289
rect 22879 4255 22885 4289
rect 22885 4255 22913 4289
rect 22951 4255 22953 4289
rect 22953 4255 22985 4289
rect 23023 4255 23055 4289
rect 23055 4255 23057 4289
rect 23095 4255 23123 4289
rect 23123 4255 23129 4289
rect 23167 4255 23191 4289
rect 23191 4255 23201 4289
rect 23239 4255 23259 4289
rect 23259 4255 23273 4289
rect 23311 4255 23327 4289
rect 23327 4255 23345 4289
rect 23383 4255 23395 4289
rect 23395 4255 23417 4289
rect 23455 4255 23463 4289
rect 23463 4255 23489 4289
rect 23527 4255 23531 4289
rect 23531 4255 23561 4289
rect 23599 4255 23633 4289
rect 23671 4255 23701 4289
rect 23701 4255 23705 4289
rect 23743 4255 23769 4289
rect 23769 4255 23777 4289
rect 23815 4255 23837 4289
rect 23837 4255 23849 4289
rect 23887 4255 23905 4289
rect 23905 4255 23921 4289
rect 23959 4255 23973 4289
rect 23973 4255 23993 4289
rect 24031 4255 24041 4289
rect 24041 4255 24065 4289
rect 24103 4255 24109 4289
rect 24109 4255 24137 4289
rect 24175 4255 24177 4289
rect 24177 4255 24209 4289
rect 24247 4255 24279 4289
rect 24279 4255 24281 4289
rect 24319 4255 24347 4289
rect 24347 4255 24353 4289
rect 24391 4255 24415 4289
rect 24415 4255 24425 4289
rect 24463 4255 24483 4289
rect 24483 4255 24497 4289
rect 24535 4255 24551 4289
rect 24551 4255 24569 4289
rect 24607 4255 24619 4289
rect 24619 4255 24641 4289
rect 24679 4255 24713 4289
rect 411 3668 445 3700
rect 411 3666 445 3668
rect 411 3600 445 3628
rect 411 3594 445 3600
rect 411 3532 445 3556
rect 411 3522 445 3532
rect 411 3464 445 3484
rect 411 3450 445 3464
rect 411 3396 445 3412
rect 411 3378 445 3396
rect 411 3328 445 3340
rect 411 3306 445 3328
rect 411 3260 445 3268
rect 411 3234 445 3260
rect 411 3192 445 3196
rect 411 3162 445 3192
rect 411 3090 445 3124
rect 411 3022 445 3052
rect 411 3018 445 3022
rect 411 2954 445 2980
rect 411 2946 445 2954
rect 411 2886 445 2908
rect 411 2874 445 2886
rect 411 2818 445 2836
rect 411 2802 445 2818
rect 411 2750 445 2764
rect 411 2730 445 2750
rect 411 2682 445 2692
rect 411 2658 445 2682
rect 411 2614 445 2620
rect 411 2586 445 2614
rect 411 2546 445 2548
rect 411 2514 445 2546
rect 411 2444 445 2476
rect 411 2442 445 2444
rect 411 2376 445 2404
rect 411 2370 445 2376
rect 411 2308 445 2332
rect 411 2298 445 2308
rect 411 2240 445 2260
rect 411 2226 445 2240
rect 411 2172 445 2188
rect 411 2154 445 2172
rect 411 2104 445 2116
rect 411 2082 445 2104
rect 411 2036 445 2044
rect 411 2010 445 2036
rect 411 1968 445 1972
rect 411 1938 445 1968
rect 411 1866 445 1900
rect 411 1798 445 1828
rect 411 1794 445 1798
rect 411 1730 445 1756
rect 411 1722 445 1730
rect 411 1662 445 1684
rect 411 1650 445 1662
rect 411 1594 445 1612
rect 411 1578 445 1594
rect 411 1526 445 1540
rect 411 1506 445 1526
rect 411 1458 445 1468
rect 411 1434 445 1458
rect 411 1390 445 1396
rect 411 1362 445 1390
rect 411 1322 445 1324
rect 411 1290 445 1322
rect 411 1220 445 1252
rect 411 1218 445 1220
rect 411 1152 445 1180
rect 411 1146 445 1152
rect 411 1084 445 1108
rect 411 1074 445 1084
rect 411 1016 445 1036
rect 411 1002 445 1016
rect 411 948 445 964
rect 411 930 445 948
rect 411 880 445 892
rect 411 858 445 880
rect 411 812 445 820
rect 411 786 445 812
rect 411 744 445 748
rect 411 714 445 744
rect 411 642 445 676
rect 411 574 445 604
rect 411 570 445 574
rect 411 506 445 532
rect 411 498 445 506
rect 411 438 445 460
rect 411 426 445 438
rect 411 370 445 388
rect 411 354 445 370
rect 411 302 445 316
rect 411 282 445 302
rect 411 234 445 244
rect 411 210 445 234
rect 411 166 445 172
rect 411 138 445 166
rect 411 98 445 100
rect 411 66 445 98
rect 411 -4 445 28
rect 411 -6 445 -4
rect 411 -72 445 -44
rect 411 -78 445 -72
rect 411 -140 445 -116
rect 411 -150 445 -140
rect 411 -208 445 -188
rect 411 -222 445 -208
rect 411 -276 445 -260
rect 411 -294 445 -276
rect 411 -344 445 -332
rect 411 -366 445 -344
rect 411 -412 445 -404
rect 411 -438 445 -412
rect 411 -480 445 -476
rect 411 -510 445 -480
rect 411 -582 445 -548
rect 411 -650 445 -620
rect 411 -654 445 -650
rect 411 -718 445 -692
rect 411 -726 445 -718
rect 411 -786 445 -764
rect 411 -798 445 -786
rect 411 -854 445 -836
rect 411 -870 445 -854
rect 411 -922 445 -908
rect 411 -942 445 -922
rect 411 -990 445 -980
rect 411 -1014 445 -990
rect 411 -1058 445 -1052
rect 411 -1086 445 -1058
rect 411 -1126 445 -1124
rect 411 -1158 445 -1126
rect 411 -1228 445 -1196
rect 411 -1230 445 -1228
rect 411 -1296 445 -1268
rect 411 -1302 445 -1296
rect 411 -1364 445 -1340
rect 411 -1374 445 -1364
rect 411 -1432 445 -1412
rect 411 -1446 445 -1432
rect 411 -1500 445 -1484
rect 411 -1518 445 -1500
rect 411 -1568 445 -1556
rect 411 -1590 445 -1568
rect 411 -1636 445 -1628
rect 411 -1662 445 -1636
rect 411 -1704 445 -1700
rect 411 -1734 445 -1704
rect 411 -1806 445 -1772
rect 411 -1874 445 -1844
rect 411 -1878 445 -1874
rect 411 -1942 445 -1916
rect 411 -1950 445 -1942
rect 411 -2010 445 -1988
rect 411 -2022 445 -2010
rect 411 -2078 445 -2060
rect 411 -2094 445 -2078
rect 411 -2146 445 -2132
rect 411 -2166 445 -2146
rect 411 -2214 445 -2204
rect 411 -2238 445 -2214
rect 411 -2282 445 -2276
rect 411 -2310 445 -2282
rect 411 -2350 445 -2348
rect 411 -2382 445 -2350
rect 411 -2452 445 -2420
rect 411 -2454 445 -2452
rect 411 -2520 445 -2492
rect 411 -2526 445 -2520
rect 411 -2588 445 -2564
rect 411 -2598 445 -2588
rect 411 -2656 445 -2636
rect 411 -2670 445 -2656
rect 411 -2724 445 -2708
rect 411 -2742 445 -2724
rect 411 -2792 445 -2780
rect 411 -2814 445 -2792
rect 411 -2860 445 -2852
rect 411 -2886 445 -2860
rect 411 -2928 445 -2924
rect 411 -2958 445 -2928
rect 411 -3030 445 -2996
rect 411 -3098 445 -3068
rect 411 -3102 445 -3098
rect 411 -3166 445 -3140
rect 411 -3174 445 -3166
rect 411 -3234 445 -3212
rect 411 -3246 445 -3234
rect 411 -3302 445 -3284
rect 411 -3318 445 -3302
rect 411 -3370 445 -3356
rect 411 -3390 445 -3370
rect 411 -3438 445 -3428
rect 411 -3462 445 -3438
rect 411 -3506 445 -3500
rect 411 -3534 445 -3506
rect 411 -3574 445 -3572
rect 411 -3606 445 -3574
rect 411 -3676 445 -3644
rect 411 -3678 445 -3676
rect 411 -3744 445 -3716
rect 411 -3750 445 -3744
rect 411 -3812 445 -3788
rect 411 -3822 445 -3812
rect 411 -3880 445 -3860
rect 411 -3894 445 -3880
rect 411 -3948 445 -3932
rect 411 -3966 445 -3948
rect 411 -4016 445 -4004
rect 411 -4038 445 -4016
rect 411 -4084 445 -4076
rect 411 -4110 445 -4084
rect 411 -4152 445 -4148
rect 411 -4182 445 -4152
rect 411 -4254 445 -4220
rect 411 -4322 445 -4292
rect 411 -4326 445 -4322
rect 411 -4390 445 -4364
rect 411 -4398 445 -4390
rect 411 -4458 445 -4436
rect 411 -4470 445 -4458
rect 411 -4526 445 -4508
rect 411 -4542 445 -4526
rect 411 -4594 445 -4580
rect 411 -4614 445 -4594
rect 411 -4662 445 -4652
rect 411 -4686 445 -4662
rect 411 -4730 445 -4724
rect 411 -4758 445 -4730
rect 411 -4798 445 -4796
rect 411 -4830 445 -4798
rect 411 -4900 445 -4868
rect 411 -4902 445 -4900
rect 411 -4968 445 -4940
rect 411 -4974 445 -4968
rect 411 -5036 445 -5012
rect 411 -5046 445 -5036
rect 411 -5104 445 -5084
rect 411 -5118 445 -5104
rect 411 -5172 445 -5156
rect 411 -5190 445 -5172
rect 411 -5240 445 -5228
rect 411 -5262 445 -5240
rect 411 -5308 445 -5300
rect 411 -5334 445 -5308
rect 411 -5376 445 -5372
rect 411 -5406 445 -5376
rect 411 -5478 445 -5444
rect 411 -5546 445 -5516
rect 411 -5550 445 -5546
rect 411 -5614 445 -5588
rect 411 -5622 445 -5614
rect 411 -5682 445 -5660
rect 411 -5694 445 -5682
rect 411 -5750 445 -5732
rect 411 -5766 445 -5750
rect 411 -5818 445 -5804
rect 411 -5838 445 -5818
rect 411 -5886 445 -5876
rect 411 -5910 445 -5886
rect 411 -5954 445 -5948
rect 411 -5982 445 -5954
rect 411 -6022 445 -6020
rect 411 -6054 445 -6022
rect 411 -6124 445 -6092
rect 411 -6126 445 -6124
rect 411 -6192 445 -6164
rect 411 -6198 445 -6192
rect 411 -6260 445 -6236
rect 411 -6270 445 -6260
rect 411 -6328 445 -6308
rect 411 -6342 445 -6328
rect 411 -6396 445 -6380
rect 411 -6414 445 -6396
rect 411 -6464 445 -6452
rect 411 -6486 445 -6464
rect 411 -6532 445 -6524
rect 411 -6558 445 -6532
rect 411 -6600 445 -6596
rect 411 -6630 445 -6600
rect 411 -6702 445 -6668
rect 411 -6770 445 -6740
rect 411 -6774 445 -6770
rect 411 -6838 445 -6812
rect 411 -6846 445 -6838
rect 411 -6906 445 -6884
rect 411 -6918 445 -6906
rect 411 -6974 445 -6956
rect 411 -6990 445 -6974
rect 411 -7042 445 -7028
rect 411 -7062 445 -7042
rect 411 -7110 445 -7100
rect 411 -7134 445 -7110
rect 411 -7178 445 -7172
rect 411 -7206 445 -7178
rect 411 -7246 445 -7244
rect 411 -7278 445 -7246
rect 411 -7348 445 -7316
rect 411 -7350 445 -7348
rect 411 -7416 445 -7388
rect 411 -7422 445 -7416
rect 411 -7484 445 -7460
rect 411 -7494 445 -7484
rect 411 -7552 445 -7532
rect 411 -7566 445 -7552
rect 411 -7620 445 -7604
rect 411 -7638 445 -7620
rect 411 -7688 445 -7676
rect 411 -7710 445 -7688
rect 411 -7756 445 -7748
rect 411 -7782 445 -7756
rect 411 -7824 445 -7820
rect 411 -7854 445 -7824
rect 411 -7926 445 -7892
rect 411 -7994 445 -7964
rect 411 -7998 445 -7994
rect 411 -8062 445 -8036
rect 411 -8070 445 -8062
rect 411 -8130 445 -8108
rect 411 -8142 445 -8130
rect 411 -8198 445 -8180
rect 411 -8214 445 -8198
rect 411 -8266 445 -8252
rect 411 -8286 445 -8266
rect 411 -8334 445 -8324
rect 411 -8358 445 -8334
rect 411 -8402 445 -8396
rect 411 -8430 445 -8402
rect 411 -8470 445 -8468
rect 411 -8502 445 -8470
rect 411 -8572 445 -8540
rect 411 -8574 445 -8572
rect 411 -8640 445 -8612
rect 411 -8646 445 -8640
rect 411 -8708 445 -8684
rect 411 -8718 445 -8708
rect 411 -8776 445 -8756
rect 411 -8790 445 -8776
rect 411 -8844 445 -8828
rect 411 -8862 445 -8844
rect 411 -8912 445 -8900
rect 411 -8934 445 -8912
rect 411 -8980 445 -8972
rect 411 -9006 445 -8980
rect 411 -9048 445 -9044
rect 411 -9078 445 -9048
rect 411 -9150 445 -9116
rect 411 -9218 445 -9188
rect 411 -9222 445 -9218
rect 411 -9286 445 -9260
rect 411 -9294 445 -9286
rect 411 -9354 445 -9332
rect 411 -9366 445 -9354
rect 411 -9422 445 -9404
rect 411 -9438 445 -9422
rect 411 -9490 445 -9476
rect 411 -9510 445 -9490
rect 411 -9558 445 -9548
rect 411 -9582 445 -9558
rect 411 -9626 445 -9620
rect 411 -9654 445 -9626
rect 411 -9694 445 -9692
rect 411 -9726 445 -9694
rect 24755 3668 24789 3700
rect 24755 3666 24789 3668
rect 24755 3600 24789 3628
rect 24755 3594 24789 3600
rect 24755 3532 24789 3556
rect 24755 3522 24789 3532
rect 24755 3464 24789 3484
rect 24755 3450 24789 3464
rect 24755 3396 24789 3412
rect 24755 3378 24789 3396
rect 24755 3328 24789 3340
rect 24755 3306 24789 3328
rect 24755 3260 24789 3268
rect 24755 3234 24789 3260
rect 24755 3192 24789 3196
rect 24755 3162 24789 3192
rect 24755 3090 24789 3124
rect 24755 3022 24789 3052
rect 24755 3018 24789 3022
rect 24755 2954 24789 2980
rect 24755 2946 24789 2954
rect 24755 2886 24789 2908
rect 24755 2874 24789 2886
rect 24755 2818 24789 2836
rect 24755 2802 24789 2818
rect 24755 2750 24789 2764
rect 24755 2730 24789 2750
rect 24755 2682 24789 2692
rect 24755 2658 24789 2682
rect 24755 2614 24789 2620
rect 24755 2586 24789 2614
rect 24755 2546 24789 2548
rect 24755 2514 24789 2546
rect 24755 2444 24789 2476
rect 24755 2442 24789 2444
rect 24755 2376 24789 2404
rect 24755 2370 24789 2376
rect 24755 2308 24789 2332
rect 24755 2298 24789 2308
rect 24755 2240 24789 2260
rect 24755 2226 24789 2240
rect 24755 2172 24789 2188
rect 24755 2154 24789 2172
rect 24755 2104 24789 2116
rect 24755 2082 24789 2104
rect 24755 2036 24789 2044
rect 24755 2010 24789 2036
rect 24755 1968 24789 1972
rect 24755 1938 24789 1968
rect 24755 1866 24789 1900
rect 24755 1798 24789 1828
rect 24755 1794 24789 1798
rect 24755 1730 24789 1756
rect 24755 1722 24789 1730
rect 24755 1662 24789 1684
rect 24755 1650 24789 1662
rect 24755 1594 24789 1612
rect 24755 1578 24789 1594
rect 24755 1526 24789 1540
rect 24755 1506 24789 1526
rect 24755 1458 24789 1468
rect 24755 1434 24789 1458
rect 24755 1390 24789 1396
rect 24755 1362 24789 1390
rect 24755 1322 24789 1324
rect 24755 1290 24789 1322
rect 24755 1220 24789 1252
rect 24755 1218 24789 1220
rect 24755 1152 24789 1180
rect 24755 1146 24789 1152
rect 24755 1084 24789 1108
rect 24755 1074 24789 1084
rect 24755 1016 24789 1036
rect 24755 1002 24789 1016
rect 24755 948 24789 964
rect 24755 930 24789 948
rect 24755 880 24789 892
rect 24755 858 24789 880
rect 24755 812 24789 820
rect 24755 786 24789 812
rect 24755 744 24789 748
rect 24755 714 24789 744
rect 24755 642 24789 676
rect 24755 574 24789 604
rect 24755 570 24789 574
rect 24755 506 24789 532
rect 24755 498 24789 506
rect 24755 438 24789 460
rect 24755 426 24789 438
rect 24755 370 24789 388
rect 24755 354 24789 370
rect 24755 302 24789 316
rect 24755 282 24789 302
rect 24755 234 24789 244
rect 24755 210 24789 234
rect 24755 166 24789 172
rect 24755 138 24789 166
rect 24755 98 24789 100
rect 24755 66 24789 98
rect 24755 -4 24789 28
rect 24755 -6 24789 -4
rect 24755 -72 24789 -44
rect 24755 -78 24789 -72
rect 24755 -140 24789 -116
rect 24755 -150 24789 -140
rect 24755 -208 24789 -188
rect 24755 -222 24789 -208
rect 24755 -276 24789 -260
rect 24755 -294 24789 -276
rect 24755 -344 24789 -332
rect 24755 -366 24789 -344
rect 24755 -412 24789 -404
rect 24755 -438 24789 -412
rect 24755 -480 24789 -476
rect 24755 -510 24789 -480
rect 24755 -582 24789 -548
rect 24755 -650 24789 -620
rect 24755 -654 24789 -650
rect 24755 -718 24789 -692
rect 24755 -726 24789 -718
rect 24755 -786 24789 -764
rect 24755 -798 24789 -786
rect 24755 -854 24789 -836
rect 24755 -870 24789 -854
rect 24755 -922 24789 -908
rect 24755 -942 24789 -922
rect 24755 -990 24789 -980
rect 24755 -1014 24789 -990
rect 24755 -1058 24789 -1052
rect 24755 -1086 24789 -1058
rect 24755 -1126 24789 -1124
rect 24755 -1158 24789 -1126
rect 24755 -1228 24789 -1196
rect 24755 -1230 24789 -1228
rect 24755 -1296 24789 -1268
rect 24755 -1302 24789 -1296
rect 24755 -1364 24789 -1340
rect 24755 -1374 24789 -1364
rect 24755 -1432 24789 -1412
rect 24755 -1446 24789 -1432
rect 24755 -1500 24789 -1484
rect 24755 -1518 24789 -1500
rect 24755 -1568 24789 -1556
rect 24755 -1590 24789 -1568
rect 24755 -1636 24789 -1628
rect 24755 -1662 24789 -1636
rect 24755 -1704 24789 -1700
rect 24755 -1734 24789 -1704
rect 24755 -1806 24789 -1772
rect 24755 -1874 24789 -1844
rect 24755 -1878 24789 -1874
rect 24755 -1942 24789 -1916
rect 24755 -1950 24789 -1942
rect 24755 -2010 24789 -1988
rect 24755 -2022 24789 -2010
rect 24755 -2078 24789 -2060
rect 24755 -2094 24789 -2078
rect 24755 -2146 24789 -2132
rect 24755 -2166 24789 -2146
rect 24755 -2214 24789 -2204
rect 24755 -2238 24789 -2214
rect 24755 -2282 24789 -2276
rect 24755 -2310 24789 -2282
rect 24755 -2350 24789 -2348
rect 24755 -2382 24789 -2350
rect 24755 -2452 24789 -2420
rect 24755 -2454 24789 -2452
rect 24755 -2520 24789 -2492
rect 24755 -2526 24789 -2520
rect 24755 -2588 24789 -2564
rect 24755 -2598 24789 -2588
rect 24755 -2656 24789 -2636
rect 24755 -2670 24789 -2656
rect 24755 -2724 24789 -2708
rect 24755 -2742 24789 -2724
rect 24755 -2792 24789 -2780
rect 24755 -2814 24789 -2792
rect 24755 -2860 24789 -2852
rect 24755 -2886 24789 -2860
rect 24755 -2928 24789 -2924
rect 24755 -2958 24789 -2928
rect 24755 -3030 24789 -2996
rect 24755 -3098 24789 -3068
rect 24755 -3102 24789 -3098
rect 24755 -3166 24789 -3140
rect 24755 -3174 24789 -3166
rect 24755 -3234 24789 -3212
rect 24755 -3246 24789 -3234
rect 24755 -3302 24789 -3284
rect 24755 -3318 24789 -3302
rect 24755 -3370 24789 -3356
rect 24755 -3390 24789 -3370
rect 24755 -3438 24789 -3428
rect 24755 -3462 24789 -3438
rect 24755 -3506 24789 -3500
rect 24755 -3534 24789 -3506
rect 24755 -3574 24789 -3572
rect 24755 -3606 24789 -3574
rect 24755 -3676 24789 -3644
rect 24755 -3678 24789 -3676
rect 24755 -3744 24789 -3716
rect 24755 -3750 24789 -3744
rect 24755 -3812 24789 -3788
rect 24755 -3822 24789 -3812
rect 24755 -3880 24789 -3860
rect 24755 -3894 24789 -3880
rect 24755 -3948 24789 -3932
rect 24755 -3966 24789 -3948
rect 24755 -4016 24789 -4004
rect 24755 -4038 24789 -4016
rect 24755 -4084 24789 -4076
rect 24755 -4110 24789 -4084
rect 24755 -4152 24789 -4148
rect 24755 -4182 24789 -4152
rect 24755 -4254 24789 -4220
rect 24755 -4322 24789 -4292
rect 24755 -4326 24789 -4322
rect 24755 -4390 24789 -4364
rect 24755 -4398 24789 -4390
rect 24755 -4458 24789 -4436
rect 24755 -4470 24789 -4458
rect 24755 -4526 24789 -4508
rect 24755 -4542 24789 -4526
rect 24755 -4594 24789 -4580
rect 24755 -4614 24789 -4594
rect 24755 -4662 24789 -4652
rect 24755 -4686 24789 -4662
rect 24755 -4730 24789 -4724
rect 24755 -4758 24789 -4730
rect 24755 -4798 24789 -4796
rect 24755 -4830 24789 -4798
rect 24755 -4900 24789 -4868
rect 24755 -4902 24789 -4900
rect 24755 -4968 24789 -4940
rect 24755 -4974 24789 -4968
rect 24755 -5036 24789 -5012
rect 24755 -5046 24789 -5036
rect 24755 -5104 24789 -5084
rect 24755 -5118 24789 -5104
rect 24755 -5172 24789 -5156
rect 24755 -5190 24789 -5172
rect 24755 -5240 24789 -5228
rect 24755 -5262 24789 -5240
rect 24755 -5308 24789 -5300
rect 24755 -5334 24789 -5308
rect 24755 -5376 24789 -5372
rect 24755 -5406 24789 -5376
rect 24755 -5478 24789 -5444
rect 24755 -5546 24789 -5516
rect 24755 -5550 24789 -5546
rect 24755 -5614 24789 -5588
rect 24755 -5622 24789 -5614
rect 24755 -5682 24789 -5660
rect 24755 -5694 24789 -5682
rect 24755 -5750 24789 -5732
rect 24755 -5766 24789 -5750
rect 24755 -5818 24789 -5804
rect 24755 -5838 24789 -5818
rect 24755 -5886 24789 -5876
rect 24755 -5910 24789 -5886
rect 24755 -5954 24789 -5948
rect 24755 -5982 24789 -5954
rect 24755 -6022 24789 -6020
rect 24755 -6054 24789 -6022
rect 24755 -6124 24789 -6092
rect 24755 -6126 24789 -6124
rect 24755 -6192 24789 -6164
rect 24755 -6198 24789 -6192
rect 24755 -6260 24789 -6236
rect 24755 -6270 24789 -6260
rect 24755 -6328 24789 -6308
rect 24755 -6342 24789 -6328
rect 24755 -6396 24789 -6380
rect 24755 -6414 24789 -6396
rect 24755 -6464 24789 -6452
rect 24755 -6486 24789 -6464
rect 24755 -6532 24789 -6524
rect 24755 -6558 24789 -6532
rect 24755 -6600 24789 -6596
rect 24755 -6630 24789 -6600
rect 24755 -6702 24789 -6668
rect 24755 -6770 24789 -6740
rect 24755 -6774 24789 -6770
rect 24755 -6838 24789 -6812
rect 24755 -6846 24789 -6838
rect 24755 -6906 24789 -6884
rect 24755 -6918 24789 -6906
rect 24755 -6974 24789 -6956
rect 24755 -6990 24789 -6974
rect 24755 -7042 24789 -7028
rect 24755 -7062 24789 -7042
rect 24755 -7110 24789 -7100
rect 24755 -7134 24789 -7110
rect 24755 -7178 24789 -7172
rect 24755 -7206 24789 -7178
rect 24755 -7246 24789 -7244
rect 24755 -7278 24789 -7246
rect 24755 -7348 24789 -7316
rect 24755 -7350 24789 -7348
rect 24755 -7416 24789 -7388
rect 24755 -7422 24789 -7416
rect 24755 -7484 24789 -7460
rect 24755 -7494 24789 -7484
rect 24755 -7552 24789 -7532
rect 24755 -7566 24789 -7552
rect 24755 -7620 24789 -7604
rect 24755 -7638 24789 -7620
rect 24755 -7688 24789 -7676
rect 24755 -7710 24789 -7688
rect 24755 -7756 24789 -7748
rect 24755 -7782 24789 -7756
rect 24755 -7824 24789 -7820
rect 24755 -7854 24789 -7824
rect 24755 -7926 24789 -7892
rect 24755 -7994 24789 -7964
rect 24755 -7998 24789 -7994
rect 24755 -8062 24789 -8036
rect 24755 -8070 24789 -8062
rect 24755 -8130 24789 -8108
rect 24755 -8142 24789 -8130
rect 24755 -8198 24789 -8180
rect 24755 -8214 24789 -8198
rect 24755 -8266 24789 -8252
rect 24755 -8286 24789 -8266
rect 24755 -8334 24789 -8324
rect 24755 -8358 24789 -8334
rect 24755 -8402 24789 -8396
rect 24755 -8430 24789 -8402
rect 24755 -8470 24789 -8468
rect 24755 -8502 24789 -8470
rect 24755 -8572 24789 -8540
rect 24755 -8574 24789 -8572
rect 24755 -8640 24789 -8612
rect 24755 -8646 24789 -8640
rect 24755 -8708 24789 -8684
rect 24755 -8718 24789 -8708
rect 24755 -8776 24789 -8756
rect 24755 -8790 24789 -8776
rect 24755 -8844 24789 -8828
rect 24755 -8862 24789 -8844
rect 24755 -8912 24789 -8900
rect 24755 -8934 24789 -8912
rect 24755 -8980 24789 -8972
rect 24755 -9006 24789 -8980
rect 24755 -9048 24789 -9044
rect 24755 -9078 24789 -9048
rect 24755 -9150 24789 -9116
rect 24755 -9218 24789 -9188
rect 24755 -9222 24789 -9218
rect 24755 -9286 24789 -9260
rect 24755 -9294 24789 -9286
rect 24755 -9354 24789 -9332
rect 24755 -9366 24789 -9354
rect 24755 -9422 24789 -9404
rect 24755 -9438 24789 -9422
rect 24755 -9490 24789 -9476
rect 24755 -9510 24789 -9490
rect 24755 -9558 24789 -9548
rect 24755 -9582 24789 -9558
rect 24755 -9626 24789 -9620
rect 24755 -9654 24789 -9626
rect 24755 -9694 24789 -9692
rect 24755 -9726 24789 -9694
rect 487 -10315 521 -10281
rect 559 -10315 581 -10281
rect 581 -10315 593 -10281
rect 631 -10315 649 -10281
rect 649 -10315 665 -10281
rect 703 -10315 717 -10281
rect 717 -10315 737 -10281
rect 775 -10315 785 -10281
rect 785 -10315 809 -10281
rect 847 -10315 853 -10281
rect 853 -10315 881 -10281
rect 919 -10315 921 -10281
rect 921 -10315 953 -10281
rect 991 -10315 1023 -10281
rect 1023 -10315 1025 -10281
rect 1063 -10315 1091 -10281
rect 1091 -10315 1097 -10281
rect 1135 -10315 1159 -10281
rect 1159 -10315 1169 -10281
rect 1207 -10315 1227 -10281
rect 1227 -10315 1241 -10281
rect 1279 -10315 1295 -10281
rect 1295 -10315 1313 -10281
rect 1351 -10315 1363 -10281
rect 1363 -10315 1385 -10281
rect 1423 -10315 1431 -10281
rect 1431 -10315 1457 -10281
rect 1495 -10315 1499 -10281
rect 1499 -10315 1529 -10281
rect 1567 -10315 1601 -10281
rect 1639 -10315 1669 -10281
rect 1669 -10315 1673 -10281
rect 1711 -10315 1737 -10281
rect 1737 -10315 1745 -10281
rect 1783 -10315 1805 -10281
rect 1805 -10315 1817 -10281
rect 1855 -10315 1873 -10281
rect 1873 -10315 1889 -10281
rect 1927 -10315 1941 -10281
rect 1941 -10315 1961 -10281
rect 1999 -10315 2009 -10281
rect 2009 -10315 2033 -10281
rect 2071 -10315 2077 -10281
rect 2077 -10315 2105 -10281
rect 2143 -10315 2145 -10281
rect 2145 -10315 2177 -10281
rect 2215 -10315 2247 -10281
rect 2247 -10315 2249 -10281
rect 2287 -10315 2315 -10281
rect 2315 -10315 2321 -10281
rect 2359 -10315 2383 -10281
rect 2383 -10315 2393 -10281
rect 2431 -10315 2451 -10281
rect 2451 -10315 2465 -10281
rect 2503 -10315 2519 -10281
rect 2519 -10315 2537 -10281
rect 2575 -10315 2587 -10281
rect 2587 -10315 2609 -10281
rect 2647 -10315 2655 -10281
rect 2655 -10315 2681 -10281
rect 2719 -10315 2723 -10281
rect 2723 -10315 2753 -10281
rect 2791 -10315 2825 -10281
rect 2863 -10315 2893 -10281
rect 2893 -10315 2897 -10281
rect 2935 -10315 2961 -10281
rect 2961 -10315 2969 -10281
rect 3007 -10315 3029 -10281
rect 3029 -10315 3041 -10281
rect 3079 -10315 3097 -10281
rect 3097 -10315 3113 -10281
rect 3151 -10315 3165 -10281
rect 3165 -10315 3185 -10281
rect 3223 -10315 3233 -10281
rect 3233 -10315 3257 -10281
rect 3295 -10315 3301 -10281
rect 3301 -10315 3329 -10281
rect 3367 -10315 3369 -10281
rect 3369 -10315 3401 -10281
rect 3439 -10315 3471 -10281
rect 3471 -10315 3473 -10281
rect 3511 -10315 3539 -10281
rect 3539 -10315 3545 -10281
rect 3583 -10315 3607 -10281
rect 3607 -10315 3617 -10281
rect 3655 -10315 3675 -10281
rect 3675 -10315 3689 -10281
rect 3727 -10315 3743 -10281
rect 3743 -10315 3761 -10281
rect 3799 -10315 3811 -10281
rect 3811 -10315 3833 -10281
rect 3871 -10315 3879 -10281
rect 3879 -10315 3905 -10281
rect 3943 -10315 3947 -10281
rect 3947 -10315 3977 -10281
rect 4015 -10315 4049 -10281
rect 4087 -10315 4117 -10281
rect 4117 -10315 4121 -10281
rect 4159 -10315 4185 -10281
rect 4185 -10315 4193 -10281
rect 4231 -10315 4253 -10281
rect 4253 -10315 4265 -10281
rect 4303 -10315 4321 -10281
rect 4321 -10315 4337 -10281
rect 4375 -10315 4389 -10281
rect 4389 -10315 4409 -10281
rect 4447 -10315 4457 -10281
rect 4457 -10315 4481 -10281
rect 4519 -10315 4525 -10281
rect 4525 -10315 4553 -10281
rect 4591 -10315 4593 -10281
rect 4593 -10315 4625 -10281
rect 4663 -10315 4695 -10281
rect 4695 -10315 4697 -10281
rect 4735 -10315 4763 -10281
rect 4763 -10315 4769 -10281
rect 4807 -10315 4831 -10281
rect 4831 -10315 4841 -10281
rect 4879 -10315 4899 -10281
rect 4899 -10315 4913 -10281
rect 4951 -10315 4967 -10281
rect 4967 -10315 4985 -10281
rect 5023 -10315 5035 -10281
rect 5035 -10315 5057 -10281
rect 5095 -10315 5103 -10281
rect 5103 -10315 5129 -10281
rect 5167 -10315 5171 -10281
rect 5171 -10315 5201 -10281
rect 5239 -10315 5273 -10281
rect 5311 -10315 5341 -10281
rect 5341 -10315 5345 -10281
rect 5383 -10315 5409 -10281
rect 5409 -10315 5417 -10281
rect 5455 -10315 5477 -10281
rect 5477 -10315 5489 -10281
rect 5527 -10315 5545 -10281
rect 5545 -10315 5561 -10281
rect 5599 -10315 5613 -10281
rect 5613 -10315 5633 -10281
rect 5671 -10315 5681 -10281
rect 5681 -10315 5705 -10281
rect 5743 -10315 5749 -10281
rect 5749 -10315 5777 -10281
rect 5815 -10315 5817 -10281
rect 5817 -10315 5849 -10281
rect 5887 -10315 5919 -10281
rect 5919 -10315 5921 -10281
rect 5959 -10315 5987 -10281
rect 5987 -10315 5993 -10281
rect 6031 -10315 6055 -10281
rect 6055 -10315 6065 -10281
rect 6103 -10315 6123 -10281
rect 6123 -10315 6137 -10281
rect 6175 -10315 6191 -10281
rect 6191 -10315 6209 -10281
rect 6247 -10315 6259 -10281
rect 6259 -10315 6281 -10281
rect 6319 -10315 6327 -10281
rect 6327 -10315 6353 -10281
rect 6391 -10315 6395 -10281
rect 6395 -10315 6425 -10281
rect 6463 -10315 6497 -10281
rect 6535 -10315 6565 -10281
rect 6565 -10315 6569 -10281
rect 6607 -10315 6633 -10281
rect 6633 -10315 6641 -10281
rect 6679 -10315 6701 -10281
rect 6701 -10315 6713 -10281
rect 6751 -10315 6769 -10281
rect 6769 -10315 6785 -10281
rect 6823 -10315 6837 -10281
rect 6837 -10315 6857 -10281
rect 6895 -10315 6905 -10281
rect 6905 -10315 6929 -10281
rect 6967 -10315 6973 -10281
rect 6973 -10315 7001 -10281
rect 7039 -10315 7041 -10281
rect 7041 -10315 7073 -10281
rect 7111 -10315 7143 -10281
rect 7143 -10315 7145 -10281
rect 7183 -10315 7211 -10281
rect 7211 -10315 7217 -10281
rect 7255 -10315 7279 -10281
rect 7279 -10315 7289 -10281
rect 7327 -10315 7347 -10281
rect 7347 -10315 7361 -10281
rect 7399 -10315 7415 -10281
rect 7415 -10315 7433 -10281
rect 7471 -10315 7483 -10281
rect 7483 -10315 7505 -10281
rect 7543 -10315 7551 -10281
rect 7551 -10315 7577 -10281
rect 7615 -10315 7619 -10281
rect 7619 -10315 7649 -10281
rect 7687 -10315 7721 -10281
rect 7759 -10315 7789 -10281
rect 7789 -10315 7793 -10281
rect 7831 -10315 7857 -10281
rect 7857 -10315 7865 -10281
rect 7903 -10315 7925 -10281
rect 7925 -10315 7937 -10281
rect 7975 -10315 7993 -10281
rect 7993 -10315 8009 -10281
rect 8047 -10315 8061 -10281
rect 8061 -10315 8081 -10281
rect 8119 -10315 8129 -10281
rect 8129 -10315 8153 -10281
rect 8191 -10315 8197 -10281
rect 8197 -10315 8225 -10281
rect 8263 -10315 8265 -10281
rect 8265 -10315 8297 -10281
rect 8335 -10315 8367 -10281
rect 8367 -10315 8369 -10281
rect 8407 -10315 8435 -10281
rect 8435 -10315 8441 -10281
rect 8479 -10315 8503 -10281
rect 8503 -10315 8513 -10281
rect 8551 -10315 8571 -10281
rect 8571 -10315 8585 -10281
rect 8623 -10315 8639 -10281
rect 8639 -10315 8657 -10281
rect 8695 -10315 8707 -10281
rect 8707 -10315 8729 -10281
rect 8767 -10315 8775 -10281
rect 8775 -10315 8801 -10281
rect 8839 -10315 8843 -10281
rect 8843 -10315 8873 -10281
rect 8911 -10315 8945 -10281
rect 8983 -10315 9013 -10281
rect 9013 -10315 9017 -10281
rect 9055 -10315 9081 -10281
rect 9081 -10315 9089 -10281
rect 9127 -10315 9149 -10281
rect 9149 -10315 9161 -10281
rect 9199 -10315 9217 -10281
rect 9217 -10315 9233 -10281
rect 9271 -10315 9285 -10281
rect 9285 -10315 9305 -10281
rect 9343 -10315 9353 -10281
rect 9353 -10315 9377 -10281
rect 9415 -10315 9421 -10281
rect 9421 -10315 9449 -10281
rect 9487 -10315 9489 -10281
rect 9489 -10315 9521 -10281
rect 9559 -10315 9591 -10281
rect 9591 -10315 9593 -10281
rect 9631 -10315 9659 -10281
rect 9659 -10315 9665 -10281
rect 9703 -10315 9727 -10281
rect 9727 -10315 9737 -10281
rect 9775 -10315 9795 -10281
rect 9795 -10315 9809 -10281
rect 9847 -10315 9863 -10281
rect 9863 -10315 9881 -10281
rect 9919 -10315 9931 -10281
rect 9931 -10315 9953 -10281
rect 9991 -10315 9999 -10281
rect 9999 -10315 10025 -10281
rect 10063 -10315 10067 -10281
rect 10067 -10315 10097 -10281
rect 10135 -10315 10169 -10281
rect 10207 -10315 10237 -10281
rect 10237 -10315 10241 -10281
rect 10279 -10315 10305 -10281
rect 10305 -10315 10313 -10281
rect 10351 -10315 10373 -10281
rect 10373 -10315 10385 -10281
rect 10423 -10315 10441 -10281
rect 10441 -10315 10457 -10281
rect 10495 -10315 10509 -10281
rect 10509 -10315 10529 -10281
rect 10567 -10315 10577 -10281
rect 10577 -10315 10601 -10281
rect 10639 -10315 10645 -10281
rect 10645 -10315 10673 -10281
rect 10711 -10315 10713 -10281
rect 10713 -10315 10745 -10281
rect 10783 -10315 10815 -10281
rect 10815 -10315 10817 -10281
rect 10855 -10315 10883 -10281
rect 10883 -10315 10889 -10281
rect 10927 -10315 10951 -10281
rect 10951 -10315 10961 -10281
rect 10999 -10315 11019 -10281
rect 11019 -10315 11033 -10281
rect 11071 -10315 11087 -10281
rect 11087 -10315 11105 -10281
rect 11143 -10315 11155 -10281
rect 11155 -10315 11177 -10281
rect 11215 -10315 11223 -10281
rect 11223 -10315 11249 -10281
rect 11287 -10315 11291 -10281
rect 11291 -10315 11321 -10281
rect 11359 -10315 11393 -10281
rect 11431 -10315 11461 -10281
rect 11461 -10315 11465 -10281
rect 11503 -10315 11529 -10281
rect 11529 -10315 11537 -10281
rect 11575 -10315 11597 -10281
rect 11597 -10315 11609 -10281
rect 11647 -10315 11665 -10281
rect 11665 -10315 11681 -10281
rect 11719 -10315 11733 -10281
rect 11733 -10315 11753 -10281
rect 11791 -10315 11801 -10281
rect 11801 -10315 11825 -10281
rect 11863 -10315 11869 -10281
rect 11869 -10315 11897 -10281
rect 11935 -10315 11937 -10281
rect 11937 -10315 11969 -10281
rect 12007 -10315 12039 -10281
rect 12039 -10315 12041 -10281
rect 12079 -10315 12107 -10281
rect 12107 -10315 12113 -10281
rect 12151 -10315 12175 -10281
rect 12175 -10315 12185 -10281
rect 12223 -10315 12243 -10281
rect 12243 -10315 12257 -10281
rect 12295 -10315 12311 -10281
rect 12311 -10315 12329 -10281
rect 12367 -10315 12379 -10281
rect 12379 -10315 12401 -10281
rect 12439 -10315 12447 -10281
rect 12447 -10315 12473 -10281
rect 12511 -10315 12515 -10281
rect 12515 -10315 12545 -10281
rect 12583 -10315 12617 -10281
rect 12655 -10315 12685 -10281
rect 12685 -10315 12689 -10281
rect 12727 -10315 12753 -10281
rect 12753 -10315 12761 -10281
rect 12799 -10315 12821 -10281
rect 12821 -10315 12833 -10281
rect 12871 -10315 12889 -10281
rect 12889 -10315 12905 -10281
rect 12943 -10315 12957 -10281
rect 12957 -10315 12977 -10281
rect 13015 -10315 13025 -10281
rect 13025 -10315 13049 -10281
rect 13087 -10315 13093 -10281
rect 13093 -10315 13121 -10281
rect 13159 -10315 13161 -10281
rect 13161 -10315 13193 -10281
rect 13231 -10315 13263 -10281
rect 13263 -10315 13265 -10281
rect 13303 -10315 13331 -10281
rect 13331 -10315 13337 -10281
rect 13375 -10315 13399 -10281
rect 13399 -10315 13409 -10281
rect 13447 -10315 13467 -10281
rect 13467 -10315 13481 -10281
rect 13519 -10315 13535 -10281
rect 13535 -10315 13553 -10281
rect 13591 -10315 13603 -10281
rect 13603 -10315 13625 -10281
rect 13663 -10315 13671 -10281
rect 13671 -10315 13697 -10281
rect 13735 -10315 13739 -10281
rect 13739 -10315 13769 -10281
rect 13807 -10315 13841 -10281
rect 13879 -10315 13909 -10281
rect 13909 -10315 13913 -10281
rect 13951 -10315 13977 -10281
rect 13977 -10315 13985 -10281
rect 14023 -10315 14045 -10281
rect 14045 -10315 14057 -10281
rect 14095 -10315 14113 -10281
rect 14113 -10315 14129 -10281
rect 14167 -10315 14181 -10281
rect 14181 -10315 14201 -10281
rect 14239 -10315 14249 -10281
rect 14249 -10315 14273 -10281
rect 14311 -10315 14317 -10281
rect 14317 -10315 14345 -10281
rect 14383 -10315 14385 -10281
rect 14385 -10315 14417 -10281
rect 14455 -10315 14487 -10281
rect 14487 -10315 14489 -10281
rect 14527 -10315 14555 -10281
rect 14555 -10315 14561 -10281
rect 14599 -10315 14623 -10281
rect 14623 -10315 14633 -10281
rect 14671 -10315 14691 -10281
rect 14691 -10315 14705 -10281
rect 14743 -10315 14759 -10281
rect 14759 -10315 14777 -10281
rect 14815 -10315 14827 -10281
rect 14827 -10315 14849 -10281
rect 14887 -10315 14895 -10281
rect 14895 -10315 14921 -10281
rect 14959 -10315 14963 -10281
rect 14963 -10315 14993 -10281
rect 15031 -10315 15065 -10281
rect 15103 -10315 15133 -10281
rect 15133 -10315 15137 -10281
rect 15175 -10315 15201 -10281
rect 15201 -10315 15209 -10281
rect 15247 -10315 15269 -10281
rect 15269 -10315 15281 -10281
rect 15319 -10315 15337 -10281
rect 15337 -10315 15353 -10281
rect 15391 -10315 15405 -10281
rect 15405 -10315 15425 -10281
rect 15463 -10315 15473 -10281
rect 15473 -10315 15497 -10281
rect 15535 -10315 15541 -10281
rect 15541 -10315 15569 -10281
rect 15607 -10315 15609 -10281
rect 15609 -10315 15641 -10281
rect 15679 -10315 15711 -10281
rect 15711 -10315 15713 -10281
rect 15751 -10315 15779 -10281
rect 15779 -10315 15785 -10281
rect 15823 -10315 15847 -10281
rect 15847 -10315 15857 -10281
rect 15895 -10315 15915 -10281
rect 15915 -10315 15929 -10281
rect 15967 -10315 15983 -10281
rect 15983 -10315 16001 -10281
rect 16039 -10315 16051 -10281
rect 16051 -10315 16073 -10281
rect 16111 -10315 16119 -10281
rect 16119 -10315 16145 -10281
rect 16183 -10315 16187 -10281
rect 16187 -10315 16217 -10281
rect 16255 -10315 16289 -10281
rect 16327 -10315 16357 -10281
rect 16357 -10315 16361 -10281
rect 16399 -10315 16425 -10281
rect 16425 -10315 16433 -10281
rect 16471 -10315 16493 -10281
rect 16493 -10315 16505 -10281
rect 16543 -10315 16561 -10281
rect 16561 -10315 16577 -10281
rect 16615 -10315 16629 -10281
rect 16629 -10315 16649 -10281
rect 16687 -10315 16697 -10281
rect 16697 -10315 16721 -10281
rect 16759 -10315 16765 -10281
rect 16765 -10315 16793 -10281
rect 16831 -10315 16833 -10281
rect 16833 -10315 16865 -10281
rect 16903 -10315 16935 -10281
rect 16935 -10315 16937 -10281
rect 16975 -10315 17003 -10281
rect 17003 -10315 17009 -10281
rect 17047 -10315 17071 -10281
rect 17071 -10315 17081 -10281
rect 17119 -10315 17139 -10281
rect 17139 -10315 17153 -10281
rect 17191 -10315 17207 -10281
rect 17207 -10315 17225 -10281
rect 17263 -10315 17275 -10281
rect 17275 -10315 17297 -10281
rect 17335 -10315 17343 -10281
rect 17343 -10315 17369 -10281
rect 17407 -10315 17411 -10281
rect 17411 -10315 17441 -10281
rect 17479 -10315 17513 -10281
rect 17551 -10315 17581 -10281
rect 17581 -10315 17585 -10281
rect 17623 -10315 17649 -10281
rect 17649 -10315 17657 -10281
rect 17695 -10315 17717 -10281
rect 17717 -10315 17729 -10281
rect 17767 -10315 17785 -10281
rect 17785 -10315 17801 -10281
rect 17839 -10315 17853 -10281
rect 17853 -10315 17873 -10281
rect 17911 -10315 17921 -10281
rect 17921 -10315 17945 -10281
rect 17983 -10315 17989 -10281
rect 17989 -10315 18017 -10281
rect 18055 -10315 18057 -10281
rect 18057 -10315 18089 -10281
rect 18127 -10315 18159 -10281
rect 18159 -10315 18161 -10281
rect 18199 -10315 18227 -10281
rect 18227 -10315 18233 -10281
rect 18271 -10315 18295 -10281
rect 18295 -10315 18305 -10281
rect 18343 -10315 18363 -10281
rect 18363 -10315 18377 -10281
rect 18415 -10315 18431 -10281
rect 18431 -10315 18449 -10281
rect 18487 -10315 18499 -10281
rect 18499 -10315 18521 -10281
rect 18559 -10315 18567 -10281
rect 18567 -10315 18593 -10281
rect 18631 -10315 18635 -10281
rect 18635 -10315 18665 -10281
rect 18703 -10315 18737 -10281
rect 18775 -10315 18805 -10281
rect 18805 -10315 18809 -10281
rect 18847 -10315 18873 -10281
rect 18873 -10315 18881 -10281
rect 18919 -10315 18941 -10281
rect 18941 -10315 18953 -10281
rect 18991 -10315 19009 -10281
rect 19009 -10315 19025 -10281
rect 19063 -10315 19077 -10281
rect 19077 -10315 19097 -10281
rect 19135 -10315 19145 -10281
rect 19145 -10315 19169 -10281
rect 19207 -10315 19213 -10281
rect 19213 -10315 19241 -10281
rect 19279 -10315 19281 -10281
rect 19281 -10315 19313 -10281
rect 19351 -10315 19383 -10281
rect 19383 -10315 19385 -10281
rect 19423 -10315 19451 -10281
rect 19451 -10315 19457 -10281
rect 19495 -10315 19519 -10281
rect 19519 -10315 19529 -10281
rect 19567 -10315 19587 -10281
rect 19587 -10315 19601 -10281
rect 19639 -10315 19655 -10281
rect 19655 -10315 19673 -10281
rect 19711 -10315 19723 -10281
rect 19723 -10315 19745 -10281
rect 19783 -10315 19791 -10281
rect 19791 -10315 19817 -10281
rect 19855 -10315 19859 -10281
rect 19859 -10315 19889 -10281
rect 19927 -10315 19961 -10281
rect 19999 -10315 20029 -10281
rect 20029 -10315 20033 -10281
rect 20071 -10315 20097 -10281
rect 20097 -10315 20105 -10281
rect 20143 -10315 20165 -10281
rect 20165 -10315 20177 -10281
rect 20215 -10315 20233 -10281
rect 20233 -10315 20249 -10281
rect 20287 -10315 20301 -10281
rect 20301 -10315 20321 -10281
rect 20359 -10315 20369 -10281
rect 20369 -10315 20393 -10281
rect 20431 -10315 20437 -10281
rect 20437 -10315 20465 -10281
rect 20503 -10315 20505 -10281
rect 20505 -10315 20537 -10281
rect 20575 -10315 20607 -10281
rect 20607 -10315 20609 -10281
rect 20647 -10315 20675 -10281
rect 20675 -10315 20681 -10281
rect 20719 -10315 20743 -10281
rect 20743 -10315 20753 -10281
rect 20791 -10315 20811 -10281
rect 20811 -10315 20825 -10281
rect 20863 -10315 20879 -10281
rect 20879 -10315 20897 -10281
rect 20935 -10315 20947 -10281
rect 20947 -10315 20969 -10281
rect 21007 -10315 21015 -10281
rect 21015 -10315 21041 -10281
rect 21079 -10315 21083 -10281
rect 21083 -10315 21113 -10281
rect 21151 -10315 21185 -10281
rect 21223 -10315 21253 -10281
rect 21253 -10315 21257 -10281
rect 21295 -10315 21321 -10281
rect 21321 -10315 21329 -10281
rect 21367 -10315 21389 -10281
rect 21389 -10315 21401 -10281
rect 21439 -10315 21457 -10281
rect 21457 -10315 21473 -10281
rect 21511 -10315 21525 -10281
rect 21525 -10315 21545 -10281
rect 21583 -10315 21593 -10281
rect 21593 -10315 21617 -10281
rect 21655 -10315 21661 -10281
rect 21661 -10315 21689 -10281
rect 21727 -10315 21729 -10281
rect 21729 -10315 21761 -10281
rect 21799 -10315 21831 -10281
rect 21831 -10315 21833 -10281
rect 21871 -10315 21899 -10281
rect 21899 -10315 21905 -10281
rect 21943 -10315 21967 -10281
rect 21967 -10315 21977 -10281
rect 22015 -10315 22035 -10281
rect 22035 -10315 22049 -10281
rect 22087 -10315 22103 -10281
rect 22103 -10315 22121 -10281
rect 22159 -10315 22171 -10281
rect 22171 -10315 22193 -10281
rect 22231 -10315 22239 -10281
rect 22239 -10315 22265 -10281
rect 22303 -10315 22307 -10281
rect 22307 -10315 22337 -10281
rect 22375 -10315 22409 -10281
rect 22447 -10315 22477 -10281
rect 22477 -10315 22481 -10281
rect 22519 -10315 22545 -10281
rect 22545 -10315 22553 -10281
rect 22591 -10315 22613 -10281
rect 22613 -10315 22625 -10281
rect 22663 -10315 22681 -10281
rect 22681 -10315 22697 -10281
rect 22735 -10315 22749 -10281
rect 22749 -10315 22769 -10281
rect 22807 -10315 22817 -10281
rect 22817 -10315 22841 -10281
rect 22879 -10315 22885 -10281
rect 22885 -10315 22913 -10281
rect 22951 -10315 22953 -10281
rect 22953 -10315 22985 -10281
rect 23023 -10315 23055 -10281
rect 23055 -10315 23057 -10281
rect 23095 -10315 23123 -10281
rect 23123 -10315 23129 -10281
rect 23167 -10315 23191 -10281
rect 23191 -10315 23201 -10281
rect 23239 -10315 23259 -10281
rect 23259 -10315 23273 -10281
rect 23311 -10315 23327 -10281
rect 23327 -10315 23345 -10281
rect 23383 -10315 23395 -10281
rect 23395 -10315 23417 -10281
rect 23455 -10315 23463 -10281
rect 23463 -10315 23489 -10281
rect 23527 -10315 23531 -10281
rect 23531 -10315 23561 -10281
rect 23599 -10315 23633 -10281
rect 23671 -10315 23701 -10281
rect 23701 -10315 23705 -10281
rect 23743 -10315 23769 -10281
rect 23769 -10315 23777 -10281
rect 23815 -10315 23837 -10281
rect 23837 -10315 23849 -10281
rect 23887 -10315 23905 -10281
rect 23905 -10315 23921 -10281
rect 23959 -10315 23973 -10281
rect 23973 -10315 23993 -10281
rect 24031 -10315 24041 -10281
rect 24041 -10315 24065 -10281
rect 24103 -10315 24109 -10281
rect 24109 -10315 24137 -10281
rect 24175 -10315 24177 -10281
rect 24177 -10315 24209 -10281
rect 24247 -10315 24279 -10281
rect 24279 -10315 24281 -10281
rect 24319 -10315 24347 -10281
rect 24347 -10315 24353 -10281
rect 24391 -10315 24415 -10281
rect 24415 -10315 24425 -10281
rect 24463 -10315 24483 -10281
rect 24483 -10315 24497 -10281
rect 24535 -10315 24551 -10281
rect 24551 -10315 24569 -10281
rect 24607 -10315 24619 -10281
rect 24619 -10315 24641 -10281
rect 24679 -10315 24713 -10281
rect -12221 -11245 -12187 -11211
rect -12149 -11245 -12145 -11211
rect -12145 -11245 -12115 -11211
rect -12077 -11245 -12043 -11211
rect -12005 -11245 -11975 -11211
rect -11975 -11245 -11971 -11211
rect -11933 -11245 -11907 -11211
rect -11907 -11245 -11899 -11211
rect -11861 -11245 -11839 -11211
rect -11839 -11245 -11827 -11211
rect -11789 -11245 -11771 -11211
rect -11771 -11245 -11755 -11211
rect -11717 -11245 -11703 -11211
rect -11703 -11245 -11683 -11211
rect -11645 -11245 -11635 -11211
rect -11635 -11245 -11611 -11211
rect -11573 -11245 -11567 -11211
rect -11567 -11245 -11539 -11211
rect -11501 -11245 -11499 -11211
rect -11499 -11245 -11467 -11211
rect -11429 -11245 -11397 -11211
rect -11397 -11245 -11395 -11211
rect -11357 -11245 -11329 -11211
rect -11329 -11245 -11323 -11211
rect -11285 -11245 -11261 -11211
rect -11261 -11245 -11251 -11211
rect -11213 -11245 -11193 -11211
rect -11193 -11245 -11179 -11211
rect -11141 -11245 -11125 -11211
rect -11125 -11245 -11107 -11211
rect -11069 -11245 -11057 -11211
rect -11057 -11245 -11035 -11211
rect -10997 -11245 -10989 -11211
rect -10989 -11245 -10963 -11211
rect -10925 -11245 -10921 -11211
rect -10921 -11245 -10891 -11211
rect -10853 -11245 -10819 -11211
rect -10781 -11245 -10751 -11211
rect -10751 -11245 -10747 -11211
rect -10709 -11245 -10683 -11211
rect -10683 -11245 -10675 -11211
rect -10637 -11245 -10615 -11211
rect -10615 -11245 -10603 -11211
rect -10565 -11245 -10547 -11211
rect -10547 -11245 -10531 -11211
rect -10493 -11245 -10479 -11211
rect -10479 -11245 -10459 -11211
rect -10421 -11245 -10411 -11211
rect -10411 -11245 -10387 -11211
rect -10349 -11245 -10343 -11211
rect -10343 -11245 -10315 -11211
rect -10277 -11245 -10275 -11211
rect -10275 -11245 -10243 -11211
rect -10205 -11245 -10173 -11211
rect -10173 -11245 -10171 -11211
rect -10133 -11245 -10105 -11211
rect -10105 -11245 -10099 -11211
rect -10061 -11245 -10037 -11211
rect -10037 -11245 -10027 -11211
rect -9989 -11245 -9969 -11211
rect -9969 -11245 -9955 -11211
rect -9917 -11245 -9901 -11211
rect -9901 -11245 -9883 -11211
rect -9845 -11245 -9833 -11211
rect -9833 -11245 -9811 -11211
rect -9773 -11245 -9765 -11211
rect -9765 -11245 -9739 -11211
rect -9701 -11245 -9697 -11211
rect -9697 -11245 -9667 -11211
rect -9629 -11245 -9595 -11211
rect -9557 -11245 -9527 -11211
rect -9527 -11245 -9523 -11211
rect -9485 -11245 -9459 -11211
rect -9459 -11245 -9451 -11211
rect -9413 -11245 -9391 -11211
rect -9391 -11245 -9379 -11211
rect -9341 -11245 -9323 -11211
rect -9323 -11245 -9307 -11211
rect -9269 -11245 -9255 -11211
rect -9255 -11245 -9235 -11211
rect -9197 -11245 -9187 -11211
rect -9187 -11245 -9163 -11211
rect -9125 -11245 -9119 -11211
rect -9119 -11245 -9091 -11211
rect -9053 -11245 -9051 -11211
rect -9051 -11245 -9019 -11211
rect -8981 -11245 -8949 -11211
rect -8949 -11245 -8947 -11211
rect -8909 -11245 -8881 -11211
rect -8881 -11245 -8875 -11211
rect -8837 -11245 -8813 -11211
rect -8813 -11245 -8803 -11211
rect -8765 -11245 -8745 -11211
rect -8745 -11245 -8731 -11211
rect -8693 -11245 -8677 -11211
rect -8677 -11245 -8659 -11211
rect -8621 -11245 -8609 -11211
rect -8609 -11245 -8587 -11211
rect -8549 -11245 -8541 -11211
rect -8541 -11245 -8515 -11211
rect -8477 -11245 -8473 -11211
rect -8473 -11245 -8443 -11211
rect -8405 -11245 -8371 -11211
rect -8333 -11245 -8303 -11211
rect -8303 -11245 -8299 -11211
rect -8261 -11245 -8235 -11211
rect -8235 -11245 -8227 -11211
rect -8189 -11245 -8167 -11211
rect -8167 -11245 -8155 -11211
rect -8117 -11245 -8099 -11211
rect -8099 -11245 -8083 -11211
rect -8045 -11245 -8031 -11211
rect -8031 -11245 -8011 -11211
rect -7973 -11245 -7963 -11211
rect -7963 -11245 -7939 -11211
rect -7901 -11245 -7895 -11211
rect -7895 -11245 -7867 -11211
rect -7829 -11245 -7827 -11211
rect -7827 -11245 -7795 -11211
rect -7757 -11245 -7725 -11211
rect -7725 -11245 -7723 -11211
rect -7685 -11245 -7657 -11211
rect -7657 -11245 -7651 -11211
rect -7613 -11245 -7589 -11211
rect -7589 -11245 -7579 -11211
rect -7541 -11245 -7521 -11211
rect -7521 -11245 -7507 -11211
rect -7469 -11245 -7453 -11211
rect -7453 -11245 -7435 -11211
rect -7397 -11245 -7385 -11211
rect -7385 -11245 -7363 -11211
rect -7325 -11245 -7317 -11211
rect -7317 -11245 -7291 -11211
rect -7253 -11245 -7249 -11211
rect -7249 -11245 -7219 -11211
rect -7181 -11245 -7147 -11211
rect -7109 -11245 -7079 -11211
rect -7079 -11245 -7075 -11211
rect -7037 -11245 -7011 -11211
rect -7011 -11245 -7003 -11211
rect -6965 -11245 -6943 -11211
rect -6943 -11245 -6931 -11211
rect -6893 -11245 -6875 -11211
rect -6875 -11245 -6859 -11211
rect -6821 -11245 -6807 -11211
rect -6807 -11245 -6787 -11211
rect -6749 -11245 -6739 -11211
rect -6739 -11245 -6715 -11211
rect -6677 -11245 -6671 -11211
rect -6671 -11245 -6643 -11211
rect -6605 -11245 -6603 -11211
rect -6603 -11245 -6571 -11211
rect -6533 -11245 -6501 -11211
rect -6501 -11245 -6499 -11211
rect -6461 -11245 -6433 -11211
rect -6433 -11245 -6427 -11211
rect -6389 -11245 -6365 -11211
rect -6365 -11245 -6355 -11211
rect -6317 -11245 -6297 -11211
rect -6297 -11245 -6283 -11211
rect -6245 -11245 -6229 -11211
rect -6229 -11245 -6211 -11211
rect -6173 -11245 -6161 -11211
rect -6161 -11245 -6139 -11211
rect -6101 -11245 -6093 -11211
rect -6093 -11245 -6067 -11211
rect -6029 -11245 -6025 -11211
rect -6025 -11245 -5995 -11211
rect -5957 -11245 -5923 -11211
rect -5885 -11245 -5855 -11211
rect -5855 -11245 -5851 -11211
rect -5813 -11245 -5787 -11211
rect -5787 -11245 -5779 -11211
rect -5741 -11245 -5719 -11211
rect -5719 -11245 -5707 -11211
rect -5669 -11245 -5651 -11211
rect -5651 -11245 -5635 -11211
rect -5597 -11245 -5583 -11211
rect -5583 -11245 -5563 -11211
rect -5525 -11245 -5515 -11211
rect -5515 -11245 -5491 -11211
rect -5453 -11245 -5447 -11211
rect -5447 -11245 -5419 -11211
rect -5381 -11245 -5379 -11211
rect -5379 -11245 -5347 -11211
rect -5309 -11245 -5277 -11211
rect -5277 -11245 -5275 -11211
rect -5237 -11245 -5209 -11211
rect -5209 -11245 -5203 -11211
rect -5165 -11245 -5141 -11211
rect -5141 -11245 -5131 -11211
rect -5093 -11245 -5073 -11211
rect -5073 -11245 -5059 -11211
rect -5021 -11245 -5005 -11211
rect -5005 -11245 -4987 -11211
rect -4949 -11245 -4937 -11211
rect -4937 -11245 -4915 -11211
rect -4877 -11245 -4869 -11211
rect -4869 -11245 -4843 -11211
rect -4805 -11245 -4801 -11211
rect -4801 -11245 -4771 -11211
rect -4733 -11245 -4699 -11211
rect -4661 -11245 -4631 -11211
rect -4631 -11245 -4627 -11211
rect -4589 -11245 -4563 -11211
rect -4563 -11245 -4555 -11211
rect -4517 -11245 -4495 -11211
rect -4495 -11245 -4483 -11211
rect -4445 -11245 -4427 -11211
rect -4427 -11245 -4411 -11211
rect -4373 -11245 -4359 -11211
rect -4359 -11245 -4339 -11211
rect -4301 -11245 -4291 -11211
rect -4291 -11245 -4267 -11211
rect -4229 -11245 -4223 -11211
rect -4223 -11245 -4195 -11211
rect -4157 -11245 -4155 -11211
rect -4155 -11245 -4123 -11211
rect -4085 -11245 -4053 -11211
rect -4053 -11245 -4051 -11211
rect -4013 -11245 -3985 -11211
rect -3985 -11245 -3979 -11211
rect -3941 -11245 -3917 -11211
rect -3917 -11245 -3907 -11211
rect -3869 -11245 -3849 -11211
rect -3849 -11245 -3835 -11211
rect -3797 -11245 -3781 -11211
rect -3781 -11245 -3763 -11211
rect -3725 -11245 -3713 -11211
rect -3713 -11245 -3691 -11211
rect -3653 -11245 -3645 -11211
rect -3645 -11245 -3619 -11211
rect -3581 -11245 -3577 -11211
rect -3577 -11245 -3547 -11211
rect -3509 -11245 -3475 -11211
rect -3437 -11245 -3407 -11211
rect -3407 -11245 -3403 -11211
rect -3365 -11245 -3339 -11211
rect -3339 -11245 -3331 -11211
rect -3293 -11245 -3271 -11211
rect -3271 -11245 -3259 -11211
rect -3221 -11245 -3203 -11211
rect -3203 -11245 -3187 -11211
rect -3149 -11245 -3135 -11211
rect -3135 -11245 -3115 -11211
rect -3077 -11245 -3067 -11211
rect -3067 -11245 -3043 -11211
rect -3005 -11245 -2999 -11211
rect -2999 -11245 -2971 -11211
rect -2933 -11245 -2931 -11211
rect -2931 -11245 -2899 -11211
rect -2861 -11245 -2829 -11211
rect -2829 -11245 -2827 -11211
rect -2789 -11245 -2761 -11211
rect -2761 -11245 -2755 -11211
rect -2717 -11245 -2693 -11211
rect -2693 -11245 -2683 -11211
rect -2645 -11245 -2625 -11211
rect -2625 -11245 -2611 -11211
rect -2573 -11245 -2557 -11211
rect -2557 -11245 -2539 -11211
rect -2501 -11245 -2489 -11211
rect -2489 -11245 -2467 -11211
rect -2429 -11245 -2421 -11211
rect -2421 -11245 -2395 -11211
rect -2357 -11245 -2353 -11211
rect -2353 -11245 -2323 -11211
rect -2285 -11245 -2251 -11211
rect -2213 -11245 -2183 -11211
rect -2183 -11245 -2179 -11211
rect -2141 -11245 -2115 -11211
rect -2115 -11245 -2107 -11211
rect -2069 -11245 -2047 -11211
rect -2047 -11245 -2035 -11211
rect -1997 -11245 -1979 -11211
rect -1979 -11245 -1963 -11211
rect -1925 -11245 -1911 -11211
rect -1911 -11245 -1891 -11211
rect -1853 -11245 -1843 -11211
rect -1843 -11245 -1819 -11211
rect -1781 -11245 -1775 -11211
rect -1775 -11245 -1747 -11211
rect -1709 -11245 -1707 -11211
rect -1707 -11245 -1675 -11211
rect -1637 -11245 -1605 -11211
rect -1605 -11245 -1603 -11211
rect -1565 -11245 -1537 -11211
rect -1537 -11245 -1531 -11211
rect -1493 -11245 -1469 -11211
rect -1469 -11245 -1459 -11211
rect -1421 -11245 -1401 -11211
rect -1401 -11245 -1387 -11211
rect -1349 -11245 -1333 -11211
rect -1333 -11245 -1315 -11211
rect -1277 -11245 -1265 -11211
rect -1265 -11245 -1243 -11211
rect -1205 -11245 -1197 -11211
rect -1197 -11245 -1171 -11211
rect -1133 -11245 -1129 -11211
rect -1129 -11245 -1099 -11211
rect -1061 -11245 -1027 -11211
rect -989 -11245 -959 -11211
rect -959 -11245 -955 -11211
rect -917 -11245 -891 -11211
rect -891 -11245 -883 -11211
rect -845 -11245 -823 -11211
rect -823 -11245 -811 -11211
rect -773 -11245 -755 -11211
rect -755 -11245 -739 -11211
rect -701 -11245 -687 -11211
rect -687 -11245 -667 -11211
rect -629 -11245 -619 -11211
rect -619 -11245 -595 -11211
rect -557 -11245 -551 -11211
rect -551 -11245 -523 -11211
rect -485 -11245 -483 -11211
rect -483 -11245 -451 -11211
rect -413 -11245 -381 -11211
rect -381 -11245 -379 -11211
rect -341 -11245 -313 -11211
rect -313 -11245 -307 -11211
rect -269 -11245 -245 -11211
rect -245 -11245 -235 -11211
rect -197 -11245 -177 -11211
rect -177 -11245 -163 -11211
rect -125 -11245 -109 -11211
rect -109 -11245 -91 -11211
rect -53 -11245 -41 -11211
rect -41 -11245 -19 -11211
rect 19 -11245 27 -11211
rect 27 -11245 53 -11211
rect 91 -11245 95 -11211
rect 95 -11245 125 -11211
rect 163 -11245 197 -11211
rect 235 -11245 265 -11211
rect 265 -11245 269 -11211
rect 307 -11245 333 -11211
rect 333 -11245 341 -11211
rect 379 -11245 401 -11211
rect 401 -11245 413 -11211
rect 451 -11245 469 -11211
rect 469 -11245 485 -11211
rect 523 -11245 537 -11211
rect 537 -11245 557 -11211
rect 595 -11245 605 -11211
rect 605 -11245 629 -11211
rect 667 -11245 673 -11211
rect 673 -11245 701 -11211
rect 739 -11245 741 -11211
rect 741 -11245 773 -11211
rect 811 -11245 843 -11211
rect 843 -11245 845 -11211
rect 883 -11245 911 -11211
rect 911 -11245 917 -11211
rect 955 -11245 979 -11211
rect 979 -11245 989 -11211
rect 1027 -11245 1047 -11211
rect 1047 -11245 1061 -11211
rect 1099 -11245 1115 -11211
rect 1115 -11245 1133 -11211
rect 1171 -11245 1183 -11211
rect 1183 -11245 1205 -11211
rect 1243 -11245 1251 -11211
rect 1251 -11245 1277 -11211
rect 1315 -11245 1319 -11211
rect 1319 -11245 1349 -11211
rect 1387 -11245 1421 -11211
rect 1459 -11245 1489 -11211
rect 1489 -11245 1493 -11211
rect 1531 -11245 1557 -11211
rect 1557 -11245 1565 -11211
rect 1603 -11245 1625 -11211
rect 1625 -11245 1637 -11211
rect 1675 -11245 1693 -11211
rect 1693 -11245 1709 -11211
rect 1747 -11245 1761 -11211
rect 1761 -11245 1781 -11211
rect 1819 -11245 1829 -11211
rect 1829 -11245 1853 -11211
rect 1891 -11245 1897 -11211
rect 1897 -11245 1925 -11211
rect 1963 -11245 1965 -11211
rect 1965 -11245 1997 -11211
rect 2035 -11245 2067 -11211
rect 2067 -11245 2069 -11211
rect 2107 -11245 2135 -11211
rect 2135 -11245 2141 -11211
rect 2179 -11245 2203 -11211
rect 2203 -11245 2213 -11211
rect 2251 -11245 2271 -11211
rect 2271 -11245 2285 -11211
rect 2323 -11245 2339 -11211
rect 2339 -11245 2357 -11211
rect 2395 -11245 2407 -11211
rect 2407 -11245 2429 -11211
rect 2467 -11245 2475 -11211
rect 2475 -11245 2501 -11211
rect 2539 -11245 2543 -11211
rect 2543 -11245 2573 -11211
rect 2611 -11245 2645 -11211
rect 2683 -11245 2713 -11211
rect 2713 -11245 2717 -11211
rect 2755 -11245 2781 -11211
rect 2781 -11245 2789 -11211
rect 2827 -11245 2849 -11211
rect 2849 -11245 2861 -11211
rect 2899 -11245 2917 -11211
rect 2917 -11245 2933 -11211
rect 2971 -11245 2985 -11211
rect 2985 -11245 3005 -11211
rect 3043 -11245 3053 -11211
rect 3053 -11245 3077 -11211
rect 3115 -11245 3121 -11211
rect 3121 -11245 3149 -11211
rect 3187 -11245 3189 -11211
rect 3189 -11245 3221 -11211
rect 3259 -11245 3291 -11211
rect 3291 -11245 3293 -11211
rect 3331 -11245 3359 -11211
rect 3359 -11245 3365 -11211
rect 3403 -11245 3427 -11211
rect 3427 -11245 3437 -11211
rect 3475 -11245 3495 -11211
rect 3495 -11245 3509 -11211
rect 3547 -11245 3563 -11211
rect 3563 -11245 3581 -11211
rect 3619 -11245 3631 -11211
rect 3631 -11245 3653 -11211
rect 3691 -11245 3699 -11211
rect 3699 -11245 3725 -11211
rect 3763 -11245 3767 -11211
rect 3767 -11245 3797 -11211
rect 3835 -11245 3869 -11211
rect 3907 -11245 3937 -11211
rect 3937 -11245 3941 -11211
rect 3979 -11245 4005 -11211
rect 4005 -11245 4013 -11211
rect 4051 -11245 4073 -11211
rect 4073 -11245 4085 -11211
rect 4123 -11245 4141 -11211
rect 4141 -11245 4157 -11211
rect 4195 -11245 4209 -11211
rect 4209 -11245 4229 -11211
rect 4267 -11245 4277 -11211
rect 4277 -11245 4301 -11211
rect 4339 -11245 4345 -11211
rect 4345 -11245 4373 -11211
rect 4411 -11245 4413 -11211
rect 4413 -11245 4445 -11211
rect 4483 -11245 4515 -11211
rect 4515 -11245 4517 -11211
rect 4555 -11245 4583 -11211
rect 4583 -11245 4589 -11211
rect 4627 -11245 4651 -11211
rect 4651 -11245 4661 -11211
rect 4699 -11245 4719 -11211
rect 4719 -11245 4733 -11211
rect 4771 -11245 4787 -11211
rect 4787 -11245 4805 -11211
rect 4843 -11245 4855 -11211
rect 4855 -11245 4877 -11211
rect 4915 -11245 4923 -11211
rect 4923 -11245 4949 -11211
rect 4987 -11245 4991 -11211
rect 4991 -11245 5021 -11211
rect 5059 -11245 5093 -11211
rect 5131 -11245 5161 -11211
rect 5161 -11245 5165 -11211
rect 5203 -11245 5229 -11211
rect 5229 -11245 5237 -11211
rect 5275 -11245 5297 -11211
rect 5297 -11245 5309 -11211
rect 5347 -11245 5365 -11211
rect 5365 -11245 5381 -11211
rect 5419 -11245 5433 -11211
rect 5433 -11245 5453 -11211
rect 5491 -11245 5501 -11211
rect 5501 -11245 5525 -11211
rect 5563 -11245 5569 -11211
rect 5569 -11245 5597 -11211
rect 5635 -11245 5637 -11211
rect 5637 -11245 5669 -11211
rect 5707 -11245 5739 -11211
rect 5739 -11245 5741 -11211
rect 5779 -11245 5807 -11211
rect 5807 -11245 5813 -11211
rect 5851 -11245 5875 -11211
rect 5875 -11245 5885 -11211
rect 5923 -11245 5943 -11211
rect 5943 -11245 5957 -11211
rect 5995 -11245 6011 -11211
rect 6011 -11245 6029 -11211
rect 6067 -11245 6079 -11211
rect 6079 -11245 6101 -11211
rect 6139 -11245 6147 -11211
rect 6147 -11245 6173 -11211
rect 6211 -11245 6215 -11211
rect 6215 -11245 6245 -11211
rect 6283 -11245 6317 -11211
rect 6355 -11245 6385 -11211
rect 6385 -11245 6389 -11211
rect 6427 -11245 6453 -11211
rect 6453 -11245 6461 -11211
rect 6499 -11245 6521 -11211
rect 6521 -11245 6533 -11211
rect 6571 -11245 6589 -11211
rect 6589 -11245 6605 -11211
rect 6643 -11245 6657 -11211
rect 6657 -11245 6677 -11211
rect 6715 -11245 6725 -11211
rect 6725 -11245 6749 -11211
rect 6787 -11245 6793 -11211
rect 6793 -11245 6821 -11211
rect 6859 -11245 6861 -11211
rect 6861 -11245 6893 -11211
rect 6931 -11245 6963 -11211
rect 6963 -11245 6965 -11211
rect 7003 -11245 7031 -11211
rect 7031 -11245 7037 -11211
rect 7075 -11245 7099 -11211
rect 7099 -11245 7109 -11211
rect 7147 -11245 7167 -11211
rect 7167 -11245 7181 -11211
rect 7219 -11245 7235 -11211
rect 7235 -11245 7253 -11211
rect 7291 -11245 7303 -11211
rect 7303 -11245 7325 -11211
rect 7363 -11245 7371 -11211
rect 7371 -11245 7397 -11211
rect 7435 -11245 7439 -11211
rect 7439 -11245 7469 -11211
rect 7507 -11245 7541 -11211
rect 7579 -11245 7609 -11211
rect 7609 -11245 7613 -11211
rect 7651 -11245 7677 -11211
rect 7677 -11245 7685 -11211
rect 7723 -11245 7745 -11211
rect 7745 -11245 7757 -11211
rect 7795 -11245 7813 -11211
rect 7813 -11245 7829 -11211
rect 7867 -11245 7881 -11211
rect 7881 -11245 7901 -11211
rect 7939 -11245 7949 -11211
rect 7949 -11245 7973 -11211
rect 8011 -11245 8017 -11211
rect 8017 -11245 8045 -11211
rect 8083 -11245 8085 -11211
rect 8085 -11245 8117 -11211
rect 8155 -11245 8187 -11211
rect 8187 -11245 8189 -11211
rect 8227 -11245 8255 -11211
rect 8255 -11245 8261 -11211
rect 8299 -11245 8323 -11211
rect 8323 -11245 8333 -11211
rect 8371 -11245 8391 -11211
rect 8391 -11245 8405 -11211
rect 8443 -11245 8459 -11211
rect 8459 -11245 8477 -11211
rect 8515 -11245 8527 -11211
rect 8527 -11245 8549 -11211
rect 8587 -11245 8595 -11211
rect 8595 -11245 8621 -11211
rect 8659 -11245 8663 -11211
rect 8663 -11245 8693 -11211
rect 8731 -11245 8765 -11211
rect 8803 -11245 8833 -11211
rect 8833 -11245 8837 -11211
rect 8875 -11245 8901 -11211
rect 8901 -11245 8909 -11211
rect 8947 -11245 8969 -11211
rect 8969 -11245 8981 -11211
rect 9019 -11245 9037 -11211
rect 9037 -11245 9053 -11211
rect 9091 -11245 9105 -11211
rect 9105 -11245 9125 -11211
rect 9163 -11245 9173 -11211
rect 9173 -11245 9197 -11211
rect 9235 -11245 9241 -11211
rect 9241 -11245 9269 -11211
rect 9307 -11245 9309 -11211
rect 9309 -11245 9341 -11211
rect 9379 -11245 9411 -11211
rect 9411 -11245 9413 -11211
rect 9451 -11245 9479 -11211
rect 9479 -11245 9485 -11211
rect 9523 -11245 9547 -11211
rect 9547 -11245 9557 -11211
rect 9595 -11245 9615 -11211
rect 9615 -11245 9629 -11211
rect 9667 -11245 9683 -11211
rect 9683 -11245 9701 -11211
rect 9739 -11245 9751 -11211
rect 9751 -11245 9773 -11211
rect 9811 -11245 9819 -11211
rect 9819 -11245 9845 -11211
rect 9883 -11245 9887 -11211
rect 9887 -11245 9917 -11211
rect 9955 -11245 9989 -11211
rect 10027 -11245 10057 -11211
rect 10057 -11245 10061 -11211
rect 10099 -11245 10125 -11211
rect 10125 -11245 10133 -11211
rect 10171 -11245 10193 -11211
rect 10193 -11245 10205 -11211
rect 10243 -11245 10261 -11211
rect 10261 -11245 10277 -11211
rect 10315 -11245 10329 -11211
rect 10329 -11245 10349 -11211
rect 10387 -11245 10397 -11211
rect 10397 -11245 10421 -11211
rect 10459 -11245 10465 -11211
rect 10465 -11245 10493 -11211
rect 10531 -11245 10533 -11211
rect 10533 -11245 10565 -11211
rect 10603 -11245 10635 -11211
rect 10635 -11245 10637 -11211
rect 10675 -11245 10703 -11211
rect 10703 -11245 10709 -11211
rect 10747 -11245 10771 -11211
rect 10771 -11245 10781 -11211
rect 10819 -11245 10839 -11211
rect 10839 -11245 10853 -11211
rect 10891 -11245 10907 -11211
rect 10907 -11245 10925 -11211
rect 10963 -11245 10975 -11211
rect 10975 -11245 10997 -11211
rect 11035 -11245 11043 -11211
rect 11043 -11245 11069 -11211
rect 11107 -11245 11111 -11211
rect 11111 -11245 11141 -11211
rect 11179 -11245 11213 -11211
rect 11251 -11245 11281 -11211
rect 11281 -11245 11285 -11211
rect 11323 -11245 11349 -11211
rect 11349 -11245 11357 -11211
rect 11395 -11245 11417 -11211
rect 11417 -11245 11429 -11211
rect 11467 -11245 11485 -11211
rect 11485 -11245 11501 -11211
rect 11539 -11245 11553 -11211
rect 11553 -11245 11573 -11211
rect 11611 -11245 11621 -11211
rect 11621 -11245 11645 -11211
rect 11683 -11245 11689 -11211
rect 11689 -11245 11717 -11211
rect 11755 -11245 11757 -11211
rect 11757 -11245 11789 -11211
rect 11827 -11245 11859 -11211
rect 11859 -11245 11861 -11211
rect 11899 -11245 11927 -11211
rect 11927 -11245 11933 -11211
rect 11971 -11245 11995 -11211
rect 11995 -11245 12005 -11211
rect 12043 -11245 12063 -11211
rect 12063 -11245 12077 -11211
rect 12115 -11245 12131 -11211
rect 12131 -11245 12149 -11211
rect 12187 -11245 12199 -11211
rect 12199 -11245 12221 -11211
rect 12259 -11245 12267 -11211
rect 12267 -11245 12293 -11211
rect 12331 -11245 12335 -11211
rect 12335 -11245 12365 -11211
rect 12403 -11245 12437 -11211
rect 12475 -11245 12505 -11211
rect 12505 -11245 12509 -11211
rect 12547 -11245 12573 -11211
rect 12573 -11245 12581 -11211
rect 12619 -11245 12641 -11211
rect 12641 -11245 12653 -11211
rect 12691 -11245 12709 -11211
rect 12709 -11245 12725 -11211
rect 12763 -11245 12777 -11211
rect 12777 -11245 12797 -11211
rect 12835 -11245 12845 -11211
rect 12845 -11245 12869 -11211
rect 12907 -11245 12913 -11211
rect 12913 -11245 12941 -11211
rect 12979 -11245 12981 -11211
rect 12981 -11245 13013 -11211
rect 13051 -11245 13083 -11211
rect 13083 -11245 13085 -11211
rect 13123 -11245 13151 -11211
rect 13151 -11245 13157 -11211
rect 13195 -11245 13219 -11211
rect 13219 -11245 13229 -11211
rect 13267 -11245 13287 -11211
rect 13287 -11245 13301 -11211
rect 13339 -11245 13355 -11211
rect 13355 -11245 13373 -11211
rect 13411 -11245 13423 -11211
rect 13423 -11245 13445 -11211
rect 13483 -11245 13491 -11211
rect 13491 -11245 13517 -11211
rect 13555 -11245 13559 -11211
rect 13559 -11245 13589 -11211
rect 13627 -11245 13661 -11211
rect 13699 -11245 13729 -11211
rect 13729 -11245 13733 -11211
rect 13771 -11245 13797 -11211
rect 13797 -11245 13805 -11211
rect 13843 -11245 13865 -11211
rect 13865 -11245 13877 -11211
rect 13915 -11245 13933 -11211
rect 13933 -11245 13949 -11211
rect 13987 -11245 14001 -11211
rect 14001 -11245 14021 -11211
rect 14059 -11245 14069 -11211
rect 14069 -11245 14093 -11211
rect 14131 -11245 14137 -11211
rect 14137 -11245 14165 -11211
rect 14203 -11245 14205 -11211
rect 14205 -11245 14237 -11211
rect 14275 -11245 14307 -11211
rect 14307 -11245 14309 -11211
rect 14347 -11245 14375 -11211
rect 14375 -11245 14381 -11211
rect 14419 -11245 14443 -11211
rect 14443 -11245 14453 -11211
rect 14491 -11245 14511 -11211
rect 14511 -11245 14525 -11211
rect 14563 -11245 14579 -11211
rect 14579 -11245 14597 -11211
rect 14635 -11245 14647 -11211
rect 14647 -11245 14669 -11211
rect 14707 -11245 14715 -11211
rect 14715 -11245 14741 -11211
rect 14779 -11245 14783 -11211
rect 14783 -11245 14813 -11211
rect 14851 -11245 14885 -11211
rect 14923 -11245 14953 -11211
rect 14953 -11245 14957 -11211
rect 14995 -11245 15021 -11211
rect 15021 -11245 15029 -11211
rect 15067 -11245 15089 -11211
rect 15089 -11245 15101 -11211
rect 15139 -11245 15157 -11211
rect 15157 -11245 15173 -11211
rect 15211 -11245 15225 -11211
rect 15225 -11245 15245 -11211
rect 15283 -11245 15293 -11211
rect 15293 -11245 15317 -11211
rect 15355 -11245 15361 -11211
rect 15361 -11245 15389 -11211
rect 15427 -11245 15429 -11211
rect 15429 -11245 15461 -11211
rect 15499 -11245 15531 -11211
rect 15531 -11245 15533 -11211
rect 15571 -11245 15599 -11211
rect 15599 -11245 15605 -11211
rect 15643 -11245 15667 -11211
rect 15667 -11245 15677 -11211
rect 15715 -11245 15735 -11211
rect 15735 -11245 15749 -11211
rect 15787 -11245 15803 -11211
rect 15803 -11245 15821 -11211
rect 15859 -11245 15871 -11211
rect 15871 -11245 15893 -11211
rect 15931 -11245 15939 -11211
rect 15939 -11245 15965 -11211
rect 16003 -11245 16007 -11211
rect 16007 -11245 16037 -11211
rect 16075 -11245 16109 -11211
rect 16147 -11245 16177 -11211
rect 16177 -11245 16181 -11211
rect 16219 -11245 16245 -11211
rect 16245 -11245 16253 -11211
rect 16291 -11245 16313 -11211
rect 16313 -11245 16325 -11211
rect 16363 -11245 16381 -11211
rect 16381 -11245 16397 -11211
rect 16435 -11245 16449 -11211
rect 16449 -11245 16469 -11211
rect 16507 -11245 16517 -11211
rect 16517 -11245 16541 -11211
rect 16579 -11245 16585 -11211
rect 16585 -11245 16613 -11211
rect 16651 -11245 16653 -11211
rect 16653 -11245 16685 -11211
rect 16723 -11245 16755 -11211
rect 16755 -11245 16757 -11211
rect 16795 -11245 16823 -11211
rect 16823 -11245 16829 -11211
rect 16867 -11245 16891 -11211
rect 16891 -11245 16901 -11211
rect 16939 -11245 16959 -11211
rect 16959 -11245 16973 -11211
rect 17011 -11245 17027 -11211
rect 17027 -11245 17045 -11211
rect 17083 -11245 17095 -11211
rect 17095 -11245 17117 -11211
rect 17155 -11245 17163 -11211
rect 17163 -11245 17189 -11211
rect 17227 -11245 17231 -11211
rect 17231 -11245 17261 -11211
rect 17299 -11245 17333 -11211
rect 17371 -11245 17401 -11211
rect 17401 -11245 17405 -11211
rect 17443 -11245 17469 -11211
rect 17469 -11245 17477 -11211
rect 17515 -11245 17537 -11211
rect 17537 -11245 17549 -11211
rect 17587 -11245 17605 -11211
rect 17605 -11245 17621 -11211
rect 17659 -11245 17673 -11211
rect 17673 -11245 17693 -11211
rect 17731 -11245 17741 -11211
rect 17741 -11245 17765 -11211
rect 17803 -11245 17809 -11211
rect 17809 -11245 17837 -11211
rect 17875 -11245 17877 -11211
rect 17877 -11245 17909 -11211
rect 17947 -11245 17979 -11211
rect 17979 -11245 17981 -11211
rect 18019 -11245 18047 -11211
rect 18047 -11245 18053 -11211
rect 18091 -11245 18115 -11211
rect 18115 -11245 18125 -11211
rect 18163 -11245 18183 -11211
rect 18183 -11245 18197 -11211
rect 18235 -11245 18251 -11211
rect 18251 -11245 18269 -11211
rect 18307 -11245 18319 -11211
rect 18319 -11245 18341 -11211
rect 18379 -11245 18387 -11211
rect 18387 -11245 18413 -11211
rect 18451 -11245 18455 -11211
rect 18455 -11245 18485 -11211
rect 18523 -11245 18557 -11211
rect 18595 -11245 18625 -11211
rect 18625 -11245 18629 -11211
rect 18667 -11245 18693 -11211
rect 18693 -11245 18701 -11211
rect 18739 -11245 18761 -11211
rect 18761 -11245 18773 -11211
rect 18811 -11245 18829 -11211
rect 18829 -11245 18845 -11211
rect 18883 -11245 18897 -11211
rect 18897 -11245 18917 -11211
rect 18955 -11245 18965 -11211
rect 18965 -11245 18989 -11211
rect 19027 -11245 19033 -11211
rect 19033 -11245 19061 -11211
rect 19099 -11245 19101 -11211
rect 19101 -11245 19133 -11211
rect 19171 -11245 19203 -11211
rect 19203 -11245 19205 -11211
rect 19243 -11245 19271 -11211
rect 19271 -11245 19277 -11211
rect 19315 -11245 19339 -11211
rect 19339 -11245 19349 -11211
rect 19387 -11245 19407 -11211
rect 19407 -11245 19421 -11211
rect 19459 -11245 19475 -11211
rect 19475 -11245 19493 -11211
rect 19531 -11245 19543 -11211
rect 19543 -11245 19565 -11211
rect 19603 -11245 19611 -11211
rect 19611 -11245 19637 -11211
rect 19675 -11245 19679 -11211
rect 19679 -11245 19709 -11211
rect 19747 -11245 19781 -11211
rect 19819 -11245 19849 -11211
rect 19849 -11245 19853 -11211
rect 19891 -11245 19917 -11211
rect 19917 -11245 19925 -11211
rect 19963 -11245 19985 -11211
rect 19985 -11245 19997 -11211
rect 20035 -11245 20053 -11211
rect 20053 -11245 20069 -11211
rect 20107 -11245 20121 -11211
rect 20121 -11245 20141 -11211
rect 20179 -11245 20189 -11211
rect 20189 -11245 20213 -11211
rect 20251 -11245 20257 -11211
rect 20257 -11245 20285 -11211
rect 20323 -11245 20325 -11211
rect 20325 -11245 20357 -11211
rect 20395 -11245 20427 -11211
rect 20427 -11245 20429 -11211
rect 20467 -11245 20495 -11211
rect 20495 -11245 20501 -11211
rect 20539 -11245 20563 -11211
rect 20563 -11245 20573 -11211
rect 20611 -11245 20631 -11211
rect 20631 -11245 20645 -11211
rect 20683 -11245 20699 -11211
rect 20699 -11245 20717 -11211
rect 20755 -11245 20767 -11211
rect 20767 -11245 20789 -11211
rect 20827 -11245 20835 -11211
rect 20835 -11245 20861 -11211
rect 20899 -11245 20903 -11211
rect 20903 -11245 20933 -11211
rect 20971 -11245 21005 -11211
rect 21043 -11245 21073 -11211
rect 21073 -11245 21077 -11211
rect 21115 -11245 21141 -11211
rect 21141 -11245 21149 -11211
rect 21187 -11245 21209 -11211
rect 21209 -11245 21221 -11211
rect 21259 -11245 21277 -11211
rect 21277 -11245 21293 -11211
rect 21331 -11245 21345 -11211
rect 21345 -11245 21365 -11211
rect 21403 -11245 21413 -11211
rect 21413 -11245 21437 -11211
rect 21475 -11245 21481 -11211
rect 21481 -11245 21509 -11211
rect 21547 -11245 21549 -11211
rect 21549 -11245 21581 -11211
rect 21619 -11245 21651 -11211
rect 21651 -11245 21653 -11211
rect 21691 -11245 21719 -11211
rect 21719 -11245 21725 -11211
rect 21763 -11245 21787 -11211
rect 21787 -11245 21797 -11211
rect 21835 -11245 21855 -11211
rect 21855 -11245 21869 -11211
rect 21907 -11245 21923 -11211
rect 21923 -11245 21941 -11211
rect 21979 -11245 21991 -11211
rect 21991 -11245 22013 -11211
rect 22051 -11245 22059 -11211
rect 22059 -11245 22085 -11211
rect 22123 -11245 22127 -11211
rect 22127 -11245 22157 -11211
rect 22195 -11245 22229 -11211
rect 22267 -11245 22297 -11211
rect 22297 -11245 22301 -11211
rect 22339 -11245 22365 -11211
rect 22365 -11245 22373 -11211
rect 22411 -11245 22433 -11211
rect 22433 -11245 22445 -11211
rect 22483 -11245 22501 -11211
rect 22501 -11245 22517 -11211
rect 22555 -11245 22569 -11211
rect 22569 -11245 22589 -11211
rect 22627 -11245 22637 -11211
rect 22637 -11245 22661 -11211
rect 22699 -11245 22705 -11211
rect 22705 -11245 22733 -11211
rect 22771 -11245 22773 -11211
rect 22773 -11245 22805 -11211
rect 22843 -11245 22875 -11211
rect 22875 -11245 22877 -11211
rect 22915 -11245 22943 -11211
rect 22943 -11245 22949 -11211
rect 22987 -11245 23011 -11211
rect 23011 -11245 23021 -11211
rect 23059 -11245 23079 -11211
rect 23079 -11245 23093 -11211
rect 23131 -11245 23147 -11211
rect 23147 -11245 23165 -11211
rect 23203 -11245 23215 -11211
rect 23215 -11245 23237 -11211
rect 23275 -11245 23283 -11211
rect 23283 -11245 23309 -11211
rect 23347 -11245 23351 -11211
rect 23351 -11245 23381 -11211
rect 23419 -11245 23453 -11211
rect 23491 -11245 23521 -11211
rect 23521 -11245 23525 -11211
rect 23563 -11245 23589 -11211
rect 23589 -11245 23597 -11211
rect 23635 -11245 23657 -11211
rect 23657 -11245 23669 -11211
rect 23707 -11245 23725 -11211
rect 23725 -11245 23741 -11211
rect 23779 -11245 23793 -11211
rect 23793 -11245 23813 -11211
rect 23851 -11245 23861 -11211
rect 23861 -11245 23885 -11211
rect 23923 -11245 23929 -11211
rect 23929 -11245 23957 -11211
rect 23995 -11245 23997 -11211
rect 23997 -11245 24029 -11211
rect 24067 -11245 24099 -11211
rect 24099 -11245 24101 -11211
rect 24139 -11245 24167 -11211
rect 24167 -11245 24173 -11211
rect 24211 -11245 24235 -11211
rect 24235 -11245 24245 -11211
rect 24283 -11245 24303 -11211
rect 24303 -11245 24317 -11211
rect 24355 -11245 24371 -11211
rect 24371 -11245 24389 -11211
rect 24427 -11245 24439 -11211
rect 24439 -11245 24461 -11211
rect 24499 -11245 24507 -11211
rect 24507 -11245 24533 -11211
rect 24571 -11245 24575 -11211
rect 24575 -11245 24605 -11211
rect 24643 -11245 24677 -11211
rect 24715 -11245 24745 -11211
rect 24745 -11245 24749 -11211
rect 24787 -11245 24821 -11211
rect -12289 -12111 -12255 -12091
rect -12289 -12125 -12255 -12111
rect -12289 -12179 -12255 -12163
rect -12289 -12197 -12255 -12179
rect -12289 -12247 -12255 -12235
rect -12289 -12269 -12255 -12247
rect -12289 -12315 -12255 -12307
rect -12289 -12341 -12255 -12315
rect -12289 -12383 -12255 -12379
rect -12289 -12413 -12255 -12383
rect 24855 -12111 24889 -12091
rect 24855 -12125 24889 -12111
rect 24855 -12179 24889 -12163
rect 24855 -12197 24889 -12179
rect 24855 -12247 24889 -12235
rect 24855 -12269 24889 -12247
rect 24855 -12315 24889 -12307
rect 24855 -12341 24889 -12315
rect 24855 -12383 24889 -12379
rect 24855 -12413 24889 -12383
rect -12289 -12485 -12255 -12451
rect -8855 -12474 -8845 -12440
rect -8845 -12474 -8821 -12440
rect -8783 -12474 -8777 -12440
rect -8777 -12474 -8749 -12440
rect -8711 -12474 -8709 -12440
rect -8709 -12474 -8677 -12440
rect -8639 -12474 -8607 -12440
rect -8607 -12474 -8605 -12440
rect -8567 -12474 -8539 -12440
rect -8539 -12474 -8533 -12440
rect -8495 -12474 -8471 -12440
rect -8471 -12474 -8461 -12440
rect -7837 -12474 -7827 -12440
rect -7827 -12474 -7803 -12440
rect -7765 -12474 -7759 -12440
rect -7759 -12474 -7731 -12440
rect -7693 -12474 -7691 -12440
rect -7691 -12474 -7659 -12440
rect -7621 -12474 -7589 -12440
rect -7589 -12474 -7587 -12440
rect -7549 -12474 -7521 -12440
rect -7521 -12474 -7515 -12440
rect -7477 -12474 -7453 -12440
rect -7453 -12474 -7443 -12440
rect -6819 -12474 -6809 -12440
rect -6809 -12474 -6785 -12440
rect -6747 -12474 -6741 -12440
rect -6741 -12474 -6713 -12440
rect -6675 -12474 -6673 -12440
rect -6673 -12474 -6641 -12440
rect -6603 -12474 -6571 -12440
rect -6571 -12474 -6569 -12440
rect -6531 -12474 -6503 -12440
rect -6503 -12474 -6497 -12440
rect -6459 -12474 -6435 -12440
rect -6435 -12474 -6425 -12440
rect -5801 -12474 -5791 -12440
rect -5791 -12474 -5767 -12440
rect -5729 -12474 -5723 -12440
rect -5723 -12474 -5695 -12440
rect -5657 -12474 -5655 -12440
rect -5655 -12474 -5623 -12440
rect -5585 -12474 -5553 -12440
rect -5553 -12474 -5551 -12440
rect -5513 -12474 -5485 -12440
rect -5485 -12474 -5479 -12440
rect -5441 -12474 -5417 -12440
rect -5417 -12474 -5407 -12440
rect -4783 -12474 -4773 -12440
rect -4773 -12474 -4749 -12440
rect -4711 -12474 -4705 -12440
rect -4705 -12474 -4677 -12440
rect -4639 -12474 -4637 -12440
rect -4637 -12474 -4605 -12440
rect -4567 -12474 -4535 -12440
rect -4535 -12474 -4533 -12440
rect -4495 -12474 -4467 -12440
rect -4467 -12474 -4461 -12440
rect -4423 -12474 -4399 -12440
rect -4399 -12474 -4389 -12440
rect -3765 -12474 -3755 -12440
rect -3755 -12474 -3731 -12440
rect -3693 -12474 -3687 -12440
rect -3687 -12474 -3659 -12440
rect -3621 -12474 -3619 -12440
rect -3619 -12474 -3587 -12440
rect -3549 -12474 -3517 -12440
rect -3517 -12474 -3515 -12440
rect -3477 -12474 -3449 -12440
rect -3449 -12474 -3443 -12440
rect -3405 -12474 -3381 -12440
rect -3381 -12474 -3371 -12440
rect -2747 -12474 -2737 -12440
rect -2737 -12474 -2713 -12440
rect -2675 -12474 -2669 -12440
rect -2669 -12474 -2641 -12440
rect -2603 -12474 -2601 -12440
rect -2601 -12474 -2569 -12440
rect -2531 -12474 -2499 -12440
rect -2499 -12474 -2497 -12440
rect -2459 -12474 -2431 -12440
rect -2431 -12474 -2425 -12440
rect -2387 -12474 -2363 -12440
rect -2363 -12474 -2353 -12440
rect -1729 -12474 -1719 -12440
rect -1719 -12474 -1695 -12440
rect -1657 -12474 -1651 -12440
rect -1651 -12474 -1623 -12440
rect -1585 -12474 -1583 -12440
rect -1583 -12474 -1551 -12440
rect -1513 -12474 -1481 -12440
rect -1481 -12474 -1479 -12440
rect -1441 -12474 -1413 -12440
rect -1413 -12474 -1407 -12440
rect -1369 -12474 -1345 -12440
rect -1345 -12474 -1335 -12440
rect -711 -12474 -701 -12440
rect -701 -12474 -677 -12440
rect -639 -12474 -633 -12440
rect -633 -12474 -605 -12440
rect -567 -12474 -565 -12440
rect -565 -12474 -533 -12440
rect -495 -12474 -463 -12440
rect -463 -12474 -461 -12440
rect -423 -12474 -395 -12440
rect -395 -12474 -389 -12440
rect -351 -12474 -327 -12440
rect -327 -12474 -317 -12440
rect 24855 -12485 24889 -12451
rect -12289 -12553 -12255 -12523
rect -12289 -12557 -12255 -12553
rect -12289 -12621 -12255 -12595
rect -12289 -12629 -12255 -12621
rect -12289 -12689 -12255 -12667
rect -12289 -12701 -12255 -12689
rect -12289 -12757 -12255 -12739
rect -12289 -12773 -12255 -12757
rect -12289 -12825 -12255 -12811
rect -12289 -12845 -12255 -12825
rect -12289 -12893 -12255 -12883
rect -12289 -12917 -12255 -12893
rect -12289 -12961 -12255 -12955
rect -12289 -12989 -12255 -12961
rect -12289 -13029 -12255 -13027
rect -12289 -13061 -12255 -13029
rect -12289 -13131 -12255 -13099
rect -12289 -13133 -12255 -13131
rect -9184 -12557 -9150 -12543
rect -9184 -12577 -9150 -12557
rect -9184 -12625 -9150 -12615
rect -9184 -12649 -9150 -12625
rect -9184 -12693 -9150 -12687
rect -9184 -12721 -9150 -12693
rect -9184 -12761 -9150 -12759
rect -9184 -12793 -9150 -12761
rect -9184 -12863 -9150 -12831
rect -9184 -12865 -9150 -12863
rect -9184 -12931 -9150 -12903
rect -9184 -12937 -9150 -12931
rect -9184 -12999 -9150 -12975
rect -9184 -13009 -9150 -12999
rect -9184 -13067 -9150 -13047
rect -9184 -13081 -9150 -13067
rect -8166 -12557 -8132 -12543
rect -8166 -12577 -8132 -12557
rect -8166 -12625 -8132 -12615
rect -8166 -12649 -8132 -12625
rect -8166 -12693 -8132 -12687
rect -8166 -12721 -8132 -12693
rect -8166 -12761 -8132 -12759
rect -8166 -12793 -8132 -12761
rect -8166 -12863 -8132 -12831
rect -8166 -12865 -8132 -12863
rect -8166 -12931 -8132 -12903
rect -8166 -12937 -8132 -12931
rect -8166 -12999 -8132 -12975
rect -8166 -13009 -8132 -12999
rect -8166 -13067 -8132 -13047
rect -8166 -13081 -8132 -13067
rect -7148 -12557 -7114 -12543
rect -7148 -12577 -7114 -12557
rect -7148 -12625 -7114 -12615
rect -7148 -12649 -7114 -12625
rect -7148 -12693 -7114 -12687
rect -7148 -12721 -7114 -12693
rect -7148 -12761 -7114 -12759
rect -7148 -12793 -7114 -12761
rect -7148 -12863 -7114 -12831
rect -7148 -12865 -7114 -12863
rect -7148 -12931 -7114 -12903
rect -7148 -12937 -7114 -12931
rect -7148 -12999 -7114 -12975
rect -7148 -13009 -7114 -12999
rect -7148 -13067 -7114 -13047
rect -7148 -13081 -7114 -13067
rect -6130 -12557 -6096 -12543
rect -6130 -12577 -6096 -12557
rect -6130 -12625 -6096 -12615
rect -6130 -12649 -6096 -12625
rect -6130 -12693 -6096 -12687
rect -6130 -12721 -6096 -12693
rect -6130 -12761 -6096 -12759
rect -6130 -12793 -6096 -12761
rect -6130 -12863 -6096 -12831
rect -6130 -12865 -6096 -12863
rect -6130 -12931 -6096 -12903
rect -6130 -12937 -6096 -12931
rect -6130 -12999 -6096 -12975
rect -6130 -13009 -6096 -12999
rect -6130 -13067 -6096 -13047
rect -6130 -13081 -6096 -13067
rect -5112 -12557 -5078 -12543
rect -5112 -12577 -5078 -12557
rect -5112 -12625 -5078 -12615
rect -5112 -12649 -5078 -12625
rect -5112 -12693 -5078 -12687
rect -5112 -12721 -5078 -12693
rect -5112 -12761 -5078 -12759
rect -5112 -12793 -5078 -12761
rect -5112 -12863 -5078 -12831
rect -5112 -12865 -5078 -12863
rect -5112 -12931 -5078 -12903
rect -5112 -12937 -5078 -12931
rect -5112 -12999 -5078 -12975
rect -5112 -13009 -5078 -12999
rect -5112 -13067 -5078 -13047
rect -5112 -13081 -5078 -13067
rect -4094 -12557 -4060 -12543
rect -4094 -12577 -4060 -12557
rect -4094 -12625 -4060 -12615
rect -4094 -12649 -4060 -12625
rect -4094 -12693 -4060 -12687
rect -4094 -12721 -4060 -12693
rect -4094 -12761 -4060 -12759
rect -4094 -12793 -4060 -12761
rect -4094 -12863 -4060 -12831
rect -4094 -12865 -4060 -12863
rect -4094 -12931 -4060 -12903
rect -4094 -12937 -4060 -12931
rect -4094 -12999 -4060 -12975
rect -4094 -13009 -4060 -12999
rect -4094 -13067 -4060 -13047
rect -4094 -13081 -4060 -13067
rect -3076 -12557 -3042 -12543
rect -3076 -12577 -3042 -12557
rect -3076 -12625 -3042 -12615
rect -3076 -12649 -3042 -12625
rect -3076 -12693 -3042 -12687
rect -3076 -12721 -3042 -12693
rect -3076 -12761 -3042 -12759
rect -3076 -12793 -3042 -12761
rect -3076 -12863 -3042 -12831
rect -3076 -12865 -3042 -12863
rect -3076 -12931 -3042 -12903
rect -3076 -12937 -3042 -12931
rect -3076 -12999 -3042 -12975
rect -3076 -13009 -3042 -12999
rect -3076 -13067 -3042 -13047
rect -3076 -13081 -3042 -13067
rect -2058 -12557 -2024 -12543
rect -2058 -12577 -2024 -12557
rect -2058 -12625 -2024 -12615
rect -2058 -12649 -2024 -12625
rect -2058 -12693 -2024 -12687
rect -2058 -12721 -2024 -12693
rect -2058 -12761 -2024 -12759
rect -2058 -12793 -2024 -12761
rect -2058 -12863 -2024 -12831
rect -2058 -12865 -2024 -12863
rect -2058 -12931 -2024 -12903
rect -2058 -12937 -2024 -12931
rect -2058 -12999 -2024 -12975
rect -2058 -13009 -2024 -12999
rect -2058 -13067 -2024 -13047
rect -2058 -13081 -2024 -13067
rect -1040 -12557 -1006 -12543
rect -1040 -12577 -1006 -12557
rect -1040 -12625 -1006 -12615
rect -1040 -12649 -1006 -12625
rect -1040 -12693 -1006 -12687
rect -1040 -12721 -1006 -12693
rect -1040 -12761 -1006 -12759
rect -1040 -12793 -1006 -12761
rect -1040 -12863 -1006 -12831
rect -1040 -12865 -1006 -12863
rect -1040 -12931 -1006 -12903
rect -1040 -12937 -1006 -12931
rect -1040 -12999 -1006 -12975
rect -1040 -13009 -1006 -12999
rect -1040 -13067 -1006 -13047
rect -1040 -13081 -1006 -13067
rect -22 -12557 12 -12543
rect -22 -12577 12 -12557
rect -22 -12625 12 -12615
rect -22 -12649 12 -12625
rect -22 -12693 12 -12687
rect -22 -12721 12 -12693
rect -22 -12761 12 -12759
rect -22 -12793 12 -12761
rect -22 -12863 12 -12831
rect -22 -12865 12 -12863
rect -22 -12931 12 -12903
rect -22 -12937 12 -12931
rect -22 -12999 12 -12975
rect -22 -13009 12 -12999
rect -22 -13067 12 -13047
rect -22 -13081 12 -13067
rect 24855 -12553 24889 -12523
rect 24855 -12557 24889 -12553
rect 24855 -12621 24889 -12595
rect 24855 -12629 24889 -12621
rect 24855 -12689 24889 -12667
rect 24855 -12701 24889 -12689
rect 24855 -12757 24889 -12739
rect 24855 -12773 24889 -12757
rect 24855 -12825 24889 -12811
rect 24855 -12845 24889 -12825
rect 24855 -12893 24889 -12883
rect 24855 -12917 24889 -12893
rect 24855 -12961 24889 -12955
rect 24855 -12989 24889 -12961
rect 24855 -13029 24889 -13027
rect 24855 -13061 24889 -13029
rect -12289 -13199 -12255 -13171
rect -12289 -13205 -12255 -13199
rect -8855 -13184 -8845 -13150
rect -8845 -13184 -8821 -13150
rect -8783 -13184 -8777 -13150
rect -8777 -13184 -8749 -13150
rect -8711 -13184 -8709 -13150
rect -8709 -13184 -8677 -13150
rect -8639 -13184 -8607 -13150
rect -8607 -13184 -8605 -13150
rect -8567 -13184 -8539 -13150
rect -8539 -13184 -8533 -13150
rect -8495 -13184 -8471 -13150
rect -8471 -13184 -8461 -13150
rect -7837 -13184 -7827 -13150
rect -7827 -13184 -7803 -13150
rect -7765 -13184 -7759 -13150
rect -7759 -13184 -7731 -13150
rect -7693 -13184 -7691 -13150
rect -7691 -13184 -7659 -13150
rect -7621 -13184 -7589 -13150
rect -7589 -13184 -7587 -13150
rect -7549 -13184 -7521 -13150
rect -7521 -13184 -7515 -13150
rect -7477 -13184 -7453 -13150
rect -7453 -13184 -7443 -13150
rect -6819 -13184 -6809 -13150
rect -6809 -13184 -6785 -13150
rect -6747 -13184 -6741 -13150
rect -6741 -13184 -6713 -13150
rect -6675 -13184 -6673 -13150
rect -6673 -13184 -6641 -13150
rect -6603 -13184 -6571 -13150
rect -6571 -13184 -6569 -13150
rect -6531 -13184 -6503 -13150
rect -6503 -13184 -6497 -13150
rect -6459 -13184 -6435 -13150
rect -6435 -13184 -6425 -13150
rect -5801 -13184 -5791 -13150
rect -5791 -13184 -5767 -13150
rect -5729 -13184 -5723 -13150
rect -5723 -13184 -5695 -13150
rect -5657 -13184 -5655 -13150
rect -5655 -13184 -5623 -13150
rect -5585 -13184 -5553 -13150
rect -5553 -13184 -5551 -13150
rect -5513 -13184 -5485 -13150
rect -5485 -13184 -5479 -13150
rect -5441 -13184 -5417 -13150
rect -5417 -13184 -5407 -13150
rect -4783 -13184 -4773 -13150
rect -4773 -13184 -4749 -13150
rect -4711 -13184 -4705 -13150
rect -4705 -13184 -4677 -13150
rect -4639 -13184 -4637 -13150
rect -4637 -13184 -4605 -13150
rect -4567 -13184 -4535 -13150
rect -4535 -13184 -4533 -13150
rect -4495 -13184 -4467 -13150
rect -4467 -13184 -4461 -13150
rect -4423 -13184 -4399 -13150
rect -4399 -13184 -4389 -13150
rect -3765 -13184 -3755 -13150
rect -3755 -13184 -3731 -13150
rect -3693 -13184 -3687 -13150
rect -3687 -13184 -3659 -13150
rect -3621 -13184 -3619 -13150
rect -3619 -13184 -3587 -13150
rect -3549 -13184 -3517 -13150
rect -3517 -13184 -3515 -13150
rect -3477 -13184 -3449 -13150
rect -3449 -13184 -3443 -13150
rect -3405 -13184 -3381 -13150
rect -3381 -13184 -3371 -13150
rect -2747 -13184 -2737 -13150
rect -2737 -13184 -2713 -13150
rect -2675 -13184 -2669 -13150
rect -2669 -13184 -2641 -13150
rect -2603 -13184 -2601 -13150
rect -2601 -13184 -2569 -13150
rect -2531 -13184 -2499 -13150
rect -2499 -13184 -2497 -13150
rect -2459 -13184 -2431 -13150
rect -2431 -13184 -2425 -13150
rect -2387 -13184 -2363 -13150
rect -2363 -13184 -2353 -13150
rect -1729 -13184 -1719 -13150
rect -1719 -13184 -1695 -13150
rect -1657 -13184 -1651 -13150
rect -1651 -13184 -1623 -13150
rect -1585 -13184 -1583 -13150
rect -1583 -13184 -1551 -13150
rect -1513 -13184 -1481 -13150
rect -1481 -13184 -1479 -13150
rect -1441 -13184 -1413 -13150
rect -1413 -13184 -1407 -13150
rect -1369 -13184 -1345 -13150
rect -1345 -13184 -1335 -13150
rect -711 -13184 -701 -13150
rect -701 -13184 -677 -13150
rect -639 -13184 -633 -13150
rect -633 -13184 -605 -13150
rect -567 -13184 -565 -13150
rect -565 -13184 -533 -13150
rect -495 -13184 -463 -13150
rect -463 -13184 -461 -13150
rect -423 -13184 -395 -13150
rect -395 -13184 -389 -13150
rect -351 -13184 -327 -13150
rect -327 -13184 -317 -13150
rect 24855 -13131 24889 -13099
rect 24855 -13133 24889 -13131
rect -12289 -13267 -12255 -13243
rect -12289 -13277 -12255 -13267
rect 24855 -13199 24889 -13171
rect 24855 -13205 24889 -13199
rect -8855 -13292 -8845 -13258
rect -8845 -13292 -8821 -13258
rect -8783 -13292 -8777 -13258
rect -8777 -13292 -8749 -13258
rect -8711 -13292 -8709 -13258
rect -8709 -13292 -8677 -13258
rect -8639 -13292 -8607 -13258
rect -8607 -13292 -8605 -13258
rect -8567 -13292 -8539 -13258
rect -8539 -13292 -8533 -13258
rect -8495 -13292 -8471 -13258
rect -8471 -13292 -8461 -13258
rect -7837 -13292 -7827 -13258
rect -7827 -13292 -7803 -13258
rect -7765 -13292 -7759 -13258
rect -7759 -13292 -7731 -13258
rect -7693 -13292 -7691 -13258
rect -7691 -13292 -7659 -13258
rect -7621 -13292 -7589 -13258
rect -7589 -13292 -7587 -13258
rect -7549 -13292 -7521 -13258
rect -7521 -13292 -7515 -13258
rect -7477 -13292 -7453 -13258
rect -7453 -13292 -7443 -13258
rect -6819 -13292 -6809 -13258
rect -6809 -13292 -6785 -13258
rect -6747 -13292 -6741 -13258
rect -6741 -13292 -6713 -13258
rect -6675 -13292 -6673 -13258
rect -6673 -13292 -6641 -13258
rect -6603 -13292 -6571 -13258
rect -6571 -13292 -6569 -13258
rect -6531 -13292 -6503 -13258
rect -6503 -13292 -6497 -13258
rect -6459 -13292 -6435 -13258
rect -6435 -13292 -6425 -13258
rect -5801 -13292 -5791 -13258
rect -5791 -13292 -5767 -13258
rect -5729 -13292 -5723 -13258
rect -5723 -13292 -5695 -13258
rect -5657 -13292 -5655 -13258
rect -5655 -13292 -5623 -13258
rect -5585 -13292 -5553 -13258
rect -5553 -13292 -5551 -13258
rect -5513 -13292 -5485 -13258
rect -5485 -13292 -5479 -13258
rect -5441 -13292 -5417 -13258
rect -5417 -13292 -5407 -13258
rect -4783 -13292 -4773 -13258
rect -4773 -13292 -4749 -13258
rect -4711 -13292 -4705 -13258
rect -4705 -13292 -4677 -13258
rect -4639 -13292 -4637 -13258
rect -4637 -13292 -4605 -13258
rect -4567 -13292 -4535 -13258
rect -4535 -13292 -4533 -13258
rect -4495 -13292 -4467 -13258
rect -4467 -13292 -4461 -13258
rect -4423 -13292 -4399 -13258
rect -4399 -13292 -4389 -13258
rect -3765 -13292 -3755 -13258
rect -3755 -13292 -3731 -13258
rect -3693 -13292 -3687 -13258
rect -3687 -13292 -3659 -13258
rect -3621 -13292 -3619 -13258
rect -3619 -13292 -3587 -13258
rect -3549 -13292 -3517 -13258
rect -3517 -13292 -3515 -13258
rect -3477 -13292 -3449 -13258
rect -3449 -13292 -3443 -13258
rect -3405 -13292 -3381 -13258
rect -3381 -13292 -3371 -13258
rect -2747 -13292 -2737 -13258
rect -2737 -13292 -2713 -13258
rect -2675 -13292 -2669 -13258
rect -2669 -13292 -2641 -13258
rect -2603 -13292 -2601 -13258
rect -2601 -13292 -2569 -13258
rect -2531 -13292 -2499 -13258
rect -2499 -13292 -2497 -13258
rect -2459 -13292 -2431 -13258
rect -2431 -13292 -2425 -13258
rect -2387 -13292 -2363 -13258
rect -2363 -13292 -2353 -13258
rect -1729 -13292 -1719 -13258
rect -1719 -13292 -1695 -13258
rect -1657 -13292 -1651 -13258
rect -1651 -13292 -1623 -13258
rect -1585 -13292 -1583 -13258
rect -1583 -13292 -1551 -13258
rect -1513 -13292 -1481 -13258
rect -1481 -13292 -1479 -13258
rect -1441 -13292 -1413 -13258
rect -1413 -13292 -1407 -13258
rect -1369 -13292 -1345 -13258
rect -1345 -13292 -1335 -13258
rect -711 -13292 -701 -13258
rect -701 -13292 -677 -13258
rect -639 -13292 -633 -13258
rect -633 -13292 -605 -13258
rect -567 -13292 -565 -13258
rect -565 -13292 -533 -13258
rect -495 -13292 -463 -13258
rect -463 -13292 -461 -13258
rect -423 -13292 -395 -13258
rect -395 -13292 -389 -13258
rect -351 -13292 -327 -13258
rect -327 -13292 -317 -13258
rect -12289 -13335 -12255 -13315
rect -12289 -13349 -12255 -13335
rect 24855 -13267 24889 -13243
rect 24855 -13277 24889 -13267
rect -12289 -13403 -12255 -13387
rect -12289 -13421 -12255 -13403
rect -12289 -13471 -12255 -13459
rect -12289 -13493 -12255 -13471
rect -12289 -13539 -12255 -13531
rect -12289 -13565 -12255 -13539
rect -12289 -13607 -12255 -13603
rect -12289 -13637 -12255 -13607
rect -12289 -13709 -12255 -13675
rect -12289 -13777 -12255 -13747
rect -12289 -13781 -12255 -13777
rect -12289 -13845 -12255 -13819
rect -12289 -13853 -12255 -13845
rect -12289 -13913 -12255 -13891
rect -12289 -13925 -12255 -13913
rect -9184 -13375 -9150 -13361
rect -9184 -13395 -9150 -13375
rect -9184 -13443 -9150 -13433
rect -9184 -13467 -9150 -13443
rect -9184 -13511 -9150 -13505
rect -9184 -13539 -9150 -13511
rect -9184 -13579 -9150 -13577
rect -9184 -13611 -9150 -13579
rect -9184 -13681 -9150 -13649
rect -9184 -13683 -9150 -13681
rect -9184 -13749 -9150 -13721
rect -9184 -13755 -9150 -13749
rect -9184 -13817 -9150 -13793
rect -9184 -13827 -9150 -13817
rect -9184 -13885 -9150 -13865
rect -9184 -13899 -9150 -13885
rect -8166 -13375 -8132 -13361
rect -8166 -13395 -8132 -13375
rect -8166 -13443 -8132 -13433
rect -8166 -13467 -8132 -13443
rect -8166 -13511 -8132 -13505
rect -8166 -13539 -8132 -13511
rect -8166 -13579 -8132 -13577
rect -8166 -13611 -8132 -13579
rect -8166 -13681 -8132 -13649
rect -8166 -13683 -8132 -13681
rect -8166 -13749 -8132 -13721
rect -8166 -13755 -8132 -13749
rect -8166 -13817 -8132 -13793
rect -8166 -13827 -8132 -13817
rect -8166 -13885 -8132 -13865
rect -8166 -13899 -8132 -13885
rect -7148 -13375 -7114 -13361
rect -7148 -13395 -7114 -13375
rect -7148 -13443 -7114 -13433
rect -7148 -13467 -7114 -13443
rect -7148 -13511 -7114 -13505
rect -7148 -13539 -7114 -13511
rect -7148 -13579 -7114 -13577
rect -7148 -13611 -7114 -13579
rect -7148 -13681 -7114 -13649
rect -7148 -13683 -7114 -13681
rect -7148 -13749 -7114 -13721
rect -7148 -13755 -7114 -13749
rect -7148 -13817 -7114 -13793
rect -7148 -13827 -7114 -13817
rect -7148 -13885 -7114 -13865
rect -7148 -13899 -7114 -13885
rect -6130 -13375 -6096 -13361
rect -6130 -13395 -6096 -13375
rect -6130 -13443 -6096 -13433
rect -6130 -13467 -6096 -13443
rect -6130 -13511 -6096 -13505
rect -6130 -13539 -6096 -13511
rect -6130 -13579 -6096 -13577
rect -6130 -13611 -6096 -13579
rect -6130 -13681 -6096 -13649
rect -6130 -13683 -6096 -13681
rect -6130 -13749 -6096 -13721
rect -6130 -13755 -6096 -13749
rect -6130 -13817 -6096 -13793
rect -6130 -13827 -6096 -13817
rect -6130 -13885 -6096 -13865
rect -6130 -13899 -6096 -13885
rect -5112 -13375 -5078 -13361
rect -5112 -13395 -5078 -13375
rect -5112 -13443 -5078 -13433
rect -5112 -13467 -5078 -13443
rect -5112 -13511 -5078 -13505
rect -5112 -13539 -5078 -13511
rect -5112 -13579 -5078 -13577
rect -5112 -13611 -5078 -13579
rect -5112 -13681 -5078 -13649
rect -5112 -13683 -5078 -13681
rect -5112 -13749 -5078 -13721
rect -5112 -13755 -5078 -13749
rect -5112 -13817 -5078 -13793
rect -5112 -13827 -5078 -13817
rect -5112 -13885 -5078 -13865
rect -5112 -13899 -5078 -13885
rect -4094 -13375 -4060 -13361
rect -4094 -13395 -4060 -13375
rect -4094 -13443 -4060 -13433
rect -4094 -13467 -4060 -13443
rect -4094 -13511 -4060 -13505
rect -4094 -13539 -4060 -13511
rect -4094 -13579 -4060 -13577
rect -4094 -13611 -4060 -13579
rect -4094 -13681 -4060 -13649
rect -4094 -13683 -4060 -13681
rect -4094 -13749 -4060 -13721
rect -4094 -13755 -4060 -13749
rect -4094 -13817 -4060 -13793
rect -4094 -13827 -4060 -13817
rect -4094 -13885 -4060 -13865
rect -4094 -13899 -4060 -13885
rect -3076 -13375 -3042 -13361
rect -3076 -13395 -3042 -13375
rect -3076 -13443 -3042 -13433
rect -3076 -13467 -3042 -13443
rect -3076 -13511 -3042 -13505
rect -3076 -13539 -3042 -13511
rect -3076 -13579 -3042 -13577
rect -3076 -13611 -3042 -13579
rect -3076 -13681 -3042 -13649
rect -3076 -13683 -3042 -13681
rect -3076 -13749 -3042 -13721
rect -3076 -13755 -3042 -13749
rect -3076 -13817 -3042 -13793
rect -3076 -13827 -3042 -13817
rect -3076 -13885 -3042 -13865
rect -3076 -13899 -3042 -13885
rect -2058 -13375 -2024 -13361
rect -2058 -13395 -2024 -13375
rect -2058 -13443 -2024 -13433
rect -2058 -13467 -2024 -13443
rect -2058 -13511 -2024 -13505
rect -2058 -13539 -2024 -13511
rect -2058 -13579 -2024 -13577
rect -2058 -13611 -2024 -13579
rect -2058 -13681 -2024 -13649
rect -2058 -13683 -2024 -13681
rect -2058 -13749 -2024 -13721
rect -2058 -13755 -2024 -13749
rect -2058 -13817 -2024 -13793
rect -2058 -13827 -2024 -13817
rect -2058 -13885 -2024 -13865
rect -2058 -13899 -2024 -13885
rect -1040 -13375 -1006 -13361
rect -1040 -13395 -1006 -13375
rect -1040 -13443 -1006 -13433
rect -1040 -13467 -1006 -13443
rect -1040 -13511 -1006 -13505
rect -1040 -13539 -1006 -13511
rect -1040 -13579 -1006 -13577
rect -1040 -13611 -1006 -13579
rect -1040 -13681 -1006 -13649
rect -1040 -13683 -1006 -13681
rect -1040 -13749 -1006 -13721
rect -1040 -13755 -1006 -13749
rect -1040 -13817 -1006 -13793
rect -1040 -13827 -1006 -13817
rect -1040 -13885 -1006 -13865
rect -1040 -13899 -1006 -13885
rect -22 -13375 12 -13361
rect -22 -13395 12 -13375
rect -22 -13443 12 -13433
rect -22 -13467 12 -13443
rect -22 -13511 12 -13505
rect -22 -13539 12 -13511
rect -22 -13579 12 -13577
rect -22 -13611 12 -13579
rect -22 -13681 12 -13649
rect -22 -13683 12 -13681
rect -22 -13749 12 -13721
rect -22 -13755 12 -13749
rect -22 -13817 12 -13793
rect -22 -13827 12 -13817
rect -22 -13885 12 -13865
rect -22 -13899 12 -13885
rect 24855 -13335 24889 -13315
rect 24855 -13349 24889 -13335
rect 24855 -13403 24889 -13387
rect 24855 -13421 24889 -13403
rect 24855 -13471 24889 -13459
rect 24855 -13493 24889 -13471
rect 24855 -13539 24889 -13531
rect 24855 -13565 24889 -13539
rect 24855 -13607 24889 -13603
rect 24855 -13637 24889 -13607
rect 24855 -13709 24889 -13675
rect 24855 -13777 24889 -13747
rect 24855 -13781 24889 -13777
rect 24855 -13845 24889 -13819
rect 24855 -13853 24889 -13845
rect 24855 -13913 24889 -13891
rect 24855 -13925 24889 -13913
rect -12289 -13981 -12255 -13963
rect -12289 -13997 -12255 -13981
rect -8855 -14002 -8845 -13968
rect -8845 -14002 -8821 -13968
rect -8783 -14002 -8777 -13968
rect -8777 -14002 -8749 -13968
rect -8711 -14002 -8709 -13968
rect -8709 -14002 -8677 -13968
rect -8639 -14002 -8607 -13968
rect -8607 -14002 -8605 -13968
rect -8567 -14002 -8539 -13968
rect -8539 -14002 -8533 -13968
rect -8495 -14002 -8471 -13968
rect -8471 -14002 -8461 -13968
rect -7837 -14002 -7827 -13968
rect -7827 -14002 -7803 -13968
rect -7765 -14002 -7759 -13968
rect -7759 -14002 -7731 -13968
rect -7693 -14002 -7691 -13968
rect -7691 -14002 -7659 -13968
rect -7621 -14002 -7589 -13968
rect -7589 -14002 -7587 -13968
rect -7549 -14002 -7521 -13968
rect -7521 -14002 -7515 -13968
rect -7477 -14002 -7453 -13968
rect -7453 -14002 -7443 -13968
rect -6819 -14002 -6809 -13968
rect -6809 -14002 -6785 -13968
rect -6747 -14002 -6741 -13968
rect -6741 -14002 -6713 -13968
rect -6675 -14002 -6673 -13968
rect -6673 -14002 -6641 -13968
rect -6603 -14002 -6571 -13968
rect -6571 -14002 -6569 -13968
rect -6531 -14002 -6503 -13968
rect -6503 -14002 -6497 -13968
rect -6459 -14002 -6435 -13968
rect -6435 -14002 -6425 -13968
rect -5801 -14002 -5791 -13968
rect -5791 -14002 -5767 -13968
rect -5729 -14002 -5723 -13968
rect -5723 -14002 -5695 -13968
rect -5657 -14002 -5655 -13968
rect -5655 -14002 -5623 -13968
rect -5585 -14002 -5553 -13968
rect -5553 -14002 -5551 -13968
rect -5513 -14002 -5485 -13968
rect -5485 -14002 -5479 -13968
rect -5441 -14002 -5417 -13968
rect -5417 -14002 -5407 -13968
rect -4783 -14002 -4773 -13968
rect -4773 -14002 -4749 -13968
rect -4711 -14002 -4705 -13968
rect -4705 -14002 -4677 -13968
rect -4639 -14002 -4637 -13968
rect -4637 -14002 -4605 -13968
rect -4567 -14002 -4535 -13968
rect -4535 -14002 -4533 -13968
rect -4495 -14002 -4467 -13968
rect -4467 -14002 -4461 -13968
rect -4423 -14002 -4399 -13968
rect -4399 -14002 -4389 -13968
rect -3765 -14002 -3755 -13968
rect -3755 -14002 -3731 -13968
rect -3693 -14002 -3687 -13968
rect -3687 -14002 -3659 -13968
rect -3621 -14002 -3619 -13968
rect -3619 -14002 -3587 -13968
rect -3549 -14002 -3517 -13968
rect -3517 -14002 -3515 -13968
rect -3477 -14002 -3449 -13968
rect -3449 -14002 -3443 -13968
rect -3405 -14002 -3381 -13968
rect -3381 -14002 -3371 -13968
rect -2747 -14002 -2737 -13968
rect -2737 -14002 -2713 -13968
rect -2675 -14002 -2669 -13968
rect -2669 -14002 -2641 -13968
rect -2603 -14002 -2601 -13968
rect -2601 -14002 -2569 -13968
rect -2531 -14002 -2499 -13968
rect -2499 -14002 -2497 -13968
rect -2459 -14002 -2431 -13968
rect -2431 -14002 -2425 -13968
rect -2387 -14002 -2363 -13968
rect -2363 -14002 -2353 -13968
rect -1729 -14002 -1719 -13968
rect -1719 -14002 -1695 -13968
rect -1657 -14002 -1651 -13968
rect -1651 -14002 -1623 -13968
rect -1585 -14002 -1583 -13968
rect -1583 -14002 -1551 -13968
rect -1513 -14002 -1481 -13968
rect -1481 -14002 -1479 -13968
rect -1441 -14002 -1413 -13968
rect -1413 -14002 -1407 -13968
rect -1369 -14002 -1345 -13968
rect -1345 -14002 -1335 -13968
rect -711 -14002 -701 -13968
rect -701 -14002 -677 -13968
rect -639 -14002 -633 -13968
rect -633 -14002 -605 -13968
rect -567 -14002 -565 -13968
rect -565 -14002 -533 -13968
rect -495 -14002 -463 -13968
rect -463 -14002 -461 -13968
rect -423 -14002 -395 -13968
rect -395 -14002 -389 -13968
rect -351 -14002 -327 -13968
rect -327 -14002 -317 -13968
rect 24855 -13981 24889 -13963
rect 24855 -13997 24889 -13981
rect -12289 -14049 -12255 -14035
rect -12289 -14069 -12255 -14049
rect 24855 -14049 24889 -14035
rect 24855 -14069 24889 -14049
rect -12289 -14117 -12255 -14107
rect -12289 -14141 -12255 -14117
rect -8855 -14110 -8845 -14076
rect -8845 -14110 -8821 -14076
rect -8783 -14110 -8777 -14076
rect -8777 -14110 -8749 -14076
rect -8711 -14110 -8709 -14076
rect -8709 -14110 -8677 -14076
rect -8639 -14110 -8607 -14076
rect -8607 -14110 -8605 -14076
rect -8567 -14110 -8539 -14076
rect -8539 -14110 -8533 -14076
rect -8495 -14110 -8471 -14076
rect -8471 -14110 -8461 -14076
rect -7837 -14110 -7827 -14076
rect -7827 -14110 -7803 -14076
rect -7765 -14110 -7759 -14076
rect -7759 -14110 -7731 -14076
rect -7693 -14110 -7691 -14076
rect -7691 -14110 -7659 -14076
rect -7621 -14110 -7589 -14076
rect -7589 -14110 -7587 -14076
rect -7549 -14110 -7521 -14076
rect -7521 -14110 -7515 -14076
rect -7477 -14110 -7453 -14076
rect -7453 -14110 -7443 -14076
rect -6819 -14110 -6809 -14076
rect -6809 -14110 -6785 -14076
rect -6747 -14110 -6741 -14076
rect -6741 -14110 -6713 -14076
rect -6675 -14110 -6673 -14076
rect -6673 -14110 -6641 -14076
rect -6603 -14110 -6571 -14076
rect -6571 -14110 -6569 -14076
rect -6531 -14110 -6503 -14076
rect -6503 -14110 -6497 -14076
rect -6459 -14110 -6435 -14076
rect -6435 -14110 -6425 -14076
rect -5801 -14110 -5791 -14076
rect -5791 -14110 -5767 -14076
rect -5729 -14110 -5723 -14076
rect -5723 -14110 -5695 -14076
rect -5657 -14110 -5655 -14076
rect -5655 -14110 -5623 -14076
rect -5585 -14110 -5553 -14076
rect -5553 -14110 -5551 -14076
rect -5513 -14110 -5485 -14076
rect -5485 -14110 -5479 -14076
rect -5441 -14110 -5417 -14076
rect -5417 -14110 -5407 -14076
rect -4783 -14110 -4773 -14076
rect -4773 -14110 -4749 -14076
rect -4711 -14110 -4705 -14076
rect -4705 -14110 -4677 -14076
rect -4639 -14110 -4637 -14076
rect -4637 -14110 -4605 -14076
rect -4567 -14110 -4535 -14076
rect -4535 -14110 -4533 -14076
rect -4495 -14110 -4467 -14076
rect -4467 -14110 -4461 -14076
rect -4423 -14110 -4399 -14076
rect -4399 -14110 -4389 -14076
rect -3765 -14110 -3755 -14076
rect -3755 -14110 -3731 -14076
rect -3693 -14110 -3687 -14076
rect -3687 -14110 -3659 -14076
rect -3621 -14110 -3619 -14076
rect -3619 -14110 -3587 -14076
rect -3549 -14110 -3517 -14076
rect -3517 -14110 -3515 -14076
rect -3477 -14110 -3449 -14076
rect -3449 -14110 -3443 -14076
rect -3405 -14110 -3381 -14076
rect -3381 -14110 -3371 -14076
rect -2747 -14110 -2737 -14076
rect -2737 -14110 -2713 -14076
rect -2675 -14110 -2669 -14076
rect -2669 -14110 -2641 -14076
rect -2603 -14110 -2601 -14076
rect -2601 -14110 -2569 -14076
rect -2531 -14110 -2499 -14076
rect -2499 -14110 -2497 -14076
rect -2459 -14110 -2431 -14076
rect -2431 -14110 -2425 -14076
rect -2387 -14110 -2363 -14076
rect -2363 -14110 -2353 -14076
rect -1729 -14110 -1719 -14076
rect -1719 -14110 -1695 -14076
rect -1657 -14110 -1651 -14076
rect -1651 -14110 -1623 -14076
rect -1585 -14110 -1583 -14076
rect -1583 -14110 -1551 -14076
rect -1513 -14110 -1481 -14076
rect -1481 -14110 -1479 -14076
rect -1441 -14110 -1413 -14076
rect -1413 -14110 -1407 -14076
rect -1369 -14110 -1345 -14076
rect -1345 -14110 -1335 -14076
rect -711 -14110 -701 -14076
rect -701 -14110 -677 -14076
rect -639 -14110 -633 -14076
rect -633 -14110 -605 -14076
rect -567 -14110 -565 -14076
rect -565 -14110 -533 -14076
rect -495 -14110 -463 -14076
rect -463 -14110 -461 -14076
rect -423 -14110 -395 -14076
rect -395 -14110 -389 -14076
rect -351 -14110 -327 -14076
rect -327 -14110 -317 -14076
rect 24855 -14117 24889 -14107
rect 24855 -14141 24889 -14117
rect -12289 -14185 -12255 -14179
rect -12289 -14213 -12255 -14185
rect -12289 -14253 -12255 -14251
rect -12289 -14285 -12255 -14253
rect -12289 -14355 -12255 -14323
rect -12289 -14357 -12255 -14355
rect -12289 -14423 -12255 -14395
rect -12289 -14429 -12255 -14423
rect -12289 -14491 -12255 -14467
rect -12289 -14501 -12255 -14491
rect -12289 -14559 -12255 -14539
rect -12289 -14573 -12255 -14559
rect -12289 -14627 -12255 -14611
rect -12289 -14645 -12255 -14627
rect -12289 -14695 -12255 -14683
rect -12289 -14717 -12255 -14695
rect -9184 -14193 -9150 -14179
rect -9184 -14213 -9150 -14193
rect -9184 -14261 -9150 -14251
rect -9184 -14285 -9150 -14261
rect -9184 -14329 -9150 -14323
rect -9184 -14357 -9150 -14329
rect -9184 -14397 -9150 -14395
rect -9184 -14429 -9150 -14397
rect -9184 -14499 -9150 -14467
rect -9184 -14501 -9150 -14499
rect -9184 -14567 -9150 -14539
rect -9184 -14573 -9150 -14567
rect -9184 -14635 -9150 -14611
rect -9184 -14645 -9150 -14635
rect -9184 -14703 -9150 -14683
rect -9184 -14717 -9150 -14703
rect -8166 -14193 -8132 -14179
rect -8166 -14213 -8132 -14193
rect -8166 -14261 -8132 -14251
rect -8166 -14285 -8132 -14261
rect -8166 -14329 -8132 -14323
rect -8166 -14357 -8132 -14329
rect -8166 -14397 -8132 -14395
rect -8166 -14429 -8132 -14397
rect -8166 -14499 -8132 -14467
rect -8166 -14501 -8132 -14499
rect -8166 -14567 -8132 -14539
rect -8166 -14573 -8132 -14567
rect -8166 -14635 -8132 -14611
rect -8166 -14645 -8132 -14635
rect -8166 -14703 -8132 -14683
rect -8166 -14717 -8132 -14703
rect -7148 -14193 -7114 -14179
rect -7148 -14213 -7114 -14193
rect -7148 -14261 -7114 -14251
rect -7148 -14285 -7114 -14261
rect -7148 -14329 -7114 -14323
rect -7148 -14357 -7114 -14329
rect -7148 -14397 -7114 -14395
rect -7148 -14429 -7114 -14397
rect -7148 -14499 -7114 -14467
rect -7148 -14501 -7114 -14499
rect -7148 -14567 -7114 -14539
rect -7148 -14573 -7114 -14567
rect -7148 -14635 -7114 -14611
rect -7148 -14645 -7114 -14635
rect -7148 -14703 -7114 -14683
rect -7148 -14717 -7114 -14703
rect -6130 -14193 -6096 -14179
rect -6130 -14213 -6096 -14193
rect -6130 -14261 -6096 -14251
rect -6130 -14285 -6096 -14261
rect -6130 -14329 -6096 -14323
rect -6130 -14357 -6096 -14329
rect -6130 -14397 -6096 -14395
rect -6130 -14429 -6096 -14397
rect -6130 -14499 -6096 -14467
rect -6130 -14501 -6096 -14499
rect -6130 -14567 -6096 -14539
rect -6130 -14573 -6096 -14567
rect -6130 -14635 -6096 -14611
rect -6130 -14645 -6096 -14635
rect -6130 -14703 -6096 -14683
rect -6130 -14717 -6096 -14703
rect -5112 -14193 -5078 -14179
rect -5112 -14213 -5078 -14193
rect -5112 -14261 -5078 -14251
rect -5112 -14285 -5078 -14261
rect -5112 -14329 -5078 -14323
rect -5112 -14357 -5078 -14329
rect -5112 -14397 -5078 -14395
rect -5112 -14429 -5078 -14397
rect -5112 -14499 -5078 -14467
rect -5112 -14501 -5078 -14499
rect -5112 -14567 -5078 -14539
rect -5112 -14573 -5078 -14567
rect -5112 -14635 -5078 -14611
rect -5112 -14645 -5078 -14635
rect -5112 -14703 -5078 -14683
rect -5112 -14717 -5078 -14703
rect -4094 -14193 -4060 -14179
rect -4094 -14213 -4060 -14193
rect -4094 -14261 -4060 -14251
rect -4094 -14285 -4060 -14261
rect -4094 -14329 -4060 -14323
rect -4094 -14357 -4060 -14329
rect -4094 -14397 -4060 -14395
rect -4094 -14429 -4060 -14397
rect -4094 -14499 -4060 -14467
rect -4094 -14501 -4060 -14499
rect -4094 -14567 -4060 -14539
rect -4094 -14573 -4060 -14567
rect -4094 -14635 -4060 -14611
rect -4094 -14645 -4060 -14635
rect -4094 -14703 -4060 -14683
rect -4094 -14717 -4060 -14703
rect -3076 -14193 -3042 -14179
rect -3076 -14213 -3042 -14193
rect -3076 -14261 -3042 -14251
rect -3076 -14285 -3042 -14261
rect -3076 -14329 -3042 -14323
rect -3076 -14357 -3042 -14329
rect -3076 -14397 -3042 -14395
rect -3076 -14429 -3042 -14397
rect -3076 -14499 -3042 -14467
rect -3076 -14501 -3042 -14499
rect -3076 -14567 -3042 -14539
rect -3076 -14573 -3042 -14567
rect -3076 -14635 -3042 -14611
rect -3076 -14645 -3042 -14635
rect -3076 -14703 -3042 -14683
rect -3076 -14717 -3042 -14703
rect -2058 -14193 -2024 -14179
rect -2058 -14213 -2024 -14193
rect -2058 -14261 -2024 -14251
rect -2058 -14285 -2024 -14261
rect -2058 -14329 -2024 -14323
rect -2058 -14357 -2024 -14329
rect -2058 -14397 -2024 -14395
rect -2058 -14429 -2024 -14397
rect -2058 -14499 -2024 -14467
rect -2058 -14501 -2024 -14499
rect -2058 -14567 -2024 -14539
rect -2058 -14573 -2024 -14567
rect -2058 -14635 -2024 -14611
rect -2058 -14645 -2024 -14635
rect -2058 -14703 -2024 -14683
rect -2058 -14717 -2024 -14703
rect -1040 -14193 -1006 -14179
rect -1040 -14213 -1006 -14193
rect -1040 -14261 -1006 -14251
rect -1040 -14285 -1006 -14261
rect -1040 -14329 -1006 -14323
rect -1040 -14357 -1006 -14329
rect -1040 -14397 -1006 -14395
rect -1040 -14429 -1006 -14397
rect -1040 -14499 -1006 -14467
rect -1040 -14501 -1006 -14499
rect -1040 -14567 -1006 -14539
rect -1040 -14573 -1006 -14567
rect -1040 -14635 -1006 -14611
rect -1040 -14645 -1006 -14635
rect -1040 -14703 -1006 -14683
rect -1040 -14717 -1006 -14703
rect -22 -14193 12 -14179
rect -22 -14213 12 -14193
rect 2911 -14194 2921 -14160
rect 2921 -14194 2945 -14160
rect 2983 -14194 2989 -14160
rect 2989 -14194 3017 -14160
rect 3055 -14194 3057 -14160
rect 3057 -14194 3089 -14160
rect 3127 -14194 3159 -14160
rect 3159 -14194 3161 -14160
rect 3199 -14194 3227 -14160
rect 3227 -14194 3233 -14160
rect 3271 -14194 3295 -14160
rect 3295 -14194 3305 -14160
rect 3929 -14194 3939 -14160
rect 3939 -14194 3963 -14160
rect 4001 -14194 4007 -14160
rect 4007 -14194 4035 -14160
rect 4073 -14194 4075 -14160
rect 4075 -14194 4107 -14160
rect 4145 -14194 4177 -14160
rect 4177 -14194 4179 -14160
rect 4217 -14194 4245 -14160
rect 4245 -14194 4251 -14160
rect 4289 -14194 4313 -14160
rect 4313 -14194 4323 -14160
rect 4947 -14194 4957 -14160
rect 4957 -14194 4981 -14160
rect 5019 -14194 5025 -14160
rect 5025 -14194 5053 -14160
rect 5091 -14194 5093 -14160
rect 5093 -14194 5125 -14160
rect 5163 -14194 5195 -14160
rect 5195 -14194 5197 -14160
rect 5235 -14194 5263 -14160
rect 5263 -14194 5269 -14160
rect 5307 -14194 5331 -14160
rect 5331 -14194 5341 -14160
rect 5965 -14194 5975 -14160
rect 5975 -14194 5999 -14160
rect 6037 -14194 6043 -14160
rect 6043 -14194 6071 -14160
rect 6109 -14194 6111 -14160
rect 6111 -14194 6143 -14160
rect 6181 -14194 6213 -14160
rect 6213 -14194 6215 -14160
rect 6253 -14194 6281 -14160
rect 6281 -14194 6287 -14160
rect 6325 -14194 6349 -14160
rect 6349 -14194 6359 -14160
rect 6983 -14194 6993 -14160
rect 6993 -14194 7017 -14160
rect 7055 -14194 7061 -14160
rect 7061 -14194 7089 -14160
rect 7127 -14194 7129 -14160
rect 7129 -14194 7161 -14160
rect 7199 -14194 7231 -14160
rect 7231 -14194 7233 -14160
rect 7271 -14194 7299 -14160
rect 7299 -14194 7305 -14160
rect 7343 -14194 7367 -14160
rect 7367 -14194 7377 -14160
rect 8001 -14194 8011 -14160
rect 8011 -14194 8035 -14160
rect 8073 -14194 8079 -14160
rect 8079 -14194 8107 -14160
rect 8145 -14194 8147 -14160
rect 8147 -14194 8179 -14160
rect 8217 -14194 8249 -14160
rect 8249 -14194 8251 -14160
rect 8289 -14194 8317 -14160
rect 8317 -14194 8323 -14160
rect 8361 -14194 8385 -14160
rect 8385 -14194 8395 -14160
rect 9019 -14194 9029 -14160
rect 9029 -14194 9053 -14160
rect 9091 -14194 9097 -14160
rect 9097 -14194 9125 -14160
rect 9163 -14194 9165 -14160
rect 9165 -14194 9197 -14160
rect 9235 -14194 9267 -14160
rect 9267 -14194 9269 -14160
rect 9307 -14194 9335 -14160
rect 9335 -14194 9341 -14160
rect 9379 -14194 9403 -14160
rect 9403 -14194 9413 -14160
rect 10037 -14194 10047 -14160
rect 10047 -14194 10071 -14160
rect 10109 -14194 10115 -14160
rect 10115 -14194 10143 -14160
rect 10181 -14194 10183 -14160
rect 10183 -14194 10215 -14160
rect 10253 -14194 10285 -14160
rect 10285 -14194 10287 -14160
rect 10325 -14194 10353 -14160
rect 10353 -14194 10359 -14160
rect 10397 -14194 10421 -14160
rect 10421 -14194 10431 -14160
rect 11055 -14194 11065 -14160
rect 11065 -14194 11089 -14160
rect 11127 -14194 11133 -14160
rect 11133 -14194 11161 -14160
rect 11199 -14194 11201 -14160
rect 11201 -14194 11233 -14160
rect 11271 -14194 11303 -14160
rect 11303 -14194 11305 -14160
rect 11343 -14194 11371 -14160
rect 11371 -14194 11377 -14160
rect 11415 -14194 11439 -14160
rect 11439 -14194 11449 -14160
rect 12073 -14194 12083 -14160
rect 12083 -14194 12107 -14160
rect 12145 -14194 12151 -14160
rect 12151 -14194 12179 -14160
rect 12217 -14194 12219 -14160
rect 12219 -14194 12251 -14160
rect 12289 -14194 12321 -14160
rect 12321 -14194 12323 -14160
rect 12361 -14194 12389 -14160
rect 12389 -14194 12395 -14160
rect 12433 -14194 12457 -14160
rect 12457 -14194 12467 -14160
rect 13091 -14194 13101 -14160
rect 13101 -14194 13125 -14160
rect 13163 -14194 13169 -14160
rect 13169 -14194 13197 -14160
rect 13235 -14194 13237 -14160
rect 13237 -14194 13269 -14160
rect 13307 -14194 13339 -14160
rect 13339 -14194 13341 -14160
rect 13379 -14194 13407 -14160
rect 13407 -14194 13413 -14160
rect 13451 -14194 13475 -14160
rect 13475 -14194 13485 -14160
rect 14109 -14194 14119 -14160
rect 14119 -14194 14143 -14160
rect 14181 -14194 14187 -14160
rect 14187 -14194 14215 -14160
rect 14253 -14194 14255 -14160
rect 14255 -14194 14287 -14160
rect 14325 -14194 14357 -14160
rect 14357 -14194 14359 -14160
rect 14397 -14194 14425 -14160
rect 14425 -14194 14431 -14160
rect 14469 -14194 14493 -14160
rect 14493 -14194 14503 -14160
rect 15127 -14194 15137 -14160
rect 15137 -14194 15161 -14160
rect 15199 -14194 15205 -14160
rect 15205 -14194 15233 -14160
rect 15271 -14194 15273 -14160
rect 15273 -14194 15305 -14160
rect 15343 -14194 15375 -14160
rect 15375 -14194 15377 -14160
rect 15415 -14194 15443 -14160
rect 15443 -14194 15449 -14160
rect 15487 -14194 15511 -14160
rect 15511 -14194 15521 -14160
rect 16145 -14194 16155 -14160
rect 16155 -14194 16179 -14160
rect 16217 -14194 16223 -14160
rect 16223 -14194 16251 -14160
rect 16289 -14194 16291 -14160
rect 16291 -14194 16323 -14160
rect 16361 -14194 16393 -14160
rect 16393 -14194 16395 -14160
rect 16433 -14194 16461 -14160
rect 16461 -14194 16467 -14160
rect 16505 -14194 16529 -14160
rect 16529 -14194 16539 -14160
rect 17163 -14194 17173 -14160
rect 17173 -14194 17197 -14160
rect 17235 -14194 17241 -14160
rect 17241 -14194 17269 -14160
rect 17307 -14194 17309 -14160
rect 17309 -14194 17341 -14160
rect 17379 -14194 17411 -14160
rect 17411 -14194 17413 -14160
rect 17451 -14194 17479 -14160
rect 17479 -14194 17485 -14160
rect 17523 -14194 17547 -14160
rect 17547 -14194 17557 -14160
rect 18181 -14194 18191 -14160
rect 18191 -14194 18215 -14160
rect 18253 -14194 18259 -14160
rect 18259 -14194 18287 -14160
rect 18325 -14194 18327 -14160
rect 18327 -14194 18359 -14160
rect 18397 -14194 18429 -14160
rect 18429 -14194 18431 -14160
rect 18469 -14194 18497 -14160
rect 18497 -14194 18503 -14160
rect 18541 -14194 18565 -14160
rect 18565 -14194 18575 -14160
rect 19199 -14194 19209 -14160
rect 19209 -14194 19233 -14160
rect 19271 -14194 19277 -14160
rect 19277 -14194 19305 -14160
rect 19343 -14194 19345 -14160
rect 19345 -14194 19377 -14160
rect 19415 -14194 19447 -14160
rect 19447 -14194 19449 -14160
rect 19487 -14194 19515 -14160
rect 19515 -14194 19521 -14160
rect 19559 -14194 19583 -14160
rect 19583 -14194 19593 -14160
rect 20217 -14194 20227 -14160
rect 20227 -14194 20251 -14160
rect 20289 -14194 20295 -14160
rect 20295 -14194 20323 -14160
rect 20361 -14194 20363 -14160
rect 20363 -14194 20395 -14160
rect 20433 -14194 20465 -14160
rect 20465 -14194 20467 -14160
rect 20505 -14194 20533 -14160
rect 20533 -14194 20539 -14160
rect 20577 -14194 20601 -14160
rect 20601 -14194 20611 -14160
rect 21235 -14194 21245 -14160
rect 21245 -14194 21269 -14160
rect 21307 -14194 21313 -14160
rect 21313 -14194 21341 -14160
rect 21379 -14194 21381 -14160
rect 21381 -14194 21413 -14160
rect 21451 -14194 21483 -14160
rect 21483 -14194 21485 -14160
rect 21523 -14194 21551 -14160
rect 21551 -14194 21557 -14160
rect 21595 -14194 21619 -14160
rect 21619 -14194 21629 -14160
rect 22253 -14194 22263 -14160
rect 22263 -14194 22287 -14160
rect 22325 -14194 22331 -14160
rect 22331 -14194 22359 -14160
rect 22397 -14194 22399 -14160
rect 22399 -14194 22431 -14160
rect 22469 -14194 22501 -14160
rect 22501 -14194 22503 -14160
rect 22541 -14194 22569 -14160
rect 22569 -14194 22575 -14160
rect 22613 -14194 22637 -14160
rect 22637 -14194 22647 -14160
rect 24855 -14185 24889 -14179
rect 24855 -14213 24889 -14185
rect -22 -14261 12 -14251
rect -22 -14285 12 -14261
rect -22 -14329 12 -14323
rect -22 -14357 12 -14329
rect -22 -14397 12 -14395
rect -22 -14429 12 -14397
rect -22 -14499 12 -14467
rect -22 -14501 12 -14499
rect -22 -14567 12 -14539
rect -22 -14573 12 -14567
rect -22 -14635 12 -14611
rect -22 -14645 12 -14635
rect -22 -14703 12 -14683
rect -22 -14717 12 -14703
rect 2582 -14277 2616 -14263
rect 2582 -14297 2616 -14277
rect 2582 -14345 2616 -14335
rect 2582 -14369 2616 -14345
rect 2582 -14413 2616 -14407
rect 2582 -14441 2616 -14413
rect 2582 -14481 2616 -14479
rect 2582 -14513 2616 -14481
rect 2582 -14583 2616 -14551
rect 2582 -14585 2616 -14583
rect 2582 -14651 2616 -14623
rect 2582 -14657 2616 -14651
rect 2582 -14719 2616 -14695
rect 2582 -14729 2616 -14719
rect -12289 -14763 -12255 -14755
rect -12289 -14789 -12255 -14763
rect -8855 -14820 -8845 -14786
rect -8845 -14820 -8821 -14786
rect -8783 -14820 -8777 -14786
rect -8777 -14820 -8749 -14786
rect -8711 -14820 -8709 -14786
rect -8709 -14820 -8677 -14786
rect -8639 -14820 -8607 -14786
rect -8607 -14820 -8605 -14786
rect -8567 -14820 -8539 -14786
rect -8539 -14820 -8533 -14786
rect -8495 -14820 -8471 -14786
rect -8471 -14820 -8461 -14786
rect -7837 -14820 -7827 -14786
rect -7827 -14820 -7803 -14786
rect -7765 -14820 -7759 -14786
rect -7759 -14820 -7731 -14786
rect -7693 -14820 -7691 -14786
rect -7691 -14820 -7659 -14786
rect -7621 -14820 -7589 -14786
rect -7589 -14820 -7587 -14786
rect -7549 -14820 -7521 -14786
rect -7521 -14820 -7515 -14786
rect -7477 -14820 -7453 -14786
rect -7453 -14820 -7443 -14786
rect -6819 -14820 -6809 -14786
rect -6809 -14820 -6785 -14786
rect -6747 -14820 -6741 -14786
rect -6741 -14820 -6713 -14786
rect -6675 -14820 -6673 -14786
rect -6673 -14820 -6641 -14786
rect -6603 -14820 -6571 -14786
rect -6571 -14820 -6569 -14786
rect -6531 -14820 -6503 -14786
rect -6503 -14820 -6497 -14786
rect -6459 -14820 -6435 -14786
rect -6435 -14820 -6425 -14786
rect -5801 -14820 -5791 -14786
rect -5791 -14820 -5767 -14786
rect -5729 -14820 -5723 -14786
rect -5723 -14820 -5695 -14786
rect -5657 -14820 -5655 -14786
rect -5655 -14820 -5623 -14786
rect -5585 -14820 -5553 -14786
rect -5553 -14820 -5551 -14786
rect -5513 -14820 -5485 -14786
rect -5485 -14820 -5479 -14786
rect -5441 -14820 -5417 -14786
rect -5417 -14820 -5407 -14786
rect -4783 -14820 -4773 -14786
rect -4773 -14820 -4749 -14786
rect -4711 -14820 -4705 -14786
rect -4705 -14820 -4677 -14786
rect -4639 -14820 -4637 -14786
rect -4637 -14820 -4605 -14786
rect -4567 -14820 -4535 -14786
rect -4535 -14820 -4533 -14786
rect -4495 -14820 -4467 -14786
rect -4467 -14820 -4461 -14786
rect -4423 -14820 -4399 -14786
rect -4399 -14820 -4389 -14786
rect -3765 -14820 -3755 -14786
rect -3755 -14820 -3731 -14786
rect -3693 -14820 -3687 -14786
rect -3687 -14820 -3659 -14786
rect -3621 -14820 -3619 -14786
rect -3619 -14820 -3587 -14786
rect -3549 -14820 -3517 -14786
rect -3517 -14820 -3515 -14786
rect -3477 -14820 -3449 -14786
rect -3449 -14820 -3443 -14786
rect -3405 -14820 -3381 -14786
rect -3381 -14820 -3371 -14786
rect -2747 -14820 -2737 -14786
rect -2737 -14820 -2713 -14786
rect -2675 -14820 -2669 -14786
rect -2669 -14820 -2641 -14786
rect -2603 -14820 -2601 -14786
rect -2601 -14820 -2569 -14786
rect -2531 -14820 -2499 -14786
rect -2499 -14820 -2497 -14786
rect -2459 -14820 -2431 -14786
rect -2431 -14820 -2425 -14786
rect -2387 -14820 -2363 -14786
rect -2363 -14820 -2353 -14786
rect -1729 -14820 -1719 -14786
rect -1719 -14820 -1695 -14786
rect -1657 -14820 -1651 -14786
rect -1651 -14820 -1623 -14786
rect -1585 -14820 -1583 -14786
rect -1583 -14820 -1551 -14786
rect -1513 -14820 -1481 -14786
rect -1481 -14820 -1479 -14786
rect -1441 -14820 -1413 -14786
rect -1413 -14820 -1407 -14786
rect -1369 -14820 -1345 -14786
rect -1345 -14820 -1335 -14786
rect -711 -14820 -701 -14786
rect -701 -14820 -677 -14786
rect -639 -14820 -633 -14786
rect -633 -14820 -605 -14786
rect -567 -14820 -565 -14786
rect -565 -14820 -533 -14786
rect -495 -14820 -463 -14786
rect -463 -14820 -461 -14786
rect -423 -14820 -395 -14786
rect -395 -14820 -389 -14786
rect -351 -14820 -327 -14786
rect -327 -14820 -317 -14786
rect 2582 -14787 2616 -14767
rect 2582 -14801 2616 -14787
rect -12289 -14831 -12255 -14827
rect -12289 -14861 -12255 -14831
rect 3600 -14277 3634 -14263
rect 3600 -14297 3634 -14277
rect 3600 -14345 3634 -14335
rect 3600 -14369 3634 -14345
rect 3600 -14413 3634 -14407
rect 3600 -14441 3634 -14413
rect 3600 -14481 3634 -14479
rect 3600 -14513 3634 -14481
rect 3600 -14583 3634 -14551
rect 3600 -14585 3634 -14583
rect 3600 -14651 3634 -14623
rect 3600 -14657 3634 -14651
rect 3600 -14719 3634 -14695
rect 3600 -14729 3634 -14719
rect 3600 -14787 3634 -14767
rect 3600 -14801 3634 -14787
rect 4618 -14277 4652 -14263
rect 4618 -14297 4652 -14277
rect 4618 -14345 4652 -14335
rect 4618 -14369 4652 -14345
rect 4618 -14413 4652 -14407
rect 4618 -14441 4652 -14413
rect 4618 -14481 4652 -14479
rect 4618 -14513 4652 -14481
rect 4618 -14583 4652 -14551
rect 4618 -14585 4652 -14583
rect 4618 -14651 4652 -14623
rect 4618 -14657 4652 -14651
rect 4618 -14719 4652 -14695
rect 4618 -14729 4652 -14719
rect 4618 -14787 4652 -14767
rect 4618 -14801 4652 -14787
rect 5636 -14277 5670 -14263
rect 5636 -14297 5670 -14277
rect 5636 -14345 5670 -14335
rect 5636 -14369 5670 -14345
rect 5636 -14413 5670 -14407
rect 5636 -14441 5670 -14413
rect 5636 -14481 5670 -14479
rect 5636 -14513 5670 -14481
rect 5636 -14583 5670 -14551
rect 5636 -14585 5670 -14583
rect 5636 -14651 5670 -14623
rect 5636 -14657 5670 -14651
rect 5636 -14719 5670 -14695
rect 5636 -14729 5670 -14719
rect 5636 -14787 5670 -14767
rect 5636 -14801 5670 -14787
rect 6654 -14277 6688 -14263
rect 6654 -14297 6688 -14277
rect 6654 -14345 6688 -14335
rect 6654 -14369 6688 -14345
rect 6654 -14413 6688 -14407
rect 6654 -14441 6688 -14413
rect 6654 -14481 6688 -14479
rect 6654 -14513 6688 -14481
rect 6654 -14583 6688 -14551
rect 6654 -14585 6688 -14583
rect 6654 -14651 6688 -14623
rect 6654 -14657 6688 -14651
rect 6654 -14719 6688 -14695
rect 6654 -14729 6688 -14719
rect 6654 -14787 6688 -14767
rect 6654 -14801 6688 -14787
rect 7672 -14277 7706 -14263
rect 7672 -14297 7706 -14277
rect 7672 -14345 7706 -14335
rect 7672 -14369 7706 -14345
rect 7672 -14413 7706 -14407
rect 7672 -14441 7706 -14413
rect 7672 -14481 7706 -14479
rect 7672 -14513 7706 -14481
rect 7672 -14583 7706 -14551
rect 7672 -14585 7706 -14583
rect 7672 -14651 7706 -14623
rect 7672 -14657 7706 -14651
rect 7672 -14719 7706 -14695
rect 7672 -14729 7706 -14719
rect 7672 -14787 7706 -14767
rect 7672 -14801 7706 -14787
rect 8690 -14277 8724 -14263
rect 8690 -14297 8724 -14277
rect 8690 -14345 8724 -14335
rect 8690 -14369 8724 -14345
rect 8690 -14413 8724 -14407
rect 8690 -14441 8724 -14413
rect 8690 -14481 8724 -14479
rect 8690 -14513 8724 -14481
rect 8690 -14583 8724 -14551
rect 8690 -14585 8724 -14583
rect 8690 -14651 8724 -14623
rect 8690 -14657 8724 -14651
rect 8690 -14719 8724 -14695
rect 8690 -14729 8724 -14719
rect 8690 -14787 8724 -14767
rect 8690 -14801 8724 -14787
rect 9708 -14277 9742 -14263
rect 9708 -14297 9742 -14277
rect 9708 -14345 9742 -14335
rect 9708 -14369 9742 -14345
rect 9708 -14413 9742 -14407
rect 9708 -14441 9742 -14413
rect 9708 -14481 9742 -14479
rect 9708 -14513 9742 -14481
rect 9708 -14583 9742 -14551
rect 9708 -14585 9742 -14583
rect 9708 -14651 9742 -14623
rect 9708 -14657 9742 -14651
rect 9708 -14719 9742 -14695
rect 9708 -14729 9742 -14719
rect 9708 -14787 9742 -14767
rect 9708 -14801 9742 -14787
rect 10726 -14277 10760 -14263
rect 10726 -14297 10760 -14277
rect 10726 -14345 10760 -14335
rect 10726 -14369 10760 -14345
rect 10726 -14413 10760 -14407
rect 10726 -14441 10760 -14413
rect 10726 -14481 10760 -14479
rect 10726 -14513 10760 -14481
rect 10726 -14583 10760 -14551
rect 10726 -14585 10760 -14583
rect 10726 -14651 10760 -14623
rect 10726 -14657 10760 -14651
rect 10726 -14719 10760 -14695
rect 10726 -14729 10760 -14719
rect 10726 -14787 10760 -14767
rect 10726 -14801 10760 -14787
rect 11744 -14277 11778 -14263
rect 11744 -14297 11778 -14277
rect 11744 -14345 11778 -14335
rect 11744 -14369 11778 -14345
rect 11744 -14413 11778 -14407
rect 11744 -14441 11778 -14413
rect 11744 -14481 11778 -14479
rect 11744 -14513 11778 -14481
rect 11744 -14583 11778 -14551
rect 11744 -14585 11778 -14583
rect 11744 -14651 11778 -14623
rect 11744 -14657 11778 -14651
rect 11744 -14719 11778 -14695
rect 11744 -14729 11778 -14719
rect 11744 -14787 11778 -14767
rect 11744 -14801 11778 -14787
rect 12762 -14277 12796 -14263
rect 12762 -14297 12796 -14277
rect 12762 -14345 12796 -14335
rect 12762 -14369 12796 -14345
rect 12762 -14413 12796 -14407
rect 12762 -14441 12796 -14413
rect 12762 -14481 12796 -14479
rect 12762 -14513 12796 -14481
rect 12762 -14583 12796 -14551
rect 12762 -14585 12796 -14583
rect 12762 -14651 12796 -14623
rect 12762 -14657 12796 -14651
rect 12762 -14719 12796 -14695
rect 12762 -14729 12796 -14719
rect 12762 -14787 12796 -14767
rect 12762 -14801 12796 -14787
rect 13780 -14277 13814 -14263
rect 13780 -14297 13814 -14277
rect 13780 -14345 13814 -14335
rect 13780 -14369 13814 -14345
rect 13780 -14413 13814 -14407
rect 13780 -14441 13814 -14413
rect 13780 -14481 13814 -14479
rect 13780 -14513 13814 -14481
rect 13780 -14583 13814 -14551
rect 13780 -14585 13814 -14583
rect 13780 -14651 13814 -14623
rect 13780 -14657 13814 -14651
rect 13780 -14719 13814 -14695
rect 13780 -14729 13814 -14719
rect 13780 -14787 13814 -14767
rect 13780 -14801 13814 -14787
rect 14798 -14277 14832 -14263
rect 14798 -14297 14832 -14277
rect 14798 -14345 14832 -14335
rect 14798 -14369 14832 -14345
rect 14798 -14413 14832 -14407
rect 14798 -14441 14832 -14413
rect 14798 -14481 14832 -14479
rect 14798 -14513 14832 -14481
rect 14798 -14583 14832 -14551
rect 14798 -14585 14832 -14583
rect 14798 -14651 14832 -14623
rect 14798 -14657 14832 -14651
rect 14798 -14719 14832 -14695
rect 14798 -14729 14832 -14719
rect 14798 -14787 14832 -14767
rect 14798 -14801 14832 -14787
rect 15816 -14277 15850 -14263
rect 15816 -14297 15850 -14277
rect 15816 -14345 15850 -14335
rect 15816 -14369 15850 -14345
rect 15816 -14413 15850 -14407
rect 15816 -14441 15850 -14413
rect 15816 -14481 15850 -14479
rect 15816 -14513 15850 -14481
rect 15816 -14583 15850 -14551
rect 15816 -14585 15850 -14583
rect 15816 -14651 15850 -14623
rect 15816 -14657 15850 -14651
rect 15816 -14719 15850 -14695
rect 15816 -14729 15850 -14719
rect 15816 -14787 15850 -14767
rect 15816 -14801 15850 -14787
rect 16834 -14277 16868 -14263
rect 16834 -14297 16868 -14277
rect 16834 -14345 16868 -14335
rect 16834 -14369 16868 -14345
rect 16834 -14413 16868 -14407
rect 16834 -14441 16868 -14413
rect 16834 -14481 16868 -14479
rect 16834 -14513 16868 -14481
rect 16834 -14583 16868 -14551
rect 16834 -14585 16868 -14583
rect 16834 -14651 16868 -14623
rect 16834 -14657 16868 -14651
rect 16834 -14719 16868 -14695
rect 16834 -14729 16868 -14719
rect 16834 -14787 16868 -14767
rect 16834 -14801 16868 -14787
rect 17852 -14277 17886 -14263
rect 17852 -14297 17886 -14277
rect 17852 -14345 17886 -14335
rect 17852 -14369 17886 -14345
rect 17852 -14413 17886 -14407
rect 17852 -14441 17886 -14413
rect 17852 -14481 17886 -14479
rect 17852 -14513 17886 -14481
rect 17852 -14583 17886 -14551
rect 17852 -14585 17886 -14583
rect 17852 -14651 17886 -14623
rect 17852 -14657 17886 -14651
rect 17852 -14719 17886 -14695
rect 17852 -14729 17886 -14719
rect 17852 -14787 17886 -14767
rect 17852 -14801 17886 -14787
rect 18870 -14277 18904 -14263
rect 18870 -14297 18904 -14277
rect 18870 -14345 18904 -14335
rect 18870 -14369 18904 -14345
rect 18870 -14413 18904 -14407
rect 18870 -14441 18904 -14413
rect 18870 -14481 18904 -14479
rect 18870 -14513 18904 -14481
rect 18870 -14583 18904 -14551
rect 18870 -14585 18904 -14583
rect 18870 -14651 18904 -14623
rect 18870 -14657 18904 -14651
rect 18870 -14719 18904 -14695
rect 18870 -14729 18904 -14719
rect 18870 -14787 18904 -14767
rect 18870 -14801 18904 -14787
rect 19888 -14277 19922 -14263
rect 19888 -14297 19922 -14277
rect 19888 -14345 19922 -14335
rect 19888 -14369 19922 -14345
rect 19888 -14413 19922 -14407
rect 19888 -14441 19922 -14413
rect 19888 -14481 19922 -14479
rect 19888 -14513 19922 -14481
rect 19888 -14583 19922 -14551
rect 19888 -14585 19922 -14583
rect 19888 -14651 19922 -14623
rect 19888 -14657 19922 -14651
rect 19888 -14719 19922 -14695
rect 19888 -14729 19922 -14719
rect 19888 -14787 19922 -14767
rect 19888 -14801 19922 -14787
rect 20906 -14277 20940 -14263
rect 20906 -14297 20940 -14277
rect 20906 -14345 20940 -14335
rect 20906 -14369 20940 -14345
rect 20906 -14413 20940 -14407
rect 20906 -14441 20940 -14413
rect 20906 -14481 20940 -14479
rect 20906 -14513 20940 -14481
rect 20906 -14583 20940 -14551
rect 20906 -14585 20940 -14583
rect 20906 -14651 20940 -14623
rect 20906 -14657 20940 -14651
rect 20906 -14719 20940 -14695
rect 20906 -14729 20940 -14719
rect 20906 -14787 20940 -14767
rect 20906 -14801 20940 -14787
rect 21924 -14277 21958 -14263
rect 21924 -14297 21958 -14277
rect 21924 -14345 21958 -14335
rect 21924 -14369 21958 -14345
rect 21924 -14413 21958 -14407
rect 21924 -14441 21958 -14413
rect 21924 -14481 21958 -14479
rect 21924 -14513 21958 -14481
rect 21924 -14583 21958 -14551
rect 21924 -14585 21958 -14583
rect 21924 -14651 21958 -14623
rect 21924 -14657 21958 -14651
rect 21924 -14719 21958 -14695
rect 21924 -14729 21958 -14719
rect 21924 -14787 21958 -14767
rect 21924 -14801 21958 -14787
rect 22942 -14277 22976 -14263
rect 22942 -14297 22976 -14277
rect 22942 -14345 22976 -14335
rect 22942 -14369 22976 -14345
rect 22942 -14413 22976 -14407
rect 22942 -14441 22976 -14413
rect 22942 -14481 22976 -14479
rect 22942 -14513 22976 -14481
rect 22942 -14583 22976 -14551
rect 22942 -14585 22976 -14583
rect 22942 -14651 22976 -14623
rect 22942 -14657 22976 -14651
rect 22942 -14719 22976 -14695
rect 22942 -14729 22976 -14719
rect 22942 -14787 22976 -14767
rect 22942 -14801 22976 -14787
rect 24855 -14253 24889 -14251
rect 24855 -14285 24889 -14253
rect 24855 -14355 24889 -14323
rect 24855 -14357 24889 -14355
rect 24855 -14423 24889 -14395
rect 24855 -14429 24889 -14423
rect 24855 -14491 24889 -14467
rect 24855 -14501 24889 -14491
rect 24855 -14559 24889 -14539
rect 24855 -14573 24889 -14559
rect 24855 -14627 24889 -14611
rect 24855 -14645 24889 -14627
rect 24855 -14695 24889 -14683
rect 24855 -14717 24889 -14695
rect 24855 -14763 24889 -14755
rect 24855 -14789 24889 -14763
rect 24855 -14831 24889 -14827
rect 24855 -14861 24889 -14831
rect -12289 -14933 -12255 -14899
rect -8855 -14928 -8845 -14894
rect -8845 -14928 -8821 -14894
rect -8783 -14928 -8777 -14894
rect -8777 -14928 -8749 -14894
rect -8711 -14928 -8709 -14894
rect -8709 -14928 -8677 -14894
rect -8639 -14928 -8607 -14894
rect -8607 -14928 -8605 -14894
rect -8567 -14928 -8539 -14894
rect -8539 -14928 -8533 -14894
rect -8495 -14928 -8471 -14894
rect -8471 -14928 -8461 -14894
rect -7837 -14928 -7827 -14894
rect -7827 -14928 -7803 -14894
rect -7765 -14928 -7759 -14894
rect -7759 -14928 -7731 -14894
rect -7693 -14928 -7691 -14894
rect -7691 -14928 -7659 -14894
rect -7621 -14928 -7589 -14894
rect -7589 -14928 -7587 -14894
rect -7549 -14928 -7521 -14894
rect -7521 -14928 -7515 -14894
rect -7477 -14928 -7453 -14894
rect -7453 -14928 -7443 -14894
rect -6819 -14928 -6809 -14894
rect -6809 -14928 -6785 -14894
rect -6747 -14928 -6741 -14894
rect -6741 -14928 -6713 -14894
rect -6675 -14928 -6673 -14894
rect -6673 -14928 -6641 -14894
rect -6603 -14928 -6571 -14894
rect -6571 -14928 -6569 -14894
rect -6531 -14928 -6503 -14894
rect -6503 -14928 -6497 -14894
rect -6459 -14928 -6435 -14894
rect -6435 -14928 -6425 -14894
rect -5801 -14928 -5791 -14894
rect -5791 -14928 -5767 -14894
rect -5729 -14928 -5723 -14894
rect -5723 -14928 -5695 -14894
rect -5657 -14928 -5655 -14894
rect -5655 -14928 -5623 -14894
rect -5585 -14928 -5553 -14894
rect -5553 -14928 -5551 -14894
rect -5513 -14928 -5485 -14894
rect -5485 -14928 -5479 -14894
rect -5441 -14928 -5417 -14894
rect -5417 -14928 -5407 -14894
rect -4783 -14928 -4773 -14894
rect -4773 -14928 -4749 -14894
rect -4711 -14928 -4705 -14894
rect -4705 -14928 -4677 -14894
rect -4639 -14928 -4637 -14894
rect -4637 -14928 -4605 -14894
rect -4567 -14928 -4535 -14894
rect -4535 -14928 -4533 -14894
rect -4495 -14928 -4467 -14894
rect -4467 -14928 -4461 -14894
rect -4423 -14928 -4399 -14894
rect -4399 -14928 -4389 -14894
rect -3765 -14928 -3755 -14894
rect -3755 -14928 -3731 -14894
rect -3693 -14928 -3687 -14894
rect -3687 -14928 -3659 -14894
rect -3621 -14928 -3619 -14894
rect -3619 -14928 -3587 -14894
rect -3549 -14928 -3517 -14894
rect -3517 -14928 -3515 -14894
rect -3477 -14928 -3449 -14894
rect -3449 -14928 -3443 -14894
rect -3405 -14928 -3381 -14894
rect -3381 -14928 -3371 -14894
rect -2747 -14928 -2737 -14894
rect -2737 -14928 -2713 -14894
rect -2675 -14928 -2669 -14894
rect -2669 -14928 -2641 -14894
rect -2603 -14928 -2601 -14894
rect -2601 -14928 -2569 -14894
rect -2531 -14928 -2499 -14894
rect -2499 -14928 -2497 -14894
rect -2459 -14928 -2431 -14894
rect -2431 -14928 -2425 -14894
rect -2387 -14928 -2363 -14894
rect -2363 -14928 -2353 -14894
rect -1729 -14928 -1719 -14894
rect -1719 -14928 -1695 -14894
rect -1657 -14928 -1651 -14894
rect -1651 -14928 -1623 -14894
rect -1585 -14928 -1583 -14894
rect -1583 -14928 -1551 -14894
rect -1513 -14928 -1481 -14894
rect -1481 -14928 -1479 -14894
rect -1441 -14928 -1413 -14894
rect -1413 -14928 -1407 -14894
rect -1369 -14928 -1345 -14894
rect -1345 -14928 -1335 -14894
rect -711 -14928 -701 -14894
rect -701 -14928 -677 -14894
rect -639 -14928 -633 -14894
rect -633 -14928 -605 -14894
rect -567 -14928 -565 -14894
rect -565 -14928 -533 -14894
rect -495 -14928 -463 -14894
rect -463 -14928 -461 -14894
rect -423 -14928 -395 -14894
rect -395 -14928 -389 -14894
rect -351 -14928 -327 -14894
rect -327 -14928 -317 -14894
rect 2911 -14904 2921 -14870
rect 2921 -14904 2945 -14870
rect 2983 -14904 2989 -14870
rect 2989 -14904 3017 -14870
rect 3055 -14904 3057 -14870
rect 3057 -14904 3089 -14870
rect 3127 -14904 3159 -14870
rect 3159 -14904 3161 -14870
rect 3199 -14904 3227 -14870
rect 3227 -14904 3233 -14870
rect 3271 -14904 3295 -14870
rect 3295 -14904 3305 -14870
rect 3929 -14904 3939 -14870
rect 3939 -14904 3963 -14870
rect 4001 -14904 4007 -14870
rect 4007 -14904 4035 -14870
rect 4073 -14904 4075 -14870
rect 4075 -14904 4107 -14870
rect 4145 -14904 4177 -14870
rect 4177 -14904 4179 -14870
rect 4217 -14904 4245 -14870
rect 4245 -14904 4251 -14870
rect 4289 -14904 4313 -14870
rect 4313 -14904 4323 -14870
rect 4947 -14904 4957 -14870
rect 4957 -14904 4981 -14870
rect 5019 -14904 5025 -14870
rect 5025 -14904 5053 -14870
rect 5091 -14904 5093 -14870
rect 5093 -14904 5125 -14870
rect 5163 -14904 5195 -14870
rect 5195 -14904 5197 -14870
rect 5235 -14904 5263 -14870
rect 5263 -14904 5269 -14870
rect 5307 -14904 5331 -14870
rect 5331 -14904 5341 -14870
rect 5965 -14904 5975 -14870
rect 5975 -14904 5999 -14870
rect 6037 -14904 6043 -14870
rect 6043 -14904 6071 -14870
rect 6109 -14904 6111 -14870
rect 6111 -14904 6143 -14870
rect 6181 -14904 6213 -14870
rect 6213 -14904 6215 -14870
rect 6253 -14904 6281 -14870
rect 6281 -14904 6287 -14870
rect 6325 -14904 6349 -14870
rect 6349 -14904 6359 -14870
rect 6983 -14904 6993 -14870
rect 6993 -14904 7017 -14870
rect 7055 -14904 7061 -14870
rect 7061 -14904 7089 -14870
rect 7127 -14904 7129 -14870
rect 7129 -14904 7161 -14870
rect 7199 -14904 7231 -14870
rect 7231 -14904 7233 -14870
rect 7271 -14904 7299 -14870
rect 7299 -14904 7305 -14870
rect 7343 -14904 7367 -14870
rect 7367 -14904 7377 -14870
rect 8001 -14904 8011 -14870
rect 8011 -14904 8035 -14870
rect 8073 -14904 8079 -14870
rect 8079 -14904 8107 -14870
rect 8145 -14904 8147 -14870
rect 8147 -14904 8179 -14870
rect 8217 -14904 8249 -14870
rect 8249 -14904 8251 -14870
rect 8289 -14904 8317 -14870
rect 8317 -14904 8323 -14870
rect 8361 -14904 8385 -14870
rect 8385 -14904 8395 -14870
rect 9019 -14904 9029 -14870
rect 9029 -14904 9053 -14870
rect 9091 -14904 9097 -14870
rect 9097 -14904 9125 -14870
rect 9163 -14904 9165 -14870
rect 9165 -14904 9197 -14870
rect 9235 -14904 9267 -14870
rect 9267 -14904 9269 -14870
rect 9307 -14904 9335 -14870
rect 9335 -14904 9341 -14870
rect 9379 -14904 9403 -14870
rect 9403 -14904 9413 -14870
rect 10037 -14904 10047 -14870
rect 10047 -14904 10071 -14870
rect 10109 -14904 10115 -14870
rect 10115 -14904 10143 -14870
rect 10181 -14904 10183 -14870
rect 10183 -14904 10215 -14870
rect 10253 -14904 10285 -14870
rect 10285 -14904 10287 -14870
rect 10325 -14904 10353 -14870
rect 10353 -14904 10359 -14870
rect 10397 -14904 10421 -14870
rect 10421 -14904 10431 -14870
rect 11055 -14904 11065 -14870
rect 11065 -14904 11089 -14870
rect 11127 -14904 11133 -14870
rect 11133 -14904 11161 -14870
rect 11199 -14904 11201 -14870
rect 11201 -14904 11233 -14870
rect 11271 -14904 11303 -14870
rect 11303 -14904 11305 -14870
rect 11343 -14904 11371 -14870
rect 11371 -14904 11377 -14870
rect 11415 -14904 11439 -14870
rect 11439 -14904 11449 -14870
rect 12073 -14904 12083 -14870
rect 12083 -14904 12107 -14870
rect 12145 -14904 12151 -14870
rect 12151 -14904 12179 -14870
rect 12217 -14904 12219 -14870
rect 12219 -14904 12251 -14870
rect 12289 -14904 12321 -14870
rect 12321 -14904 12323 -14870
rect 12361 -14904 12389 -14870
rect 12389 -14904 12395 -14870
rect 12433 -14904 12457 -14870
rect 12457 -14904 12467 -14870
rect 13091 -14904 13101 -14870
rect 13101 -14904 13125 -14870
rect 13163 -14904 13169 -14870
rect 13169 -14904 13197 -14870
rect 13235 -14904 13237 -14870
rect 13237 -14904 13269 -14870
rect 13307 -14904 13339 -14870
rect 13339 -14904 13341 -14870
rect 13379 -14904 13407 -14870
rect 13407 -14904 13413 -14870
rect 13451 -14904 13475 -14870
rect 13475 -14904 13485 -14870
rect 14109 -14904 14119 -14870
rect 14119 -14904 14143 -14870
rect 14181 -14904 14187 -14870
rect 14187 -14904 14215 -14870
rect 14253 -14904 14255 -14870
rect 14255 -14904 14287 -14870
rect 14325 -14904 14357 -14870
rect 14357 -14904 14359 -14870
rect 14397 -14904 14425 -14870
rect 14425 -14904 14431 -14870
rect 14469 -14904 14493 -14870
rect 14493 -14904 14503 -14870
rect 15127 -14904 15137 -14870
rect 15137 -14904 15161 -14870
rect 15199 -14904 15205 -14870
rect 15205 -14904 15233 -14870
rect 15271 -14904 15273 -14870
rect 15273 -14904 15305 -14870
rect 15343 -14904 15375 -14870
rect 15375 -14904 15377 -14870
rect 15415 -14904 15443 -14870
rect 15443 -14904 15449 -14870
rect 15487 -14904 15511 -14870
rect 15511 -14904 15521 -14870
rect 16145 -14904 16155 -14870
rect 16155 -14904 16179 -14870
rect 16217 -14904 16223 -14870
rect 16223 -14904 16251 -14870
rect 16289 -14904 16291 -14870
rect 16291 -14904 16323 -14870
rect 16361 -14904 16393 -14870
rect 16393 -14904 16395 -14870
rect 16433 -14904 16461 -14870
rect 16461 -14904 16467 -14870
rect 16505 -14904 16529 -14870
rect 16529 -14904 16539 -14870
rect 17163 -14904 17173 -14870
rect 17173 -14904 17197 -14870
rect 17235 -14904 17241 -14870
rect 17241 -14904 17269 -14870
rect 17307 -14904 17309 -14870
rect 17309 -14904 17341 -14870
rect 17379 -14904 17411 -14870
rect 17411 -14904 17413 -14870
rect 17451 -14904 17479 -14870
rect 17479 -14904 17485 -14870
rect 17523 -14904 17547 -14870
rect 17547 -14904 17557 -14870
rect 18181 -14904 18191 -14870
rect 18191 -14904 18215 -14870
rect 18253 -14904 18259 -14870
rect 18259 -14904 18287 -14870
rect 18325 -14904 18327 -14870
rect 18327 -14904 18359 -14870
rect 18397 -14904 18429 -14870
rect 18429 -14904 18431 -14870
rect 18469 -14904 18497 -14870
rect 18497 -14904 18503 -14870
rect 18541 -14904 18565 -14870
rect 18565 -14904 18575 -14870
rect 19199 -14904 19209 -14870
rect 19209 -14904 19233 -14870
rect 19271 -14904 19277 -14870
rect 19277 -14904 19305 -14870
rect 19343 -14904 19345 -14870
rect 19345 -14904 19377 -14870
rect 19415 -14904 19447 -14870
rect 19447 -14904 19449 -14870
rect 19487 -14904 19515 -14870
rect 19515 -14904 19521 -14870
rect 19559 -14904 19583 -14870
rect 19583 -14904 19593 -14870
rect 20217 -14904 20227 -14870
rect 20227 -14904 20251 -14870
rect 20289 -14904 20295 -14870
rect 20295 -14904 20323 -14870
rect 20361 -14904 20363 -14870
rect 20363 -14904 20395 -14870
rect 20433 -14904 20465 -14870
rect 20465 -14904 20467 -14870
rect 20505 -14904 20533 -14870
rect 20533 -14904 20539 -14870
rect 20577 -14904 20601 -14870
rect 20601 -14904 20611 -14870
rect 21235 -14904 21245 -14870
rect 21245 -14904 21269 -14870
rect 21307 -14904 21313 -14870
rect 21313 -14904 21341 -14870
rect 21379 -14904 21381 -14870
rect 21381 -14904 21413 -14870
rect 21451 -14904 21483 -14870
rect 21483 -14904 21485 -14870
rect 21523 -14904 21551 -14870
rect 21551 -14904 21557 -14870
rect 21595 -14904 21619 -14870
rect 21619 -14904 21629 -14870
rect 22253 -14904 22263 -14870
rect 22263 -14904 22287 -14870
rect 22325 -14904 22331 -14870
rect 22331 -14904 22359 -14870
rect 22397 -14904 22399 -14870
rect 22399 -14904 22431 -14870
rect 22469 -14904 22501 -14870
rect 22501 -14904 22503 -14870
rect 22541 -14904 22569 -14870
rect 22569 -14904 22575 -14870
rect 22613 -14904 22637 -14870
rect 22637 -14904 22647 -14870
rect 24855 -14933 24889 -14899
rect -12289 -15001 -12255 -14971
rect -12289 -15005 -12255 -15001
rect -12289 -15069 -12255 -15043
rect -12289 -15077 -12255 -15069
rect -12289 -15137 -12255 -15115
rect -12289 -15149 -12255 -15137
rect -12289 -15205 -12255 -15187
rect -12289 -15221 -12255 -15205
rect -12289 -15273 -12255 -15259
rect -12289 -15293 -12255 -15273
rect -12289 -15341 -12255 -15331
rect -12289 -15365 -12255 -15341
rect -12289 -15409 -12255 -15403
rect -12289 -15437 -12255 -15409
rect -12289 -15477 -12255 -15475
rect -12289 -15509 -12255 -15477
rect -12289 -15579 -12255 -15547
rect -12289 -15581 -12255 -15579
rect -9184 -15011 -9150 -14997
rect -9184 -15031 -9150 -15011
rect -9184 -15079 -9150 -15069
rect -9184 -15103 -9150 -15079
rect -9184 -15147 -9150 -15141
rect -9184 -15175 -9150 -15147
rect -9184 -15215 -9150 -15213
rect -9184 -15247 -9150 -15215
rect -9184 -15317 -9150 -15285
rect -9184 -15319 -9150 -15317
rect -9184 -15385 -9150 -15357
rect -9184 -15391 -9150 -15385
rect -9184 -15453 -9150 -15429
rect -9184 -15463 -9150 -15453
rect -9184 -15521 -9150 -15501
rect -9184 -15535 -9150 -15521
rect -8166 -15011 -8132 -14997
rect -8166 -15031 -8132 -15011
rect -8166 -15079 -8132 -15069
rect -8166 -15103 -8132 -15079
rect -8166 -15147 -8132 -15141
rect -8166 -15175 -8132 -15147
rect -8166 -15215 -8132 -15213
rect -8166 -15247 -8132 -15215
rect -8166 -15317 -8132 -15285
rect -8166 -15319 -8132 -15317
rect -8166 -15385 -8132 -15357
rect -8166 -15391 -8132 -15385
rect -8166 -15453 -8132 -15429
rect -8166 -15463 -8132 -15453
rect -8166 -15521 -8132 -15501
rect -8166 -15535 -8132 -15521
rect -7148 -15011 -7114 -14997
rect -7148 -15031 -7114 -15011
rect -7148 -15079 -7114 -15069
rect -7148 -15103 -7114 -15079
rect -7148 -15147 -7114 -15141
rect -7148 -15175 -7114 -15147
rect -7148 -15215 -7114 -15213
rect -7148 -15247 -7114 -15215
rect -7148 -15317 -7114 -15285
rect -7148 -15319 -7114 -15317
rect -7148 -15385 -7114 -15357
rect -7148 -15391 -7114 -15385
rect -7148 -15453 -7114 -15429
rect -7148 -15463 -7114 -15453
rect -7148 -15521 -7114 -15501
rect -7148 -15535 -7114 -15521
rect -6130 -15011 -6096 -14997
rect -6130 -15031 -6096 -15011
rect -6130 -15079 -6096 -15069
rect -6130 -15103 -6096 -15079
rect -6130 -15147 -6096 -15141
rect -6130 -15175 -6096 -15147
rect -6130 -15215 -6096 -15213
rect -6130 -15247 -6096 -15215
rect -6130 -15317 -6096 -15285
rect -6130 -15319 -6096 -15317
rect -6130 -15385 -6096 -15357
rect -6130 -15391 -6096 -15385
rect -6130 -15453 -6096 -15429
rect -6130 -15463 -6096 -15453
rect -6130 -15521 -6096 -15501
rect -6130 -15535 -6096 -15521
rect -5112 -15011 -5078 -14997
rect -5112 -15031 -5078 -15011
rect -5112 -15079 -5078 -15069
rect -5112 -15103 -5078 -15079
rect -5112 -15147 -5078 -15141
rect -5112 -15175 -5078 -15147
rect -5112 -15215 -5078 -15213
rect -5112 -15247 -5078 -15215
rect -5112 -15317 -5078 -15285
rect -5112 -15319 -5078 -15317
rect -5112 -15385 -5078 -15357
rect -5112 -15391 -5078 -15385
rect -5112 -15453 -5078 -15429
rect -5112 -15463 -5078 -15453
rect -5112 -15521 -5078 -15501
rect -5112 -15535 -5078 -15521
rect -4094 -15011 -4060 -14997
rect -4094 -15031 -4060 -15011
rect -4094 -15079 -4060 -15069
rect -4094 -15103 -4060 -15079
rect -4094 -15147 -4060 -15141
rect -4094 -15175 -4060 -15147
rect -4094 -15215 -4060 -15213
rect -4094 -15247 -4060 -15215
rect -4094 -15317 -4060 -15285
rect -4094 -15319 -4060 -15317
rect -4094 -15385 -4060 -15357
rect -4094 -15391 -4060 -15385
rect -4094 -15453 -4060 -15429
rect -4094 -15463 -4060 -15453
rect -4094 -15521 -4060 -15501
rect -4094 -15535 -4060 -15521
rect -3076 -15011 -3042 -14997
rect -3076 -15031 -3042 -15011
rect -3076 -15079 -3042 -15069
rect -3076 -15103 -3042 -15079
rect -3076 -15147 -3042 -15141
rect -3076 -15175 -3042 -15147
rect -3076 -15215 -3042 -15213
rect -3076 -15247 -3042 -15215
rect -3076 -15317 -3042 -15285
rect -3076 -15319 -3042 -15317
rect -3076 -15385 -3042 -15357
rect -3076 -15391 -3042 -15385
rect -3076 -15453 -3042 -15429
rect -3076 -15463 -3042 -15453
rect -3076 -15521 -3042 -15501
rect -3076 -15535 -3042 -15521
rect -2058 -15011 -2024 -14997
rect -2058 -15031 -2024 -15011
rect -2058 -15079 -2024 -15069
rect -2058 -15103 -2024 -15079
rect -2058 -15147 -2024 -15141
rect -2058 -15175 -2024 -15147
rect -2058 -15215 -2024 -15213
rect -2058 -15247 -2024 -15215
rect -2058 -15317 -2024 -15285
rect -2058 -15319 -2024 -15317
rect -2058 -15385 -2024 -15357
rect -2058 -15391 -2024 -15385
rect -2058 -15453 -2024 -15429
rect -2058 -15463 -2024 -15453
rect -2058 -15521 -2024 -15501
rect -2058 -15535 -2024 -15521
rect -1040 -15011 -1006 -14997
rect -1040 -15031 -1006 -15011
rect -1040 -15079 -1006 -15069
rect -1040 -15103 -1006 -15079
rect -1040 -15147 -1006 -15141
rect -1040 -15175 -1006 -15147
rect -1040 -15215 -1006 -15213
rect -1040 -15247 -1006 -15215
rect -1040 -15317 -1006 -15285
rect -1040 -15319 -1006 -15317
rect -1040 -15385 -1006 -15357
rect -1040 -15391 -1006 -15385
rect -1040 -15453 -1006 -15429
rect -1040 -15463 -1006 -15453
rect -1040 -15521 -1006 -15501
rect -1040 -15535 -1006 -15521
rect -22 -15011 12 -14997
rect -22 -15031 12 -15011
rect -22 -15079 12 -15069
rect -22 -15103 12 -15079
rect -22 -15147 12 -15141
rect -22 -15175 12 -15147
rect -22 -15215 12 -15213
rect -22 -15247 12 -15215
rect -22 -15317 12 -15285
rect -22 -15319 12 -15317
rect -22 -15385 12 -15357
rect -22 -15391 12 -15385
rect 24855 -15001 24889 -14971
rect 24855 -15005 24889 -15001
rect 24855 -15069 24889 -15043
rect 24855 -15077 24889 -15069
rect 24855 -15137 24889 -15115
rect 24855 -15149 24889 -15137
rect 24855 -15205 24889 -15187
rect 24855 -15221 24889 -15205
rect 24855 -15273 24889 -15259
rect 24855 -15293 24889 -15273
rect 24855 -15341 24889 -15331
rect 24855 -15365 24889 -15341
rect 2911 -15426 2921 -15392
rect 2921 -15426 2945 -15392
rect 2983 -15426 2989 -15392
rect 2989 -15426 3017 -15392
rect 3055 -15426 3057 -15392
rect 3057 -15426 3089 -15392
rect 3127 -15426 3159 -15392
rect 3159 -15426 3161 -15392
rect 3199 -15426 3227 -15392
rect 3227 -15426 3233 -15392
rect 3271 -15426 3295 -15392
rect 3295 -15426 3305 -15392
rect 3929 -15426 3939 -15392
rect 3939 -15426 3963 -15392
rect 4001 -15426 4007 -15392
rect 4007 -15426 4035 -15392
rect 4073 -15426 4075 -15392
rect 4075 -15426 4107 -15392
rect 4145 -15426 4177 -15392
rect 4177 -15426 4179 -15392
rect 4217 -15426 4245 -15392
rect 4245 -15426 4251 -15392
rect 4289 -15426 4313 -15392
rect 4313 -15426 4323 -15392
rect 4947 -15426 4957 -15392
rect 4957 -15426 4981 -15392
rect 5019 -15426 5025 -15392
rect 5025 -15426 5053 -15392
rect 5091 -15426 5093 -15392
rect 5093 -15426 5125 -15392
rect 5163 -15426 5195 -15392
rect 5195 -15426 5197 -15392
rect 5235 -15426 5263 -15392
rect 5263 -15426 5269 -15392
rect 5307 -15426 5331 -15392
rect 5331 -15426 5341 -15392
rect 5965 -15426 5975 -15392
rect 5975 -15426 5999 -15392
rect 6037 -15426 6043 -15392
rect 6043 -15426 6071 -15392
rect 6109 -15426 6111 -15392
rect 6111 -15426 6143 -15392
rect 6181 -15426 6213 -15392
rect 6213 -15426 6215 -15392
rect 6253 -15426 6281 -15392
rect 6281 -15426 6287 -15392
rect 6325 -15426 6349 -15392
rect 6349 -15426 6359 -15392
rect 6983 -15426 6993 -15392
rect 6993 -15426 7017 -15392
rect 7055 -15426 7061 -15392
rect 7061 -15426 7089 -15392
rect 7127 -15426 7129 -15392
rect 7129 -15426 7161 -15392
rect 7199 -15426 7231 -15392
rect 7231 -15426 7233 -15392
rect 7271 -15426 7299 -15392
rect 7299 -15426 7305 -15392
rect 7343 -15426 7367 -15392
rect 7367 -15426 7377 -15392
rect 8001 -15426 8011 -15392
rect 8011 -15426 8035 -15392
rect 8073 -15426 8079 -15392
rect 8079 -15426 8107 -15392
rect 8145 -15426 8147 -15392
rect 8147 -15426 8179 -15392
rect 8217 -15426 8249 -15392
rect 8249 -15426 8251 -15392
rect 8289 -15426 8317 -15392
rect 8317 -15426 8323 -15392
rect 8361 -15426 8385 -15392
rect 8385 -15426 8395 -15392
rect 9019 -15426 9029 -15392
rect 9029 -15426 9053 -15392
rect 9091 -15426 9097 -15392
rect 9097 -15426 9125 -15392
rect 9163 -15426 9165 -15392
rect 9165 -15426 9197 -15392
rect 9235 -15426 9267 -15392
rect 9267 -15426 9269 -15392
rect 9307 -15426 9335 -15392
rect 9335 -15426 9341 -15392
rect 9379 -15426 9403 -15392
rect 9403 -15426 9413 -15392
rect 10037 -15426 10047 -15392
rect 10047 -15426 10071 -15392
rect 10109 -15426 10115 -15392
rect 10115 -15426 10143 -15392
rect 10181 -15426 10183 -15392
rect 10183 -15426 10215 -15392
rect 10253 -15426 10285 -15392
rect 10285 -15426 10287 -15392
rect 10325 -15426 10353 -15392
rect 10353 -15426 10359 -15392
rect 10397 -15426 10421 -15392
rect 10421 -15426 10431 -15392
rect 11055 -15426 11065 -15392
rect 11065 -15426 11089 -15392
rect 11127 -15426 11133 -15392
rect 11133 -15426 11161 -15392
rect 11199 -15426 11201 -15392
rect 11201 -15426 11233 -15392
rect 11271 -15426 11303 -15392
rect 11303 -15426 11305 -15392
rect 11343 -15426 11371 -15392
rect 11371 -15426 11377 -15392
rect 11415 -15426 11439 -15392
rect 11439 -15426 11449 -15392
rect 12073 -15426 12083 -15392
rect 12083 -15426 12107 -15392
rect 12145 -15426 12151 -15392
rect 12151 -15426 12179 -15392
rect 12217 -15426 12219 -15392
rect 12219 -15426 12251 -15392
rect 12289 -15426 12321 -15392
rect 12321 -15426 12323 -15392
rect 12361 -15426 12389 -15392
rect 12389 -15426 12395 -15392
rect 12433 -15426 12457 -15392
rect 12457 -15426 12467 -15392
rect 13091 -15426 13101 -15392
rect 13101 -15426 13125 -15392
rect 13163 -15426 13169 -15392
rect 13169 -15426 13197 -15392
rect 13235 -15426 13237 -15392
rect 13237 -15426 13269 -15392
rect 13307 -15426 13339 -15392
rect 13339 -15426 13341 -15392
rect 13379 -15426 13407 -15392
rect 13407 -15426 13413 -15392
rect 13451 -15426 13475 -15392
rect 13475 -15426 13485 -15392
rect 14109 -15426 14119 -15392
rect 14119 -15426 14143 -15392
rect 14181 -15426 14187 -15392
rect 14187 -15426 14215 -15392
rect 14253 -15426 14255 -15392
rect 14255 -15426 14287 -15392
rect 14325 -15426 14357 -15392
rect 14357 -15426 14359 -15392
rect 14397 -15426 14425 -15392
rect 14425 -15426 14431 -15392
rect 14469 -15426 14493 -15392
rect 14493 -15426 14503 -15392
rect 15127 -15426 15137 -15392
rect 15137 -15426 15161 -15392
rect 15199 -15426 15205 -15392
rect 15205 -15426 15233 -15392
rect 15271 -15426 15273 -15392
rect 15273 -15426 15305 -15392
rect 15343 -15426 15375 -15392
rect 15375 -15426 15377 -15392
rect 15415 -15426 15443 -15392
rect 15443 -15426 15449 -15392
rect 15487 -15426 15511 -15392
rect 15511 -15426 15521 -15392
rect 16145 -15426 16155 -15392
rect 16155 -15426 16179 -15392
rect 16217 -15426 16223 -15392
rect 16223 -15426 16251 -15392
rect 16289 -15426 16291 -15392
rect 16291 -15426 16323 -15392
rect 16361 -15426 16393 -15392
rect 16393 -15426 16395 -15392
rect 16433 -15426 16461 -15392
rect 16461 -15426 16467 -15392
rect 16505 -15426 16529 -15392
rect 16529 -15426 16539 -15392
rect 17163 -15426 17173 -15392
rect 17173 -15426 17197 -15392
rect 17235 -15426 17241 -15392
rect 17241 -15426 17269 -15392
rect 17307 -15426 17309 -15392
rect 17309 -15426 17341 -15392
rect 17379 -15426 17411 -15392
rect 17411 -15426 17413 -15392
rect 17451 -15426 17479 -15392
rect 17479 -15426 17485 -15392
rect 17523 -15426 17547 -15392
rect 17547 -15426 17557 -15392
rect 18181 -15426 18191 -15392
rect 18191 -15426 18215 -15392
rect 18253 -15426 18259 -15392
rect 18259 -15426 18287 -15392
rect 18325 -15426 18327 -15392
rect 18327 -15426 18359 -15392
rect 18397 -15426 18429 -15392
rect 18429 -15426 18431 -15392
rect 18469 -15426 18497 -15392
rect 18497 -15426 18503 -15392
rect 18541 -15426 18565 -15392
rect 18565 -15426 18575 -15392
rect 19199 -15426 19209 -15392
rect 19209 -15426 19233 -15392
rect 19271 -15426 19277 -15392
rect 19277 -15426 19305 -15392
rect 19343 -15426 19345 -15392
rect 19345 -15426 19377 -15392
rect 19415 -15426 19447 -15392
rect 19447 -15426 19449 -15392
rect 19487 -15426 19515 -15392
rect 19515 -15426 19521 -15392
rect 19559 -15426 19583 -15392
rect 19583 -15426 19593 -15392
rect 20217 -15426 20227 -15392
rect 20227 -15426 20251 -15392
rect 20289 -15426 20295 -15392
rect 20295 -15426 20323 -15392
rect 20361 -15426 20363 -15392
rect 20363 -15426 20395 -15392
rect 20433 -15426 20465 -15392
rect 20465 -15426 20467 -15392
rect 20505 -15426 20533 -15392
rect 20533 -15426 20539 -15392
rect 20577 -15426 20601 -15392
rect 20601 -15426 20611 -15392
rect 21235 -15426 21245 -15392
rect 21245 -15426 21269 -15392
rect 21307 -15426 21313 -15392
rect 21313 -15426 21341 -15392
rect 21379 -15426 21381 -15392
rect 21381 -15426 21413 -15392
rect 21451 -15426 21483 -15392
rect 21483 -15426 21485 -15392
rect 21523 -15426 21551 -15392
rect 21551 -15426 21557 -15392
rect 21595 -15426 21619 -15392
rect 21619 -15426 21629 -15392
rect 22253 -15426 22263 -15392
rect 22263 -15426 22287 -15392
rect 22325 -15426 22331 -15392
rect 22331 -15426 22359 -15392
rect 22397 -15426 22399 -15392
rect 22399 -15426 22431 -15392
rect 22469 -15426 22501 -15392
rect 22501 -15426 22503 -15392
rect 22541 -15426 22569 -15392
rect 22569 -15426 22575 -15392
rect 22613 -15426 22637 -15392
rect 22637 -15426 22647 -15392
rect -22 -15453 12 -15429
rect -22 -15463 12 -15453
rect 24855 -15409 24889 -15403
rect 24855 -15437 24889 -15409
rect -22 -15521 12 -15501
rect -22 -15535 12 -15521
rect 2582 -15509 2616 -15495
rect 2582 -15529 2616 -15509
rect 2582 -15577 2616 -15567
rect 2582 -15601 2616 -15577
rect -12289 -15647 -12255 -15619
rect -12289 -15653 -12255 -15647
rect -8855 -15638 -8845 -15604
rect -8845 -15638 -8821 -15604
rect -8783 -15638 -8777 -15604
rect -8777 -15638 -8749 -15604
rect -8711 -15638 -8709 -15604
rect -8709 -15638 -8677 -15604
rect -8639 -15638 -8607 -15604
rect -8607 -15638 -8605 -15604
rect -8567 -15638 -8539 -15604
rect -8539 -15638 -8533 -15604
rect -8495 -15638 -8471 -15604
rect -8471 -15638 -8461 -15604
rect -7837 -15638 -7827 -15604
rect -7827 -15638 -7803 -15604
rect -7765 -15638 -7759 -15604
rect -7759 -15638 -7731 -15604
rect -7693 -15638 -7691 -15604
rect -7691 -15638 -7659 -15604
rect -7621 -15638 -7589 -15604
rect -7589 -15638 -7587 -15604
rect -7549 -15638 -7521 -15604
rect -7521 -15638 -7515 -15604
rect -7477 -15638 -7453 -15604
rect -7453 -15638 -7443 -15604
rect -6819 -15638 -6809 -15604
rect -6809 -15638 -6785 -15604
rect -6747 -15638 -6741 -15604
rect -6741 -15638 -6713 -15604
rect -6675 -15638 -6673 -15604
rect -6673 -15638 -6641 -15604
rect -6603 -15638 -6571 -15604
rect -6571 -15638 -6569 -15604
rect -6531 -15638 -6503 -15604
rect -6503 -15638 -6497 -15604
rect -6459 -15638 -6435 -15604
rect -6435 -15638 -6425 -15604
rect -5801 -15638 -5791 -15604
rect -5791 -15638 -5767 -15604
rect -5729 -15638 -5723 -15604
rect -5723 -15638 -5695 -15604
rect -5657 -15638 -5655 -15604
rect -5655 -15638 -5623 -15604
rect -5585 -15638 -5553 -15604
rect -5553 -15638 -5551 -15604
rect -5513 -15638 -5485 -15604
rect -5485 -15638 -5479 -15604
rect -5441 -15638 -5417 -15604
rect -5417 -15638 -5407 -15604
rect -4783 -15638 -4773 -15604
rect -4773 -15638 -4749 -15604
rect -4711 -15638 -4705 -15604
rect -4705 -15638 -4677 -15604
rect -4639 -15638 -4637 -15604
rect -4637 -15638 -4605 -15604
rect -4567 -15638 -4535 -15604
rect -4535 -15638 -4533 -15604
rect -4495 -15638 -4467 -15604
rect -4467 -15638 -4461 -15604
rect -4423 -15638 -4399 -15604
rect -4399 -15638 -4389 -15604
rect -3765 -15638 -3755 -15604
rect -3755 -15638 -3731 -15604
rect -3693 -15638 -3687 -15604
rect -3687 -15638 -3659 -15604
rect -3621 -15638 -3619 -15604
rect -3619 -15638 -3587 -15604
rect -3549 -15638 -3517 -15604
rect -3517 -15638 -3515 -15604
rect -3477 -15638 -3449 -15604
rect -3449 -15638 -3443 -15604
rect -3405 -15638 -3381 -15604
rect -3381 -15638 -3371 -15604
rect -2747 -15638 -2737 -15604
rect -2737 -15638 -2713 -15604
rect -2675 -15638 -2669 -15604
rect -2669 -15638 -2641 -15604
rect -2603 -15638 -2601 -15604
rect -2601 -15638 -2569 -15604
rect -2531 -15638 -2499 -15604
rect -2499 -15638 -2497 -15604
rect -2459 -15638 -2431 -15604
rect -2431 -15638 -2425 -15604
rect -2387 -15638 -2363 -15604
rect -2363 -15638 -2353 -15604
rect -1729 -15638 -1719 -15604
rect -1719 -15638 -1695 -15604
rect -1657 -15638 -1651 -15604
rect -1651 -15638 -1623 -15604
rect -1585 -15638 -1583 -15604
rect -1583 -15638 -1551 -15604
rect -1513 -15638 -1481 -15604
rect -1481 -15638 -1479 -15604
rect -1441 -15638 -1413 -15604
rect -1413 -15638 -1407 -15604
rect -1369 -15638 -1345 -15604
rect -1345 -15638 -1335 -15604
rect -711 -15638 -701 -15604
rect -701 -15638 -677 -15604
rect -639 -15638 -633 -15604
rect -633 -15638 -605 -15604
rect -567 -15638 -565 -15604
rect -565 -15638 -533 -15604
rect -495 -15638 -463 -15604
rect -463 -15638 -461 -15604
rect -423 -15638 -395 -15604
rect -395 -15638 -389 -15604
rect -351 -15638 -327 -15604
rect -327 -15638 -317 -15604
rect -12289 -15715 -12255 -15691
rect -12289 -15725 -12255 -15715
rect 2582 -15645 2616 -15639
rect 2582 -15673 2616 -15645
rect -8855 -15746 -8845 -15712
rect -8845 -15746 -8821 -15712
rect -8783 -15746 -8777 -15712
rect -8777 -15746 -8749 -15712
rect -8711 -15746 -8709 -15712
rect -8709 -15746 -8677 -15712
rect -8639 -15746 -8607 -15712
rect -8607 -15746 -8605 -15712
rect -8567 -15746 -8539 -15712
rect -8539 -15746 -8533 -15712
rect -8495 -15746 -8471 -15712
rect -8471 -15746 -8461 -15712
rect -7837 -15746 -7827 -15712
rect -7827 -15746 -7803 -15712
rect -7765 -15746 -7759 -15712
rect -7759 -15746 -7731 -15712
rect -7693 -15746 -7691 -15712
rect -7691 -15746 -7659 -15712
rect -7621 -15746 -7589 -15712
rect -7589 -15746 -7587 -15712
rect -7549 -15746 -7521 -15712
rect -7521 -15746 -7515 -15712
rect -7477 -15746 -7453 -15712
rect -7453 -15746 -7443 -15712
rect -6819 -15746 -6809 -15712
rect -6809 -15746 -6785 -15712
rect -6747 -15746 -6741 -15712
rect -6741 -15746 -6713 -15712
rect -6675 -15746 -6673 -15712
rect -6673 -15746 -6641 -15712
rect -6603 -15746 -6571 -15712
rect -6571 -15746 -6569 -15712
rect -6531 -15746 -6503 -15712
rect -6503 -15746 -6497 -15712
rect -6459 -15746 -6435 -15712
rect -6435 -15746 -6425 -15712
rect -5801 -15746 -5791 -15712
rect -5791 -15746 -5767 -15712
rect -5729 -15746 -5723 -15712
rect -5723 -15746 -5695 -15712
rect -5657 -15746 -5655 -15712
rect -5655 -15746 -5623 -15712
rect -5585 -15746 -5553 -15712
rect -5553 -15746 -5551 -15712
rect -5513 -15746 -5485 -15712
rect -5485 -15746 -5479 -15712
rect -5441 -15746 -5417 -15712
rect -5417 -15746 -5407 -15712
rect -4783 -15746 -4773 -15712
rect -4773 -15746 -4749 -15712
rect -4711 -15746 -4705 -15712
rect -4705 -15746 -4677 -15712
rect -4639 -15746 -4637 -15712
rect -4637 -15746 -4605 -15712
rect -4567 -15746 -4535 -15712
rect -4535 -15746 -4533 -15712
rect -4495 -15746 -4467 -15712
rect -4467 -15746 -4461 -15712
rect -4423 -15746 -4399 -15712
rect -4399 -15746 -4389 -15712
rect -3765 -15746 -3755 -15712
rect -3755 -15746 -3731 -15712
rect -3693 -15746 -3687 -15712
rect -3687 -15746 -3659 -15712
rect -3621 -15746 -3619 -15712
rect -3619 -15746 -3587 -15712
rect -3549 -15746 -3517 -15712
rect -3517 -15746 -3515 -15712
rect -3477 -15746 -3449 -15712
rect -3449 -15746 -3443 -15712
rect -3405 -15746 -3381 -15712
rect -3381 -15746 -3371 -15712
rect -2747 -15746 -2737 -15712
rect -2737 -15746 -2713 -15712
rect -2675 -15746 -2669 -15712
rect -2669 -15746 -2641 -15712
rect -2603 -15746 -2601 -15712
rect -2601 -15746 -2569 -15712
rect -2531 -15746 -2499 -15712
rect -2499 -15746 -2497 -15712
rect -2459 -15746 -2431 -15712
rect -2431 -15746 -2425 -15712
rect -2387 -15746 -2363 -15712
rect -2363 -15746 -2353 -15712
rect -1729 -15746 -1719 -15712
rect -1719 -15746 -1695 -15712
rect -1657 -15746 -1651 -15712
rect -1651 -15746 -1623 -15712
rect -1585 -15746 -1583 -15712
rect -1583 -15746 -1551 -15712
rect -1513 -15746 -1481 -15712
rect -1481 -15746 -1479 -15712
rect -1441 -15746 -1413 -15712
rect -1413 -15746 -1407 -15712
rect -1369 -15746 -1345 -15712
rect -1345 -15746 -1335 -15712
rect -711 -15746 -701 -15712
rect -701 -15746 -677 -15712
rect -639 -15746 -633 -15712
rect -633 -15746 -605 -15712
rect -567 -15746 -565 -15712
rect -565 -15746 -533 -15712
rect -495 -15746 -463 -15712
rect -463 -15746 -461 -15712
rect -423 -15746 -395 -15712
rect -395 -15746 -389 -15712
rect -351 -15746 -327 -15712
rect -327 -15746 -317 -15712
rect 2582 -15713 2616 -15711
rect 2582 -15745 2616 -15713
rect -12289 -15783 -12255 -15763
rect -12289 -15797 -12255 -15783
rect -12289 -15851 -12255 -15835
rect -12289 -15869 -12255 -15851
rect -12289 -15919 -12255 -15907
rect -12289 -15941 -12255 -15919
rect -12289 -15987 -12255 -15979
rect -12289 -16013 -12255 -15987
rect -12289 -16055 -12255 -16051
rect -12289 -16085 -12255 -16055
rect -12289 -16157 -12255 -16123
rect -12289 -16225 -12255 -16195
rect -12289 -16229 -12255 -16225
rect -12289 -16293 -12255 -16267
rect -12289 -16301 -12255 -16293
rect -12289 -16361 -12255 -16339
rect -12289 -16373 -12255 -16361
rect -9184 -15829 -9150 -15815
rect -9184 -15849 -9150 -15829
rect -9184 -15897 -9150 -15887
rect -9184 -15921 -9150 -15897
rect -9184 -15965 -9150 -15959
rect -9184 -15993 -9150 -15965
rect -9184 -16033 -9150 -16031
rect -9184 -16065 -9150 -16033
rect -9184 -16135 -9150 -16103
rect -9184 -16137 -9150 -16135
rect -9184 -16203 -9150 -16175
rect -9184 -16209 -9150 -16203
rect -9184 -16271 -9150 -16247
rect -9184 -16281 -9150 -16271
rect -9184 -16339 -9150 -16319
rect -9184 -16353 -9150 -16339
rect -8166 -15829 -8132 -15815
rect -8166 -15849 -8132 -15829
rect -8166 -15897 -8132 -15887
rect -8166 -15921 -8132 -15897
rect -8166 -15965 -8132 -15959
rect -8166 -15993 -8132 -15965
rect -8166 -16033 -8132 -16031
rect -8166 -16065 -8132 -16033
rect -8166 -16135 -8132 -16103
rect -8166 -16137 -8132 -16135
rect -8166 -16203 -8132 -16175
rect -8166 -16209 -8132 -16203
rect -8166 -16271 -8132 -16247
rect -8166 -16281 -8132 -16271
rect -8166 -16339 -8132 -16319
rect -8166 -16353 -8132 -16339
rect -7148 -15829 -7114 -15815
rect -7148 -15849 -7114 -15829
rect -7148 -15897 -7114 -15887
rect -7148 -15921 -7114 -15897
rect -7148 -15965 -7114 -15959
rect -7148 -15993 -7114 -15965
rect -7148 -16033 -7114 -16031
rect -7148 -16065 -7114 -16033
rect -7148 -16135 -7114 -16103
rect -7148 -16137 -7114 -16135
rect -7148 -16203 -7114 -16175
rect -7148 -16209 -7114 -16203
rect -7148 -16271 -7114 -16247
rect -7148 -16281 -7114 -16271
rect -7148 -16339 -7114 -16319
rect -7148 -16353 -7114 -16339
rect -6130 -15829 -6096 -15815
rect -6130 -15849 -6096 -15829
rect -6130 -15897 -6096 -15887
rect -6130 -15921 -6096 -15897
rect -6130 -15965 -6096 -15959
rect -6130 -15993 -6096 -15965
rect -6130 -16033 -6096 -16031
rect -6130 -16065 -6096 -16033
rect -6130 -16135 -6096 -16103
rect -6130 -16137 -6096 -16135
rect -6130 -16203 -6096 -16175
rect -6130 -16209 -6096 -16203
rect -6130 -16271 -6096 -16247
rect -6130 -16281 -6096 -16271
rect -6130 -16339 -6096 -16319
rect -6130 -16353 -6096 -16339
rect -5112 -15829 -5078 -15815
rect -5112 -15849 -5078 -15829
rect -5112 -15897 -5078 -15887
rect -5112 -15921 -5078 -15897
rect -5112 -15965 -5078 -15959
rect -5112 -15993 -5078 -15965
rect -5112 -16033 -5078 -16031
rect -5112 -16065 -5078 -16033
rect -5112 -16135 -5078 -16103
rect -5112 -16137 -5078 -16135
rect -5112 -16203 -5078 -16175
rect -5112 -16209 -5078 -16203
rect -5112 -16271 -5078 -16247
rect -5112 -16281 -5078 -16271
rect -5112 -16339 -5078 -16319
rect -5112 -16353 -5078 -16339
rect -4094 -15829 -4060 -15815
rect -4094 -15849 -4060 -15829
rect -4094 -15897 -4060 -15887
rect -4094 -15921 -4060 -15897
rect -4094 -15965 -4060 -15959
rect -4094 -15993 -4060 -15965
rect -4094 -16033 -4060 -16031
rect -4094 -16065 -4060 -16033
rect -4094 -16135 -4060 -16103
rect -4094 -16137 -4060 -16135
rect -4094 -16203 -4060 -16175
rect -4094 -16209 -4060 -16203
rect -4094 -16271 -4060 -16247
rect -4094 -16281 -4060 -16271
rect -4094 -16339 -4060 -16319
rect -4094 -16353 -4060 -16339
rect -3076 -15829 -3042 -15815
rect -3076 -15849 -3042 -15829
rect -3076 -15897 -3042 -15887
rect -3076 -15921 -3042 -15897
rect -3076 -15965 -3042 -15959
rect -3076 -15993 -3042 -15965
rect -3076 -16033 -3042 -16031
rect -3076 -16065 -3042 -16033
rect -3076 -16135 -3042 -16103
rect -3076 -16137 -3042 -16135
rect -3076 -16203 -3042 -16175
rect -3076 -16209 -3042 -16203
rect -3076 -16271 -3042 -16247
rect -3076 -16281 -3042 -16271
rect -3076 -16339 -3042 -16319
rect -3076 -16353 -3042 -16339
rect -2058 -15829 -2024 -15815
rect -2058 -15849 -2024 -15829
rect -2058 -15897 -2024 -15887
rect -2058 -15921 -2024 -15897
rect -2058 -15965 -2024 -15959
rect -2058 -15993 -2024 -15965
rect -2058 -16033 -2024 -16031
rect -2058 -16065 -2024 -16033
rect -2058 -16135 -2024 -16103
rect -2058 -16137 -2024 -16135
rect -2058 -16203 -2024 -16175
rect -2058 -16209 -2024 -16203
rect -2058 -16271 -2024 -16247
rect -2058 -16281 -2024 -16271
rect -2058 -16339 -2024 -16319
rect -2058 -16353 -2024 -16339
rect -1040 -15829 -1006 -15815
rect -1040 -15849 -1006 -15829
rect -1040 -15897 -1006 -15887
rect -1040 -15921 -1006 -15897
rect -1040 -15965 -1006 -15959
rect -1040 -15993 -1006 -15965
rect -1040 -16033 -1006 -16031
rect -1040 -16065 -1006 -16033
rect -1040 -16135 -1006 -16103
rect -1040 -16137 -1006 -16135
rect -1040 -16203 -1006 -16175
rect -1040 -16209 -1006 -16203
rect -1040 -16271 -1006 -16247
rect -1040 -16281 -1006 -16271
rect -1040 -16339 -1006 -16319
rect -1040 -16353 -1006 -16339
rect -22 -15829 12 -15815
rect -22 -15849 12 -15829
rect -22 -15897 12 -15887
rect -22 -15921 12 -15897
rect -22 -15965 12 -15959
rect -22 -15993 12 -15965
rect -22 -16033 12 -16031
rect -22 -16065 12 -16033
rect 2582 -15815 2616 -15783
rect 2582 -15817 2616 -15815
rect 2582 -15883 2616 -15855
rect 2582 -15889 2616 -15883
rect 2582 -15951 2616 -15927
rect 2582 -15961 2616 -15951
rect 2582 -16019 2616 -15999
rect 2582 -16033 2616 -16019
rect 3600 -15509 3634 -15495
rect 3600 -15529 3634 -15509
rect 3600 -15577 3634 -15567
rect 3600 -15601 3634 -15577
rect 3600 -15645 3634 -15639
rect 3600 -15673 3634 -15645
rect 3600 -15713 3634 -15711
rect 3600 -15745 3634 -15713
rect 3600 -15815 3634 -15783
rect 3600 -15817 3634 -15815
rect 3600 -15883 3634 -15855
rect 3600 -15889 3634 -15883
rect 3600 -15951 3634 -15927
rect 3600 -15961 3634 -15951
rect 3600 -16019 3634 -15999
rect 3600 -16033 3634 -16019
rect 4618 -15509 4652 -15495
rect 4618 -15529 4652 -15509
rect 4618 -15577 4652 -15567
rect 4618 -15601 4652 -15577
rect 4618 -15645 4652 -15639
rect 4618 -15673 4652 -15645
rect 4618 -15713 4652 -15711
rect 4618 -15745 4652 -15713
rect 4618 -15815 4652 -15783
rect 4618 -15817 4652 -15815
rect 4618 -15883 4652 -15855
rect 4618 -15889 4652 -15883
rect 4618 -15951 4652 -15927
rect 4618 -15961 4652 -15951
rect 4618 -16019 4652 -15999
rect 4618 -16033 4652 -16019
rect 5636 -15509 5670 -15495
rect 5636 -15529 5670 -15509
rect 5636 -15577 5670 -15567
rect 5636 -15601 5670 -15577
rect 5636 -15645 5670 -15639
rect 5636 -15673 5670 -15645
rect 5636 -15713 5670 -15711
rect 5636 -15745 5670 -15713
rect 5636 -15815 5670 -15783
rect 5636 -15817 5670 -15815
rect 5636 -15883 5670 -15855
rect 5636 -15889 5670 -15883
rect 5636 -15951 5670 -15927
rect 5636 -15961 5670 -15951
rect 5636 -16019 5670 -15999
rect 5636 -16033 5670 -16019
rect 6654 -15509 6688 -15495
rect 6654 -15529 6688 -15509
rect 6654 -15577 6688 -15567
rect 6654 -15601 6688 -15577
rect 6654 -15645 6688 -15639
rect 6654 -15673 6688 -15645
rect 6654 -15713 6688 -15711
rect 6654 -15745 6688 -15713
rect 6654 -15815 6688 -15783
rect 6654 -15817 6688 -15815
rect 6654 -15883 6688 -15855
rect 6654 -15889 6688 -15883
rect 6654 -15951 6688 -15927
rect 6654 -15961 6688 -15951
rect 6654 -16019 6688 -15999
rect 6654 -16033 6688 -16019
rect 7672 -15509 7706 -15495
rect 7672 -15529 7706 -15509
rect 7672 -15577 7706 -15567
rect 7672 -15601 7706 -15577
rect 7672 -15645 7706 -15639
rect 7672 -15673 7706 -15645
rect 7672 -15713 7706 -15711
rect 7672 -15745 7706 -15713
rect 7672 -15815 7706 -15783
rect 7672 -15817 7706 -15815
rect 7672 -15883 7706 -15855
rect 7672 -15889 7706 -15883
rect 7672 -15951 7706 -15927
rect 7672 -15961 7706 -15951
rect 7672 -16019 7706 -15999
rect 7672 -16033 7706 -16019
rect 8690 -15509 8724 -15495
rect 8690 -15529 8724 -15509
rect 8690 -15577 8724 -15567
rect 8690 -15601 8724 -15577
rect 8690 -15645 8724 -15639
rect 8690 -15673 8724 -15645
rect 8690 -15713 8724 -15711
rect 8690 -15745 8724 -15713
rect 8690 -15815 8724 -15783
rect 8690 -15817 8724 -15815
rect 8690 -15883 8724 -15855
rect 8690 -15889 8724 -15883
rect 8690 -15951 8724 -15927
rect 8690 -15961 8724 -15951
rect 8690 -16019 8724 -15999
rect 8690 -16033 8724 -16019
rect 9708 -15509 9742 -15495
rect 9708 -15529 9742 -15509
rect 9708 -15577 9742 -15567
rect 9708 -15601 9742 -15577
rect 9708 -15645 9742 -15639
rect 9708 -15673 9742 -15645
rect 9708 -15713 9742 -15711
rect 9708 -15745 9742 -15713
rect 9708 -15815 9742 -15783
rect 9708 -15817 9742 -15815
rect 9708 -15883 9742 -15855
rect 9708 -15889 9742 -15883
rect 9708 -15951 9742 -15927
rect 9708 -15961 9742 -15951
rect 9708 -16019 9742 -15999
rect 9708 -16033 9742 -16019
rect 10726 -15509 10760 -15495
rect 10726 -15529 10760 -15509
rect 10726 -15577 10760 -15567
rect 10726 -15601 10760 -15577
rect 10726 -15645 10760 -15639
rect 10726 -15673 10760 -15645
rect 10726 -15713 10760 -15711
rect 10726 -15745 10760 -15713
rect 10726 -15815 10760 -15783
rect 10726 -15817 10760 -15815
rect 10726 -15883 10760 -15855
rect 10726 -15889 10760 -15883
rect 10726 -15951 10760 -15927
rect 10726 -15961 10760 -15951
rect 10726 -16019 10760 -15999
rect 10726 -16033 10760 -16019
rect 11744 -15509 11778 -15495
rect 11744 -15529 11778 -15509
rect 11744 -15577 11778 -15567
rect 11744 -15601 11778 -15577
rect 11744 -15645 11778 -15639
rect 11744 -15673 11778 -15645
rect 11744 -15713 11778 -15711
rect 11744 -15745 11778 -15713
rect 11744 -15815 11778 -15783
rect 11744 -15817 11778 -15815
rect 11744 -15883 11778 -15855
rect 11744 -15889 11778 -15883
rect 11744 -15951 11778 -15927
rect 11744 -15961 11778 -15951
rect 11744 -16019 11778 -15999
rect 11744 -16033 11778 -16019
rect 12762 -15509 12796 -15495
rect 12762 -15529 12796 -15509
rect 12762 -15577 12796 -15567
rect 12762 -15601 12796 -15577
rect 12762 -15645 12796 -15639
rect 12762 -15673 12796 -15645
rect 12762 -15713 12796 -15711
rect 12762 -15745 12796 -15713
rect 12762 -15815 12796 -15783
rect 12762 -15817 12796 -15815
rect 12762 -15883 12796 -15855
rect 12762 -15889 12796 -15883
rect 12762 -15951 12796 -15927
rect 12762 -15961 12796 -15951
rect 12762 -16019 12796 -15999
rect 12762 -16033 12796 -16019
rect 13780 -15509 13814 -15495
rect 13780 -15529 13814 -15509
rect 13780 -15577 13814 -15567
rect 13780 -15601 13814 -15577
rect 13780 -15645 13814 -15639
rect 13780 -15673 13814 -15645
rect 13780 -15713 13814 -15711
rect 13780 -15745 13814 -15713
rect 13780 -15815 13814 -15783
rect 13780 -15817 13814 -15815
rect 13780 -15883 13814 -15855
rect 13780 -15889 13814 -15883
rect 13780 -15951 13814 -15927
rect 13780 -15961 13814 -15951
rect 13780 -16019 13814 -15999
rect 13780 -16033 13814 -16019
rect 14798 -15509 14832 -15495
rect 14798 -15529 14832 -15509
rect 14798 -15577 14832 -15567
rect 14798 -15601 14832 -15577
rect 14798 -15645 14832 -15639
rect 14798 -15673 14832 -15645
rect 14798 -15713 14832 -15711
rect 14798 -15745 14832 -15713
rect 14798 -15815 14832 -15783
rect 14798 -15817 14832 -15815
rect 14798 -15883 14832 -15855
rect 14798 -15889 14832 -15883
rect 14798 -15951 14832 -15927
rect 14798 -15961 14832 -15951
rect 14798 -16019 14832 -15999
rect 14798 -16033 14832 -16019
rect 15816 -15509 15850 -15495
rect 15816 -15529 15850 -15509
rect 15816 -15577 15850 -15567
rect 15816 -15601 15850 -15577
rect 15816 -15645 15850 -15639
rect 15816 -15673 15850 -15645
rect 15816 -15713 15850 -15711
rect 15816 -15745 15850 -15713
rect 15816 -15815 15850 -15783
rect 15816 -15817 15850 -15815
rect 15816 -15883 15850 -15855
rect 15816 -15889 15850 -15883
rect 15816 -15951 15850 -15927
rect 15816 -15961 15850 -15951
rect 15816 -16019 15850 -15999
rect 15816 -16033 15850 -16019
rect 16834 -15509 16868 -15495
rect 16834 -15529 16868 -15509
rect 16834 -15577 16868 -15567
rect 16834 -15601 16868 -15577
rect 16834 -15645 16868 -15639
rect 16834 -15673 16868 -15645
rect 16834 -15713 16868 -15711
rect 16834 -15745 16868 -15713
rect 16834 -15815 16868 -15783
rect 16834 -15817 16868 -15815
rect 16834 -15883 16868 -15855
rect 16834 -15889 16868 -15883
rect 16834 -15951 16868 -15927
rect 16834 -15961 16868 -15951
rect 16834 -16019 16868 -15999
rect 16834 -16033 16868 -16019
rect 17852 -15509 17886 -15495
rect 17852 -15529 17886 -15509
rect 17852 -15577 17886 -15567
rect 17852 -15601 17886 -15577
rect 17852 -15645 17886 -15639
rect 17852 -15673 17886 -15645
rect 17852 -15713 17886 -15711
rect 17852 -15745 17886 -15713
rect 17852 -15815 17886 -15783
rect 17852 -15817 17886 -15815
rect 17852 -15883 17886 -15855
rect 17852 -15889 17886 -15883
rect 17852 -15951 17886 -15927
rect 17852 -15961 17886 -15951
rect 17852 -16019 17886 -15999
rect 17852 -16033 17886 -16019
rect 18870 -15509 18904 -15495
rect 18870 -15529 18904 -15509
rect 18870 -15577 18904 -15567
rect 18870 -15601 18904 -15577
rect 18870 -15645 18904 -15639
rect 18870 -15673 18904 -15645
rect 18870 -15713 18904 -15711
rect 18870 -15745 18904 -15713
rect 18870 -15815 18904 -15783
rect 18870 -15817 18904 -15815
rect 18870 -15883 18904 -15855
rect 18870 -15889 18904 -15883
rect 18870 -15951 18904 -15927
rect 18870 -15961 18904 -15951
rect 18870 -16019 18904 -15999
rect 18870 -16033 18904 -16019
rect 19888 -15509 19922 -15495
rect 19888 -15529 19922 -15509
rect 19888 -15577 19922 -15567
rect 19888 -15601 19922 -15577
rect 19888 -15645 19922 -15639
rect 19888 -15673 19922 -15645
rect 19888 -15713 19922 -15711
rect 19888 -15745 19922 -15713
rect 19888 -15815 19922 -15783
rect 19888 -15817 19922 -15815
rect 19888 -15883 19922 -15855
rect 19888 -15889 19922 -15883
rect 19888 -15951 19922 -15927
rect 19888 -15961 19922 -15951
rect 19888 -16019 19922 -15999
rect 19888 -16033 19922 -16019
rect 20906 -15509 20940 -15495
rect 20906 -15529 20940 -15509
rect 20906 -15577 20940 -15567
rect 20906 -15601 20940 -15577
rect 20906 -15645 20940 -15639
rect 20906 -15673 20940 -15645
rect 20906 -15713 20940 -15711
rect 20906 -15745 20940 -15713
rect 20906 -15815 20940 -15783
rect 20906 -15817 20940 -15815
rect 20906 -15883 20940 -15855
rect 20906 -15889 20940 -15883
rect 20906 -15951 20940 -15927
rect 20906 -15961 20940 -15951
rect 20906 -16019 20940 -15999
rect 20906 -16033 20940 -16019
rect 21924 -15509 21958 -15495
rect 21924 -15529 21958 -15509
rect 21924 -15577 21958 -15567
rect 21924 -15601 21958 -15577
rect 21924 -15645 21958 -15639
rect 21924 -15673 21958 -15645
rect 21924 -15713 21958 -15711
rect 21924 -15745 21958 -15713
rect 21924 -15815 21958 -15783
rect 21924 -15817 21958 -15815
rect 21924 -15883 21958 -15855
rect 21924 -15889 21958 -15883
rect 21924 -15951 21958 -15927
rect 21924 -15961 21958 -15951
rect 21924 -16019 21958 -15999
rect 21924 -16033 21958 -16019
rect 22942 -15509 22976 -15495
rect 22942 -15529 22976 -15509
rect 22942 -15577 22976 -15567
rect 22942 -15601 22976 -15577
rect 22942 -15645 22976 -15639
rect 22942 -15673 22976 -15645
rect 22942 -15713 22976 -15711
rect 22942 -15745 22976 -15713
rect 22942 -15815 22976 -15783
rect 22942 -15817 22976 -15815
rect 22942 -15883 22976 -15855
rect 22942 -15889 22976 -15883
rect 22942 -15951 22976 -15927
rect 22942 -15961 22976 -15951
rect 22942 -16019 22976 -15999
rect 24855 -15477 24889 -15475
rect 24855 -15509 24889 -15477
rect 24855 -15579 24889 -15547
rect 24855 -15581 24889 -15579
rect 24855 -15647 24889 -15619
rect 24855 -15653 24889 -15647
rect 24855 -15715 24889 -15691
rect 24855 -15725 24889 -15715
rect 24855 -15783 24889 -15763
rect 24855 -15797 24889 -15783
rect 24855 -15851 24889 -15835
rect 24855 -15869 24889 -15851
rect 24855 -15919 24889 -15907
rect 24855 -15941 24889 -15919
rect 22942 -16033 22976 -16019
rect 24855 -15987 24889 -15979
rect 24855 -16013 24889 -15987
rect 24855 -16055 24889 -16051
rect 24855 -16085 24889 -16055
rect -22 -16135 12 -16103
rect -22 -16137 12 -16135
rect 2911 -16136 2921 -16102
rect 2921 -16136 2945 -16102
rect 2983 -16136 2989 -16102
rect 2989 -16136 3017 -16102
rect 3055 -16136 3057 -16102
rect 3057 -16136 3089 -16102
rect 3127 -16136 3159 -16102
rect 3159 -16136 3161 -16102
rect 3199 -16136 3227 -16102
rect 3227 -16136 3233 -16102
rect 3271 -16136 3295 -16102
rect 3295 -16136 3305 -16102
rect 3929 -16136 3939 -16102
rect 3939 -16136 3963 -16102
rect 4001 -16136 4007 -16102
rect 4007 -16136 4035 -16102
rect 4073 -16136 4075 -16102
rect 4075 -16136 4107 -16102
rect 4145 -16136 4177 -16102
rect 4177 -16136 4179 -16102
rect 4217 -16136 4245 -16102
rect 4245 -16136 4251 -16102
rect 4289 -16136 4313 -16102
rect 4313 -16136 4323 -16102
rect 4947 -16136 4957 -16102
rect 4957 -16136 4981 -16102
rect 5019 -16136 5025 -16102
rect 5025 -16136 5053 -16102
rect 5091 -16136 5093 -16102
rect 5093 -16136 5125 -16102
rect 5163 -16136 5195 -16102
rect 5195 -16136 5197 -16102
rect 5235 -16136 5263 -16102
rect 5263 -16136 5269 -16102
rect 5307 -16136 5331 -16102
rect 5331 -16136 5341 -16102
rect 5965 -16136 5975 -16102
rect 5975 -16136 5999 -16102
rect 6037 -16136 6043 -16102
rect 6043 -16136 6071 -16102
rect 6109 -16136 6111 -16102
rect 6111 -16136 6143 -16102
rect 6181 -16136 6213 -16102
rect 6213 -16136 6215 -16102
rect 6253 -16136 6281 -16102
rect 6281 -16136 6287 -16102
rect 6325 -16136 6349 -16102
rect 6349 -16136 6359 -16102
rect 6983 -16136 6993 -16102
rect 6993 -16136 7017 -16102
rect 7055 -16136 7061 -16102
rect 7061 -16136 7089 -16102
rect 7127 -16136 7129 -16102
rect 7129 -16136 7161 -16102
rect 7199 -16136 7231 -16102
rect 7231 -16136 7233 -16102
rect 7271 -16136 7299 -16102
rect 7299 -16136 7305 -16102
rect 7343 -16136 7367 -16102
rect 7367 -16136 7377 -16102
rect 8001 -16136 8011 -16102
rect 8011 -16136 8035 -16102
rect 8073 -16136 8079 -16102
rect 8079 -16136 8107 -16102
rect 8145 -16136 8147 -16102
rect 8147 -16136 8179 -16102
rect 8217 -16136 8249 -16102
rect 8249 -16136 8251 -16102
rect 8289 -16136 8317 -16102
rect 8317 -16136 8323 -16102
rect 8361 -16136 8385 -16102
rect 8385 -16136 8395 -16102
rect 9019 -16136 9029 -16102
rect 9029 -16136 9053 -16102
rect 9091 -16136 9097 -16102
rect 9097 -16136 9125 -16102
rect 9163 -16136 9165 -16102
rect 9165 -16136 9197 -16102
rect 9235 -16136 9267 -16102
rect 9267 -16136 9269 -16102
rect 9307 -16136 9335 -16102
rect 9335 -16136 9341 -16102
rect 9379 -16136 9403 -16102
rect 9403 -16136 9413 -16102
rect 10037 -16136 10047 -16102
rect 10047 -16136 10071 -16102
rect 10109 -16136 10115 -16102
rect 10115 -16136 10143 -16102
rect 10181 -16136 10183 -16102
rect 10183 -16136 10215 -16102
rect 10253 -16136 10285 -16102
rect 10285 -16136 10287 -16102
rect 10325 -16136 10353 -16102
rect 10353 -16136 10359 -16102
rect 10397 -16136 10421 -16102
rect 10421 -16136 10431 -16102
rect 11055 -16136 11065 -16102
rect 11065 -16136 11089 -16102
rect 11127 -16136 11133 -16102
rect 11133 -16136 11161 -16102
rect 11199 -16136 11201 -16102
rect 11201 -16136 11233 -16102
rect 11271 -16136 11303 -16102
rect 11303 -16136 11305 -16102
rect 11343 -16136 11371 -16102
rect 11371 -16136 11377 -16102
rect 11415 -16136 11439 -16102
rect 11439 -16136 11449 -16102
rect 12073 -16136 12083 -16102
rect 12083 -16136 12107 -16102
rect 12145 -16136 12151 -16102
rect 12151 -16136 12179 -16102
rect 12217 -16136 12219 -16102
rect 12219 -16136 12251 -16102
rect 12289 -16136 12321 -16102
rect 12321 -16136 12323 -16102
rect 12361 -16136 12389 -16102
rect 12389 -16136 12395 -16102
rect 12433 -16136 12457 -16102
rect 12457 -16136 12467 -16102
rect 13091 -16136 13101 -16102
rect 13101 -16136 13125 -16102
rect 13163 -16136 13169 -16102
rect 13169 -16136 13197 -16102
rect 13235 -16136 13237 -16102
rect 13237 -16136 13269 -16102
rect 13307 -16136 13339 -16102
rect 13339 -16136 13341 -16102
rect 13379 -16136 13407 -16102
rect 13407 -16136 13413 -16102
rect 13451 -16136 13475 -16102
rect 13475 -16136 13485 -16102
rect 14109 -16136 14119 -16102
rect 14119 -16136 14143 -16102
rect 14181 -16136 14187 -16102
rect 14187 -16136 14215 -16102
rect 14253 -16136 14255 -16102
rect 14255 -16136 14287 -16102
rect 14325 -16136 14357 -16102
rect 14357 -16136 14359 -16102
rect 14397 -16136 14425 -16102
rect 14425 -16136 14431 -16102
rect 14469 -16136 14493 -16102
rect 14493 -16136 14503 -16102
rect 15127 -16136 15137 -16102
rect 15137 -16136 15161 -16102
rect 15199 -16136 15205 -16102
rect 15205 -16136 15233 -16102
rect 15271 -16136 15273 -16102
rect 15273 -16136 15305 -16102
rect 15343 -16136 15375 -16102
rect 15375 -16136 15377 -16102
rect 15415 -16136 15443 -16102
rect 15443 -16136 15449 -16102
rect 15487 -16136 15511 -16102
rect 15511 -16136 15521 -16102
rect 16145 -16136 16155 -16102
rect 16155 -16136 16179 -16102
rect 16217 -16136 16223 -16102
rect 16223 -16136 16251 -16102
rect 16289 -16136 16291 -16102
rect 16291 -16136 16323 -16102
rect 16361 -16136 16393 -16102
rect 16393 -16136 16395 -16102
rect 16433 -16136 16461 -16102
rect 16461 -16136 16467 -16102
rect 16505 -16136 16529 -16102
rect 16529 -16136 16539 -16102
rect 17163 -16136 17173 -16102
rect 17173 -16136 17197 -16102
rect 17235 -16136 17241 -16102
rect 17241 -16136 17269 -16102
rect 17379 -16136 17411 -16102
rect 17411 -16136 17413 -16102
rect 17451 -16136 17479 -16102
rect 17479 -16136 17485 -16102
rect 17523 -16136 17547 -16102
rect 17547 -16136 17557 -16102
rect 18181 -16136 18191 -16102
rect 18191 -16136 18215 -16102
rect 18253 -16136 18259 -16102
rect 18259 -16136 18287 -16102
rect 18469 -16136 18497 -16102
rect 18497 -16136 18503 -16102
rect 18541 -16136 18565 -16102
rect 18565 -16136 18575 -16102
rect 19199 -16136 19209 -16102
rect 19209 -16136 19233 -16102
rect 19271 -16136 19277 -16102
rect 19277 -16136 19305 -16102
rect 19343 -16136 19345 -16102
rect 19345 -16136 19377 -16102
rect 19415 -16136 19447 -16102
rect 19447 -16136 19449 -16102
rect 19487 -16136 19515 -16102
rect 19515 -16136 19521 -16102
rect 19559 -16136 19583 -16102
rect 19583 -16136 19593 -16102
rect 20217 -16136 20227 -16102
rect 20227 -16136 20251 -16102
rect 20289 -16136 20295 -16102
rect 20295 -16136 20323 -16102
rect 20361 -16136 20363 -16102
rect 20363 -16136 20395 -16102
rect 20433 -16136 20465 -16102
rect 20465 -16136 20467 -16102
rect 20505 -16136 20533 -16102
rect 20533 -16136 20539 -16102
rect 20577 -16136 20601 -16102
rect 20601 -16136 20611 -16102
rect 21235 -16136 21245 -16102
rect 21245 -16136 21269 -16102
rect 21307 -16136 21313 -16102
rect 21313 -16136 21341 -16102
rect 21379 -16136 21381 -16102
rect 21381 -16136 21413 -16102
rect 21451 -16136 21483 -16102
rect 21483 -16136 21485 -16102
rect 21523 -16136 21551 -16102
rect 21551 -16136 21557 -16102
rect 21595 -16136 21619 -16102
rect 21619 -16136 21629 -16102
rect 22253 -16136 22263 -16102
rect 22263 -16136 22287 -16102
rect 22325 -16136 22331 -16102
rect 22331 -16136 22359 -16102
rect 22397 -16136 22399 -16102
rect 22399 -16136 22431 -16102
rect 22469 -16136 22501 -16102
rect 22501 -16136 22503 -16102
rect 22541 -16136 22569 -16102
rect 22569 -16136 22575 -16102
rect 22613 -16136 22637 -16102
rect 22637 -16136 22647 -16102
rect -22 -16203 12 -16175
rect -22 -16209 12 -16203
rect -22 -16271 12 -16247
rect -22 -16281 12 -16271
rect -22 -16339 12 -16319
rect -22 -16353 12 -16339
rect 24855 -16157 24889 -16123
rect 24855 -16225 24889 -16195
rect 24855 -16229 24889 -16225
rect 24855 -16293 24889 -16267
rect 24855 -16301 24889 -16293
rect 24855 -16361 24889 -16339
rect 24855 -16373 24889 -16361
rect -12289 -16429 -12255 -16411
rect -12289 -16445 -12255 -16429
rect -8855 -16456 -8845 -16422
rect -8845 -16456 -8821 -16422
rect -8783 -16456 -8777 -16422
rect -8777 -16456 -8749 -16422
rect -8711 -16456 -8709 -16422
rect -8709 -16456 -8677 -16422
rect -8639 -16456 -8607 -16422
rect -8607 -16456 -8605 -16422
rect -8567 -16456 -8539 -16422
rect -8539 -16456 -8533 -16422
rect -8495 -16456 -8471 -16422
rect -8471 -16456 -8461 -16422
rect -7837 -16456 -7827 -16422
rect -7827 -16456 -7803 -16422
rect -7765 -16456 -7759 -16422
rect -7759 -16456 -7731 -16422
rect -7693 -16456 -7691 -16422
rect -7691 -16456 -7659 -16422
rect -7621 -16456 -7589 -16422
rect -7589 -16456 -7587 -16422
rect -7549 -16456 -7521 -16422
rect -7521 -16456 -7515 -16422
rect -7477 -16456 -7453 -16422
rect -7453 -16456 -7443 -16422
rect -6819 -16456 -6809 -16422
rect -6809 -16456 -6785 -16422
rect -6747 -16456 -6741 -16422
rect -6741 -16456 -6713 -16422
rect -6675 -16456 -6673 -16422
rect -6673 -16456 -6641 -16422
rect -6603 -16456 -6571 -16422
rect -6571 -16456 -6569 -16422
rect -6531 -16456 -6503 -16422
rect -6503 -16456 -6497 -16422
rect -6459 -16456 -6435 -16422
rect -6435 -16456 -6425 -16422
rect -5801 -16456 -5791 -16422
rect -5791 -16456 -5767 -16422
rect -5729 -16456 -5723 -16422
rect -5723 -16456 -5695 -16422
rect -5657 -16456 -5655 -16422
rect -5655 -16456 -5623 -16422
rect -5585 -16456 -5553 -16422
rect -5553 -16456 -5551 -16422
rect -5513 -16456 -5485 -16422
rect -5485 -16456 -5479 -16422
rect -5441 -16456 -5417 -16422
rect -5417 -16456 -5407 -16422
rect -4783 -16456 -4773 -16422
rect -4773 -16456 -4749 -16422
rect -4711 -16456 -4705 -16422
rect -4705 -16456 -4677 -16422
rect -4639 -16456 -4637 -16422
rect -4637 -16456 -4605 -16422
rect -4567 -16456 -4535 -16422
rect -4535 -16456 -4533 -16422
rect -4495 -16456 -4467 -16422
rect -4467 -16456 -4461 -16422
rect -4423 -16456 -4399 -16422
rect -4399 -16456 -4389 -16422
rect -3765 -16456 -3755 -16422
rect -3755 -16456 -3731 -16422
rect -3693 -16456 -3687 -16422
rect -3687 -16456 -3659 -16422
rect -3621 -16456 -3619 -16422
rect -3619 -16456 -3587 -16422
rect -3549 -16456 -3517 -16422
rect -3517 -16456 -3515 -16422
rect -3477 -16456 -3449 -16422
rect -3449 -16456 -3443 -16422
rect -3405 -16456 -3381 -16422
rect -3381 -16456 -3371 -16422
rect -2747 -16456 -2737 -16422
rect -2737 -16456 -2713 -16422
rect -2675 -16456 -2669 -16422
rect -2669 -16456 -2641 -16422
rect -2603 -16456 -2601 -16422
rect -2601 -16456 -2569 -16422
rect -2531 -16456 -2499 -16422
rect -2499 -16456 -2497 -16422
rect -2459 -16456 -2431 -16422
rect -2431 -16456 -2425 -16422
rect -2387 -16456 -2363 -16422
rect -2363 -16456 -2353 -16422
rect -1729 -16456 -1719 -16422
rect -1719 -16456 -1695 -16422
rect -1657 -16456 -1651 -16422
rect -1651 -16456 -1623 -16422
rect -1585 -16456 -1583 -16422
rect -1583 -16456 -1551 -16422
rect -1513 -16456 -1481 -16422
rect -1481 -16456 -1479 -16422
rect -1441 -16456 -1413 -16422
rect -1413 -16456 -1407 -16422
rect -1369 -16456 -1345 -16422
rect -1345 -16456 -1335 -16422
rect -711 -16456 -701 -16422
rect -701 -16456 -677 -16422
rect -639 -16456 -633 -16422
rect -633 -16456 -605 -16422
rect -567 -16456 -565 -16422
rect -565 -16456 -533 -16422
rect -495 -16456 -463 -16422
rect -463 -16456 -461 -16422
rect -423 -16456 -395 -16422
rect -395 -16456 -389 -16422
rect -351 -16456 -327 -16422
rect -327 -16456 -317 -16422
rect 24855 -16429 24889 -16411
rect 24855 -16445 24889 -16429
rect -12289 -16497 -12255 -16483
rect -12289 -16517 -12255 -16497
rect 24855 -16497 24889 -16483
rect 24855 -16517 24889 -16497
rect -12289 -16565 -12255 -16555
rect -12289 -16589 -12255 -16565
rect -8855 -16564 -8845 -16530
rect -8845 -16564 -8821 -16530
rect -8783 -16564 -8777 -16530
rect -8777 -16564 -8749 -16530
rect -8711 -16564 -8709 -16530
rect -8709 -16564 -8677 -16530
rect -8639 -16564 -8607 -16530
rect -8607 -16564 -8605 -16530
rect -8567 -16564 -8539 -16530
rect -8539 -16564 -8533 -16530
rect -8495 -16564 -8471 -16530
rect -8471 -16564 -8461 -16530
rect -7837 -16564 -7827 -16530
rect -7827 -16564 -7803 -16530
rect -7765 -16564 -7759 -16530
rect -7759 -16564 -7731 -16530
rect -7693 -16564 -7691 -16530
rect -7691 -16564 -7659 -16530
rect -7621 -16564 -7589 -16530
rect -7589 -16564 -7587 -16530
rect -7549 -16564 -7521 -16530
rect -7521 -16564 -7515 -16530
rect -7477 -16564 -7453 -16530
rect -7453 -16564 -7443 -16530
rect -6819 -16564 -6809 -16530
rect -6809 -16564 -6785 -16530
rect -6747 -16564 -6741 -16530
rect -6741 -16564 -6713 -16530
rect -6675 -16564 -6673 -16530
rect -6673 -16564 -6641 -16530
rect -6603 -16564 -6571 -16530
rect -6571 -16564 -6569 -16530
rect -6531 -16564 -6503 -16530
rect -6503 -16564 -6497 -16530
rect -6459 -16564 -6435 -16530
rect -6435 -16564 -6425 -16530
rect -5801 -16564 -5791 -16530
rect -5791 -16564 -5767 -16530
rect -5729 -16564 -5723 -16530
rect -5723 -16564 -5695 -16530
rect -5657 -16564 -5655 -16530
rect -5655 -16564 -5623 -16530
rect -5585 -16564 -5553 -16530
rect -5553 -16564 -5551 -16530
rect -5513 -16564 -5485 -16530
rect -5485 -16564 -5479 -16530
rect -5441 -16564 -5417 -16530
rect -5417 -16564 -5407 -16530
rect -4783 -16564 -4773 -16530
rect -4773 -16564 -4749 -16530
rect -4711 -16564 -4705 -16530
rect -4705 -16564 -4677 -16530
rect -4639 -16564 -4637 -16530
rect -4637 -16564 -4605 -16530
rect -4567 -16564 -4535 -16530
rect -4535 -16564 -4533 -16530
rect -4495 -16564 -4467 -16530
rect -4467 -16564 -4461 -16530
rect -4423 -16564 -4399 -16530
rect -4399 -16564 -4389 -16530
rect -3765 -16564 -3755 -16530
rect -3755 -16564 -3731 -16530
rect -3693 -16564 -3687 -16530
rect -3687 -16564 -3659 -16530
rect -3621 -16564 -3619 -16530
rect -3619 -16564 -3587 -16530
rect -3549 -16564 -3517 -16530
rect -3517 -16564 -3515 -16530
rect -3477 -16564 -3449 -16530
rect -3449 -16564 -3443 -16530
rect -3405 -16564 -3381 -16530
rect -3381 -16564 -3371 -16530
rect -2747 -16564 -2737 -16530
rect -2737 -16564 -2713 -16530
rect -2675 -16564 -2669 -16530
rect -2669 -16564 -2641 -16530
rect -2603 -16564 -2601 -16530
rect -2601 -16564 -2569 -16530
rect -2531 -16564 -2499 -16530
rect -2499 -16564 -2497 -16530
rect -2459 -16564 -2431 -16530
rect -2431 -16564 -2425 -16530
rect -2387 -16564 -2363 -16530
rect -2363 -16564 -2353 -16530
rect -1729 -16564 -1719 -16530
rect -1719 -16564 -1695 -16530
rect -1657 -16564 -1651 -16530
rect -1651 -16564 -1623 -16530
rect -1585 -16564 -1583 -16530
rect -1583 -16564 -1551 -16530
rect -1513 -16564 -1481 -16530
rect -1481 -16564 -1479 -16530
rect -1441 -16564 -1413 -16530
rect -1413 -16564 -1407 -16530
rect -1369 -16564 -1345 -16530
rect -1345 -16564 -1335 -16530
rect -711 -16564 -701 -16530
rect -701 -16564 -677 -16530
rect -639 -16564 -633 -16530
rect -633 -16564 -605 -16530
rect -567 -16564 -565 -16530
rect -565 -16564 -533 -16530
rect -495 -16564 -463 -16530
rect -463 -16564 -461 -16530
rect -423 -16564 -395 -16530
rect -395 -16564 -389 -16530
rect -351 -16564 -327 -16530
rect -327 -16564 -317 -16530
rect 24855 -16565 24889 -16555
rect 24855 -16589 24889 -16565
rect -12289 -16633 -12255 -16627
rect -12289 -16661 -12255 -16633
rect -12289 -16701 -12255 -16699
rect -12289 -16733 -12255 -16701
rect -12289 -16803 -12255 -16771
rect -12289 -16805 -12255 -16803
rect -12289 -16871 -12255 -16843
rect -12289 -16877 -12255 -16871
rect -12289 -16939 -12255 -16915
rect -12289 -16949 -12255 -16939
rect -12289 -17007 -12255 -16987
rect -12289 -17021 -12255 -17007
rect -12289 -17075 -12255 -17059
rect -12289 -17093 -12255 -17075
rect -12289 -17143 -12255 -17131
rect -12289 -17165 -12255 -17143
rect -12289 -17211 -12255 -17203
rect -12289 -17237 -12255 -17211
rect -9184 -16647 -9150 -16633
rect -9184 -16667 -9150 -16647
rect -9184 -16715 -9150 -16705
rect -9184 -16739 -9150 -16715
rect -9184 -16783 -9150 -16777
rect -9184 -16811 -9150 -16783
rect -9184 -16851 -9150 -16849
rect -9184 -16883 -9150 -16851
rect -9184 -16953 -9150 -16921
rect -9184 -16955 -9150 -16953
rect -9184 -17021 -9150 -16993
rect -9184 -17027 -9150 -17021
rect -9184 -17089 -9150 -17065
rect -9184 -17099 -9150 -17089
rect -9184 -17157 -9150 -17137
rect -9184 -17171 -9150 -17157
rect -8166 -16647 -8132 -16633
rect -8166 -16667 -8132 -16647
rect -8166 -16715 -8132 -16705
rect -8166 -16739 -8132 -16715
rect -8166 -16783 -8132 -16777
rect -8166 -16811 -8132 -16783
rect -8166 -16851 -8132 -16849
rect -8166 -16883 -8132 -16851
rect -8166 -16953 -8132 -16921
rect -8166 -16955 -8132 -16953
rect -8166 -17021 -8132 -16993
rect -8166 -17027 -8132 -17021
rect -8166 -17089 -8132 -17065
rect -8166 -17099 -8132 -17089
rect -8166 -17157 -8132 -17137
rect -8166 -17171 -8132 -17157
rect -7148 -16647 -7114 -16633
rect -7148 -16667 -7114 -16647
rect -7148 -16715 -7114 -16705
rect -7148 -16739 -7114 -16715
rect -7148 -16783 -7114 -16777
rect -7148 -16811 -7114 -16783
rect -7148 -16851 -7114 -16849
rect -7148 -16883 -7114 -16851
rect -7148 -16953 -7114 -16921
rect -7148 -16955 -7114 -16953
rect -7148 -17021 -7114 -16993
rect -7148 -17027 -7114 -17021
rect -7148 -17089 -7114 -17065
rect -7148 -17099 -7114 -17089
rect -7148 -17157 -7114 -17137
rect -7148 -17171 -7114 -17157
rect -6130 -16647 -6096 -16633
rect -6130 -16667 -6096 -16647
rect -6130 -16715 -6096 -16705
rect -6130 -16739 -6096 -16715
rect -6130 -16783 -6096 -16777
rect -6130 -16811 -6096 -16783
rect -6130 -16851 -6096 -16849
rect -6130 -16883 -6096 -16851
rect -6130 -16953 -6096 -16921
rect -6130 -16955 -6096 -16953
rect -6130 -17021 -6096 -16993
rect -6130 -17027 -6096 -17021
rect -6130 -17089 -6096 -17065
rect -6130 -17099 -6096 -17089
rect -6130 -17157 -6096 -17137
rect -6130 -17171 -6096 -17157
rect -5112 -16647 -5078 -16633
rect -5112 -16667 -5078 -16647
rect -5112 -16715 -5078 -16705
rect -5112 -16739 -5078 -16715
rect -5112 -16783 -5078 -16777
rect -5112 -16811 -5078 -16783
rect -5112 -16851 -5078 -16849
rect -5112 -16883 -5078 -16851
rect -5112 -16953 -5078 -16921
rect -5112 -16955 -5078 -16953
rect -5112 -17021 -5078 -16993
rect -5112 -17027 -5078 -17021
rect -5112 -17089 -5078 -17065
rect -5112 -17099 -5078 -17089
rect -5112 -17157 -5078 -17137
rect -5112 -17171 -5078 -17157
rect -4094 -16647 -4060 -16633
rect -4094 -16667 -4060 -16647
rect -4094 -16715 -4060 -16705
rect -4094 -16739 -4060 -16715
rect -4094 -16783 -4060 -16777
rect -4094 -16811 -4060 -16783
rect -4094 -16851 -4060 -16849
rect -4094 -16883 -4060 -16851
rect -4094 -16953 -4060 -16921
rect -4094 -16955 -4060 -16953
rect -4094 -17021 -4060 -16993
rect -4094 -17027 -4060 -17021
rect -4094 -17089 -4060 -17065
rect -4094 -17099 -4060 -17089
rect -4094 -17157 -4060 -17137
rect -4094 -17171 -4060 -17157
rect -3076 -16647 -3042 -16633
rect -3076 -16667 -3042 -16647
rect -3076 -16715 -3042 -16705
rect -3076 -16739 -3042 -16715
rect -3076 -16783 -3042 -16777
rect -3076 -16811 -3042 -16783
rect -3076 -16851 -3042 -16849
rect -3076 -16883 -3042 -16851
rect -3076 -16953 -3042 -16921
rect -3076 -16955 -3042 -16953
rect -3076 -17021 -3042 -16993
rect -3076 -17027 -3042 -17021
rect -3076 -17089 -3042 -17065
rect -3076 -17099 -3042 -17089
rect -3076 -17157 -3042 -17137
rect -3076 -17171 -3042 -17157
rect -2058 -16647 -2024 -16633
rect -2058 -16667 -2024 -16647
rect -2058 -16715 -2024 -16705
rect -2058 -16739 -2024 -16715
rect -2058 -16783 -2024 -16777
rect -2058 -16811 -2024 -16783
rect -2058 -16851 -2024 -16849
rect -2058 -16883 -2024 -16851
rect -2058 -16953 -2024 -16921
rect -2058 -16955 -2024 -16953
rect -2058 -17021 -2024 -16993
rect -2058 -17027 -2024 -17021
rect -2058 -17089 -2024 -17065
rect -2058 -17099 -2024 -17089
rect -2058 -17157 -2024 -17137
rect -2058 -17171 -2024 -17157
rect -1040 -16647 -1006 -16633
rect -1040 -16667 -1006 -16647
rect -1040 -16715 -1006 -16705
rect -1040 -16739 -1006 -16715
rect -1040 -16783 -1006 -16777
rect -1040 -16811 -1006 -16783
rect -1040 -16851 -1006 -16849
rect -1040 -16883 -1006 -16851
rect -1040 -16953 -1006 -16921
rect -1040 -16955 -1006 -16953
rect -1040 -17021 -1006 -16993
rect -1040 -17027 -1006 -17021
rect -1040 -17089 -1006 -17065
rect -1040 -17099 -1006 -17089
rect -1040 -17157 -1006 -17137
rect -1040 -17171 -1006 -17157
rect -22 -16647 12 -16633
rect -22 -16667 12 -16647
rect 2909 -16660 2919 -16626
rect 2919 -16660 2943 -16626
rect 2981 -16660 2987 -16626
rect 2987 -16660 3015 -16626
rect 3053 -16660 3055 -16626
rect 3055 -16660 3087 -16626
rect 3125 -16660 3157 -16626
rect 3157 -16660 3159 -16626
rect 3197 -16660 3225 -16626
rect 3225 -16660 3231 -16626
rect 3269 -16660 3293 -16626
rect 3293 -16660 3303 -16626
rect 3927 -16660 3937 -16626
rect 3937 -16660 3961 -16626
rect 3999 -16660 4005 -16626
rect 4005 -16660 4033 -16626
rect 4071 -16660 4073 -16626
rect 4073 -16660 4105 -16626
rect 4143 -16660 4175 -16626
rect 4175 -16660 4177 -16626
rect 4215 -16660 4243 -16626
rect 4243 -16660 4249 -16626
rect 4287 -16660 4311 -16626
rect 4311 -16660 4321 -16626
rect 4945 -16660 4955 -16626
rect 4955 -16660 4979 -16626
rect 5017 -16660 5023 -16626
rect 5023 -16660 5051 -16626
rect 5089 -16660 5091 -16626
rect 5091 -16660 5123 -16626
rect 5161 -16660 5193 -16626
rect 5193 -16660 5195 -16626
rect 5233 -16660 5261 -16626
rect 5261 -16660 5267 -16626
rect 5305 -16660 5329 -16626
rect 5329 -16660 5339 -16626
rect 5963 -16660 5973 -16626
rect 5973 -16660 5997 -16626
rect 6035 -16660 6041 -16626
rect 6041 -16660 6069 -16626
rect 6107 -16660 6109 -16626
rect 6109 -16660 6141 -16626
rect 6179 -16660 6211 -16626
rect 6211 -16660 6213 -16626
rect 6251 -16660 6279 -16626
rect 6279 -16660 6285 -16626
rect 6323 -16660 6347 -16626
rect 6347 -16660 6357 -16626
rect 6981 -16660 6991 -16626
rect 6991 -16660 7015 -16626
rect 7053 -16660 7059 -16626
rect 7059 -16660 7087 -16626
rect 7125 -16660 7127 -16626
rect 7127 -16660 7159 -16626
rect 7197 -16660 7229 -16626
rect 7229 -16660 7231 -16626
rect 7269 -16660 7297 -16626
rect 7297 -16660 7303 -16626
rect 7341 -16660 7365 -16626
rect 7365 -16660 7375 -16626
rect 7999 -16660 8009 -16626
rect 8009 -16660 8033 -16626
rect 8071 -16660 8077 -16626
rect 8077 -16660 8105 -16626
rect 8143 -16660 8145 -16626
rect 8145 -16660 8177 -16626
rect 8215 -16660 8247 -16626
rect 8247 -16660 8249 -16626
rect 8287 -16660 8315 -16626
rect 8315 -16660 8321 -16626
rect 8359 -16660 8383 -16626
rect 8383 -16660 8393 -16626
rect 9017 -16660 9027 -16626
rect 9027 -16660 9051 -16626
rect 9089 -16660 9095 -16626
rect 9095 -16660 9123 -16626
rect 9161 -16660 9163 -16626
rect 9163 -16660 9195 -16626
rect 9233 -16660 9265 -16626
rect 9265 -16660 9267 -16626
rect 9305 -16660 9333 -16626
rect 9333 -16660 9339 -16626
rect 9377 -16660 9401 -16626
rect 9401 -16660 9411 -16626
rect 10035 -16660 10045 -16626
rect 10045 -16660 10069 -16626
rect 10107 -16660 10113 -16626
rect 10113 -16660 10141 -16626
rect 10179 -16660 10181 -16626
rect 10181 -16660 10213 -16626
rect 10251 -16660 10283 -16626
rect 10283 -16660 10285 -16626
rect 10323 -16660 10351 -16626
rect 10351 -16660 10357 -16626
rect 10395 -16660 10419 -16626
rect 10419 -16660 10429 -16626
rect 11053 -16660 11063 -16626
rect 11063 -16660 11087 -16626
rect 11125 -16660 11131 -16626
rect 11131 -16660 11159 -16626
rect 11197 -16660 11199 -16626
rect 11199 -16660 11231 -16626
rect 11269 -16660 11301 -16626
rect 11301 -16660 11303 -16626
rect 11341 -16660 11369 -16626
rect 11369 -16660 11375 -16626
rect 11413 -16660 11437 -16626
rect 11437 -16660 11447 -16626
rect 12071 -16660 12081 -16626
rect 12081 -16660 12105 -16626
rect 12143 -16660 12149 -16626
rect 12149 -16660 12177 -16626
rect 12215 -16660 12217 -16626
rect 12217 -16660 12249 -16626
rect 12287 -16660 12319 -16626
rect 12319 -16660 12321 -16626
rect 12359 -16660 12387 -16626
rect 12387 -16660 12393 -16626
rect 12431 -16660 12455 -16626
rect 12455 -16660 12465 -16626
rect 13089 -16660 13099 -16626
rect 13099 -16660 13123 -16626
rect 13161 -16660 13167 -16626
rect 13167 -16660 13195 -16626
rect 13233 -16660 13235 -16626
rect 13235 -16660 13267 -16626
rect 13305 -16660 13337 -16626
rect 13337 -16660 13339 -16626
rect 13377 -16660 13405 -16626
rect 13405 -16660 13411 -16626
rect 13449 -16660 13473 -16626
rect 13473 -16660 13483 -16626
rect 14107 -16660 14117 -16626
rect 14117 -16660 14141 -16626
rect 14179 -16660 14185 -16626
rect 14185 -16660 14213 -16626
rect 14251 -16660 14253 -16626
rect 14253 -16660 14285 -16626
rect 14323 -16660 14355 -16626
rect 14355 -16660 14357 -16626
rect 14395 -16660 14423 -16626
rect 14423 -16660 14429 -16626
rect 14467 -16660 14491 -16626
rect 14491 -16660 14501 -16626
rect 15125 -16660 15135 -16626
rect 15135 -16660 15159 -16626
rect 15197 -16660 15203 -16626
rect 15203 -16660 15231 -16626
rect 15269 -16660 15271 -16626
rect 15271 -16660 15303 -16626
rect 15341 -16660 15373 -16626
rect 15373 -16660 15375 -16626
rect 15413 -16660 15441 -16626
rect 15441 -16660 15447 -16626
rect 15485 -16660 15509 -16626
rect 15509 -16660 15519 -16626
rect 16143 -16660 16153 -16626
rect 16153 -16660 16177 -16626
rect 16215 -16660 16221 -16626
rect 16221 -16660 16249 -16626
rect 16287 -16660 16289 -16626
rect 16289 -16660 16321 -16626
rect 16359 -16660 16391 -16626
rect 16391 -16660 16393 -16626
rect 16431 -16660 16459 -16626
rect 16459 -16660 16465 -16626
rect 16503 -16660 16527 -16626
rect 16527 -16660 16537 -16626
rect 17161 -16660 17171 -16626
rect 17171 -16660 17195 -16626
rect 17233 -16660 17239 -16626
rect 17239 -16660 17267 -16626
rect 17305 -16660 17307 -16626
rect 17307 -16660 17339 -16626
rect 17377 -16660 17409 -16626
rect 17409 -16660 17411 -16626
rect 17449 -16660 17477 -16626
rect 17477 -16660 17483 -16626
rect 17521 -16660 17545 -16626
rect 17545 -16660 17555 -16626
rect 18179 -16660 18189 -16626
rect 18189 -16660 18213 -16626
rect 18251 -16660 18257 -16626
rect 18257 -16660 18285 -16626
rect 18323 -16660 18325 -16626
rect 18325 -16660 18357 -16626
rect 18395 -16660 18427 -16626
rect 18427 -16660 18429 -16626
rect 18467 -16660 18495 -16626
rect 18495 -16660 18501 -16626
rect 18539 -16660 18563 -16626
rect 18563 -16660 18573 -16626
rect 19197 -16660 19207 -16626
rect 19207 -16660 19231 -16626
rect 19269 -16660 19275 -16626
rect 19275 -16660 19303 -16626
rect 19341 -16660 19343 -16626
rect 19343 -16660 19375 -16626
rect 19413 -16660 19445 -16626
rect 19445 -16660 19447 -16626
rect 19485 -16660 19513 -16626
rect 19513 -16660 19519 -16626
rect 19557 -16660 19581 -16626
rect 19581 -16660 19591 -16626
rect 20215 -16660 20225 -16626
rect 20225 -16660 20249 -16626
rect 20287 -16660 20293 -16626
rect 20293 -16660 20321 -16626
rect 20359 -16660 20361 -16626
rect 20361 -16660 20393 -16626
rect 20431 -16660 20463 -16626
rect 20463 -16660 20465 -16626
rect 20503 -16660 20531 -16626
rect 20531 -16660 20537 -16626
rect 20575 -16660 20599 -16626
rect 20599 -16660 20609 -16626
rect 21233 -16660 21243 -16626
rect 21243 -16660 21267 -16626
rect 21305 -16660 21311 -16626
rect 21311 -16660 21339 -16626
rect 21377 -16660 21379 -16626
rect 21379 -16660 21411 -16626
rect 21449 -16660 21481 -16626
rect 21481 -16660 21483 -16626
rect 21521 -16660 21549 -16626
rect 21549 -16660 21555 -16626
rect 21593 -16660 21617 -16626
rect 21617 -16660 21627 -16626
rect 22251 -16660 22261 -16626
rect 22261 -16660 22285 -16626
rect 22323 -16660 22329 -16626
rect 22329 -16660 22357 -16626
rect 22395 -16660 22397 -16626
rect 22397 -16660 22429 -16626
rect 22467 -16660 22499 -16626
rect 22499 -16660 22501 -16626
rect 22539 -16660 22567 -16626
rect 22567 -16660 22573 -16626
rect 22611 -16660 22635 -16626
rect 22635 -16660 22645 -16626
rect 24855 -16633 24889 -16627
rect 24855 -16661 24889 -16633
rect -22 -16715 12 -16705
rect -22 -16739 12 -16715
rect -22 -16783 12 -16777
rect -22 -16811 12 -16783
rect -22 -16851 12 -16849
rect -22 -16883 12 -16851
rect -22 -16953 12 -16921
rect -22 -16955 12 -16953
rect -22 -17021 12 -16993
rect -22 -17027 12 -17021
rect -22 -17089 12 -17065
rect -22 -17099 12 -17089
rect -22 -17157 12 -17137
rect -22 -17171 12 -17157
rect 2580 -16743 2614 -16729
rect 2580 -16763 2614 -16743
rect 2580 -16811 2614 -16801
rect 2580 -16835 2614 -16811
rect 2580 -16879 2614 -16873
rect 2580 -16907 2614 -16879
rect 2580 -16947 2614 -16945
rect 2580 -16979 2614 -16947
rect 2580 -17049 2614 -17017
rect 2580 -17051 2614 -17049
rect 2580 -17117 2614 -17089
rect 2580 -17123 2614 -17117
rect 2580 -17185 2614 -17161
rect 2580 -17195 2614 -17185
rect -8855 -17274 -8845 -17240
rect -8845 -17274 -8821 -17240
rect -8783 -17274 -8777 -17240
rect -8777 -17274 -8749 -17240
rect -8711 -17274 -8709 -17240
rect -8709 -17274 -8677 -17240
rect -8639 -17274 -8607 -17240
rect -8607 -17274 -8605 -17240
rect -8567 -17274 -8539 -17240
rect -8539 -17274 -8533 -17240
rect -8495 -17274 -8471 -17240
rect -8471 -17274 -8461 -17240
rect -7837 -17274 -7827 -17240
rect -7827 -17274 -7803 -17240
rect -7765 -17274 -7759 -17240
rect -7759 -17274 -7731 -17240
rect -7693 -17274 -7691 -17240
rect -7691 -17274 -7659 -17240
rect -7621 -17274 -7589 -17240
rect -7589 -17274 -7587 -17240
rect -7549 -17274 -7521 -17240
rect -7521 -17274 -7515 -17240
rect -7477 -17274 -7453 -17240
rect -7453 -17274 -7443 -17240
rect -6819 -17274 -6809 -17240
rect -6809 -17274 -6785 -17240
rect -6747 -17274 -6741 -17240
rect -6741 -17274 -6713 -17240
rect -6675 -17274 -6673 -17240
rect -6673 -17274 -6641 -17240
rect -6603 -17274 -6571 -17240
rect -6571 -17274 -6569 -17240
rect -6531 -17274 -6503 -17240
rect -6503 -17274 -6497 -17240
rect -6459 -17274 -6435 -17240
rect -6435 -17274 -6425 -17240
rect -5801 -17274 -5791 -17240
rect -5791 -17274 -5767 -17240
rect -5729 -17274 -5723 -17240
rect -5723 -17274 -5695 -17240
rect -5657 -17274 -5655 -17240
rect -5655 -17274 -5623 -17240
rect -5585 -17274 -5553 -17240
rect -5553 -17274 -5551 -17240
rect -5513 -17274 -5485 -17240
rect -5485 -17274 -5479 -17240
rect -5441 -17274 -5417 -17240
rect -5417 -17274 -5407 -17240
rect -4783 -17274 -4773 -17240
rect -4773 -17274 -4749 -17240
rect -4711 -17274 -4705 -17240
rect -4705 -17274 -4677 -17240
rect -4639 -17274 -4637 -17240
rect -4637 -17274 -4605 -17240
rect -4567 -17274 -4535 -17240
rect -4535 -17274 -4533 -17240
rect -4495 -17274 -4467 -17240
rect -4467 -17274 -4461 -17240
rect -4423 -17274 -4399 -17240
rect -4399 -17274 -4389 -17240
rect -3765 -17274 -3755 -17240
rect -3755 -17274 -3731 -17240
rect -3693 -17274 -3687 -17240
rect -3687 -17274 -3659 -17240
rect -3621 -17274 -3619 -17240
rect -3619 -17274 -3587 -17240
rect -3549 -17274 -3517 -17240
rect -3517 -17274 -3515 -17240
rect -3477 -17274 -3449 -17240
rect -3449 -17274 -3443 -17240
rect -3405 -17274 -3381 -17240
rect -3381 -17274 -3371 -17240
rect -2747 -17274 -2737 -17240
rect -2737 -17274 -2713 -17240
rect -2675 -17274 -2669 -17240
rect -2669 -17274 -2641 -17240
rect -2603 -17274 -2601 -17240
rect -2601 -17274 -2569 -17240
rect -2531 -17274 -2499 -17240
rect -2499 -17274 -2497 -17240
rect -2459 -17274 -2431 -17240
rect -2431 -17274 -2425 -17240
rect -2387 -17274 -2363 -17240
rect -2363 -17274 -2353 -17240
rect -1729 -17274 -1719 -17240
rect -1719 -17274 -1695 -17240
rect -1657 -17274 -1651 -17240
rect -1651 -17274 -1623 -17240
rect -1585 -17274 -1583 -17240
rect -1583 -17274 -1551 -17240
rect -1513 -17274 -1481 -17240
rect -1481 -17274 -1479 -17240
rect -1441 -17274 -1413 -17240
rect -1413 -17274 -1407 -17240
rect -1369 -17274 -1345 -17240
rect -1345 -17274 -1335 -17240
rect -711 -17274 -701 -17240
rect -701 -17274 -677 -17240
rect -639 -17274 -633 -17240
rect -633 -17274 -605 -17240
rect -567 -17274 -565 -17240
rect -565 -17274 -533 -17240
rect -495 -17274 -463 -17240
rect -463 -17274 -461 -17240
rect -423 -17274 -395 -17240
rect -395 -17274 -389 -17240
rect -351 -17274 -327 -17240
rect -327 -17274 -317 -17240
rect 2580 -17253 2614 -17233
rect 2580 -17267 2614 -17253
rect -12289 -17279 -12255 -17275
rect -12289 -17309 -12255 -17279
rect 3598 -16743 3632 -16729
rect 3598 -16763 3632 -16743
rect 3598 -16811 3632 -16801
rect 3598 -16835 3632 -16811
rect 3598 -16879 3632 -16873
rect 3598 -16907 3632 -16879
rect 3598 -16947 3632 -16945
rect 3598 -16979 3632 -16947
rect 3598 -17049 3632 -17017
rect 3598 -17051 3632 -17049
rect 3598 -17117 3632 -17089
rect 3598 -17123 3632 -17117
rect 3598 -17185 3632 -17161
rect 3598 -17195 3632 -17185
rect 3598 -17253 3632 -17233
rect 3598 -17267 3632 -17253
rect 4616 -16743 4650 -16729
rect 4616 -16763 4650 -16743
rect 4616 -16811 4650 -16801
rect 4616 -16835 4650 -16811
rect 4616 -16879 4650 -16873
rect 4616 -16907 4650 -16879
rect 4616 -16947 4650 -16945
rect 4616 -16979 4650 -16947
rect 4616 -17049 4650 -17017
rect 4616 -17051 4650 -17049
rect 4616 -17117 4650 -17089
rect 4616 -17123 4650 -17117
rect 4616 -17185 4650 -17161
rect 4616 -17195 4650 -17185
rect 4616 -17253 4650 -17233
rect 4616 -17267 4650 -17253
rect 5634 -16743 5668 -16729
rect 5634 -16763 5668 -16743
rect 5634 -16811 5668 -16801
rect 5634 -16835 5668 -16811
rect 5634 -16879 5668 -16873
rect 5634 -16907 5668 -16879
rect 5634 -16947 5668 -16945
rect 5634 -16979 5668 -16947
rect 5634 -17049 5668 -17017
rect 5634 -17051 5668 -17049
rect 5634 -17117 5668 -17089
rect 5634 -17123 5668 -17117
rect 5634 -17185 5668 -17161
rect 5634 -17195 5668 -17185
rect 5634 -17253 5668 -17233
rect 5634 -17267 5668 -17253
rect 6652 -16743 6686 -16729
rect 6652 -16763 6686 -16743
rect 6652 -16811 6686 -16801
rect 6652 -16835 6686 -16811
rect 6652 -16879 6686 -16873
rect 6652 -16907 6686 -16879
rect 6652 -16947 6686 -16945
rect 6652 -16979 6686 -16947
rect 6652 -17049 6686 -17017
rect 6652 -17051 6686 -17049
rect 6652 -17117 6686 -17089
rect 6652 -17123 6686 -17117
rect 6652 -17185 6686 -17161
rect 6652 -17195 6686 -17185
rect 6652 -17253 6686 -17233
rect 6652 -17267 6686 -17253
rect 7670 -16743 7704 -16729
rect 7670 -16763 7704 -16743
rect 7670 -16811 7704 -16801
rect 7670 -16835 7704 -16811
rect 7670 -16879 7704 -16873
rect 7670 -16907 7704 -16879
rect 7670 -16947 7704 -16945
rect 7670 -16979 7704 -16947
rect 7670 -17049 7704 -17017
rect 7670 -17051 7704 -17049
rect 7670 -17117 7704 -17089
rect 7670 -17123 7704 -17117
rect 7670 -17185 7704 -17161
rect 7670 -17195 7704 -17185
rect 7670 -17253 7704 -17233
rect 7670 -17267 7704 -17253
rect 8688 -16743 8722 -16729
rect 8688 -16763 8722 -16743
rect 8688 -16811 8722 -16801
rect 8688 -16835 8722 -16811
rect 8688 -16879 8722 -16873
rect 8688 -16907 8722 -16879
rect 8688 -16947 8722 -16945
rect 8688 -16979 8722 -16947
rect 8688 -17049 8722 -17017
rect 8688 -17051 8722 -17049
rect 8688 -17117 8722 -17089
rect 8688 -17123 8722 -17117
rect 8688 -17185 8722 -17161
rect 8688 -17195 8722 -17185
rect 8688 -17253 8722 -17233
rect 8688 -17267 8722 -17253
rect 9706 -16743 9740 -16729
rect 9706 -16763 9740 -16743
rect 9706 -16811 9740 -16801
rect 9706 -16835 9740 -16811
rect 9706 -16879 9740 -16873
rect 9706 -16907 9740 -16879
rect 9706 -16947 9740 -16945
rect 9706 -16979 9740 -16947
rect 9706 -17049 9740 -17017
rect 9706 -17051 9740 -17049
rect 9706 -17117 9740 -17089
rect 9706 -17123 9740 -17117
rect 9706 -17185 9740 -17161
rect 9706 -17195 9740 -17185
rect 9706 -17253 9740 -17233
rect 9706 -17267 9740 -17253
rect 10724 -16743 10758 -16729
rect 10724 -16763 10758 -16743
rect 10724 -16811 10758 -16801
rect 10724 -16835 10758 -16811
rect 10724 -16879 10758 -16873
rect 10724 -16907 10758 -16879
rect 10724 -16947 10758 -16945
rect 10724 -16979 10758 -16947
rect 10724 -17049 10758 -17017
rect 10724 -17051 10758 -17049
rect 10724 -17117 10758 -17089
rect 10724 -17123 10758 -17117
rect 10724 -17185 10758 -17161
rect 10724 -17195 10758 -17185
rect 10724 -17253 10758 -17233
rect 10724 -17267 10758 -17253
rect 11742 -16743 11776 -16729
rect 11742 -16763 11776 -16743
rect 11742 -16811 11776 -16801
rect 11742 -16835 11776 -16811
rect 11742 -16879 11776 -16873
rect 11742 -16907 11776 -16879
rect 11742 -16947 11776 -16945
rect 11742 -16979 11776 -16947
rect 11742 -17049 11776 -17017
rect 11742 -17051 11776 -17049
rect 11742 -17117 11776 -17089
rect 11742 -17123 11776 -17117
rect 11742 -17185 11776 -17161
rect 11742 -17195 11776 -17185
rect 11742 -17253 11776 -17233
rect 11742 -17267 11776 -17253
rect 12760 -16743 12794 -16729
rect 12760 -16763 12794 -16743
rect 12760 -16811 12794 -16801
rect 12760 -16835 12794 -16811
rect 12760 -16879 12794 -16873
rect 12760 -16907 12794 -16879
rect 12760 -16947 12794 -16945
rect 12760 -16979 12794 -16947
rect 12760 -17049 12794 -17017
rect 12760 -17051 12794 -17049
rect 12760 -17117 12794 -17089
rect 12760 -17123 12794 -17117
rect 12760 -17185 12794 -17161
rect 12760 -17195 12794 -17185
rect 12760 -17253 12794 -17233
rect 12760 -17267 12794 -17253
rect 13778 -16743 13812 -16729
rect 13778 -16763 13812 -16743
rect 13778 -16811 13812 -16801
rect 13778 -16835 13812 -16811
rect 13778 -16879 13812 -16873
rect 13778 -16907 13812 -16879
rect 13778 -16947 13812 -16945
rect 13778 -16979 13812 -16947
rect 13778 -17049 13812 -17017
rect 13778 -17051 13812 -17049
rect 13778 -17117 13812 -17089
rect 13778 -17123 13812 -17117
rect 13778 -17185 13812 -17161
rect 13778 -17195 13812 -17185
rect 13778 -17253 13812 -17233
rect 13778 -17267 13812 -17253
rect 14796 -16743 14830 -16729
rect 14796 -16763 14830 -16743
rect 14796 -16811 14830 -16801
rect 14796 -16835 14830 -16811
rect 14796 -16879 14830 -16873
rect 14796 -16907 14830 -16879
rect 14796 -16947 14830 -16945
rect 14796 -16979 14830 -16947
rect 14796 -17049 14830 -17017
rect 14796 -17051 14830 -17049
rect 14796 -17117 14830 -17089
rect 14796 -17123 14830 -17117
rect 14796 -17185 14830 -17161
rect 14796 -17195 14830 -17185
rect 14796 -17253 14830 -17233
rect 14796 -17267 14830 -17253
rect 15814 -16743 15848 -16729
rect 15814 -16763 15848 -16743
rect 15814 -16811 15848 -16801
rect 15814 -16835 15848 -16811
rect 15814 -16879 15848 -16873
rect 15814 -16907 15848 -16879
rect 15814 -16947 15848 -16945
rect 15814 -16979 15848 -16947
rect 15814 -17049 15848 -17017
rect 15814 -17051 15848 -17049
rect 15814 -17117 15848 -17089
rect 15814 -17123 15848 -17117
rect 15814 -17185 15848 -17161
rect 15814 -17195 15848 -17185
rect 15814 -17253 15848 -17233
rect 15814 -17267 15848 -17253
rect 16832 -16743 16866 -16729
rect 16832 -16763 16866 -16743
rect 16832 -16811 16866 -16801
rect 16832 -16835 16866 -16811
rect 16832 -16879 16866 -16873
rect 16832 -16907 16866 -16879
rect 16832 -16947 16866 -16945
rect 16832 -16979 16866 -16947
rect 16832 -17049 16866 -17017
rect 16832 -17051 16866 -17049
rect 16832 -17117 16866 -17089
rect 16832 -17123 16866 -17117
rect 16832 -17185 16866 -17161
rect 16832 -17195 16866 -17185
rect 16832 -17253 16866 -17233
rect 16832 -17267 16866 -17253
rect 17850 -16743 17884 -16729
rect 17850 -16763 17884 -16743
rect 17850 -16811 17884 -16801
rect 17850 -16835 17884 -16811
rect 17850 -16879 17884 -16873
rect 17850 -16907 17884 -16879
rect 17850 -16947 17884 -16945
rect 17850 -16979 17884 -16947
rect 17850 -17049 17884 -17017
rect 17850 -17051 17884 -17049
rect 17850 -17117 17884 -17089
rect 17850 -17123 17884 -17117
rect 17850 -17185 17884 -17161
rect 17850 -17195 17884 -17185
rect 17850 -17253 17884 -17233
rect 17850 -17267 17884 -17253
rect 18868 -16743 18902 -16729
rect 18868 -16763 18902 -16743
rect 18868 -16811 18902 -16801
rect 18868 -16835 18902 -16811
rect 18868 -16879 18902 -16873
rect 18868 -16907 18902 -16879
rect 18868 -16947 18902 -16945
rect 18868 -16979 18902 -16947
rect 18868 -17049 18902 -17017
rect 18868 -17051 18902 -17049
rect 18868 -17117 18902 -17089
rect 18868 -17123 18902 -17117
rect 18868 -17185 18902 -17161
rect 18868 -17195 18902 -17185
rect 18868 -17253 18902 -17233
rect 18868 -17267 18902 -17253
rect 19886 -16743 19920 -16729
rect 19886 -16763 19920 -16743
rect 19886 -16811 19920 -16801
rect 19886 -16835 19920 -16811
rect 19886 -16879 19920 -16873
rect 19886 -16907 19920 -16879
rect 19886 -16947 19920 -16945
rect 19886 -16979 19920 -16947
rect 19886 -17049 19920 -17017
rect 19886 -17051 19920 -17049
rect 19886 -17117 19920 -17089
rect 19886 -17123 19920 -17117
rect 19886 -17185 19920 -17161
rect 19886 -17195 19920 -17185
rect 19886 -17253 19920 -17233
rect 19886 -17267 19920 -17253
rect 20904 -16743 20938 -16729
rect 20904 -16763 20938 -16743
rect 20904 -16811 20938 -16801
rect 20904 -16835 20938 -16811
rect 20904 -16879 20938 -16873
rect 20904 -16907 20938 -16879
rect 20904 -16947 20938 -16945
rect 20904 -16979 20938 -16947
rect 20904 -17049 20938 -17017
rect 20904 -17051 20938 -17049
rect 20904 -17117 20938 -17089
rect 20904 -17123 20938 -17117
rect 20904 -17185 20938 -17161
rect 20904 -17195 20938 -17185
rect 20904 -17253 20938 -17233
rect 20904 -17267 20938 -17253
rect 21922 -16743 21956 -16729
rect 21922 -16763 21956 -16743
rect 21922 -16811 21956 -16801
rect 21922 -16835 21956 -16811
rect 21922 -16879 21956 -16873
rect 21922 -16907 21956 -16879
rect 21922 -16947 21956 -16945
rect 21922 -16979 21956 -16947
rect 21922 -17049 21956 -17017
rect 21922 -17051 21956 -17049
rect 21922 -17117 21956 -17089
rect 21922 -17123 21956 -17117
rect 21922 -17185 21956 -17161
rect 21922 -17195 21956 -17185
rect 21922 -17253 21956 -17233
rect 21922 -17267 21956 -17253
rect 22940 -16743 22974 -16729
rect 22940 -16763 22974 -16743
rect 22940 -16811 22974 -16801
rect 22940 -16835 22974 -16811
rect 22940 -16879 22974 -16873
rect 22940 -16907 22974 -16879
rect 22940 -16947 22974 -16945
rect 22940 -16979 22974 -16947
rect 22940 -17049 22974 -17017
rect 22940 -17051 22974 -17049
rect 22940 -17117 22974 -17089
rect 22940 -17123 22974 -17117
rect 22940 -17185 22974 -17161
rect 22940 -17195 22974 -17185
rect 22940 -17253 22974 -17233
rect 22940 -17267 22974 -17253
rect 24855 -16701 24889 -16699
rect 24855 -16733 24889 -16701
rect 24855 -16803 24889 -16771
rect 24855 -16805 24889 -16803
rect 24855 -16871 24889 -16843
rect 24855 -16877 24889 -16871
rect 24855 -16939 24889 -16915
rect 24855 -16949 24889 -16939
rect 24855 -17007 24889 -16987
rect 24855 -17021 24889 -17007
rect 24855 -17075 24889 -17059
rect 24855 -17093 24889 -17075
rect 24855 -17143 24889 -17131
rect 24855 -17165 24889 -17143
rect 24855 -17211 24889 -17203
rect 24855 -17237 24889 -17211
rect 24855 -17279 24889 -17275
rect 24855 -17309 24889 -17279
rect -12289 -17381 -12255 -17347
rect -8855 -17382 -8845 -17348
rect -8845 -17382 -8821 -17348
rect -8783 -17382 -8777 -17348
rect -8777 -17382 -8749 -17348
rect -8711 -17382 -8709 -17348
rect -8709 -17382 -8677 -17348
rect -8639 -17382 -8607 -17348
rect -8607 -17382 -8605 -17348
rect -8567 -17382 -8539 -17348
rect -8539 -17382 -8533 -17348
rect -8495 -17382 -8471 -17348
rect -8471 -17382 -8461 -17348
rect -7837 -17382 -7827 -17348
rect -7827 -17382 -7803 -17348
rect -7765 -17382 -7759 -17348
rect -7759 -17382 -7731 -17348
rect -7693 -17382 -7691 -17348
rect -7691 -17382 -7659 -17348
rect -7621 -17382 -7589 -17348
rect -7589 -17382 -7587 -17348
rect -7549 -17382 -7521 -17348
rect -7521 -17382 -7515 -17348
rect -7477 -17382 -7453 -17348
rect -7453 -17382 -7443 -17348
rect -6819 -17382 -6809 -17348
rect -6809 -17382 -6785 -17348
rect -6747 -17382 -6741 -17348
rect -6741 -17382 -6713 -17348
rect -6675 -17382 -6673 -17348
rect -6673 -17382 -6641 -17348
rect -6603 -17382 -6571 -17348
rect -6571 -17382 -6569 -17348
rect -6531 -17382 -6503 -17348
rect -6503 -17382 -6497 -17348
rect -6459 -17382 -6435 -17348
rect -6435 -17382 -6425 -17348
rect -5801 -17382 -5791 -17348
rect -5791 -17382 -5767 -17348
rect -5729 -17382 -5723 -17348
rect -5723 -17382 -5695 -17348
rect -5657 -17382 -5655 -17348
rect -5655 -17382 -5623 -17348
rect -5585 -17382 -5553 -17348
rect -5553 -17382 -5551 -17348
rect -5513 -17382 -5485 -17348
rect -5485 -17382 -5479 -17348
rect -5441 -17382 -5417 -17348
rect -5417 -17382 -5407 -17348
rect -4783 -17382 -4773 -17348
rect -4773 -17382 -4749 -17348
rect -4711 -17382 -4705 -17348
rect -4705 -17382 -4677 -17348
rect -4639 -17382 -4637 -17348
rect -4637 -17382 -4605 -17348
rect -4567 -17382 -4535 -17348
rect -4535 -17382 -4533 -17348
rect -4495 -17382 -4467 -17348
rect -4467 -17382 -4461 -17348
rect -4423 -17382 -4399 -17348
rect -4399 -17382 -4389 -17348
rect -3765 -17382 -3755 -17348
rect -3755 -17382 -3731 -17348
rect -3693 -17382 -3687 -17348
rect -3687 -17382 -3659 -17348
rect -3621 -17382 -3619 -17348
rect -3619 -17382 -3587 -17348
rect -3549 -17382 -3517 -17348
rect -3517 -17382 -3515 -17348
rect -3477 -17382 -3449 -17348
rect -3449 -17382 -3443 -17348
rect -3405 -17382 -3381 -17348
rect -3381 -17382 -3371 -17348
rect -2747 -17382 -2737 -17348
rect -2737 -17382 -2713 -17348
rect -2675 -17382 -2669 -17348
rect -2669 -17382 -2641 -17348
rect -2603 -17382 -2601 -17348
rect -2601 -17382 -2569 -17348
rect -2531 -17382 -2499 -17348
rect -2499 -17382 -2497 -17348
rect -2459 -17382 -2431 -17348
rect -2431 -17382 -2425 -17348
rect -2387 -17382 -2363 -17348
rect -2363 -17382 -2353 -17348
rect -1729 -17382 -1719 -17348
rect -1719 -17382 -1695 -17348
rect -1657 -17382 -1651 -17348
rect -1651 -17382 -1623 -17348
rect -1585 -17382 -1583 -17348
rect -1583 -17382 -1551 -17348
rect -1513 -17382 -1481 -17348
rect -1481 -17382 -1479 -17348
rect -1441 -17382 -1413 -17348
rect -1413 -17382 -1407 -17348
rect -1369 -17382 -1345 -17348
rect -1345 -17382 -1335 -17348
rect -711 -17382 -701 -17348
rect -701 -17382 -677 -17348
rect -639 -17382 -633 -17348
rect -633 -17382 -605 -17348
rect -567 -17382 -565 -17348
rect -565 -17382 -533 -17348
rect -495 -17382 -463 -17348
rect -463 -17382 -461 -17348
rect -423 -17382 -395 -17348
rect -395 -17382 -389 -17348
rect -351 -17382 -327 -17348
rect -327 -17382 -317 -17348
rect 2909 -17370 2919 -17336
rect 2919 -17370 2943 -17336
rect 2981 -17370 2987 -17336
rect 2987 -17370 3015 -17336
rect 3053 -17370 3055 -17336
rect 3055 -17370 3087 -17336
rect 3125 -17370 3157 -17336
rect 3157 -17370 3159 -17336
rect 3197 -17370 3225 -17336
rect 3225 -17370 3231 -17336
rect 3269 -17370 3293 -17336
rect 3293 -17370 3303 -17336
rect 3927 -17370 3937 -17336
rect 3937 -17370 3961 -17336
rect 3999 -17370 4005 -17336
rect 4005 -17370 4033 -17336
rect 4071 -17370 4073 -17336
rect 4073 -17370 4105 -17336
rect 4143 -17370 4175 -17336
rect 4175 -17370 4177 -17336
rect 4215 -17370 4243 -17336
rect 4243 -17370 4249 -17336
rect 4287 -17370 4311 -17336
rect 4311 -17370 4321 -17336
rect 4945 -17370 4955 -17336
rect 4955 -17370 4979 -17336
rect 5017 -17370 5023 -17336
rect 5023 -17370 5051 -17336
rect 5089 -17370 5091 -17336
rect 5091 -17370 5123 -17336
rect 5161 -17370 5193 -17336
rect 5193 -17370 5195 -17336
rect 5233 -17370 5261 -17336
rect 5261 -17370 5267 -17336
rect 5305 -17370 5329 -17336
rect 5329 -17370 5339 -17336
rect 5963 -17370 5973 -17336
rect 5973 -17370 5997 -17336
rect 6035 -17370 6041 -17336
rect 6041 -17370 6069 -17336
rect 6107 -17370 6109 -17336
rect 6109 -17370 6141 -17336
rect 6179 -17370 6211 -17336
rect 6211 -17370 6213 -17336
rect 6251 -17370 6279 -17336
rect 6279 -17370 6285 -17336
rect 6323 -17370 6347 -17336
rect 6347 -17370 6357 -17336
rect 6981 -17370 6991 -17336
rect 6991 -17370 7015 -17336
rect 7053 -17370 7059 -17336
rect 7059 -17370 7087 -17336
rect 7125 -17370 7127 -17336
rect 7127 -17370 7159 -17336
rect 7197 -17370 7229 -17336
rect 7229 -17370 7231 -17336
rect 7269 -17370 7297 -17336
rect 7297 -17370 7303 -17336
rect 7341 -17370 7365 -17336
rect 7365 -17370 7375 -17336
rect 7999 -17370 8009 -17336
rect 8009 -17370 8033 -17336
rect 8071 -17370 8077 -17336
rect 8077 -17370 8105 -17336
rect 8143 -17370 8145 -17336
rect 8145 -17370 8177 -17336
rect 8215 -17370 8247 -17336
rect 8247 -17370 8249 -17336
rect 8287 -17370 8315 -17336
rect 8315 -17370 8321 -17336
rect 8359 -17370 8383 -17336
rect 8383 -17370 8393 -17336
rect 9017 -17370 9027 -17336
rect 9027 -17370 9051 -17336
rect 9089 -17370 9095 -17336
rect 9095 -17370 9123 -17336
rect 9161 -17370 9163 -17336
rect 9163 -17370 9195 -17336
rect 9233 -17370 9265 -17336
rect 9265 -17370 9267 -17336
rect 9305 -17370 9333 -17336
rect 9333 -17370 9339 -17336
rect 9377 -17370 9401 -17336
rect 9401 -17370 9411 -17336
rect 10035 -17370 10045 -17336
rect 10045 -17370 10069 -17336
rect 10107 -17370 10113 -17336
rect 10113 -17370 10141 -17336
rect 10179 -17370 10181 -17336
rect 10181 -17370 10213 -17336
rect 10251 -17370 10283 -17336
rect 10283 -17370 10285 -17336
rect 10323 -17370 10351 -17336
rect 10351 -17370 10357 -17336
rect 10395 -17370 10419 -17336
rect 10419 -17370 10429 -17336
rect 11053 -17370 11063 -17336
rect 11063 -17370 11087 -17336
rect 11125 -17370 11131 -17336
rect 11131 -17370 11159 -17336
rect 11197 -17370 11199 -17336
rect 11199 -17370 11231 -17336
rect 11269 -17370 11301 -17336
rect 11301 -17370 11303 -17336
rect 11341 -17370 11369 -17336
rect 11369 -17370 11375 -17336
rect 11413 -17370 11437 -17336
rect 11437 -17370 11447 -17336
rect 12071 -17370 12081 -17336
rect 12081 -17370 12105 -17336
rect 12143 -17370 12149 -17336
rect 12149 -17370 12177 -17336
rect 12215 -17370 12217 -17336
rect 12217 -17370 12249 -17336
rect 12287 -17370 12319 -17336
rect 12319 -17370 12321 -17336
rect 12359 -17370 12387 -17336
rect 12387 -17370 12393 -17336
rect 12431 -17370 12455 -17336
rect 12455 -17370 12465 -17336
rect 13089 -17370 13099 -17336
rect 13099 -17370 13123 -17336
rect 13161 -17370 13167 -17336
rect 13167 -17370 13195 -17336
rect 13233 -17370 13235 -17336
rect 13235 -17370 13267 -17336
rect 13305 -17370 13337 -17336
rect 13337 -17370 13339 -17336
rect 13377 -17370 13405 -17336
rect 13405 -17370 13411 -17336
rect 13449 -17370 13473 -17336
rect 13473 -17370 13483 -17336
rect 14107 -17370 14117 -17336
rect 14117 -17370 14141 -17336
rect 14179 -17370 14185 -17336
rect 14185 -17370 14213 -17336
rect 14251 -17370 14253 -17336
rect 14253 -17370 14285 -17336
rect 14323 -17370 14355 -17336
rect 14355 -17370 14357 -17336
rect 14395 -17370 14423 -17336
rect 14423 -17370 14429 -17336
rect 14467 -17370 14491 -17336
rect 14491 -17370 14501 -17336
rect 15125 -17370 15135 -17336
rect 15135 -17370 15159 -17336
rect 15197 -17370 15203 -17336
rect 15203 -17370 15231 -17336
rect 15269 -17370 15271 -17336
rect 15271 -17370 15303 -17336
rect 15341 -17370 15373 -17336
rect 15373 -17370 15375 -17336
rect 15413 -17370 15441 -17336
rect 15441 -17370 15447 -17336
rect 15485 -17370 15509 -17336
rect 15509 -17370 15519 -17336
rect 16143 -17370 16153 -17336
rect 16153 -17370 16177 -17336
rect 16215 -17370 16221 -17336
rect 16221 -17370 16249 -17336
rect 16287 -17370 16289 -17336
rect 16289 -17370 16321 -17336
rect 16359 -17370 16391 -17336
rect 16391 -17370 16393 -17336
rect 16431 -17370 16459 -17336
rect 16459 -17370 16465 -17336
rect 16503 -17370 16527 -17336
rect 16527 -17370 16537 -17336
rect 17161 -17370 17171 -17336
rect 17171 -17370 17195 -17336
rect 17233 -17370 17239 -17336
rect 17239 -17370 17267 -17336
rect 17305 -17370 17307 -17336
rect 17307 -17370 17339 -17336
rect 17377 -17370 17409 -17336
rect 17409 -17370 17411 -17336
rect 17449 -17370 17477 -17336
rect 17477 -17370 17483 -17336
rect 17521 -17370 17545 -17336
rect 17545 -17370 17555 -17336
rect 18179 -17370 18189 -17336
rect 18189 -17370 18213 -17336
rect 18251 -17370 18257 -17336
rect 18257 -17370 18285 -17336
rect 18323 -17370 18325 -17336
rect 18325 -17370 18357 -17336
rect 18395 -17370 18427 -17336
rect 18427 -17370 18429 -17336
rect 18467 -17370 18495 -17336
rect 18495 -17370 18501 -17336
rect 18539 -17370 18563 -17336
rect 18563 -17370 18573 -17336
rect 19197 -17370 19207 -17336
rect 19207 -17370 19231 -17336
rect 19269 -17370 19275 -17336
rect 19275 -17370 19303 -17336
rect 19341 -17370 19343 -17336
rect 19343 -17370 19375 -17336
rect 19413 -17370 19445 -17336
rect 19445 -17370 19447 -17336
rect 19485 -17370 19513 -17336
rect 19513 -17370 19519 -17336
rect 19557 -17370 19581 -17336
rect 19581 -17370 19591 -17336
rect 20215 -17370 20225 -17336
rect 20225 -17370 20249 -17336
rect 20287 -17370 20293 -17336
rect 20293 -17370 20321 -17336
rect 20359 -17370 20361 -17336
rect 20361 -17370 20393 -17336
rect 20431 -17370 20463 -17336
rect 20463 -17370 20465 -17336
rect 20503 -17370 20531 -17336
rect 20531 -17370 20537 -17336
rect 20575 -17370 20599 -17336
rect 20599 -17370 20609 -17336
rect 21233 -17370 21243 -17336
rect 21243 -17370 21267 -17336
rect 21305 -17370 21311 -17336
rect 21311 -17370 21339 -17336
rect 21377 -17370 21379 -17336
rect 21379 -17370 21411 -17336
rect 21449 -17370 21481 -17336
rect 21481 -17370 21483 -17336
rect 21521 -17370 21549 -17336
rect 21549 -17370 21555 -17336
rect 21593 -17370 21617 -17336
rect 21617 -17370 21627 -17336
rect 22251 -17370 22261 -17336
rect 22261 -17370 22285 -17336
rect 22323 -17370 22329 -17336
rect 22329 -17370 22357 -17336
rect 22395 -17370 22397 -17336
rect 22397 -17370 22429 -17336
rect 22467 -17370 22499 -17336
rect 22499 -17370 22501 -17336
rect 22539 -17370 22567 -17336
rect 22567 -17370 22573 -17336
rect 22611 -17370 22635 -17336
rect 22635 -17370 22645 -17336
rect 24855 -17381 24889 -17347
rect -12289 -17449 -12255 -17419
rect -12289 -17453 -12255 -17449
rect -12289 -17517 -12255 -17491
rect -12289 -17525 -12255 -17517
rect -12289 -17585 -12255 -17563
rect -12289 -17597 -12255 -17585
rect -12289 -17653 -12255 -17635
rect -12289 -17669 -12255 -17653
rect -12289 -17721 -12255 -17707
rect -12289 -17741 -12255 -17721
rect -12289 -17789 -12255 -17779
rect -12289 -17813 -12255 -17789
rect -12289 -17857 -12255 -17851
rect -12289 -17885 -12255 -17857
rect -12289 -17925 -12255 -17923
rect -12289 -17957 -12255 -17925
rect -12289 -18027 -12255 -17995
rect -12289 -18029 -12255 -18027
rect -9184 -17465 -9150 -17451
rect -9184 -17485 -9150 -17465
rect -9184 -17533 -9150 -17523
rect -9184 -17557 -9150 -17533
rect -9184 -17601 -9150 -17595
rect -9184 -17629 -9150 -17601
rect -9184 -17669 -9150 -17667
rect -9184 -17701 -9150 -17669
rect -9184 -17771 -9150 -17739
rect -9184 -17773 -9150 -17771
rect -9184 -17839 -9150 -17811
rect -9184 -17845 -9150 -17839
rect -9184 -17907 -9150 -17883
rect -9184 -17917 -9150 -17907
rect -9184 -17975 -9150 -17955
rect -9184 -17989 -9150 -17975
rect -8166 -17465 -8132 -17451
rect -8166 -17485 -8132 -17465
rect -8166 -17533 -8132 -17523
rect -8166 -17557 -8132 -17533
rect -8166 -17601 -8132 -17595
rect -8166 -17629 -8132 -17601
rect -8166 -17669 -8132 -17667
rect -8166 -17701 -8132 -17669
rect -8166 -17771 -8132 -17739
rect -8166 -17773 -8132 -17771
rect -8166 -17839 -8132 -17811
rect -8166 -17845 -8132 -17839
rect -8166 -17907 -8132 -17883
rect -8166 -17917 -8132 -17907
rect -8166 -17975 -8132 -17955
rect -8166 -17989 -8132 -17975
rect -7148 -17465 -7114 -17451
rect -7148 -17485 -7114 -17465
rect -7148 -17533 -7114 -17523
rect -7148 -17557 -7114 -17533
rect -7148 -17601 -7114 -17595
rect -7148 -17629 -7114 -17601
rect -7148 -17669 -7114 -17667
rect -7148 -17701 -7114 -17669
rect -7148 -17771 -7114 -17739
rect -7148 -17773 -7114 -17771
rect -7148 -17839 -7114 -17811
rect -7148 -17845 -7114 -17839
rect -7148 -17907 -7114 -17883
rect -7148 -17917 -7114 -17907
rect -7148 -17975 -7114 -17955
rect -7148 -17989 -7114 -17975
rect -6130 -17465 -6096 -17451
rect -6130 -17485 -6096 -17465
rect -6130 -17533 -6096 -17523
rect -6130 -17557 -6096 -17533
rect -6130 -17601 -6096 -17595
rect -6130 -17629 -6096 -17601
rect -6130 -17669 -6096 -17667
rect -6130 -17701 -6096 -17669
rect -6130 -17771 -6096 -17739
rect -6130 -17773 -6096 -17771
rect -6130 -17839 -6096 -17811
rect -6130 -17845 -6096 -17839
rect -6130 -17907 -6096 -17883
rect -6130 -17917 -6096 -17907
rect -6130 -17975 -6096 -17955
rect -6130 -17989 -6096 -17975
rect -5112 -17465 -5078 -17451
rect -5112 -17485 -5078 -17465
rect -5112 -17533 -5078 -17523
rect -5112 -17557 -5078 -17533
rect -5112 -17601 -5078 -17595
rect -5112 -17629 -5078 -17601
rect -5112 -17669 -5078 -17667
rect -5112 -17701 -5078 -17669
rect -5112 -17771 -5078 -17739
rect -5112 -17773 -5078 -17771
rect -5112 -17839 -5078 -17811
rect -5112 -17845 -5078 -17839
rect -5112 -17907 -5078 -17883
rect -5112 -17917 -5078 -17907
rect -5112 -17975 -5078 -17955
rect -5112 -17989 -5078 -17975
rect -4094 -17465 -4060 -17451
rect -4094 -17485 -4060 -17465
rect -4094 -17533 -4060 -17523
rect -4094 -17557 -4060 -17533
rect -4094 -17601 -4060 -17595
rect -4094 -17629 -4060 -17601
rect -4094 -17669 -4060 -17667
rect -4094 -17701 -4060 -17669
rect -4094 -17771 -4060 -17739
rect -4094 -17773 -4060 -17771
rect -4094 -17839 -4060 -17811
rect -4094 -17845 -4060 -17839
rect -4094 -17907 -4060 -17883
rect -4094 -17917 -4060 -17907
rect -4094 -17975 -4060 -17955
rect -4094 -17989 -4060 -17975
rect -3076 -17465 -3042 -17451
rect -3076 -17485 -3042 -17465
rect -3076 -17533 -3042 -17523
rect -3076 -17557 -3042 -17533
rect -3076 -17601 -3042 -17595
rect -3076 -17629 -3042 -17601
rect -3076 -17669 -3042 -17667
rect -3076 -17701 -3042 -17669
rect -3076 -17771 -3042 -17739
rect -3076 -17773 -3042 -17771
rect -3076 -17839 -3042 -17811
rect -3076 -17845 -3042 -17839
rect -3076 -17907 -3042 -17883
rect -3076 -17917 -3042 -17907
rect -3076 -17975 -3042 -17955
rect -3076 -17989 -3042 -17975
rect -2058 -17465 -2024 -17451
rect -2058 -17485 -2024 -17465
rect -2058 -17533 -2024 -17523
rect -2058 -17557 -2024 -17533
rect -2058 -17601 -2024 -17595
rect -2058 -17629 -2024 -17601
rect -2058 -17669 -2024 -17667
rect -2058 -17701 -2024 -17669
rect -2058 -17771 -2024 -17739
rect -2058 -17773 -2024 -17771
rect -2058 -17839 -2024 -17811
rect -2058 -17845 -2024 -17839
rect -2058 -17907 -2024 -17883
rect -2058 -17917 -2024 -17907
rect -2058 -17975 -2024 -17955
rect -2058 -17989 -2024 -17975
rect -1040 -17465 -1006 -17451
rect -1040 -17485 -1006 -17465
rect -1040 -17533 -1006 -17523
rect -1040 -17557 -1006 -17533
rect -1040 -17601 -1006 -17595
rect -1040 -17629 -1006 -17601
rect -1040 -17669 -1006 -17667
rect -1040 -17701 -1006 -17669
rect -1040 -17771 -1006 -17739
rect -1040 -17773 -1006 -17771
rect -1040 -17839 -1006 -17811
rect -1040 -17845 -1006 -17839
rect -1040 -17907 -1006 -17883
rect -1040 -17917 -1006 -17907
rect -1040 -17975 -1006 -17955
rect -1040 -17989 -1006 -17975
rect -22 -17465 12 -17451
rect -22 -17485 12 -17465
rect -22 -17533 12 -17523
rect -22 -17557 12 -17533
rect -22 -17601 12 -17595
rect -22 -17629 12 -17601
rect -22 -17669 12 -17667
rect -22 -17701 12 -17669
rect -22 -17771 12 -17739
rect -22 -17773 12 -17771
rect -22 -17839 12 -17811
rect -22 -17845 12 -17839
rect 24855 -17449 24889 -17419
rect 24855 -17453 24889 -17449
rect 24855 -17517 24889 -17491
rect 24855 -17525 24889 -17517
rect 24855 -17585 24889 -17563
rect 24855 -17597 24889 -17585
rect 24855 -17653 24889 -17635
rect 24855 -17669 24889 -17653
rect 24855 -17721 24889 -17707
rect 24855 -17741 24889 -17721
rect 24855 -17789 24889 -17779
rect 24855 -17813 24889 -17789
rect -22 -17907 12 -17883
rect 2909 -17894 2919 -17860
rect 2919 -17894 2943 -17860
rect 2981 -17894 2987 -17860
rect 2987 -17894 3015 -17860
rect 3053 -17894 3055 -17860
rect 3055 -17894 3087 -17860
rect 3125 -17894 3157 -17860
rect 3157 -17894 3159 -17860
rect 3197 -17894 3225 -17860
rect 3225 -17894 3231 -17860
rect 3269 -17894 3293 -17860
rect 3293 -17894 3303 -17860
rect 3927 -17894 3937 -17860
rect 3937 -17894 3961 -17860
rect 3999 -17894 4005 -17860
rect 4005 -17894 4033 -17860
rect 4071 -17894 4073 -17860
rect 4073 -17894 4105 -17860
rect 4143 -17894 4175 -17860
rect 4175 -17894 4177 -17860
rect 4215 -17894 4243 -17860
rect 4243 -17894 4249 -17860
rect 4287 -17894 4311 -17860
rect 4311 -17894 4321 -17860
rect 4945 -17894 4955 -17860
rect 4955 -17894 4979 -17860
rect 5017 -17894 5023 -17860
rect 5023 -17894 5051 -17860
rect 5089 -17894 5091 -17860
rect 5091 -17894 5123 -17860
rect 5161 -17894 5193 -17860
rect 5193 -17894 5195 -17860
rect 5233 -17894 5261 -17860
rect 5261 -17894 5267 -17860
rect 5305 -17894 5329 -17860
rect 5329 -17894 5339 -17860
rect 5963 -17894 5973 -17860
rect 5973 -17894 5997 -17860
rect 6035 -17894 6041 -17860
rect 6041 -17894 6069 -17860
rect 6107 -17894 6109 -17860
rect 6109 -17894 6141 -17860
rect 6179 -17894 6211 -17860
rect 6211 -17894 6213 -17860
rect 6251 -17894 6279 -17860
rect 6279 -17894 6285 -17860
rect 6323 -17894 6347 -17860
rect 6347 -17894 6357 -17860
rect 6981 -17894 6991 -17860
rect 6991 -17894 7015 -17860
rect 7053 -17894 7059 -17860
rect 7059 -17894 7087 -17860
rect 7125 -17894 7127 -17860
rect 7127 -17894 7159 -17860
rect 7197 -17894 7229 -17860
rect 7229 -17894 7231 -17860
rect 7269 -17894 7297 -17860
rect 7297 -17894 7303 -17860
rect 7341 -17894 7365 -17860
rect 7365 -17894 7375 -17860
rect 7999 -17894 8009 -17860
rect 8009 -17894 8033 -17860
rect 8071 -17894 8077 -17860
rect 8077 -17894 8105 -17860
rect 8143 -17894 8145 -17860
rect 8145 -17894 8177 -17860
rect 8215 -17894 8247 -17860
rect 8247 -17894 8249 -17860
rect 8287 -17894 8315 -17860
rect 8315 -17894 8321 -17860
rect 8359 -17894 8383 -17860
rect 8383 -17894 8393 -17860
rect 9017 -17894 9027 -17860
rect 9027 -17894 9051 -17860
rect 9089 -17894 9095 -17860
rect 9095 -17894 9123 -17860
rect 9161 -17894 9163 -17860
rect 9163 -17894 9195 -17860
rect 9233 -17894 9265 -17860
rect 9265 -17894 9267 -17860
rect 9305 -17894 9333 -17860
rect 9333 -17894 9339 -17860
rect 9377 -17894 9401 -17860
rect 9401 -17894 9411 -17860
rect 10035 -17894 10045 -17860
rect 10045 -17894 10069 -17860
rect 10107 -17894 10113 -17860
rect 10113 -17894 10141 -17860
rect 10179 -17894 10181 -17860
rect 10181 -17894 10213 -17860
rect 10251 -17894 10283 -17860
rect 10283 -17894 10285 -17860
rect 10323 -17894 10351 -17860
rect 10351 -17894 10357 -17860
rect 10395 -17894 10419 -17860
rect 10419 -17894 10429 -17860
rect 11053 -17894 11063 -17860
rect 11063 -17894 11087 -17860
rect 11125 -17894 11131 -17860
rect 11131 -17894 11159 -17860
rect 11197 -17894 11199 -17860
rect 11199 -17894 11231 -17860
rect 11269 -17894 11301 -17860
rect 11301 -17894 11303 -17860
rect 11341 -17894 11369 -17860
rect 11369 -17894 11375 -17860
rect 11413 -17894 11437 -17860
rect 11437 -17894 11447 -17860
rect 12071 -17894 12081 -17860
rect 12081 -17894 12105 -17860
rect 12143 -17894 12149 -17860
rect 12149 -17894 12177 -17860
rect 12215 -17894 12217 -17860
rect 12217 -17894 12249 -17860
rect 12287 -17894 12319 -17860
rect 12319 -17894 12321 -17860
rect 12359 -17894 12387 -17860
rect 12387 -17894 12393 -17860
rect 12431 -17894 12455 -17860
rect 12455 -17894 12465 -17860
rect 13089 -17894 13099 -17860
rect 13099 -17894 13123 -17860
rect 13161 -17894 13167 -17860
rect 13167 -17894 13195 -17860
rect 13233 -17894 13235 -17860
rect 13235 -17894 13267 -17860
rect 13305 -17894 13337 -17860
rect 13337 -17894 13339 -17860
rect 13377 -17894 13405 -17860
rect 13405 -17894 13411 -17860
rect 13449 -17894 13473 -17860
rect 13473 -17894 13483 -17860
rect 14107 -17894 14117 -17860
rect 14117 -17894 14141 -17860
rect 14179 -17894 14185 -17860
rect 14185 -17894 14213 -17860
rect 14251 -17894 14253 -17860
rect 14253 -17894 14285 -17860
rect 14323 -17894 14355 -17860
rect 14355 -17894 14357 -17860
rect 14395 -17894 14423 -17860
rect 14423 -17894 14429 -17860
rect 14467 -17894 14491 -17860
rect 14491 -17894 14501 -17860
rect 15125 -17894 15135 -17860
rect 15135 -17894 15159 -17860
rect 15197 -17894 15203 -17860
rect 15203 -17894 15231 -17860
rect 15269 -17894 15271 -17860
rect 15271 -17894 15303 -17860
rect 15341 -17894 15373 -17860
rect 15373 -17894 15375 -17860
rect 15413 -17894 15441 -17860
rect 15441 -17894 15447 -17860
rect 15485 -17894 15509 -17860
rect 15509 -17894 15519 -17860
rect 16143 -17894 16153 -17860
rect 16153 -17894 16177 -17860
rect 16215 -17894 16221 -17860
rect 16221 -17894 16249 -17860
rect 16287 -17894 16289 -17860
rect 16289 -17894 16321 -17860
rect 16359 -17894 16391 -17860
rect 16391 -17894 16393 -17860
rect 16431 -17894 16459 -17860
rect 16459 -17894 16465 -17860
rect 16503 -17894 16527 -17860
rect 16527 -17894 16537 -17860
rect 17161 -17894 17171 -17860
rect 17171 -17894 17195 -17860
rect 17233 -17894 17239 -17860
rect 17239 -17894 17267 -17860
rect 17305 -17894 17307 -17860
rect 17307 -17894 17339 -17860
rect 17377 -17894 17409 -17860
rect 17409 -17894 17411 -17860
rect 17449 -17894 17477 -17860
rect 17477 -17894 17483 -17860
rect 17521 -17894 17545 -17860
rect 17545 -17894 17555 -17860
rect 18179 -17894 18189 -17860
rect 18189 -17894 18213 -17860
rect 18251 -17894 18257 -17860
rect 18257 -17894 18285 -17860
rect 18323 -17894 18325 -17860
rect 18325 -17894 18357 -17860
rect 18395 -17894 18427 -17860
rect 18427 -17894 18429 -17860
rect 18467 -17894 18495 -17860
rect 18495 -17894 18501 -17860
rect 18539 -17894 18563 -17860
rect 18563 -17894 18573 -17860
rect 19197 -17894 19207 -17860
rect 19207 -17894 19231 -17860
rect 19269 -17894 19275 -17860
rect 19275 -17894 19303 -17860
rect 19341 -17894 19343 -17860
rect 19343 -17894 19375 -17860
rect 19413 -17894 19445 -17860
rect 19445 -17894 19447 -17860
rect 19485 -17894 19513 -17860
rect 19513 -17894 19519 -17860
rect 19557 -17894 19581 -17860
rect 19581 -17894 19591 -17860
rect 20215 -17894 20225 -17860
rect 20225 -17894 20249 -17860
rect 20287 -17894 20293 -17860
rect 20293 -17894 20321 -17860
rect 20359 -17894 20361 -17860
rect 20361 -17894 20393 -17860
rect 20431 -17894 20463 -17860
rect 20463 -17894 20465 -17860
rect 20503 -17894 20531 -17860
rect 20531 -17894 20537 -17860
rect 20575 -17894 20599 -17860
rect 20599 -17894 20609 -17860
rect 21233 -17894 21243 -17860
rect 21243 -17894 21267 -17860
rect 21305 -17894 21311 -17860
rect 21311 -17894 21339 -17860
rect 21377 -17894 21379 -17860
rect 21379 -17894 21411 -17860
rect 21449 -17894 21481 -17860
rect 21481 -17894 21483 -17860
rect 21521 -17894 21549 -17860
rect 21549 -17894 21555 -17860
rect 21593 -17894 21617 -17860
rect 21617 -17894 21627 -17860
rect 22251 -17894 22261 -17860
rect 22261 -17894 22285 -17860
rect 22323 -17894 22329 -17860
rect 22329 -17894 22357 -17860
rect 22395 -17894 22397 -17860
rect 22397 -17894 22429 -17860
rect 22467 -17894 22499 -17860
rect 22499 -17894 22501 -17860
rect 22539 -17894 22567 -17860
rect 22567 -17894 22573 -17860
rect 22611 -17894 22635 -17860
rect 22635 -17894 22645 -17860
rect 24855 -17857 24889 -17851
rect 24855 -17885 24889 -17857
rect -22 -17917 12 -17907
rect -22 -17975 12 -17955
rect -22 -17989 12 -17975
rect 2580 -17977 2614 -17963
rect 2580 -17997 2614 -17977
rect 2580 -18045 2614 -18035
rect -12289 -18095 -12255 -18067
rect -12289 -18101 -12255 -18095
rect -8855 -18092 -8845 -18058
rect -8845 -18092 -8821 -18058
rect -8783 -18092 -8777 -18058
rect -8777 -18092 -8749 -18058
rect -8711 -18092 -8709 -18058
rect -8709 -18092 -8677 -18058
rect -8639 -18092 -8607 -18058
rect -8607 -18092 -8605 -18058
rect -8567 -18092 -8539 -18058
rect -8539 -18092 -8533 -18058
rect -8495 -18092 -8471 -18058
rect -8471 -18092 -8461 -18058
rect -7837 -18092 -7827 -18058
rect -7827 -18092 -7803 -18058
rect -7765 -18092 -7759 -18058
rect -7759 -18092 -7731 -18058
rect -7693 -18092 -7691 -18058
rect -7691 -18092 -7659 -18058
rect -7621 -18092 -7589 -18058
rect -7589 -18092 -7587 -18058
rect -7549 -18092 -7521 -18058
rect -7521 -18092 -7515 -18058
rect -7477 -18092 -7453 -18058
rect -7453 -18092 -7443 -18058
rect -6819 -18092 -6809 -18058
rect -6809 -18092 -6785 -18058
rect -6747 -18092 -6741 -18058
rect -6741 -18092 -6713 -18058
rect -6675 -18092 -6673 -18058
rect -6673 -18092 -6641 -18058
rect -6603 -18092 -6571 -18058
rect -6571 -18092 -6569 -18058
rect -6531 -18092 -6503 -18058
rect -6503 -18092 -6497 -18058
rect -6459 -18092 -6435 -18058
rect -6435 -18092 -6425 -18058
rect -5801 -18092 -5791 -18058
rect -5791 -18092 -5767 -18058
rect -5729 -18092 -5723 -18058
rect -5723 -18092 -5695 -18058
rect -5657 -18092 -5655 -18058
rect -5655 -18092 -5623 -18058
rect -5585 -18092 -5553 -18058
rect -5553 -18092 -5551 -18058
rect -5513 -18092 -5485 -18058
rect -5485 -18092 -5479 -18058
rect -5441 -18092 -5417 -18058
rect -5417 -18092 -5407 -18058
rect -4783 -18092 -4773 -18058
rect -4773 -18092 -4749 -18058
rect -4711 -18092 -4705 -18058
rect -4705 -18092 -4677 -18058
rect -4639 -18092 -4637 -18058
rect -4637 -18092 -4605 -18058
rect -4567 -18092 -4535 -18058
rect -4535 -18092 -4533 -18058
rect -4495 -18092 -4467 -18058
rect -4467 -18092 -4461 -18058
rect -4423 -18092 -4399 -18058
rect -4399 -18092 -4389 -18058
rect -3765 -18092 -3755 -18058
rect -3755 -18092 -3731 -18058
rect -3693 -18092 -3687 -18058
rect -3687 -18092 -3659 -18058
rect -3621 -18092 -3619 -18058
rect -3619 -18092 -3587 -18058
rect -3549 -18092 -3517 -18058
rect -3517 -18092 -3515 -18058
rect -3477 -18092 -3449 -18058
rect -3449 -18092 -3443 -18058
rect -3405 -18092 -3381 -18058
rect -3381 -18092 -3371 -18058
rect -2747 -18092 -2737 -18058
rect -2737 -18092 -2713 -18058
rect -2675 -18092 -2669 -18058
rect -2669 -18092 -2641 -18058
rect -2603 -18092 -2601 -18058
rect -2601 -18092 -2569 -18058
rect -2531 -18092 -2499 -18058
rect -2499 -18092 -2497 -18058
rect -2459 -18092 -2431 -18058
rect -2431 -18092 -2425 -18058
rect -2387 -18092 -2363 -18058
rect -2363 -18092 -2353 -18058
rect -1729 -18092 -1719 -18058
rect -1719 -18092 -1695 -18058
rect -1657 -18092 -1651 -18058
rect -1651 -18092 -1623 -18058
rect -1585 -18092 -1583 -18058
rect -1583 -18092 -1551 -18058
rect -1513 -18092 -1481 -18058
rect -1481 -18092 -1479 -18058
rect -1441 -18092 -1413 -18058
rect -1413 -18092 -1407 -18058
rect -1369 -18092 -1345 -18058
rect -1345 -18092 -1335 -18058
rect -711 -18092 -701 -18058
rect -701 -18092 -677 -18058
rect -639 -18092 -633 -18058
rect -633 -18092 -605 -18058
rect -567 -18092 -565 -18058
rect -565 -18092 -533 -18058
rect -495 -18092 -463 -18058
rect -463 -18092 -461 -18058
rect -423 -18092 -395 -18058
rect -395 -18092 -389 -18058
rect -351 -18092 -327 -18058
rect -327 -18092 -317 -18058
rect 2580 -18069 2614 -18045
rect -12289 -18163 -12255 -18139
rect -12289 -18173 -12255 -18163
rect 2580 -18113 2614 -18107
rect 2580 -18141 2614 -18113
rect -8855 -18200 -8845 -18166
rect -8845 -18200 -8821 -18166
rect -8783 -18200 -8777 -18166
rect -8777 -18200 -8749 -18166
rect -8711 -18200 -8709 -18166
rect -8709 -18200 -8677 -18166
rect -8639 -18200 -8607 -18166
rect -8607 -18200 -8605 -18166
rect -8567 -18200 -8539 -18166
rect -8539 -18200 -8533 -18166
rect -8495 -18200 -8471 -18166
rect -8471 -18200 -8461 -18166
rect -7837 -18200 -7827 -18166
rect -7827 -18200 -7803 -18166
rect -7765 -18200 -7759 -18166
rect -7759 -18200 -7731 -18166
rect -7693 -18200 -7691 -18166
rect -7691 -18200 -7659 -18166
rect -7621 -18200 -7589 -18166
rect -7589 -18200 -7587 -18166
rect -7549 -18200 -7521 -18166
rect -7521 -18200 -7515 -18166
rect -7477 -18200 -7453 -18166
rect -7453 -18200 -7443 -18166
rect -6819 -18200 -6809 -18166
rect -6809 -18200 -6785 -18166
rect -6747 -18200 -6741 -18166
rect -6741 -18200 -6713 -18166
rect -6675 -18200 -6673 -18166
rect -6673 -18200 -6641 -18166
rect -6603 -18200 -6571 -18166
rect -6571 -18200 -6569 -18166
rect -6531 -18200 -6503 -18166
rect -6503 -18200 -6497 -18166
rect -6459 -18200 -6435 -18166
rect -6435 -18200 -6425 -18166
rect -5801 -18200 -5791 -18166
rect -5791 -18200 -5767 -18166
rect -5729 -18200 -5723 -18166
rect -5723 -18200 -5695 -18166
rect -5657 -18200 -5655 -18166
rect -5655 -18200 -5623 -18166
rect -5585 -18200 -5553 -18166
rect -5553 -18200 -5551 -18166
rect -5513 -18200 -5485 -18166
rect -5485 -18200 -5479 -18166
rect -5441 -18200 -5417 -18166
rect -5417 -18200 -5407 -18166
rect -4783 -18200 -4773 -18166
rect -4773 -18200 -4749 -18166
rect -4711 -18200 -4705 -18166
rect -4705 -18200 -4677 -18166
rect -4639 -18200 -4637 -18166
rect -4637 -18200 -4605 -18166
rect -4567 -18200 -4535 -18166
rect -4535 -18200 -4533 -18166
rect -4495 -18200 -4467 -18166
rect -4467 -18200 -4461 -18166
rect -4423 -18200 -4399 -18166
rect -4399 -18200 -4389 -18166
rect -3765 -18200 -3755 -18166
rect -3755 -18200 -3731 -18166
rect -3693 -18200 -3687 -18166
rect -3687 -18200 -3659 -18166
rect -3621 -18200 -3619 -18166
rect -3619 -18200 -3587 -18166
rect -3549 -18200 -3517 -18166
rect -3517 -18200 -3515 -18166
rect -3477 -18200 -3449 -18166
rect -3449 -18200 -3443 -18166
rect -3405 -18200 -3381 -18166
rect -3381 -18200 -3371 -18166
rect -2747 -18200 -2737 -18166
rect -2737 -18200 -2713 -18166
rect -2675 -18200 -2669 -18166
rect -2669 -18200 -2641 -18166
rect -2603 -18200 -2601 -18166
rect -2601 -18200 -2569 -18166
rect -2531 -18200 -2499 -18166
rect -2499 -18200 -2497 -18166
rect -2459 -18200 -2431 -18166
rect -2431 -18200 -2425 -18166
rect -2387 -18200 -2363 -18166
rect -2363 -18200 -2353 -18166
rect -1729 -18200 -1719 -18166
rect -1719 -18200 -1695 -18166
rect -1657 -18200 -1651 -18166
rect -1651 -18200 -1623 -18166
rect -1585 -18200 -1583 -18166
rect -1583 -18200 -1551 -18166
rect -1513 -18200 -1481 -18166
rect -1481 -18200 -1479 -18166
rect -1441 -18200 -1413 -18166
rect -1413 -18200 -1407 -18166
rect -1369 -18200 -1345 -18166
rect -1345 -18200 -1335 -18166
rect -711 -18200 -701 -18166
rect -701 -18200 -677 -18166
rect -639 -18200 -633 -18166
rect -633 -18200 -605 -18166
rect -567 -18200 -565 -18166
rect -565 -18200 -533 -18166
rect -495 -18200 -463 -18166
rect -463 -18200 -461 -18166
rect -423 -18200 -395 -18166
rect -395 -18200 -389 -18166
rect -351 -18200 -327 -18166
rect -327 -18200 -317 -18166
rect 2580 -18181 2614 -18179
rect -12289 -18231 -12255 -18211
rect -12289 -18245 -12255 -18231
rect 2580 -18213 2614 -18181
rect -12289 -18299 -12255 -18283
rect -12289 -18317 -12255 -18299
rect -12289 -18367 -12255 -18355
rect -12289 -18389 -12255 -18367
rect -12289 -18435 -12255 -18427
rect -12289 -18461 -12255 -18435
rect -12289 -18503 -12255 -18499
rect -12289 -18533 -12255 -18503
rect -12289 -18605 -12255 -18571
rect -12289 -18673 -12255 -18643
rect -12289 -18677 -12255 -18673
rect -12289 -18741 -12255 -18715
rect -12289 -18749 -12255 -18741
rect -12289 -18809 -12255 -18787
rect -12289 -18821 -12255 -18809
rect -9184 -18283 -9150 -18269
rect -9184 -18303 -9150 -18283
rect -9184 -18351 -9150 -18341
rect -9184 -18375 -9150 -18351
rect -9184 -18419 -9150 -18413
rect -9184 -18447 -9150 -18419
rect -9184 -18487 -9150 -18485
rect -9184 -18519 -9150 -18487
rect -9184 -18589 -9150 -18557
rect -9184 -18591 -9150 -18589
rect -9184 -18657 -9150 -18629
rect -9184 -18663 -9150 -18657
rect -9184 -18725 -9150 -18701
rect -9184 -18735 -9150 -18725
rect -9184 -18793 -9150 -18773
rect -9184 -18807 -9150 -18793
rect -8166 -18283 -8132 -18269
rect -8166 -18303 -8132 -18283
rect -8166 -18351 -8132 -18341
rect -8166 -18375 -8132 -18351
rect -8166 -18419 -8132 -18413
rect -8166 -18447 -8132 -18419
rect -8166 -18487 -8132 -18485
rect -8166 -18519 -8132 -18487
rect -8166 -18589 -8132 -18557
rect -8166 -18591 -8132 -18589
rect -8166 -18657 -8132 -18629
rect -8166 -18663 -8132 -18657
rect -8166 -18725 -8132 -18701
rect -8166 -18735 -8132 -18725
rect -8166 -18793 -8132 -18773
rect -8166 -18807 -8132 -18793
rect -7148 -18283 -7114 -18269
rect -7148 -18303 -7114 -18283
rect -7148 -18351 -7114 -18341
rect -7148 -18375 -7114 -18351
rect -7148 -18419 -7114 -18413
rect -7148 -18447 -7114 -18419
rect -7148 -18487 -7114 -18485
rect -7148 -18519 -7114 -18487
rect -7148 -18589 -7114 -18557
rect -7148 -18591 -7114 -18589
rect -7148 -18657 -7114 -18629
rect -7148 -18663 -7114 -18657
rect -7148 -18725 -7114 -18701
rect -7148 -18735 -7114 -18725
rect -7148 -18793 -7114 -18773
rect -7148 -18807 -7114 -18793
rect -6130 -18283 -6096 -18269
rect -6130 -18303 -6096 -18283
rect -6130 -18351 -6096 -18341
rect -6130 -18375 -6096 -18351
rect -6130 -18419 -6096 -18413
rect -6130 -18447 -6096 -18419
rect -6130 -18487 -6096 -18485
rect -6130 -18519 -6096 -18487
rect -6130 -18589 -6096 -18557
rect -6130 -18591 -6096 -18589
rect -6130 -18657 -6096 -18629
rect -6130 -18663 -6096 -18657
rect -6130 -18725 -6096 -18701
rect -6130 -18735 -6096 -18725
rect -6130 -18793 -6096 -18773
rect -6130 -18807 -6096 -18793
rect -5112 -18283 -5078 -18269
rect -5112 -18303 -5078 -18283
rect -5112 -18351 -5078 -18341
rect -5112 -18375 -5078 -18351
rect -5112 -18419 -5078 -18413
rect -5112 -18447 -5078 -18419
rect -5112 -18487 -5078 -18485
rect -5112 -18519 -5078 -18487
rect -5112 -18589 -5078 -18557
rect -5112 -18591 -5078 -18589
rect -5112 -18657 -5078 -18629
rect -5112 -18663 -5078 -18657
rect -5112 -18725 -5078 -18701
rect -5112 -18735 -5078 -18725
rect -5112 -18793 -5078 -18773
rect -5112 -18807 -5078 -18793
rect -4094 -18283 -4060 -18269
rect -4094 -18303 -4060 -18283
rect -4094 -18351 -4060 -18341
rect -4094 -18375 -4060 -18351
rect -4094 -18419 -4060 -18413
rect -4094 -18447 -4060 -18419
rect -4094 -18487 -4060 -18485
rect -4094 -18519 -4060 -18487
rect -4094 -18589 -4060 -18557
rect -4094 -18591 -4060 -18589
rect -4094 -18657 -4060 -18629
rect -4094 -18663 -4060 -18657
rect -4094 -18725 -4060 -18701
rect -4094 -18735 -4060 -18725
rect -4094 -18793 -4060 -18773
rect -4094 -18807 -4060 -18793
rect -3076 -18283 -3042 -18269
rect -3076 -18303 -3042 -18283
rect -3076 -18351 -3042 -18341
rect -3076 -18375 -3042 -18351
rect -3076 -18419 -3042 -18413
rect -3076 -18447 -3042 -18419
rect -3076 -18487 -3042 -18485
rect -3076 -18519 -3042 -18487
rect -3076 -18589 -3042 -18557
rect -3076 -18591 -3042 -18589
rect -3076 -18657 -3042 -18629
rect -3076 -18663 -3042 -18657
rect -3076 -18725 -3042 -18701
rect -3076 -18735 -3042 -18725
rect -3076 -18793 -3042 -18773
rect -3076 -18807 -3042 -18793
rect -2058 -18283 -2024 -18269
rect -2058 -18303 -2024 -18283
rect -2058 -18351 -2024 -18341
rect -2058 -18375 -2024 -18351
rect -2058 -18419 -2024 -18413
rect -2058 -18447 -2024 -18419
rect -2058 -18487 -2024 -18485
rect -2058 -18519 -2024 -18487
rect -2058 -18589 -2024 -18557
rect -2058 -18591 -2024 -18589
rect -2058 -18657 -2024 -18629
rect -2058 -18663 -2024 -18657
rect -2058 -18725 -2024 -18701
rect -2058 -18735 -2024 -18725
rect -2058 -18793 -2024 -18773
rect -2058 -18807 -2024 -18793
rect -1040 -18283 -1006 -18269
rect -1040 -18303 -1006 -18283
rect -1040 -18351 -1006 -18341
rect -1040 -18375 -1006 -18351
rect -1040 -18419 -1006 -18413
rect -1040 -18447 -1006 -18419
rect -1040 -18487 -1006 -18485
rect -1040 -18519 -1006 -18487
rect -1040 -18589 -1006 -18557
rect -1040 -18591 -1006 -18589
rect -1040 -18657 -1006 -18629
rect -1040 -18663 -1006 -18657
rect -1040 -18725 -1006 -18701
rect -1040 -18735 -1006 -18725
rect -1040 -18793 -1006 -18773
rect -1040 -18807 -1006 -18793
rect -22 -18283 12 -18269
rect -22 -18303 12 -18283
rect -22 -18351 12 -18341
rect -22 -18375 12 -18351
rect -22 -18419 12 -18413
rect -22 -18447 12 -18419
rect -22 -18487 12 -18485
rect -22 -18519 12 -18487
rect 2580 -18283 2614 -18251
rect 2580 -18285 2614 -18283
rect 2580 -18351 2614 -18323
rect 2580 -18357 2614 -18351
rect 2580 -18419 2614 -18395
rect 2580 -18429 2614 -18419
rect 2580 -18487 2614 -18467
rect 2580 -18501 2614 -18487
rect 3598 -17977 3632 -17963
rect 3598 -17997 3632 -17977
rect 3598 -18045 3632 -18035
rect 3598 -18069 3632 -18045
rect 3598 -18113 3632 -18107
rect 3598 -18141 3632 -18113
rect 3598 -18181 3632 -18179
rect 3598 -18213 3632 -18181
rect 3598 -18283 3632 -18251
rect 3598 -18285 3632 -18283
rect 3598 -18351 3632 -18323
rect 3598 -18357 3632 -18351
rect 3598 -18419 3632 -18395
rect 3598 -18429 3632 -18419
rect 3598 -18487 3632 -18467
rect 3598 -18501 3632 -18487
rect 4616 -17977 4650 -17963
rect 4616 -17997 4650 -17977
rect 4616 -18045 4650 -18035
rect 4616 -18069 4650 -18045
rect 4616 -18113 4650 -18107
rect 4616 -18141 4650 -18113
rect 4616 -18181 4650 -18179
rect 4616 -18213 4650 -18181
rect 4616 -18283 4650 -18251
rect 4616 -18285 4650 -18283
rect 4616 -18351 4650 -18323
rect 4616 -18357 4650 -18351
rect 4616 -18419 4650 -18395
rect 4616 -18429 4650 -18419
rect 4616 -18487 4650 -18467
rect 4616 -18501 4650 -18487
rect 5634 -17977 5668 -17963
rect 5634 -17997 5668 -17977
rect 5634 -18045 5668 -18035
rect 5634 -18069 5668 -18045
rect 5634 -18113 5668 -18107
rect 5634 -18141 5668 -18113
rect 5634 -18181 5668 -18179
rect 5634 -18213 5668 -18181
rect 5634 -18283 5668 -18251
rect 5634 -18285 5668 -18283
rect 5634 -18351 5668 -18323
rect 5634 -18357 5668 -18351
rect 5634 -18419 5668 -18395
rect 5634 -18429 5668 -18419
rect 5634 -18487 5668 -18467
rect 5634 -18501 5668 -18487
rect 6652 -17977 6686 -17963
rect 6652 -17997 6686 -17977
rect 6652 -18045 6686 -18035
rect 6652 -18069 6686 -18045
rect 6652 -18113 6686 -18107
rect 6652 -18141 6686 -18113
rect 6652 -18181 6686 -18179
rect 6652 -18213 6686 -18181
rect 6652 -18283 6686 -18251
rect 6652 -18285 6686 -18283
rect 6652 -18351 6686 -18323
rect 6652 -18357 6686 -18351
rect 6652 -18419 6686 -18395
rect 6652 -18429 6686 -18419
rect 6652 -18487 6686 -18467
rect 6652 -18501 6686 -18487
rect 7670 -17977 7704 -17963
rect 7670 -17997 7704 -17977
rect 7670 -18045 7704 -18035
rect 7670 -18069 7704 -18045
rect 7670 -18113 7704 -18107
rect 7670 -18141 7704 -18113
rect 7670 -18181 7704 -18179
rect 7670 -18213 7704 -18181
rect 7670 -18283 7704 -18251
rect 7670 -18285 7704 -18283
rect 7670 -18351 7704 -18323
rect 7670 -18357 7704 -18351
rect 7670 -18419 7704 -18395
rect 7670 -18429 7704 -18419
rect 7670 -18487 7704 -18467
rect 7670 -18501 7704 -18487
rect 8688 -17977 8722 -17963
rect 8688 -17997 8722 -17977
rect 8688 -18045 8722 -18035
rect 8688 -18069 8722 -18045
rect 8688 -18113 8722 -18107
rect 8688 -18141 8722 -18113
rect 8688 -18181 8722 -18179
rect 8688 -18213 8722 -18181
rect 8688 -18283 8722 -18251
rect 8688 -18285 8722 -18283
rect 8688 -18351 8722 -18323
rect 8688 -18357 8722 -18351
rect 8688 -18419 8722 -18395
rect 8688 -18429 8722 -18419
rect 8688 -18487 8722 -18467
rect 8688 -18501 8722 -18487
rect 9706 -17977 9740 -17963
rect 9706 -17997 9740 -17977
rect 9706 -18045 9740 -18035
rect 9706 -18069 9740 -18045
rect 9706 -18113 9740 -18107
rect 9706 -18141 9740 -18113
rect 9706 -18181 9740 -18179
rect 9706 -18213 9740 -18181
rect 9706 -18283 9740 -18251
rect 9706 -18285 9740 -18283
rect 9706 -18351 9740 -18323
rect 9706 -18357 9740 -18351
rect 9706 -18419 9740 -18395
rect 9706 -18429 9740 -18419
rect 9706 -18487 9740 -18467
rect 9706 -18501 9740 -18487
rect 10724 -17977 10758 -17963
rect 10724 -17997 10758 -17977
rect 10724 -18045 10758 -18035
rect 10724 -18069 10758 -18045
rect 10724 -18113 10758 -18107
rect 10724 -18141 10758 -18113
rect 10724 -18181 10758 -18179
rect 10724 -18213 10758 -18181
rect 10724 -18283 10758 -18251
rect 10724 -18285 10758 -18283
rect 10724 -18351 10758 -18323
rect 10724 -18357 10758 -18351
rect 10724 -18419 10758 -18395
rect 10724 -18429 10758 -18419
rect 10724 -18487 10758 -18467
rect 10724 -18501 10758 -18487
rect 11742 -17977 11776 -17963
rect 11742 -17997 11776 -17977
rect 11742 -18045 11776 -18035
rect 11742 -18069 11776 -18045
rect 11742 -18113 11776 -18107
rect 11742 -18141 11776 -18113
rect 11742 -18181 11776 -18179
rect 11742 -18213 11776 -18181
rect 11742 -18283 11776 -18251
rect 11742 -18285 11776 -18283
rect 11742 -18351 11776 -18323
rect 11742 -18357 11776 -18351
rect 11742 -18419 11776 -18395
rect 11742 -18429 11776 -18419
rect 11742 -18487 11776 -18467
rect 11742 -18501 11776 -18487
rect 12760 -17977 12794 -17963
rect 12760 -17997 12794 -17977
rect 12760 -18045 12794 -18035
rect 12760 -18069 12794 -18045
rect 12760 -18113 12794 -18107
rect 12760 -18141 12794 -18113
rect 12760 -18181 12794 -18179
rect 12760 -18213 12794 -18181
rect 12760 -18283 12794 -18251
rect 12760 -18285 12794 -18283
rect 12760 -18351 12794 -18323
rect 12760 -18357 12794 -18351
rect 12760 -18419 12794 -18395
rect 12760 -18429 12794 -18419
rect 12760 -18487 12794 -18467
rect 12760 -18501 12794 -18487
rect 13778 -17977 13812 -17963
rect 13778 -17997 13812 -17977
rect 13778 -18045 13812 -18035
rect 13778 -18069 13812 -18045
rect 13778 -18113 13812 -18107
rect 13778 -18141 13812 -18113
rect 13778 -18181 13812 -18179
rect 13778 -18213 13812 -18181
rect 13778 -18283 13812 -18251
rect 13778 -18285 13812 -18283
rect 13778 -18351 13812 -18323
rect 13778 -18357 13812 -18351
rect 13778 -18419 13812 -18395
rect 13778 -18429 13812 -18419
rect 13778 -18487 13812 -18467
rect 13778 -18501 13812 -18487
rect 14796 -17977 14830 -17963
rect 14796 -17997 14830 -17977
rect 14796 -18045 14830 -18035
rect 14796 -18069 14830 -18045
rect 14796 -18113 14830 -18107
rect 14796 -18141 14830 -18113
rect 14796 -18181 14830 -18179
rect 14796 -18213 14830 -18181
rect 14796 -18283 14830 -18251
rect 14796 -18285 14830 -18283
rect 14796 -18351 14830 -18323
rect 14796 -18357 14830 -18351
rect 14796 -18419 14830 -18395
rect 14796 -18429 14830 -18419
rect 14796 -18487 14830 -18467
rect 14796 -18501 14830 -18487
rect 15814 -17977 15848 -17963
rect 15814 -17997 15848 -17977
rect 15814 -18045 15848 -18035
rect 15814 -18069 15848 -18045
rect 15814 -18113 15848 -18107
rect 15814 -18141 15848 -18113
rect 15814 -18181 15848 -18179
rect 15814 -18213 15848 -18181
rect 15814 -18283 15848 -18251
rect 15814 -18285 15848 -18283
rect 15814 -18351 15848 -18323
rect 15814 -18357 15848 -18351
rect 15814 -18419 15848 -18395
rect 15814 -18429 15848 -18419
rect 15814 -18487 15848 -18467
rect 15814 -18501 15848 -18487
rect 16832 -17977 16866 -17963
rect 16832 -17997 16866 -17977
rect 16832 -18045 16866 -18035
rect 16832 -18069 16866 -18045
rect 16832 -18113 16866 -18107
rect 16832 -18141 16866 -18113
rect 16832 -18181 16866 -18179
rect 16832 -18213 16866 -18181
rect 16832 -18283 16866 -18251
rect 16832 -18285 16866 -18283
rect 16832 -18351 16866 -18323
rect 16832 -18357 16866 -18351
rect 16832 -18419 16866 -18395
rect 16832 -18429 16866 -18419
rect 16832 -18487 16866 -18467
rect 16832 -18501 16866 -18487
rect 17850 -17977 17884 -17963
rect 17850 -17997 17884 -17977
rect 17850 -18045 17884 -18035
rect 17850 -18069 17884 -18045
rect 17850 -18113 17884 -18107
rect 17850 -18141 17884 -18113
rect 17850 -18181 17884 -18179
rect 17850 -18213 17884 -18181
rect 17850 -18283 17884 -18251
rect 17850 -18285 17884 -18283
rect 17850 -18351 17884 -18323
rect 17850 -18357 17884 -18351
rect 17850 -18419 17884 -18395
rect 17850 -18429 17884 -18419
rect 17850 -18487 17884 -18467
rect 17850 -18501 17884 -18487
rect 18868 -17977 18902 -17963
rect 18868 -17997 18902 -17977
rect 18868 -18045 18902 -18035
rect 18868 -18069 18902 -18045
rect 18868 -18113 18902 -18107
rect 18868 -18141 18902 -18113
rect 18868 -18181 18902 -18179
rect 18868 -18213 18902 -18181
rect 18868 -18283 18902 -18251
rect 18868 -18285 18902 -18283
rect 18868 -18351 18902 -18323
rect 18868 -18357 18902 -18351
rect 18868 -18419 18902 -18395
rect 18868 -18429 18902 -18419
rect 18868 -18487 18902 -18467
rect 18868 -18501 18902 -18487
rect 19886 -17977 19920 -17963
rect 19886 -17997 19920 -17977
rect 19886 -18045 19920 -18035
rect 19886 -18069 19920 -18045
rect 19886 -18113 19920 -18107
rect 19886 -18141 19920 -18113
rect 19886 -18181 19920 -18179
rect 19886 -18213 19920 -18181
rect 19886 -18283 19920 -18251
rect 19886 -18285 19920 -18283
rect 19886 -18351 19920 -18323
rect 19886 -18357 19920 -18351
rect 19886 -18419 19920 -18395
rect 19886 -18429 19920 -18419
rect 19886 -18487 19920 -18467
rect 19886 -18501 19920 -18487
rect 20904 -17977 20938 -17963
rect 20904 -17997 20938 -17977
rect 20904 -18045 20938 -18035
rect 20904 -18069 20938 -18045
rect 20904 -18113 20938 -18107
rect 20904 -18141 20938 -18113
rect 20904 -18181 20938 -18179
rect 20904 -18213 20938 -18181
rect 20904 -18283 20938 -18251
rect 20904 -18285 20938 -18283
rect 20904 -18351 20938 -18323
rect 20904 -18357 20938 -18351
rect 20904 -18419 20938 -18395
rect 20904 -18429 20938 -18419
rect 20904 -18487 20938 -18467
rect 20904 -18501 20938 -18487
rect 21922 -17977 21956 -17963
rect 21922 -17997 21956 -17977
rect 21922 -18045 21956 -18035
rect 21922 -18069 21956 -18045
rect 21922 -18113 21956 -18107
rect 21922 -18141 21956 -18113
rect 21922 -18181 21956 -18179
rect 21922 -18213 21956 -18181
rect 21922 -18283 21956 -18251
rect 21922 -18285 21956 -18283
rect 21922 -18351 21956 -18323
rect 21922 -18357 21956 -18351
rect 21922 -18419 21956 -18395
rect 21922 -18429 21956 -18419
rect 21922 -18487 21956 -18467
rect 21922 -18501 21956 -18487
rect 22940 -17977 22974 -17963
rect 22940 -17997 22974 -17977
rect 22940 -18045 22974 -18035
rect 22940 -18069 22974 -18045
rect 22940 -18113 22974 -18107
rect 22940 -18141 22974 -18113
rect 22940 -18181 22974 -18179
rect 22940 -18213 22974 -18181
rect 22940 -18283 22974 -18251
rect 22940 -18285 22974 -18283
rect 22940 -18351 22974 -18323
rect 22940 -18357 22974 -18351
rect 22940 -18419 22974 -18395
rect 22940 -18429 22974 -18419
rect 22940 -18487 22974 -18467
rect 22940 -18501 22974 -18487
rect 24855 -17925 24889 -17923
rect 24855 -17957 24889 -17925
rect 24855 -18027 24889 -17995
rect 24855 -18029 24889 -18027
rect 24855 -18095 24889 -18067
rect 24855 -18101 24889 -18095
rect 24855 -18163 24889 -18139
rect 24855 -18173 24889 -18163
rect 24855 -18231 24889 -18211
rect 24855 -18245 24889 -18231
rect 24855 -18299 24889 -18283
rect 24855 -18317 24889 -18299
rect 24855 -18367 24889 -18355
rect 24855 -18389 24889 -18367
rect 24855 -18435 24889 -18427
rect 24855 -18461 24889 -18435
rect -22 -18589 12 -18557
rect 24855 -18503 24889 -18499
rect 24855 -18533 24889 -18503
rect -22 -18591 12 -18589
rect 2909 -18604 2919 -18570
rect 2919 -18604 2943 -18570
rect 2981 -18604 2987 -18570
rect 2987 -18604 3015 -18570
rect 3053 -18604 3055 -18570
rect 3055 -18604 3087 -18570
rect 3125 -18604 3157 -18570
rect 3157 -18604 3159 -18570
rect 3197 -18604 3225 -18570
rect 3225 -18604 3231 -18570
rect 3269 -18604 3293 -18570
rect 3293 -18604 3303 -18570
rect 3927 -18604 3937 -18570
rect 3937 -18604 3961 -18570
rect 3999 -18604 4005 -18570
rect 4005 -18604 4033 -18570
rect 4071 -18604 4073 -18570
rect 4073 -18604 4105 -18570
rect 4143 -18604 4175 -18570
rect 4175 -18604 4177 -18570
rect 4215 -18604 4243 -18570
rect 4243 -18604 4249 -18570
rect 4287 -18604 4311 -18570
rect 4311 -18604 4321 -18570
rect 4945 -18604 4955 -18570
rect 4955 -18604 4979 -18570
rect 5017 -18604 5023 -18570
rect 5023 -18604 5051 -18570
rect 5089 -18604 5091 -18570
rect 5091 -18604 5123 -18570
rect 5161 -18604 5193 -18570
rect 5193 -18604 5195 -18570
rect 5233 -18604 5261 -18570
rect 5261 -18604 5267 -18570
rect 5305 -18604 5329 -18570
rect 5329 -18604 5339 -18570
rect 5963 -18604 5973 -18570
rect 5973 -18604 5997 -18570
rect 6035 -18604 6041 -18570
rect 6041 -18604 6069 -18570
rect 6107 -18604 6109 -18570
rect 6109 -18604 6141 -18570
rect 6179 -18604 6211 -18570
rect 6211 -18604 6213 -18570
rect 6251 -18604 6279 -18570
rect 6279 -18604 6285 -18570
rect 6323 -18604 6347 -18570
rect 6347 -18604 6357 -18570
rect 6981 -18604 6991 -18570
rect 6991 -18604 7015 -18570
rect 7053 -18604 7059 -18570
rect 7059 -18604 7087 -18570
rect 7125 -18604 7127 -18570
rect 7127 -18604 7159 -18570
rect 7197 -18604 7229 -18570
rect 7229 -18604 7231 -18570
rect 7269 -18604 7297 -18570
rect 7297 -18604 7303 -18570
rect 7341 -18604 7365 -18570
rect 7365 -18604 7375 -18570
rect 7999 -18604 8009 -18570
rect 8009 -18604 8033 -18570
rect 8071 -18604 8077 -18570
rect 8077 -18604 8105 -18570
rect 8143 -18604 8145 -18570
rect 8145 -18604 8177 -18570
rect 8215 -18604 8247 -18570
rect 8247 -18604 8249 -18570
rect 8287 -18604 8315 -18570
rect 8315 -18604 8321 -18570
rect 8359 -18604 8383 -18570
rect 8383 -18604 8393 -18570
rect 9017 -18604 9027 -18570
rect 9027 -18604 9051 -18570
rect 9089 -18604 9095 -18570
rect 9095 -18604 9123 -18570
rect 9161 -18604 9163 -18570
rect 9163 -18604 9195 -18570
rect 9233 -18604 9265 -18570
rect 9265 -18604 9267 -18570
rect 9305 -18604 9333 -18570
rect 9333 -18604 9339 -18570
rect 9377 -18604 9401 -18570
rect 9401 -18604 9411 -18570
rect 10035 -18604 10045 -18570
rect 10045 -18604 10069 -18570
rect 10107 -18604 10113 -18570
rect 10113 -18604 10141 -18570
rect 10179 -18604 10181 -18570
rect 10181 -18604 10213 -18570
rect 10251 -18604 10283 -18570
rect 10283 -18604 10285 -18570
rect 10323 -18604 10351 -18570
rect 10351 -18604 10357 -18570
rect 10395 -18604 10419 -18570
rect 10419 -18604 10429 -18570
rect 11053 -18604 11063 -18570
rect 11063 -18604 11087 -18570
rect 11125 -18604 11131 -18570
rect 11131 -18604 11159 -18570
rect 11197 -18604 11199 -18570
rect 11199 -18604 11231 -18570
rect 11269 -18604 11301 -18570
rect 11301 -18604 11303 -18570
rect 11341 -18604 11369 -18570
rect 11369 -18604 11375 -18570
rect 11413 -18604 11437 -18570
rect 11437 -18604 11447 -18570
rect 12071 -18604 12081 -18570
rect 12081 -18604 12105 -18570
rect 12143 -18604 12149 -18570
rect 12149 -18604 12177 -18570
rect 12215 -18604 12217 -18570
rect 12217 -18604 12249 -18570
rect 12287 -18604 12319 -18570
rect 12319 -18604 12321 -18570
rect 12359 -18604 12387 -18570
rect 12387 -18604 12393 -18570
rect 12431 -18604 12455 -18570
rect 12455 -18604 12465 -18570
rect 13089 -18604 13099 -18570
rect 13099 -18604 13123 -18570
rect 13161 -18604 13167 -18570
rect 13167 -18604 13195 -18570
rect 13233 -18604 13235 -18570
rect 13235 -18604 13267 -18570
rect 13305 -18604 13337 -18570
rect 13337 -18604 13339 -18570
rect 13377 -18604 13405 -18570
rect 13405 -18604 13411 -18570
rect 13449 -18604 13473 -18570
rect 13473 -18604 13483 -18570
rect 14107 -18604 14117 -18570
rect 14117 -18604 14141 -18570
rect 14179 -18604 14185 -18570
rect 14185 -18604 14213 -18570
rect 14251 -18604 14253 -18570
rect 14253 -18604 14285 -18570
rect 14323 -18604 14355 -18570
rect 14355 -18604 14357 -18570
rect 14395 -18604 14423 -18570
rect 14423 -18604 14429 -18570
rect 14467 -18604 14491 -18570
rect 14491 -18604 14501 -18570
rect 15125 -18604 15135 -18570
rect 15135 -18604 15159 -18570
rect 15197 -18604 15203 -18570
rect 15203 -18604 15231 -18570
rect 15269 -18604 15271 -18570
rect 15271 -18604 15303 -18570
rect 15341 -18604 15373 -18570
rect 15373 -18604 15375 -18570
rect 15413 -18604 15441 -18570
rect 15441 -18604 15447 -18570
rect 15485 -18604 15509 -18570
rect 15509 -18604 15519 -18570
rect 16143 -18604 16153 -18570
rect 16153 -18604 16177 -18570
rect 16215 -18604 16221 -18570
rect 16221 -18604 16249 -18570
rect 16287 -18604 16289 -18570
rect 16289 -18604 16321 -18570
rect 16359 -18604 16391 -18570
rect 16391 -18604 16393 -18570
rect 16431 -18604 16459 -18570
rect 16459 -18604 16465 -18570
rect 16503 -18604 16527 -18570
rect 16527 -18604 16537 -18570
rect 17161 -18604 17171 -18570
rect 17171 -18604 17195 -18570
rect 17233 -18604 17239 -18570
rect 17239 -18604 17267 -18570
rect 17305 -18604 17307 -18570
rect 17307 -18604 17339 -18570
rect 17377 -18604 17409 -18570
rect 17409 -18604 17411 -18570
rect 17449 -18604 17477 -18570
rect 17477 -18604 17483 -18570
rect 17521 -18604 17545 -18570
rect 17545 -18604 17555 -18570
rect 18179 -18604 18189 -18570
rect 18189 -18604 18213 -18570
rect 18251 -18604 18257 -18570
rect 18257 -18604 18285 -18570
rect 18323 -18604 18325 -18570
rect 18325 -18604 18357 -18570
rect 18395 -18604 18427 -18570
rect 18427 -18604 18429 -18570
rect 18467 -18604 18495 -18570
rect 18495 -18604 18501 -18570
rect 18539 -18604 18563 -18570
rect 18563 -18604 18573 -18570
rect 19197 -18604 19207 -18570
rect 19207 -18604 19231 -18570
rect 19269 -18604 19275 -18570
rect 19275 -18604 19303 -18570
rect 19341 -18604 19343 -18570
rect 19343 -18604 19375 -18570
rect 19413 -18604 19445 -18570
rect 19445 -18604 19447 -18570
rect 19485 -18604 19513 -18570
rect 19513 -18604 19519 -18570
rect 19557 -18604 19581 -18570
rect 19581 -18604 19591 -18570
rect 20215 -18604 20225 -18570
rect 20225 -18604 20249 -18570
rect 20287 -18604 20293 -18570
rect 20293 -18604 20321 -18570
rect 20359 -18604 20361 -18570
rect 20361 -18604 20393 -18570
rect 20431 -18604 20463 -18570
rect 20463 -18604 20465 -18570
rect 20503 -18604 20531 -18570
rect 20531 -18604 20537 -18570
rect 20575 -18604 20599 -18570
rect 20599 -18604 20609 -18570
rect 21233 -18604 21243 -18570
rect 21243 -18604 21267 -18570
rect 21305 -18604 21311 -18570
rect 21311 -18604 21339 -18570
rect 21377 -18604 21379 -18570
rect 21379 -18604 21411 -18570
rect 21449 -18604 21481 -18570
rect 21481 -18604 21483 -18570
rect 21521 -18604 21549 -18570
rect 21549 -18604 21555 -18570
rect 21593 -18604 21617 -18570
rect 21617 -18604 21627 -18570
rect 22251 -18604 22261 -18570
rect 22261 -18604 22285 -18570
rect 22323 -18604 22329 -18570
rect 22329 -18604 22357 -18570
rect 22395 -18604 22397 -18570
rect 22397 -18604 22429 -18570
rect 22467 -18604 22499 -18570
rect 22499 -18604 22501 -18570
rect 22539 -18604 22567 -18570
rect 22567 -18604 22573 -18570
rect 22611 -18604 22635 -18570
rect 22635 -18604 22645 -18570
rect -22 -18657 12 -18629
rect -22 -18663 12 -18657
rect -22 -18725 12 -18701
rect -22 -18735 12 -18725
rect -22 -18793 12 -18773
rect -22 -18807 12 -18793
rect 24855 -18605 24889 -18571
rect 24855 -18673 24889 -18643
rect 24855 -18677 24889 -18673
rect 24855 -18741 24889 -18715
rect 24855 -18749 24889 -18741
rect 24855 -18809 24889 -18787
rect 24855 -18821 24889 -18809
rect -12289 -18877 -12255 -18859
rect -12289 -18893 -12255 -18877
rect -8855 -18910 -8845 -18876
rect -8845 -18910 -8821 -18876
rect -8783 -18910 -8777 -18876
rect -8777 -18910 -8749 -18876
rect -8711 -18910 -8709 -18876
rect -8709 -18910 -8677 -18876
rect -8639 -18910 -8607 -18876
rect -8607 -18910 -8605 -18876
rect -8567 -18910 -8539 -18876
rect -8539 -18910 -8533 -18876
rect -8495 -18910 -8471 -18876
rect -8471 -18910 -8461 -18876
rect -7837 -18910 -7827 -18876
rect -7827 -18910 -7803 -18876
rect -7765 -18910 -7759 -18876
rect -7759 -18910 -7731 -18876
rect -7693 -18910 -7691 -18876
rect -7691 -18910 -7659 -18876
rect -7621 -18910 -7589 -18876
rect -7589 -18910 -7587 -18876
rect -7549 -18910 -7521 -18876
rect -7521 -18910 -7515 -18876
rect -7477 -18910 -7453 -18876
rect -7453 -18910 -7443 -18876
rect -6819 -18910 -6809 -18876
rect -6809 -18910 -6785 -18876
rect -6747 -18910 -6741 -18876
rect -6741 -18910 -6713 -18876
rect -6675 -18910 -6673 -18876
rect -6673 -18910 -6641 -18876
rect -6603 -18910 -6571 -18876
rect -6571 -18910 -6569 -18876
rect -6531 -18910 -6503 -18876
rect -6503 -18910 -6497 -18876
rect -6459 -18910 -6435 -18876
rect -6435 -18910 -6425 -18876
rect -5801 -18910 -5791 -18876
rect -5791 -18910 -5767 -18876
rect -5729 -18910 -5723 -18876
rect -5723 -18910 -5695 -18876
rect -5657 -18910 -5655 -18876
rect -5655 -18910 -5623 -18876
rect -5585 -18910 -5553 -18876
rect -5553 -18910 -5551 -18876
rect -5513 -18910 -5485 -18876
rect -5485 -18910 -5479 -18876
rect -5441 -18910 -5417 -18876
rect -5417 -18910 -5407 -18876
rect -4783 -18910 -4773 -18876
rect -4773 -18910 -4749 -18876
rect -4711 -18910 -4705 -18876
rect -4705 -18910 -4677 -18876
rect -4639 -18910 -4637 -18876
rect -4637 -18910 -4605 -18876
rect -4567 -18910 -4535 -18876
rect -4535 -18910 -4533 -18876
rect -4495 -18910 -4467 -18876
rect -4467 -18910 -4461 -18876
rect -4423 -18910 -4399 -18876
rect -4399 -18910 -4389 -18876
rect -3765 -18910 -3755 -18876
rect -3755 -18910 -3731 -18876
rect -3693 -18910 -3687 -18876
rect -3687 -18910 -3659 -18876
rect -3621 -18910 -3619 -18876
rect -3619 -18910 -3587 -18876
rect -3549 -18910 -3517 -18876
rect -3517 -18910 -3515 -18876
rect -3477 -18910 -3449 -18876
rect -3449 -18910 -3443 -18876
rect -3405 -18910 -3381 -18876
rect -3381 -18910 -3371 -18876
rect -2747 -18910 -2737 -18876
rect -2737 -18910 -2713 -18876
rect -2675 -18910 -2669 -18876
rect -2669 -18910 -2641 -18876
rect -2603 -18910 -2601 -18876
rect -2601 -18910 -2569 -18876
rect -2531 -18910 -2499 -18876
rect -2499 -18910 -2497 -18876
rect -2459 -18910 -2431 -18876
rect -2431 -18910 -2425 -18876
rect -2387 -18910 -2363 -18876
rect -2363 -18910 -2353 -18876
rect -1729 -18910 -1719 -18876
rect -1719 -18910 -1695 -18876
rect -1657 -18910 -1651 -18876
rect -1651 -18910 -1623 -18876
rect -1585 -18910 -1583 -18876
rect -1583 -18910 -1551 -18876
rect -1513 -18910 -1481 -18876
rect -1481 -18910 -1479 -18876
rect -1441 -18910 -1413 -18876
rect -1413 -18910 -1407 -18876
rect -1369 -18910 -1345 -18876
rect -1345 -18910 -1335 -18876
rect -711 -18910 -701 -18876
rect -701 -18910 -677 -18876
rect -639 -18910 -633 -18876
rect -633 -18910 -605 -18876
rect -567 -18910 -565 -18876
rect -565 -18910 -533 -18876
rect -495 -18910 -463 -18876
rect -463 -18910 -461 -18876
rect -423 -18910 -395 -18876
rect -395 -18910 -389 -18876
rect -351 -18910 -327 -18876
rect -327 -18910 -317 -18876
rect 24855 -18877 24889 -18859
rect 24855 -18893 24889 -18877
rect -12289 -18945 -12255 -18931
rect -12289 -18965 -12255 -18945
rect -12289 -19013 -12255 -19003
rect -12289 -19037 -12255 -19013
rect -12289 -19081 -12255 -19075
rect -12289 -19109 -12255 -19081
rect 24855 -18945 24889 -18931
rect 24855 -18965 24889 -18945
rect 24855 -19013 24889 -19003
rect 24855 -19037 24889 -19013
rect -12289 -19149 -12255 -19147
rect -12289 -19181 -12255 -19149
rect 2909 -19126 2919 -19092
rect 2919 -19126 2943 -19092
rect 2981 -19126 2987 -19092
rect 2987 -19126 3015 -19092
rect 3053 -19126 3055 -19092
rect 3055 -19126 3087 -19092
rect 3125 -19126 3157 -19092
rect 3157 -19126 3159 -19092
rect 3197 -19126 3225 -19092
rect 3225 -19126 3231 -19092
rect 3269 -19126 3293 -19092
rect 3293 -19126 3303 -19092
rect 3927 -19126 3937 -19092
rect 3937 -19126 3961 -19092
rect 3999 -19126 4005 -19092
rect 4005 -19126 4033 -19092
rect 4071 -19126 4073 -19092
rect 4073 -19126 4105 -19092
rect 4143 -19126 4175 -19092
rect 4175 -19126 4177 -19092
rect 4215 -19126 4243 -19092
rect 4243 -19126 4249 -19092
rect 4287 -19126 4311 -19092
rect 4311 -19126 4321 -19092
rect 4945 -19126 4955 -19092
rect 4955 -19126 4979 -19092
rect 5017 -19126 5023 -19092
rect 5023 -19126 5051 -19092
rect 5089 -19126 5091 -19092
rect 5091 -19126 5123 -19092
rect 5161 -19126 5193 -19092
rect 5193 -19126 5195 -19092
rect 5233 -19126 5261 -19092
rect 5261 -19126 5267 -19092
rect 5305 -19126 5329 -19092
rect 5329 -19126 5339 -19092
rect 5963 -19126 5973 -19092
rect 5973 -19126 5997 -19092
rect 6035 -19126 6041 -19092
rect 6041 -19126 6069 -19092
rect 6107 -19126 6109 -19092
rect 6109 -19126 6141 -19092
rect 6179 -19126 6211 -19092
rect 6211 -19126 6213 -19092
rect 6251 -19126 6279 -19092
rect 6279 -19126 6285 -19092
rect 6323 -19126 6347 -19092
rect 6347 -19126 6357 -19092
rect 6981 -19126 6991 -19092
rect 6991 -19126 7015 -19092
rect 7053 -19126 7059 -19092
rect 7059 -19126 7087 -19092
rect 7125 -19126 7127 -19092
rect 7127 -19126 7159 -19092
rect 7197 -19126 7229 -19092
rect 7229 -19126 7231 -19092
rect 7269 -19126 7297 -19092
rect 7297 -19126 7303 -19092
rect 7341 -19126 7365 -19092
rect 7365 -19126 7375 -19092
rect 7999 -19126 8009 -19092
rect 8009 -19126 8033 -19092
rect 8071 -19126 8077 -19092
rect 8077 -19126 8105 -19092
rect 8143 -19126 8145 -19092
rect 8145 -19126 8177 -19092
rect 8215 -19126 8247 -19092
rect 8247 -19126 8249 -19092
rect 8287 -19126 8315 -19092
rect 8315 -19126 8321 -19092
rect 8359 -19126 8383 -19092
rect 8383 -19126 8393 -19092
rect 9017 -19126 9027 -19092
rect 9027 -19126 9051 -19092
rect 9089 -19126 9095 -19092
rect 9095 -19126 9123 -19092
rect 9161 -19126 9163 -19092
rect 9163 -19126 9195 -19092
rect 9233 -19126 9265 -19092
rect 9265 -19126 9267 -19092
rect 9305 -19126 9333 -19092
rect 9333 -19126 9339 -19092
rect 9377 -19126 9401 -19092
rect 9401 -19126 9411 -19092
rect 10035 -19126 10045 -19092
rect 10045 -19126 10069 -19092
rect 10107 -19126 10113 -19092
rect 10113 -19126 10141 -19092
rect 10179 -19126 10181 -19092
rect 10181 -19126 10213 -19092
rect 10251 -19126 10283 -19092
rect 10283 -19126 10285 -19092
rect 10323 -19126 10351 -19092
rect 10351 -19126 10357 -19092
rect 10395 -19126 10419 -19092
rect 10419 -19126 10429 -19092
rect 11053 -19126 11063 -19092
rect 11063 -19126 11087 -19092
rect 11125 -19126 11131 -19092
rect 11131 -19126 11159 -19092
rect 11197 -19126 11199 -19092
rect 11199 -19126 11231 -19092
rect 11269 -19126 11301 -19092
rect 11301 -19126 11303 -19092
rect 11341 -19126 11369 -19092
rect 11369 -19126 11375 -19092
rect 11413 -19126 11437 -19092
rect 11437 -19126 11447 -19092
rect 12071 -19126 12081 -19092
rect 12081 -19126 12105 -19092
rect 12143 -19126 12149 -19092
rect 12149 -19126 12177 -19092
rect 12215 -19126 12217 -19092
rect 12217 -19126 12249 -19092
rect 12287 -19126 12319 -19092
rect 12319 -19126 12321 -19092
rect 12359 -19126 12387 -19092
rect 12387 -19126 12393 -19092
rect 12431 -19126 12455 -19092
rect 12455 -19126 12465 -19092
rect 13089 -19126 13099 -19092
rect 13099 -19126 13123 -19092
rect 13161 -19126 13167 -19092
rect 13167 -19126 13195 -19092
rect 13233 -19126 13235 -19092
rect 13235 -19126 13267 -19092
rect 13305 -19126 13337 -19092
rect 13337 -19126 13339 -19092
rect 13377 -19126 13405 -19092
rect 13405 -19126 13411 -19092
rect 13449 -19126 13473 -19092
rect 13473 -19126 13483 -19092
rect 14107 -19126 14117 -19092
rect 14117 -19126 14141 -19092
rect 14179 -19126 14185 -19092
rect 14185 -19126 14213 -19092
rect 14251 -19126 14253 -19092
rect 14253 -19126 14285 -19092
rect 14323 -19126 14355 -19092
rect 14355 -19126 14357 -19092
rect 14395 -19126 14423 -19092
rect 14423 -19126 14429 -19092
rect 14467 -19126 14491 -19092
rect 14491 -19126 14501 -19092
rect 15125 -19126 15135 -19092
rect 15135 -19126 15159 -19092
rect 15197 -19126 15203 -19092
rect 15203 -19126 15231 -19092
rect 15269 -19126 15271 -19092
rect 15271 -19126 15303 -19092
rect 15341 -19126 15373 -19092
rect 15373 -19126 15375 -19092
rect 15413 -19126 15441 -19092
rect 15441 -19126 15447 -19092
rect 15485 -19126 15509 -19092
rect 15509 -19126 15519 -19092
rect 16143 -19126 16153 -19092
rect 16153 -19126 16177 -19092
rect 16215 -19126 16221 -19092
rect 16221 -19126 16249 -19092
rect 16287 -19126 16289 -19092
rect 16289 -19126 16321 -19092
rect 16359 -19126 16391 -19092
rect 16391 -19126 16393 -19092
rect 16431 -19126 16459 -19092
rect 16459 -19126 16465 -19092
rect 16503 -19126 16527 -19092
rect 16527 -19126 16537 -19092
rect 17161 -19126 17171 -19092
rect 17171 -19126 17195 -19092
rect 17233 -19126 17239 -19092
rect 17239 -19126 17267 -19092
rect 17305 -19126 17307 -19092
rect 17307 -19126 17339 -19092
rect 17377 -19126 17409 -19092
rect 17409 -19126 17411 -19092
rect 17449 -19126 17477 -19092
rect 17477 -19126 17483 -19092
rect 17521 -19126 17545 -19092
rect 17545 -19126 17555 -19092
rect 18179 -19126 18189 -19092
rect 18189 -19126 18213 -19092
rect 18251 -19126 18257 -19092
rect 18257 -19126 18285 -19092
rect 18323 -19126 18325 -19092
rect 18325 -19126 18357 -19092
rect 18395 -19126 18427 -19092
rect 18427 -19126 18429 -19092
rect 18467 -19126 18495 -19092
rect 18495 -19126 18501 -19092
rect 18539 -19126 18563 -19092
rect 18563 -19126 18573 -19092
rect 19197 -19126 19207 -19092
rect 19207 -19126 19231 -19092
rect 19269 -19126 19275 -19092
rect 19275 -19126 19303 -19092
rect 19341 -19126 19343 -19092
rect 19343 -19126 19375 -19092
rect 19413 -19126 19445 -19092
rect 19445 -19126 19447 -19092
rect 19485 -19126 19513 -19092
rect 19513 -19126 19519 -19092
rect 19557 -19126 19581 -19092
rect 19581 -19126 19591 -19092
rect 20215 -19126 20225 -19092
rect 20225 -19126 20249 -19092
rect 20287 -19126 20293 -19092
rect 20293 -19126 20321 -19092
rect 20359 -19126 20361 -19092
rect 20361 -19126 20393 -19092
rect 20431 -19126 20463 -19092
rect 20463 -19126 20465 -19092
rect 20503 -19126 20531 -19092
rect 20531 -19126 20537 -19092
rect 20575 -19126 20599 -19092
rect 20599 -19126 20609 -19092
rect 21233 -19126 21243 -19092
rect 21243 -19126 21267 -19092
rect 21305 -19126 21311 -19092
rect 21311 -19126 21339 -19092
rect 21377 -19126 21379 -19092
rect 21379 -19126 21411 -19092
rect 21449 -19126 21481 -19092
rect 21481 -19126 21483 -19092
rect 21521 -19126 21549 -19092
rect 21549 -19126 21555 -19092
rect 21593 -19126 21617 -19092
rect 21617 -19126 21627 -19092
rect 22251 -19126 22261 -19092
rect 22261 -19126 22285 -19092
rect 22323 -19126 22329 -19092
rect 22329 -19126 22357 -19092
rect 22395 -19126 22397 -19092
rect 22397 -19126 22429 -19092
rect 22467 -19126 22499 -19092
rect 22499 -19126 22501 -19092
rect 22539 -19126 22567 -19092
rect 22567 -19126 22573 -19092
rect 22611 -19126 22635 -19092
rect 22635 -19126 22645 -19092
rect 24855 -19081 24889 -19075
rect 24855 -19109 24889 -19081
rect -12289 -19251 -12255 -19219
rect -12289 -19253 -12255 -19251
rect -12289 -19319 -12255 -19291
rect -12289 -19325 -12255 -19319
rect -12289 -19387 -12255 -19363
rect -12289 -19397 -12255 -19387
rect -12289 -19455 -12255 -19435
rect -12289 -19469 -12255 -19455
rect -12289 -19523 -12255 -19507
rect -12289 -19541 -12255 -19523
rect -12289 -19591 -12255 -19579
rect -12289 -19613 -12255 -19591
rect -12289 -19659 -12255 -19651
rect -12289 -19685 -12255 -19659
rect -12289 -19727 -12255 -19723
rect -12289 -19757 -12255 -19727
rect 2580 -19209 2614 -19195
rect 2580 -19229 2614 -19209
rect 2580 -19277 2614 -19267
rect 2580 -19301 2614 -19277
rect 2580 -19345 2614 -19339
rect 2580 -19373 2614 -19345
rect 2580 -19413 2614 -19411
rect 2580 -19445 2614 -19413
rect 2580 -19515 2614 -19483
rect 2580 -19517 2614 -19515
rect 2580 -19583 2614 -19555
rect 2580 -19589 2614 -19583
rect 2580 -19651 2614 -19627
rect 2580 -19661 2614 -19651
rect 2580 -19719 2614 -19699
rect 2580 -19733 2614 -19719
rect 3598 -19209 3632 -19195
rect 3598 -19229 3632 -19209
rect 3598 -19277 3632 -19267
rect 3598 -19301 3632 -19277
rect 3598 -19345 3632 -19339
rect 3598 -19373 3632 -19345
rect 3598 -19413 3632 -19411
rect 3598 -19445 3632 -19413
rect 3598 -19515 3632 -19483
rect 3598 -19517 3632 -19515
rect 3598 -19583 3632 -19555
rect 3598 -19589 3632 -19583
rect 3598 -19651 3632 -19627
rect 3598 -19661 3632 -19651
rect 3598 -19719 3632 -19699
rect 3598 -19733 3632 -19719
rect 4616 -19209 4650 -19195
rect 4616 -19229 4650 -19209
rect 4616 -19277 4650 -19267
rect 4616 -19301 4650 -19277
rect 4616 -19345 4650 -19339
rect 4616 -19373 4650 -19345
rect 4616 -19413 4650 -19411
rect 4616 -19445 4650 -19413
rect 4616 -19515 4650 -19483
rect 4616 -19517 4650 -19515
rect 4616 -19583 4650 -19555
rect 4616 -19589 4650 -19583
rect 4616 -19651 4650 -19627
rect 4616 -19661 4650 -19651
rect 4616 -19719 4650 -19699
rect 4616 -19733 4650 -19719
rect 5634 -19209 5668 -19195
rect 5634 -19229 5668 -19209
rect 5634 -19277 5668 -19267
rect 5634 -19301 5668 -19277
rect 5634 -19345 5668 -19339
rect 5634 -19373 5668 -19345
rect 5634 -19413 5668 -19411
rect 5634 -19445 5668 -19413
rect 5634 -19515 5668 -19483
rect 5634 -19517 5668 -19515
rect 5634 -19583 5668 -19555
rect 5634 -19589 5668 -19583
rect 5634 -19651 5668 -19627
rect 5634 -19661 5668 -19651
rect 5634 -19719 5668 -19699
rect 5634 -19733 5668 -19719
rect 6652 -19209 6686 -19195
rect 6652 -19229 6686 -19209
rect 6652 -19277 6686 -19267
rect 6652 -19301 6686 -19277
rect 6652 -19345 6686 -19339
rect 6652 -19373 6686 -19345
rect 6652 -19413 6686 -19411
rect 6652 -19445 6686 -19413
rect 6652 -19515 6686 -19483
rect 6652 -19517 6686 -19515
rect 6652 -19583 6686 -19555
rect 6652 -19589 6686 -19583
rect 6652 -19651 6686 -19627
rect 6652 -19661 6686 -19651
rect 6652 -19719 6686 -19699
rect 6652 -19733 6686 -19719
rect 7670 -19209 7704 -19195
rect 7670 -19229 7704 -19209
rect 7670 -19277 7704 -19267
rect 7670 -19301 7704 -19277
rect 7670 -19345 7704 -19339
rect 7670 -19373 7704 -19345
rect 7670 -19413 7704 -19411
rect 7670 -19445 7704 -19413
rect 7670 -19515 7704 -19483
rect 7670 -19517 7704 -19515
rect 7670 -19583 7704 -19555
rect 7670 -19589 7704 -19583
rect 7670 -19651 7704 -19627
rect 7670 -19661 7704 -19651
rect 7670 -19719 7704 -19699
rect 7670 -19733 7704 -19719
rect 8688 -19209 8722 -19195
rect 8688 -19229 8722 -19209
rect 8688 -19277 8722 -19267
rect 8688 -19301 8722 -19277
rect 8688 -19345 8722 -19339
rect 8688 -19373 8722 -19345
rect 8688 -19413 8722 -19411
rect 8688 -19445 8722 -19413
rect 8688 -19515 8722 -19483
rect 8688 -19517 8722 -19515
rect 8688 -19583 8722 -19555
rect 8688 -19589 8722 -19583
rect 8688 -19651 8722 -19627
rect 8688 -19661 8722 -19651
rect 8688 -19719 8722 -19699
rect 8688 -19733 8722 -19719
rect 9706 -19209 9740 -19195
rect 9706 -19229 9740 -19209
rect 9706 -19277 9740 -19267
rect 9706 -19301 9740 -19277
rect 9706 -19345 9740 -19339
rect 9706 -19373 9740 -19345
rect 9706 -19413 9740 -19411
rect 9706 -19445 9740 -19413
rect 9706 -19515 9740 -19483
rect 9706 -19517 9740 -19515
rect 9706 -19583 9740 -19555
rect 9706 -19589 9740 -19583
rect 9706 -19651 9740 -19627
rect 9706 -19661 9740 -19651
rect 9706 -19719 9740 -19699
rect 9706 -19733 9740 -19719
rect 10724 -19209 10758 -19195
rect 10724 -19229 10758 -19209
rect 10724 -19277 10758 -19267
rect 10724 -19301 10758 -19277
rect 10724 -19345 10758 -19339
rect 10724 -19373 10758 -19345
rect 10724 -19413 10758 -19411
rect 10724 -19445 10758 -19413
rect 10724 -19515 10758 -19483
rect 10724 -19517 10758 -19515
rect 10724 -19583 10758 -19555
rect 10724 -19589 10758 -19583
rect 10724 -19651 10758 -19627
rect 10724 -19661 10758 -19651
rect 10724 -19719 10758 -19699
rect 10724 -19733 10758 -19719
rect 11742 -19209 11776 -19195
rect 11742 -19229 11776 -19209
rect 11742 -19277 11776 -19267
rect 11742 -19301 11776 -19277
rect 11742 -19345 11776 -19339
rect 11742 -19373 11776 -19345
rect 11742 -19413 11776 -19411
rect 11742 -19445 11776 -19413
rect 11742 -19515 11776 -19483
rect 11742 -19517 11776 -19515
rect 11742 -19583 11776 -19555
rect 11742 -19589 11776 -19583
rect 11742 -19651 11776 -19627
rect 11742 -19661 11776 -19651
rect 11742 -19719 11776 -19699
rect 11742 -19733 11776 -19719
rect 12760 -19209 12794 -19195
rect 12760 -19229 12794 -19209
rect 12760 -19277 12794 -19267
rect 12760 -19301 12794 -19277
rect 12760 -19345 12794 -19339
rect 12760 -19373 12794 -19345
rect 12760 -19413 12794 -19411
rect 12760 -19445 12794 -19413
rect 12760 -19515 12794 -19483
rect 12760 -19517 12794 -19515
rect 12760 -19583 12794 -19555
rect 12760 -19589 12794 -19583
rect 12760 -19651 12794 -19627
rect 12760 -19661 12794 -19651
rect 12760 -19719 12794 -19699
rect 12760 -19733 12794 -19719
rect 13778 -19209 13812 -19195
rect 13778 -19229 13812 -19209
rect 13778 -19277 13812 -19267
rect 13778 -19301 13812 -19277
rect 13778 -19345 13812 -19339
rect 13778 -19373 13812 -19345
rect 13778 -19413 13812 -19411
rect 13778 -19445 13812 -19413
rect 13778 -19515 13812 -19483
rect 13778 -19517 13812 -19515
rect 13778 -19583 13812 -19555
rect 13778 -19589 13812 -19583
rect 13778 -19651 13812 -19627
rect 13778 -19661 13812 -19651
rect 13778 -19719 13812 -19699
rect 13778 -19733 13812 -19719
rect 14796 -19209 14830 -19195
rect 14796 -19229 14830 -19209
rect 14796 -19277 14830 -19267
rect 14796 -19301 14830 -19277
rect 14796 -19345 14830 -19339
rect 14796 -19373 14830 -19345
rect 14796 -19413 14830 -19411
rect 14796 -19445 14830 -19413
rect 14796 -19515 14830 -19483
rect 14796 -19517 14830 -19515
rect 14796 -19583 14830 -19555
rect 14796 -19589 14830 -19583
rect 14796 -19651 14830 -19627
rect 14796 -19661 14830 -19651
rect 14796 -19719 14830 -19699
rect 14796 -19733 14830 -19719
rect 15814 -19209 15848 -19195
rect 15814 -19229 15848 -19209
rect 15814 -19277 15848 -19267
rect 15814 -19301 15848 -19277
rect 15814 -19345 15848 -19339
rect 15814 -19373 15848 -19345
rect 15814 -19413 15848 -19411
rect 15814 -19445 15848 -19413
rect 15814 -19515 15848 -19483
rect 15814 -19517 15848 -19515
rect 15814 -19583 15848 -19555
rect 15814 -19589 15848 -19583
rect 15814 -19651 15848 -19627
rect 15814 -19661 15848 -19651
rect 15814 -19719 15848 -19699
rect 15814 -19733 15848 -19719
rect 16832 -19209 16866 -19195
rect 16832 -19229 16866 -19209
rect 16832 -19277 16866 -19267
rect 16832 -19301 16866 -19277
rect 16832 -19345 16866 -19339
rect 16832 -19373 16866 -19345
rect 16832 -19413 16866 -19411
rect 16832 -19445 16866 -19413
rect 16832 -19515 16866 -19483
rect 16832 -19517 16866 -19515
rect 16832 -19583 16866 -19555
rect 16832 -19589 16866 -19583
rect 16832 -19651 16866 -19627
rect 16832 -19661 16866 -19651
rect 16832 -19719 16866 -19699
rect 16832 -19733 16866 -19719
rect 17850 -19209 17884 -19195
rect 17850 -19229 17884 -19209
rect 17850 -19277 17884 -19267
rect 17850 -19301 17884 -19277
rect 17850 -19345 17884 -19339
rect 17850 -19373 17884 -19345
rect 17850 -19413 17884 -19411
rect 17850 -19445 17884 -19413
rect 17850 -19515 17884 -19483
rect 17850 -19517 17884 -19515
rect 17850 -19583 17884 -19555
rect 17850 -19589 17884 -19583
rect 17850 -19651 17884 -19627
rect 17850 -19661 17884 -19651
rect 17850 -19719 17884 -19699
rect 17850 -19733 17884 -19719
rect 18868 -19209 18902 -19195
rect 18868 -19229 18902 -19209
rect 18868 -19277 18902 -19267
rect 18868 -19301 18902 -19277
rect 18868 -19345 18902 -19339
rect 18868 -19373 18902 -19345
rect 18868 -19413 18902 -19411
rect 18868 -19445 18902 -19413
rect 18868 -19515 18902 -19483
rect 18868 -19517 18902 -19515
rect 18868 -19583 18902 -19555
rect 18868 -19589 18902 -19583
rect 18868 -19651 18902 -19627
rect 18868 -19661 18902 -19651
rect 18868 -19719 18902 -19699
rect 18868 -19733 18902 -19719
rect 19886 -19209 19920 -19195
rect 19886 -19229 19920 -19209
rect 19886 -19277 19920 -19267
rect 19886 -19301 19920 -19277
rect 19886 -19345 19920 -19339
rect 19886 -19373 19920 -19345
rect 19886 -19413 19920 -19411
rect 19886 -19445 19920 -19413
rect 19886 -19515 19920 -19483
rect 19886 -19517 19920 -19515
rect 19886 -19583 19920 -19555
rect 19886 -19589 19920 -19583
rect 19886 -19651 19920 -19627
rect 19886 -19661 19920 -19651
rect 19886 -19719 19920 -19699
rect 19886 -19733 19920 -19719
rect 20904 -19209 20938 -19195
rect 20904 -19229 20938 -19209
rect 20904 -19277 20938 -19267
rect 20904 -19301 20938 -19277
rect 20904 -19345 20938 -19339
rect 20904 -19373 20938 -19345
rect 20904 -19413 20938 -19411
rect 20904 -19445 20938 -19413
rect 20904 -19515 20938 -19483
rect 20904 -19517 20938 -19515
rect 20904 -19583 20938 -19555
rect 20904 -19589 20938 -19583
rect 20904 -19651 20938 -19627
rect 20904 -19661 20938 -19651
rect 20904 -19719 20938 -19699
rect 20904 -19733 20938 -19719
rect 21922 -19209 21956 -19195
rect 21922 -19229 21956 -19209
rect 21922 -19277 21956 -19267
rect 21922 -19301 21956 -19277
rect 21922 -19345 21956 -19339
rect 21922 -19373 21956 -19345
rect 21922 -19413 21956 -19411
rect 21922 -19445 21956 -19413
rect 21922 -19515 21956 -19483
rect 21922 -19517 21956 -19515
rect 21922 -19583 21956 -19555
rect 21922 -19589 21956 -19583
rect 21922 -19651 21956 -19627
rect 21922 -19661 21956 -19651
rect 21922 -19719 21956 -19699
rect 21922 -19733 21956 -19719
rect 22940 -19209 22974 -19195
rect 22940 -19229 22974 -19209
rect 22940 -19277 22974 -19267
rect 22940 -19301 22974 -19277
rect 22940 -19345 22974 -19339
rect 22940 -19373 22974 -19345
rect 22940 -19413 22974 -19411
rect 22940 -19445 22974 -19413
rect 22940 -19515 22974 -19483
rect 22940 -19517 22974 -19515
rect 22940 -19583 22974 -19555
rect 22940 -19589 22974 -19583
rect 22940 -19651 22974 -19627
rect 22940 -19661 22974 -19651
rect 22940 -19719 22974 -19699
rect 22940 -19733 22974 -19719
rect 24855 -19149 24889 -19147
rect 24855 -19181 24889 -19149
rect 24855 -19251 24889 -19219
rect 24855 -19253 24889 -19251
rect 24855 -19319 24889 -19291
rect 24855 -19325 24889 -19319
rect 24855 -19387 24889 -19363
rect 24855 -19397 24889 -19387
rect 24855 -19455 24889 -19435
rect 24855 -19469 24889 -19455
rect 24855 -19523 24889 -19507
rect 24855 -19541 24889 -19523
rect 24855 -19591 24889 -19579
rect 24855 -19613 24889 -19591
rect 24855 -19659 24889 -19651
rect 24855 -19685 24889 -19659
rect 24855 -19727 24889 -19723
rect 24855 -19757 24889 -19727
rect -12289 -19829 -12255 -19795
rect 2909 -19836 2919 -19802
rect 2919 -19836 2943 -19802
rect 2981 -19836 2987 -19802
rect 2987 -19836 3015 -19802
rect 3053 -19836 3055 -19802
rect 3055 -19836 3087 -19802
rect 3125 -19836 3157 -19802
rect 3157 -19836 3159 -19802
rect 3197 -19836 3225 -19802
rect 3225 -19836 3231 -19802
rect 3269 -19836 3293 -19802
rect 3293 -19836 3303 -19802
rect 3927 -19836 3937 -19802
rect 3937 -19836 3961 -19802
rect 3999 -19836 4005 -19802
rect 4005 -19836 4033 -19802
rect 4071 -19836 4073 -19802
rect 4073 -19836 4105 -19802
rect 4143 -19836 4175 -19802
rect 4175 -19836 4177 -19802
rect 4215 -19836 4243 -19802
rect 4243 -19836 4249 -19802
rect 4287 -19836 4311 -19802
rect 4311 -19836 4321 -19802
rect 4945 -19836 4955 -19802
rect 4955 -19836 4979 -19802
rect 5017 -19836 5023 -19802
rect 5023 -19836 5051 -19802
rect 5089 -19836 5091 -19802
rect 5091 -19836 5123 -19802
rect 5161 -19836 5193 -19802
rect 5193 -19836 5195 -19802
rect 5233 -19836 5261 -19802
rect 5261 -19836 5267 -19802
rect 5305 -19836 5329 -19802
rect 5329 -19836 5339 -19802
rect 5963 -19836 5973 -19802
rect 5973 -19836 5997 -19802
rect 6035 -19836 6041 -19802
rect 6041 -19836 6069 -19802
rect 6107 -19836 6109 -19802
rect 6109 -19836 6141 -19802
rect 6179 -19836 6211 -19802
rect 6211 -19836 6213 -19802
rect 6251 -19836 6279 -19802
rect 6279 -19836 6285 -19802
rect 6323 -19836 6347 -19802
rect 6347 -19836 6357 -19802
rect 6981 -19836 6991 -19802
rect 6991 -19836 7015 -19802
rect 7053 -19836 7059 -19802
rect 7059 -19836 7087 -19802
rect 7125 -19836 7127 -19802
rect 7127 -19836 7159 -19802
rect 7197 -19836 7229 -19802
rect 7229 -19836 7231 -19802
rect 7269 -19836 7297 -19802
rect 7297 -19836 7303 -19802
rect 7341 -19836 7365 -19802
rect 7365 -19836 7375 -19802
rect 7999 -19836 8009 -19802
rect 8009 -19836 8033 -19802
rect 8071 -19836 8077 -19802
rect 8077 -19836 8105 -19802
rect 8143 -19836 8145 -19802
rect 8145 -19836 8177 -19802
rect 8215 -19836 8247 -19802
rect 8247 -19836 8249 -19802
rect 8287 -19836 8315 -19802
rect 8315 -19836 8321 -19802
rect 8359 -19836 8383 -19802
rect 8383 -19836 8393 -19802
rect 9017 -19836 9027 -19802
rect 9027 -19836 9051 -19802
rect 9089 -19836 9095 -19802
rect 9095 -19836 9123 -19802
rect 9161 -19836 9163 -19802
rect 9163 -19836 9195 -19802
rect 9233 -19836 9265 -19802
rect 9265 -19836 9267 -19802
rect 9305 -19836 9333 -19802
rect 9333 -19836 9339 -19802
rect 9377 -19836 9401 -19802
rect 9401 -19836 9411 -19802
rect 10035 -19836 10045 -19802
rect 10045 -19836 10069 -19802
rect 10107 -19836 10113 -19802
rect 10113 -19836 10141 -19802
rect 10179 -19836 10181 -19802
rect 10181 -19836 10213 -19802
rect 10251 -19836 10283 -19802
rect 10283 -19836 10285 -19802
rect 10323 -19836 10351 -19802
rect 10351 -19836 10357 -19802
rect 10395 -19836 10419 -19802
rect 10419 -19836 10429 -19802
rect 11053 -19836 11063 -19802
rect 11063 -19836 11087 -19802
rect 11125 -19836 11131 -19802
rect 11131 -19836 11159 -19802
rect 11197 -19836 11199 -19802
rect 11199 -19836 11231 -19802
rect 11269 -19836 11301 -19802
rect 11301 -19836 11303 -19802
rect 11341 -19836 11369 -19802
rect 11369 -19836 11375 -19802
rect 11413 -19836 11437 -19802
rect 11437 -19836 11447 -19802
rect 12071 -19836 12081 -19802
rect 12081 -19836 12105 -19802
rect 12143 -19836 12149 -19802
rect 12149 -19836 12177 -19802
rect 12215 -19836 12217 -19802
rect 12217 -19836 12249 -19802
rect 12287 -19836 12319 -19802
rect 12319 -19836 12321 -19802
rect 12359 -19836 12387 -19802
rect 12387 -19836 12393 -19802
rect 12431 -19836 12455 -19802
rect 12455 -19836 12465 -19802
rect 13089 -19836 13099 -19802
rect 13099 -19836 13123 -19802
rect 13161 -19836 13167 -19802
rect 13167 -19836 13195 -19802
rect 13233 -19836 13235 -19802
rect 13235 -19836 13267 -19802
rect 13305 -19836 13337 -19802
rect 13337 -19836 13339 -19802
rect 13377 -19836 13405 -19802
rect 13405 -19836 13411 -19802
rect 13449 -19836 13473 -19802
rect 13473 -19836 13483 -19802
rect 14107 -19836 14117 -19802
rect 14117 -19836 14141 -19802
rect 14179 -19836 14185 -19802
rect 14185 -19836 14213 -19802
rect 14251 -19836 14253 -19802
rect 14253 -19836 14285 -19802
rect 14323 -19836 14355 -19802
rect 14355 -19836 14357 -19802
rect 14395 -19836 14423 -19802
rect 14423 -19836 14429 -19802
rect 14467 -19836 14491 -19802
rect 14491 -19836 14501 -19802
rect 15125 -19836 15135 -19802
rect 15135 -19836 15159 -19802
rect 15197 -19836 15203 -19802
rect 15203 -19836 15231 -19802
rect 15269 -19836 15271 -19802
rect 15271 -19836 15303 -19802
rect 15341 -19836 15373 -19802
rect 15373 -19836 15375 -19802
rect 15413 -19836 15441 -19802
rect 15441 -19836 15447 -19802
rect 15485 -19836 15509 -19802
rect 15509 -19836 15519 -19802
rect 16143 -19836 16153 -19802
rect 16153 -19836 16177 -19802
rect 16215 -19836 16221 -19802
rect 16221 -19836 16249 -19802
rect 16287 -19836 16289 -19802
rect 16289 -19836 16321 -19802
rect 16359 -19836 16391 -19802
rect 16391 -19836 16393 -19802
rect 16431 -19836 16459 -19802
rect 16459 -19836 16465 -19802
rect 16503 -19836 16527 -19802
rect 16527 -19836 16537 -19802
rect 17161 -19836 17171 -19802
rect 17171 -19836 17195 -19802
rect 17233 -19836 17239 -19802
rect 17239 -19836 17267 -19802
rect 17305 -19836 17307 -19802
rect 17307 -19836 17339 -19802
rect 17377 -19836 17409 -19802
rect 17409 -19836 17411 -19802
rect 17449 -19836 17477 -19802
rect 17477 -19836 17483 -19802
rect 17521 -19836 17545 -19802
rect 17545 -19836 17555 -19802
rect 18179 -19836 18189 -19802
rect 18189 -19836 18213 -19802
rect 18251 -19836 18257 -19802
rect 18257 -19836 18285 -19802
rect 18323 -19836 18325 -19802
rect 18325 -19836 18357 -19802
rect 18395 -19836 18427 -19802
rect 18427 -19836 18429 -19802
rect 18467 -19836 18495 -19802
rect 18495 -19836 18501 -19802
rect 18539 -19836 18563 -19802
rect 18563 -19836 18573 -19802
rect 19197 -19836 19207 -19802
rect 19207 -19836 19231 -19802
rect 19269 -19836 19275 -19802
rect 19275 -19836 19303 -19802
rect 19341 -19836 19343 -19802
rect 19343 -19836 19375 -19802
rect 19413 -19836 19445 -19802
rect 19445 -19836 19447 -19802
rect 19485 -19836 19513 -19802
rect 19513 -19836 19519 -19802
rect 19557 -19836 19581 -19802
rect 19581 -19836 19591 -19802
rect 20215 -19836 20225 -19802
rect 20225 -19836 20249 -19802
rect 20287 -19836 20293 -19802
rect 20293 -19836 20321 -19802
rect 20359 -19836 20361 -19802
rect 20361 -19836 20393 -19802
rect 20431 -19836 20463 -19802
rect 20463 -19836 20465 -19802
rect 20503 -19836 20531 -19802
rect 20531 -19836 20537 -19802
rect 20575 -19836 20599 -19802
rect 20599 -19836 20609 -19802
rect 21233 -19836 21243 -19802
rect 21243 -19836 21267 -19802
rect 21305 -19836 21311 -19802
rect 21311 -19836 21339 -19802
rect 21377 -19836 21379 -19802
rect 21379 -19836 21411 -19802
rect 21449 -19836 21481 -19802
rect 21481 -19836 21483 -19802
rect 21521 -19836 21549 -19802
rect 21549 -19836 21555 -19802
rect 21593 -19836 21617 -19802
rect 21617 -19836 21627 -19802
rect 22251 -19836 22261 -19802
rect 22261 -19836 22285 -19802
rect 22323 -19836 22329 -19802
rect 22329 -19836 22357 -19802
rect 22395 -19836 22397 -19802
rect 22397 -19836 22429 -19802
rect 22467 -19836 22499 -19802
rect 22499 -19836 22501 -19802
rect 22539 -19836 22567 -19802
rect 22567 -19836 22573 -19802
rect 22611 -19836 22635 -19802
rect 22635 -19836 22645 -19802
rect 24855 -19829 24889 -19795
rect -12289 -19897 -12255 -19867
rect -12289 -19901 -12255 -19897
rect -12289 -19965 -12255 -19939
rect -12289 -19973 -12255 -19965
rect -12289 -20033 -12255 -20011
rect -12289 -20045 -12255 -20033
rect -12289 -20101 -12255 -20083
rect -12289 -20117 -12255 -20101
rect -12289 -20169 -12255 -20155
rect -12289 -20189 -12255 -20169
rect -12289 -20237 -12255 -20227
rect -12289 -20261 -12255 -20237
rect -12289 -20305 -12255 -20299
rect -12289 -20333 -12255 -20305
rect 24855 -19897 24889 -19867
rect 24855 -19901 24889 -19897
rect 24855 -19965 24889 -19939
rect 24855 -19973 24889 -19965
rect 24855 -20033 24889 -20011
rect 24855 -20045 24889 -20033
rect 24855 -20101 24889 -20083
rect 24855 -20117 24889 -20101
rect 24855 -20169 24889 -20155
rect 24855 -20189 24889 -20169
rect 24855 -20237 24889 -20227
rect 24855 -20261 24889 -20237
rect -12289 -20373 -12255 -20371
rect -12289 -20405 -12255 -20373
rect 2909 -20360 2919 -20326
rect 2919 -20360 2943 -20326
rect 2981 -20360 2987 -20326
rect 2987 -20360 3015 -20326
rect 3053 -20360 3055 -20326
rect 3055 -20360 3087 -20326
rect 3125 -20360 3157 -20326
rect 3157 -20360 3159 -20326
rect 3197 -20360 3225 -20326
rect 3225 -20360 3231 -20326
rect 3269 -20360 3293 -20326
rect 3293 -20360 3303 -20326
rect 3927 -20360 3937 -20326
rect 3937 -20360 3961 -20326
rect 3999 -20360 4005 -20326
rect 4005 -20360 4033 -20326
rect 4071 -20360 4073 -20326
rect 4073 -20360 4105 -20326
rect 4143 -20360 4175 -20326
rect 4175 -20360 4177 -20326
rect 4215 -20360 4243 -20326
rect 4243 -20360 4249 -20326
rect 4287 -20360 4311 -20326
rect 4311 -20360 4321 -20326
rect 4945 -20360 4955 -20326
rect 4955 -20360 4979 -20326
rect 5017 -20360 5023 -20326
rect 5023 -20360 5051 -20326
rect 5089 -20360 5091 -20326
rect 5091 -20360 5123 -20326
rect 5161 -20360 5193 -20326
rect 5193 -20360 5195 -20326
rect 5233 -20360 5261 -20326
rect 5261 -20360 5267 -20326
rect 5305 -20360 5329 -20326
rect 5329 -20360 5339 -20326
rect 5963 -20360 5973 -20326
rect 5973 -20360 5997 -20326
rect 6035 -20360 6041 -20326
rect 6041 -20360 6069 -20326
rect 6107 -20360 6109 -20326
rect 6109 -20360 6141 -20326
rect 6179 -20360 6211 -20326
rect 6211 -20360 6213 -20326
rect 6251 -20360 6279 -20326
rect 6279 -20360 6285 -20326
rect 6323 -20360 6347 -20326
rect 6347 -20360 6357 -20326
rect 6981 -20360 6991 -20326
rect 6991 -20360 7015 -20326
rect 7053 -20360 7059 -20326
rect 7059 -20360 7087 -20326
rect 7125 -20360 7127 -20326
rect 7127 -20360 7159 -20326
rect 7197 -20360 7229 -20326
rect 7229 -20360 7231 -20326
rect 7269 -20360 7297 -20326
rect 7297 -20360 7303 -20326
rect 7341 -20360 7365 -20326
rect 7365 -20360 7375 -20326
rect 7999 -20360 8009 -20326
rect 8009 -20360 8033 -20326
rect 8071 -20360 8077 -20326
rect 8077 -20360 8105 -20326
rect 8143 -20360 8145 -20326
rect 8145 -20360 8177 -20326
rect 8215 -20360 8247 -20326
rect 8247 -20360 8249 -20326
rect 8287 -20360 8315 -20326
rect 8315 -20360 8321 -20326
rect 8359 -20360 8383 -20326
rect 8383 -20360 8393 -20326
rect 9017 -20360 9027 -20326
rect 9027 -20360 9051 -20326
rect 9089 -20360 9095 -20326
rect 9095 -20360 9123 -20326
rect 9161 -20360 9163 -20326
rect 9163 -20360 9195 -20326
rect 9233 -20360 9265 -20326
rect 9265 -20360 9267 -20326
rect 9305 -20360 9333 -20326
rect 9333 -20360 9339 -20326
rect 9377 -20360 9401 -20326
rect 9401 -20360 9411 -20326
rect 10035 -20360 10045 -20326
rect 10045 -20360 10069 -20326
rect 10107 -20360 10113 -20326
rect 10113 -20360 10141 -20326
rect 10179 -20360 10181 -20326
rect 10181 -20360 10213 -20326
rect 10251 -20360 10283 -20326
rect 10283 -20360 10285 -20326
rect 10323 -20360 10351 -20326
rect 10351 -20360 10357 -20326
rect 10395 -20360 10419 -20326
rect 10419 -20360 10429 -20326
rect 11053 -20360 11063 -20326
rect 11063 -20360 11087 -20326
rect 11125 -20360 11131 -20326
rect 11131 -20360 11159 -20326
rect 11197 -20360 11199 -20326
rect 11199 -20360 11231 -20326
rect 11269 -20360 11301 -20326
rect 11301 -20360 11303 -20326
rect 11341 -20360 11369 -20326
rect 11369 -20360 11375 -20326
rect 11413 -20360 11437 -20326
rect 11437 -20360 11447 -20326
rect 12071 -20360 12081 -20326
rect 12081 -20360 12105 -20326
rect 12143 -20360 12149 -20326
rect 12149 -20360 12177 -20326
rect 12215 -20360 12217 -20326
rect 12217 -20360 12249 -20326
rect 12287 -20360 12319 -20326
rect 12319 -20360 12321 -20326
rect 12359 -20360 12387 -20326
rect 12387 -20360 12393 -20326
rect 12431 -20360 12455 -20326
rect 12455 -20360 12465 -20326
rect 13089 -20360 13099 -20326
rect 13099 -20360 13123 -20326
rect 13161 -20360 13167 -20326
rect 13167 -20360 13195 -20326
rect 13233 -20360 13235 -20326
rect 13235 -20360 13267 -20326
rect 13305 -20360 13337 -20326
rect 13337 -20360 13339 -20326
rect 13377 -20360 13405 -20326
rect 13405 -20360 13411 -20326
rect 13449 -20360 13473 -20326
rect 13473 -20360 13483 -20326
rect 14107 -20360 14117 -20326
rect 14117 -20360 14141 -20326
rect 14179 -20360 14185 -20326
rect 14185 -20360 14213 -20326
rect 14251 -20360 14253 -20326
rect 14253 -20360 14285 -20326
rect 14323 -20360 14355 -20326
rect 14355 -20360 14357 -20326
rect 14395 -20360 14423 -20326
rect 14423 -20360 14429 -20326
rect 14467 -20360 14491 -20326
rect 14491 -20360 14501 -20326
rect 15125 -20360 15135 -20326
rect 15135 -20360 15159 -20326
rect 15197 -20360 15203 -20326
rect 15203 -20360 15231 -20326
rect 15269 -20360 15271 -20326
rect 15271 -20360 15303 -20326
rect 15341 -20360 15373 -20326
rect 15373 -20360 15375 -20326
rect 15413 -20360 15441 -20326
rect 15441 -20360 15447 -20326
rect 15485 -20360 15509 -20326
rect 15509 -20360 15519 -20326
rect 16143 -20360 16153 -20326
rect 16153 -20360 16177 -20326
rect 16215 -20360 16221 -20326
rect 16221 -20360 16249 -20326
rect 16287 -20360 16289 -20326
rect 16289 -20360 16321 -20326
rect 16359 -20360 16391 -20326
rect 16391 -20360 16393 -20326
rect 16431 -20360 16459 -20326
rect 16459 -20360 16465 -20326
rect 16503 -20360 16527 -20326
rect 16527 -20360 16537 -20326
rect 17161 -20360 17171 -20326
rect 17171 -20360 17195 -20326
rect 17233 -20360 17239 -20326
rect 17239 -20360 17267 -20326
rect 17305 -20360 17307 -20326
rect 17307 -20360 17339 -20326
rect 17377 -20360 17409 -20326
rect 17409 -20360 17411 -20326
rect 17449 -20360 17477 -20326
rect 17477 -20360 17483 -20326
rect 17521 -20360 17545 -20326
rect 17545 -20360 17555 -20326
rect 18179 -20360 18189 -20326
rect 18189 -20360 18213 -20326
rect 18251 -20360 18257 -20326
rect 18257 -20360 18285 -20326
rect 18323 -20360 18325 -20326
rect 18325 -20360 18357 -20326
rect 18395 -20360 18427 -20326
rect 18427 -20360 18429 -20326
rect 18467 -20360 18495 -20326
rect 18495 -20360 18501 -20326
rect 18539 -20360 18563 -20326
rect 18563 -20360 18573 -20326
rect 19197 -20360 19207 -20326
rect 19207 -20360 19231 -20326
rect 19269 -20360 19275 -20326
rect 19275 -20360 19303 -20326
rect 19341 -20360 19343 -20326
rect 19343 -20360 19375 -20326
rect 19413 -20360 19445 -20326
rect 19445 -20360 19447 -20326
rect 19485 -20360 19513 -20326
rect 19513 -20360 19519 -20326
rect 19557 -20360 19581 -20326
rect 19581 -20360 19591 -20326
rect 20215 -20360 20225 -20326
rect 20225 -20360 20249 -20326
rect 20287 -20360 20293 -20326
rect 20293 -20360 20321 -20326
rect 20359 -20360 20361 -20326
rect 20361 -20360 20393 -20326
rect 20431 -20360 20463 -20326
rect 20463 -20360 20465 -20326
rect 20503 -20360 20531 -20326
rect 20531 -20360 20537 -20326
rect 20575 -20360 20599 -20326
rect 20599 -20360 20609 -20326
rect 21233 -20360 21243 -20326
rect 21243 -20360 21267 -20326
rect 21305 -20360 21311 -20326
rect 21311 -20360 21339 -20326
rect 21377 -20360 21379 -20326
rect 21379 -20360 21411 -20326
rect 21449 -20360 21481 -20326
rect 21481 -20360 21483 -20326
rect 21521 -20360 21549 -20326
rect 21549 -20360 21555 -20326
rect 21593 -20360 21617 -20326
rect 21617 -20360 21627 -20326
rect 22251 -20360 22261 -20326
rect 22261 -20360 22285 -20326
rect 22323 -20360 22329 -20326
rect 22329 -20360 22357 -20326
rect 22395 -20360 22397 -20326
rect 22397 -20360 22429 -20326
rect 22467 -20360 22499 -20326
rect 22499 -20360 22501 -20326
rect 22539 -20360 22567 -20326
rect 22567 -20360 22573 -20326
rect 22611 -20360 22635 -20326
rect 22635 -20360 22645 -20326
rect 24855 -20305 24889 -20299
rect 24855 -20333 24889 -20305
rect -12289 -20475 -12255 -20443
rect -12289 -20477 -12255 -20475
rect -12289 -20543 -12255 -20515
rect -12289 -20549 -12255 -20543
rect -12289 -20611 -12255 -20587
rect -12289 -20621 -12255 -20611
rect -12289 -20679 -12255 -20659
rect -12289 -20693 -12255 -20679
rect -12289 -20747 -12255 -20731
rect -12289 -20765 -12255 -20747
rect -12289 -20815 -12255 -20803
rect -12289 -20837 -12255 -20815
rect -12289 -20883 -12255 -20875
rect -12289 -20909 -12255 -20883
rect -12289 -20951 -12255 -20947
rect -12289 -20981 -12255 -20951
rect 2580 -20443 2614 -20429
rect 2580 -20463 2614 -20443
rect 2580 -20511 2614 -20501
rect 2580 -20535 2614 -20511
rect 2580 -20579 2614 -20573
rect 2580 -20607 2614 -20579
rect 2580 -20647 2614 -20645
rect 2580 -20679 2614 -20647
rect 2580 -20749 2614 -20717
rect 2580 -20751 2614 -20749
rect 2580 -20817 2614 -20789
rect 2580 -20823 2614 -20817
rect 2580 -20885 2614 -20861
rect 2580 -20895 2614 -20885
rect 2580 -20953 2614 -20933
rect 2580 -20967 2614 -20953
rect 3598 -20443 3632 -20429
rect 3598 -20463 3632 -20443
rect 3598 -20511 3632 -20501
rect 3598 -20535 3632 -20511
rect 3598 -20579 3632 -20573
rect 3598 -20607 3632 -20579
rect 3598 -20647 3632 -20645
rect 3598 -20679 3632 -20647
rect 3598 -20749 3632 -20717
rect 3598 -20751 3632 -20749
rect 3598 -20817 3632 -20789
rect 3598 -20823 3632 -20817
rect 3598 -20885 3632 -20861
rect 3598 -20895 3632 -20885
rect 3598 -20953 3632 -20933
rect 3598 -20967 3632 -20953
rect 4616 -20443 4650 -20429
rect 4616 -20463 4650 -20443
rect 4616 -20511 4650 -20501
rect 4616 -20535 4650 -20511
rect 4616 -20579 4650 -20573
rect 4616 -20607 4650 -20579
rect 4616 -20647 4650 -20645
rect 4616 -20679 4650 -20647
rect 4616 -20749 4650 -20717
rect 4616 -20751 4650 -20749
rect 4616 -20817 4650 -20789
rect 4616 -20823 4650 -20817
rect 4616 -20885 4650 -20861
rect 4616 -20895 4650 -20885
rect 4616 -20953 4650 -20933
rect 4616 -20967 4650 -20953
rect 5634 -20443 5668 -20429
rect 5634 -20463 5668 -20443
rect 5634 -20511 5668 -20501
rect 5634 -20535 5668 -20511
rect 5634 -20579 5668 -20573
rect 5634 -20607 5668 -20579
rect 5634 -20647 5668 -20645
rect 5634 -20679 5668 -20647
rect 5634 -20749 5668 -20717
rect 5634 -20751 5668 -20749
rect 5634 -20817 5668 -20789
rect 5634 -20823 5668 -20817
rect 5634 -20885 5668 -20861
rect 5634 -20895 5668 -20885
rect 5634 -20953 5668 -20933
rect 5634 -20967 5668 -20953
rect 6652 -20443 6686 -20429
rect 6652 -20463 6686 -20443
rect 6652 -20511 6686 -20501
rect 6652 -20535 6686 -20511
rect 6652 -20579 6686 -20573
rect 6652 -20607 6686 -20579
rect 6652 -20647 6686 -20645
rect 6652 -20679 6686 -20647
rect 6652 -20749 6686 -20717
rect 6652 -20751 6686 -20749
rect 6652 -20817 6686 -20789
rect 6652 -20823 6686 -20817
rect 6652 -20885 6686 -20861
rect 6652 -20895 6686 -20885
rect 6652 -20953 6686 -20933
rect 6652 -20967 6686 -20953
rect 7670 -20443 7704 -20429
rect 7670 -20463 7704 -20443
rect 7670 -20511 7704 -20501
rect 7670 -20535 7704 -20511
rect 7670 -20579 7704 -20573
rect 7670 -20607 7704 -20579
rect 7670 -20647 7704 -20645
rect 7670 -20679 7704 -20647
rect 7670 -20749 7704 -20717
rect 7670 -20751 7704 -20749
rect 7670 -20817 7704 -20789
rect 7670 -20823 7704 -20817
rect 7670 -20885 7704 -20861
rect 7670 -20895 7704 -20885
rect 7670 -20953 7704 -20933
rect 7670 -20967 7704 -20953
rect 8688 -20443 8722 -20429
rect 8688 -20463 8722 -20443
rect 8688 -20511 8722 -20501
rect 8688 -20535 8722 -20511
rect 8688 -20579 8722 -20573
rect 8688 -20607 8722 -20579
rect 8688 -20647 8722 -20645
rect 8688 -20679 8722 -20647
rect 8688 -20749 8722 -20717
rect 8688 -20751 8722 -20749
rect 8688 -20817 8722 -20789
rect 8688 -20823 8722 -20817
rect 8688 -20885 8722 -20861
rect 8688 -20895 8722 -20885
rect 8688 -20953 8722 -20933
rect 8688 -20967 8722 -20953
rect 9706 -20443 9740 -20429
rect 9706 -20463 9740 -20443
rect 9706 -20511 9740 -20501
rect 9706 -20535 9740 -20511
rect 9706 -20579 9740 -20573
rect 9706 -20607 9740 -20579
rect 9706 -20647 9740 -20645
rect 9706 -20679 9740 -20647
rect 9706 -20749 9740 -20717
rect 9706 -20751 9740 -20749
rect 9706 -20817 9740 -20789
rect 9706 -20823 9740 -20817
rect 9706 -20885 9740 -20861
rect 9706 -20895 9740 -20885
rect 9706 -20953 9740 -20933
rect 9706 -20967 9740 -20953
rect 10724 -20443 10758 -20429
rect 10724 -20463 10758 -20443
rect 10724 -20511 10758 -20501
rect 10724 -20535 10758 -20511
rect 10724 -20579 10758 -20573
rect 10724 -20607 10758 -20579
rect 10724 -20647 10758 -20645
rect 10724 -20679 10758 -20647
rect 10724 -20749 10758 -20717
rect 10724 -20751 10758 -20749
rect 10724 -20817 10758 -20789
rect 10724 -20823 10758 -20817
rect 10724 -20885 10758 -20861
rect 10724 -20895 10758 -20885
rect 10724 -20953 10758 -20933
rect 10724 -20967 10758 -20953
rect 11742 -20443 11776 -20429
rect 11742 -20463 11776 -20443
rect 11742 -20511 11776 -20501
rect 11742 -20535 11776 -20511
rect 11742 -20579 11776 -20573
rect 11742 -20607 11776 -20579
rect 11742 -20647 11776 -20645
rect 11742 -20679 11776 -20647
rect 11742 -20749 11776 -20717
rect 11742 -20751 11776 -20749
rect 11742 -20817 11776 -20789
rect 11742 -20823 11776 -20817
rect 11742 -20885 11776 -20861
rect 11742 -20895 11776 -20885
rect 11742 -20953 11776 -20933
rect 11742 -20967 11776 -20953
rect 12760 -20443 12794 -20429
rect 12760 -20463 12794 -20443
rect 12760 -20511 12794 -20501
rect 12760 -20535 12794 -20511
rect 12760 -20579 12794 -20573
rect 12760 -20607 12794 -20579
rect 12760 -20647 12794 -20645
rect 12760 -20679 12794 -20647
rect 12760 -20749 12794 -20717
rect 12760 -20751 12794 -20749
rect 12760 -20817 12794 -20789
rect 12760 -20823 12794 -20817
rect 12760 -20885 12794 -20861
rect 12760 -20895 12794 -20885
rect 12760 -20953 12794 -20933
rect 12760 -20967 12794 -20953
rect 13778 -20443 13812 -20429
rect 13778 -20463 13812 -20443
rect 13778 -20511 13812 -20501
rect 13778 -20535 13812 -20511
rect 13778 -20579 13812 -20573
rect 13778 -20607 13812 -20579
rect 13778 -20647 13812 -20645
rect 13778 -20679 13812 -20647
rect 13778 -20749 13812 -20717
rect 13778 -20751 13812 -20749
rect 13778 -20817 13812 -20789
rect 13778 -20823 13812 -20817
rect 13778 -20885 13812 -20861
rect 13778 -20895 13812 -20885
rect 13778 -20953 13812 -20933
rect 13778 -20967 13812 -20953
rect 14796 -20443 14830 -20429
rect 14796 -20463 14830 -20443
rect 14796 -20511 14830 -20501
rect 14796 -20535 14830 -20511
rect 14796 -20579 14830 -20573
rect 14796 -20607 14830 -20579
rect 14796 -20647 14830 -20645
rect 14796 -20679 14830 -20647
rect 14796 -20749 14830 -20717
rect 14796 -20751 14830 -20749
rect 14796 -20817 14830 -20789
rect 14796 -20823 14830 -20817
rect 14796 -20885 14830 -20861
rect 14796 -20895 14830 -20885
rect 14796 -20953 14830 -20933
rect 14796 -20967 14830 -20953
rect 15814 -20443 15848 -20429
rect 15814 -20463 15848 -20443
rect 15814 -20511 15848 -20501
rect 15814 -20535 15848 -20511
rect 15814 -20579 15848 -20573
rect 15814 -20607 15848 -20579
rect 15814 -20647 15848 -20645
rect 15814 -20679 15848 -20647
rect 15814 -20749 15848 -20717
rect 15814 -20751 15848 -20749
rect 15814 -20817 15848 -20789
rect 15814 -20823 15848 -20817
rect 15814 -20885 15848 -20861
rect 15814 -20895 15848 -20885
rect 15814 -20953 15848 -20933
rect 15814 -20967 15848 -20953
rect 16832 -20443 16866 -20429
rect 16832 -20463 16866 -20443
rect 16832 -20511 16866 -20501
rect 16832 -20535 16866 -20511
rect 16832 -20579 16866 -20573
rect 16832 -20607 16866 -20579
rect 16832 -20647 16866 -20645
rect 16832 -20679 16866 -20647
rect 16832 -20749 16866 -20717
rect 16832 -20751 16866 -20749
rect 16832 -20817 16866 -20789
rect 16832 -20823 16866 -20817
rect 16832 -20885 16866 -20861
rect 16832 -20895 16866 -20885
rect 16832 -20953 16866 -20933
rect 16832 -20967 16866 -20953
rect 17850 -20443 17884 -20429
rect 17850 -20463 17884 -20443
rect 17850 -20511 17884 -20501
rect 17850 -20535 17884 -20511
rect 17850 -20579 17884 -20573
rect 17850 -20607 17884 -20579
rect 17850 -20647 17884 -20645
rect 17850 -20679 17884 -20647
rect 17850 -20749 17884 -20717
rect 17850 -20751 17884 -20749
rect 17850 -20817 17884 -20789
rect 17850 -20823 17884 -20817
rect 17850 -20885 17884 -20861
rect 17850 -20895 17884 -20885
rect 17850 -20953 17884 -20933
rect 17850 -20967 17884 -20953
rect 18868 -20443 18902 -20429
rect 18868 -20463 18902 -20443
rect 18868 -20511 18902 -20501
rect 18868 -20535 18902 -20511
rect 18868 -20579 18902 -20573
rect 18868 -20607 18902 -20579
rect 18868 -20647 18902 -20645
rect 18868 -20679 18902 -20647
rect 18868 -20749 18902 -20717
rect 18868 -20751 18902 -20749
rect 18868 -20817 18902 -20789
rect 18868 -20823 18902 -20817
rect 18868 -20885 18902 -20861
rect 18868 -20895 18902 -20885
rect 18868 -20953 18902 -20933
rect 18868 -20967 18902 -20953
rect 19886 -20443 19920 -20429
rect 19886 -20463 19920 -20443
rect 19886 -20511 19920 -20501
rect 19886 -20535 19920 -20511
rect 19886 -20579 19920 -20573
rect 19886 -20607 19920 -20579
rect 19886 -20647 19920 -20645
rect 19886 -20679 19920 -20647
rect 19886 -20749 19920 -20717
rect 19886 -20751 19920 -20749
rect 19886 -20817 19920 -20789
rect 19886 -20823 19920 -20817
rect 19886 -20885 19920 -20861
rect 19886 -20895 19920 -20885
rect 19886 -20953 19920 -20933
rect 19886 -20967 19920 -20953
rect 20904 -20443 20938 -20429
rect 20904 -20463 20938 -20443
rect 20904 -20511 20938 -20501
rect 20904 -20535 20938 -20511
rect 20904 -20579 20938 -20573
rect 20904 -20607 20938 -20579
rect 20904 -20647 20938 -20645
rect 20904 -20679 20938 -20647
rect 20904 -20749 20938 -20717
rect 20904 -20751 20938 -20749
rect 20904 -20817 20938 -20789
rect 20904 -20823 20938 -20817
rect 20904 -20885 20938 -20861
rect 20904 -20895 20938 -20885
rect 20904 -20953 20938 -20933
rect 20904 -20967 20938 -20953
rect 21922 -20443 21956 -20429
rect 21922 -20463 21956 -20443
rect 21922 -20511 21956 -20501
rect 21922 -20535 21956 -20511
rect 21922 -20579 21956 -20573
rect 21922 -20607 21956 -20579
rect 21922 -20647 21956 -20645
rect 21922 -20679 21956 -20647
rect 21922 -20749 21956 -20717
rect 21922 -20751 21956 -20749
rect 21922 -20817 21956 -20789
rect 21922 -20823 21956 -20817
rect 21922 -20885 21956 -20861
rect 21922 -20895 21956 -20885
rect 21922 -20953 21956 -20933
rect 21922 -20967 21956 -20953
rect 22940 -20443 22974 -20429
rect 22940 -20463 22974 -20443
rect 22940 -20511 22974 -20501
rect 22940 -20535 22974 -20511
rect 22940 -20579 22974 -20573
rect 22940 -20607 22974 -20579
rect 22940 -20647 22974 -20645
rect 22940 -20679 22974 -20647
rect 22940 -20749 22974 -20717
rect 22940 -20751 22974 -20749
rect 22940 -20817 22974 -20789
rect 22940 -20823 22974 -20817
rect 22940 -20885 22974 -20861
rect 22940 -20895 22974 -20885
rect 22940 -20953 22974 -20933
rect 22940 -20967 22974 -20953
rect 24855 -20373 24889 -20371
rect 24855 -20405 24889 -20373
rect 24855 -20475 24889 -20443
rect 24855 -20477 24889 -20475
rect 24855 -20543 24889 -20515
rect 24855 -20549 24889 -20543
rect 24855 -20611 24889 -20587
rect 24855 -20621 24889 -20611
rect 24855 -20679 24889 -20659
rect 24855 -20693 24889 -20679
rect 24855 -20747 24889 -20731
rect 24855 -20765 24889 -20747
rect 24855 -20815 24889 -20803
rect 24855 -20837 24889 -20815
rect 24855 -20883 24889 -20875
rect 24855 -20909 24889 -20883
rect 24855 -20951 24889 -20947
rect 24855 -20981 24889 -20951
rect -12289 -21053 -12255 -21019
rect 2909 -21070 2919 -21036
rect 2919 -21070 2943 -21036
rect 2981 -21070 2987 -21036
rect 2987 -21070 3015 -21036
rect 3053 -21070 3055 -21036
rect 3055 -21070 3087 -21036
rect 3125 -21070 3157 -21036
rect 3157 -21070 3159 -21036
rect 3197 -21070 3225 -21036
rect 3225 -21070 3231 -21036
rect 3269 -21070 3293 -21036
rect 3293 -21070 3303 -21036
rect 3927 -21070 3937 -21036
rect 3937 -21070 3961 -21036
rect 3999 -21070 4005 -21036
rect 4005 -21070 4033 -21036
rect 4071 -21070 4073 -21036
rect 4073 -21070 4105 -21036
rect 4143 -21070 4175 -21036
rect 4175 -21070 4177 -21036
rect 4215 -21070 4243 -21036
rect 4243 -21070 4249 -21036
rect 4287 -21070 4311 -21036
rect 4311 -21070 4321 -21036
rect 4945 -21070 4955 -21036
rect 4955 -21070 4979 -21036
rect 5017 -21070 5023 -21036
rect 5023 -21070 5051 -21036
rect 5089 -21070 5091 -21036
rect 5091 -21070 5123 -21036
rect 5161 -21070 5193 -21036
rect 5193 -21070 5195 -21036
rect 5233 -21070 5261 -21036
rect 5261 -21070 5267 -21036
rect 5305 -21070 5329 -21036
rect 5329 -21070 5339 -21036
rect 5963 -21070 5973 -21036
rect 5973 -21070 5997 -21036
rect 6035 -21070 6041 -21036
rect 6041 -21070 6069 -21036
rect 6107 -21070 6109 -21036
rect 6109 -21070 6141 -21036
rect 6179 -21070 6211 -21036
rect 6211 -21070 6213 -21036
rect 6251 -21070 6279 -21036
rect 6279 -21070 6285 -21036
rect 6323 -21070 6347 -21036
rect 6347 -21070 6357 -21036
rect 6981 -21070 6991 -21036
rect 6991 -21070 7015 -21036
rect 7053 -21070 7059 -21036
rect 7059 -21070 7087 -21036
rect 7125 -21070 7127 -21036
rect 7127 -21070 7159 -21036
rect 7197 -21070 7229 -21036
rect 7229 -21070 7231 -21036
rect 7269 -21070 7297 -21036
rect 7297 -21070 7303 -21036
rect 7341 -21070 7365 -21036
rect 7365 -21070 7375 -21036
rect 7999 -21070 8009 -21036
rect 8009 -21070 8033 -21036
rect 8071 -21070 8077 -21036
rect 8077 -21070 8105 -21036
rect 8143 -21070 8145 -21036
rect 8145 -21070 8177 -21036
rect 8215 -21070 8247 -21036
rect 8247 -21070 8249 -21036
rect 8287 -21070 8315 -21036
rect 8315 -21070 8321 -21036
rect 8359 -21070 8383 -21036
rect 8383 -21070 8393 -21036
rect 9017 -21070 9027 -21036
rect 9027 -21070 9051 -21036
rect 9089 -21070 9095 -21036
rect 9095 -21070 9123 -21036
rect 9161 -21070 9163 -21036
rect 9163 -21070 9195 -21036
rect 9233 -21070 9265 -21036
rect 9265 -21070 9267 -21036
rect 9305 -21070 9333 -21036
rect 9333 -21070 9339 -21036
rect 9377 -21070 9401 -21036
rect 9401 -21070 9411 -21036
rect 10035 -21070 10045 -21036
rect 10045 -21070 10069 -21036
rect 10107 -21070 10113 -21036
rect 10113 -21070 10141 -21036
rect 10179 -21070 10181 -21036
rect 10181 -21070 10213 -21036
rect 10251 -21070 10283 -21036
rect 10283 -21070 10285 -21036
rect 10323 -21070 10351 -21036
rect 10351 -21070 10357 -21036
rect 10395 -21070 10419 -21036
rect 10419 -21070 10429 -21036
rect 11053 -21070 11063 -21036
rect 11063 -21070 11087 -21036
rect 11125 -21070 11131 -21036
rect 11131 -21070 11159 -21036
rect 11197 -21070 11199 -21036
rect 11199 -21070 11231 -21036
rect 11269 -21070 11301 -21036
rect 11301 -21070 11303 -21036
rect 11341 -21070 11369 -21036
rect 11369 -21070 11375 -21036
rect 11413 -21070 11437 -21036
rect 11437 -21070 11447 -21036
rect 12071 -21070 12081 -21036
rect 12081 -21070 12105 -21036
rect 12143 -21070 12149 -21036
rect 12149 -21070 12177 -21036
rect 12215 -21070 12217 -21036
rect 12217 -21070 12249 -21036
rect 12287 -21070 12319 -21036
rect 12319 -21070 12321 -21036
rect 12359 -21070 12387 -21036
rect 12387 -21070 12393 -21036
rect 12431 -21070 12455 -21036
rect 12455 -21070 12465 -21036
rect 13089 -21070 13099 -21036
rect 13099 -21070 13123 -21036
rect 13161 -21070 13167 -21036
rect 13167 -21070 13195 -21036
rect 13233 -21070 13235 -21036
rect 13235 -21070 13267 -21036
rect 13305 -21070 13337 -21036
rect 13337 -21070 13339 -21036
rect 13377 -21070 13405 -21036
rect 13405 -21070 13411 -21036
rect 13449 -21070 13473 -21036
rect 13473 -21070 13483 -21036
rect 14107 -21070 14117 -21036
rect 14117 -21070 14141 -21036
rect 14179 -21070 14185 -21036
rect 14185 -21070 14213 -21036
rect 14251 -21070 14253 -21036
rect 14253 -21070 14285 -21036
rect 14323 -21070 14355 -21036
rect 14355 -21070 14357 -21036
rect 14395 -21070 14423 -21036
rect 14423 -21070 14429 -21036
rect 14467 -21070 14491 -21036
rect 14491 -21070 14501 -21036
rect 15125 -21070 15135 -21036
rect 15135 -21070 15159 -21036
rect 15197 -21070 15203 -21036
rect 15203 -21070 15231 -21036
rect 15269 -21070 15271 -21036
rect 15271 -21070 15303 -21036
rect 15341 -21070 15373 -21036
rect 15373 -21070 15375 -21036
rect 15413 -21070 15441 -21036
rect 15441 -21070 15447 -21036
rect 15485 -21070 15509 -21036
rect 15509 -21070 15519 -21036
rect 16143 -21070 16153 -21036
rect 16153 -21070 16177 -21036
rect 16215 -21070 16221 -21036
rect 16221 -21070 16249 -21036
rect 16287 -21070 16289 -21036
rect 16289 -21070 16321 -21036
rect 16359 -21070 16391 -21036
rect 16391 -21070 16393 -21036
rect 16431 -21070 16459 -21036
rect 16459 -21070 16465 -21036
rect 16503 -21070 16527 -21036
rect 16527 -21070 16537 -21036
rect 17161 -21070 17171 -21036
rect 17171 -21070 17195 -21036
rect 17233 -21070 17239 -21036
rect 17239 -21070 17267 -21036
rect 17305 -21070 17307 -21036
rect 17307 -21070 17339 -21036
rect 17377 -21070 17409 -21036
rect 17409 -21070 17411 -21036
rect 17449 -21070 17477 -21036
rect 17477 -21070 17483 -21036
rect 17521 -21070 17545 -21036
rect 17545 -21070 17555 -21036
rect 18179 -21070 18189 -21036
rect 18189 -21070 18213 -21036
rect 18251 -21070 18257 -21036
rect 18257 -21070 18285 -21036
rect 18323 -21070 18325 -21036
rect 18325 -21070 18357 -21036
rect 18395 -21070 18427 -21036
rect 18427 -21070 18429 -21036
rect 18467 -21070 18495 -21036
rect 18495 -21070 18501 -21036
rect 18539 -21070 18563 -21036
rect 18563 -21070 18573 -21036
rect 19197 -21070 19207 -21036
rect 19207 -21070 19231 -21036
rect 19269 -21070 19275 -21036
rect 19275 -21070 19303 -21036
rect 19341 -21070 19343 -21036
rect 19343 -21070 19375 -21036
rect 19413 -21070 19445 -21036
rect 19445 -21070 19447 -21036
rect 19485 -21070 19513 -21036
rect 19513 -21070 19519 -21036
rect 19557 -21070 19581 -21036
rect 19581 -21070 19591 -21036
rect 20215 -21070 20225 -21036
rect 20225 -21070 20249 -21036
rect 20287 -21070 20293 -21036
rect 20293 -21070 20321 -21036
rect 20359 -21070 20361 -21036
rect 20361 -21070 20393 -21036
rect 20431 -21070 20463 -21036
rect 20463 -21070 20465 -21036
rect 20503 -21070 20531 -21036
rect 20531 -21070 20537 -21036
rect 20575 -21070 20599 -21036
rect 20599 -21070 20609 -21036
rect 21233 -21070 21243 -21036
rect 21243 -21070 21267 -21036
rect 21305 -21070 21311 -21036
rect 21311 -21070 21339 -21036
rect 21377 -21070 21379 -21036
rect 21379 -21070 21411 -21036
rect 21449 -21070 21481 -21036
rect 21481 -21070 21483 -21036
rect 21521 -21070 21549 -21036
rect 21549 -21070 21555 -21036
rect 21593 -21070 21617 -21036
rect 21617 -21070 21627 -21036
rect 22251 -21070 22261 -21036
rect 22261 -21070 22285 -21036
rect 22323 -21070 22329 -21036
rect 22329 -21070 22357 -21036
rect 22395 -21070 22397 -21036
rect 22397 -21070 22429 -21036
rect 22467 -21070 22499 -21036
rect 22499 -21070 22501 -21036
rect 22539 -21070 22567 -21036
rect 22567 -21070 22573 -21036
rect 22611 -21070 22635 -21036
rect 22635 -21070 22645 -21036
rect 24855 -21053 24889 -21019
rect -12289 -21121 -12255 -21091
rect -12289 -21125 -12255 -21121
rect -12289 -21189 -12255 -21163
rect -12289 -21197 -12255 -21189
rect -12289 -21257 -12255 -21235
rect -12289 -21269 -12255 -21257
rect -12289 -21325 -12255 -21307
rect -12289 -21341 -12255 -21325
rect -12289 -21393 -12255 -21379
rect -12289 -21413 -12255 -21393
rect -12289 -21461 -12255 -21451
rect -12289 -21485 -12255 -21461
rect -12289 -21529 -12255 -21523
rect -12289 -21557 -12255 -21529
rect 24855 -21121 24889 -21091
rect 24855 -21125 24889 -21121
rect 24855 -21189 24889 -21163
rect 24855 -21197 24889 -21189
rect 24855 -21257 24889 -21235
rect 24855 -21269 24889 -21257
rect 24855 -21325 24889 -21307
rect 24855 -21341 24889 -21325
rect 24855 -21393 24889 -21379
rect 24855 -21413 24889 -21393
rect 24855 -21461 24889 -21451
rect 24855 -21485 24889 -21461
rect 24855 -21529 24889 -21523
rect 24855 -21557 24889 -21529
rect -12289 -21597 -12255 -21595
rect -12289 -21629 -12255 -21597
rect 2909 -21594 2919 -21560
rect 2919 -21594 2943 -21560
rect 2981 -21594 2987 -21560
rect 2987 -21594 3015 -21560
rect 3053 -21594 3055 -21560
rect 3055 -21594 3087 -21560
rect 3125 -21594 3157 -21560
rect 3157 -21594 3159 -21560
rect 3197 -21594 3225 -21560
rect 3225 -21594 3231 -21560
rect 3269 -21594 3293 -21560
rect 3293 -21594 3303 -21560
rect 3927 -21594 3937 -21560
rect 3937 -21594 3961 -21560
rect 3999 -21594 4005 -21560
rect 4005 -21594 4033 -21560
rect 4071 -21594 4073 -21560
rect 4073 -21594 4105 -21560
rect 4143 -21594 4175 -21560
rect 4175 -21594 4177 -21560
rect 4215 -21594 4243 -21560
rect 4243 -21594 4249 -21560
rect 4287 -21594 4311 -21560
rect 4311 -21594 4321 -21560
rect 4945 -21594 4955 -21560
rect 4955 -21594 4979 -21560
rect 5017 -21594 5023 -21560
rect 5023 -21594 5051 -21560
rect 5089 -21594 5091 -21560
rect 5091 -21594 5123 -21560
rect 5161 -21594 5193 -21560
rect 5193 -21594 5195 -21560
rect 5233 -21594 5261 -21560
rect 5261 -21594 5267 -21560
rect 5305 -21594 5329 -21560
rect 5329 -21594 5339 -21560
rect 5963 -21594 5973 -21560
rect 5973 -21594 5997 -21560
rect 6035 -21594 6041 -21560
rect 6041 -21594 6069 -21560
rect 6107 -21594 6109 -21560
rect 6109 -21594 6141 -21560
rect 6179 -21594 6211 -21560
rect 6211 -21594 6213 -21560
rect 6251 -21594 6279 -21560
rect 6279 -21594 6285 -21560
rect 6323 -21594 6347 -21560
rect 6347 -21594 6357 -21560
rect 6981 -21594 6991 -21560
rect 6991 -21594 7015 -21560
rect 7053 -21594 7059 -21560
rect 7059 -21594 7087 -21560
rect 7125 -21594 7127 -21560
rect 7127 -21594 7159 -21560
rect 7197 -21594 7229 -21560
rect 7229 -21594 7231 -21560
rect 7269 -21594 7297 -21560
rect 7297 -21594 7303 -21560
rect 7341 -21594 7365 -21560
rect 7365 -21594 7375 -21560
rect 7999 -21594 8009 -21560
rect 8009 -21594 8033 -21560
rect 8071 -21594 8077 -21560
rect 8077 -21594 8105 -21560
rect 8143 -21594 8145 -21560
rect 8145 -21594 8177 -21560
rect 8215 -21594 8247 -21560
rect 8247 -21594 8249 -21560
rect 8287 -21594 8315 -21560
rect 8315 -21594 8321 -21560
rect 8359 -21594 8383 -21560
rect 8383 -21594 8393 -21560
rect 9017 -21594 9027 -21560
rect 9027 -21594 9051 -21560
rect 9089 -21594 9095 -21560
rect 9095 -21594 9123 -21560
rect 9161 -21594 9163 -21560
rect 9163 -21594 9195 -21560
rect 9233 -21594 9265 -21560
rect 9265 -21594 9267 -21560
rect 9305 -21594 9333 -21560
rect 9333 -21594 9339 -21560
rect 9377 -21594 9401 -21560
rect 9401 -21594 9411 -21560
rect 10035 -21594 10045 -21560
rect 10045 -21594 10069 -21560
rect 10107 -21594 10113 -21560
rect 10113 -21594 10141 -21560
rect 10179 -21594 10181 -21560
rect 10181 -21594 10213 -21560
rect 10251 -21594 10283 -21560
rect 10283 -21594 10285 -21560
rect 10323 -21594 10351 -21560
rect 10351 -21594 10357 -21560
rect 10395 -21594 10419 -21560
rect 10419 -21594 10429 -21560
rect 11053 -21594 11063 -21560
rect 11063 -21594 11087 -21560
rect 11125 -21594 11131 -21560
rect 11131 -21594 11159 -21560
rect 11197 -21594 11199 -21560
rect 11199 -21594 11231 -21560
rect 11269 -21594 11301 -21560
rect 11301 -21594 11303 -21560
rect 11341 -21594 11369 -21560
rect 11369 -21594 11375 -21560
rect 11413 -21594 11437 -21560
rect 11437 -21594 11447 -21560
rect 12071 -21594 12081 -21560
rect 12081 -21594 12105 -21560
rect 12143 -21594 12149 -21560
rect 12149 -21594 12177 -21560
rect 12215 -21594 12217 -21560
rect 12217 -21594 12249 -21560
rect 12287 -21594 12319 -21560
rect 12319 -21594 12321 -21560
rect 12359 -21594 12387 -21560
rect 12387 -21594 12393 -21560
rect 12431 -21594 12455 -21560
rect 12455 -21594 12465 -21560
rect 13089 -21594 13099 -21560
rect 13099 -21594 13123 -21560
rect 13161 -21594 13167 -21560
rect 13167 -21594 13195 -21560
rect 13233 -21594 13235 -21560
rect 13235 -21594 13267 -21560
rect 13305 -21594 13337 -21560
rect 13337 -21594 13339 -21560
rect 13377 -21594 13405 -21560
rect 13405 -21594 13411 -21560
rect 13449 -21594 13473 -21560
rect 13473 -21594 13483 -21560
rect 14107 -21594 14117 -21560
rect 14117 -21594 14141 -21560
rect 14179 -21594 14185 -21560
rect 14185 -21594 14213 -21560
rect 14251 -21594 14253 -21560
rect 14253 -21594 14285 -21560
rect 14323 -21594 14355 -21560
rect 14355 -21594 14357 -21560
rect 14395 -21594 14423 -21560
rect 14423 -21594 14429 -21560
rect 14467 -21594 14491 -21560
rect 14491 -21594 14501 -21560
rect 15125 -21594 15135 -21560
rect 15135 -21594 15159 -21560
rect 15197 -21594 15203 -21560
rect 15203 -21594 15231 -21560
rect 15269 -21594 15271 -21560
rect 15271 -21594 15303 -21560
rect 15341 -21594 15373 -21560
rect 15373 -21594 15375 -21560
rect 15413 -21594 15441 -21560
rect 15441 -21594 15447 -21560
rect 15485 -21594 15509 -21560
rect 15509 -21594 15519 -21560
rect 16143 -21594 16153 -21560
rect 16153 -21594 16177 -21560
rect 16215 -21594 16221 -21560
rect 16221 -21594 16249 -21560
rect 16287 -21594 16289 -21560
rect 16289 -21594 16321 -21560
rect 16359 -21594 16391 -21560
rect 16391 -21594 16393 -21560
rect 16431 -21594 16459 -21560
rect 16459 -21594 16465 -21560
rect 16503 -21594 16527 -21560
rect 16527 -21594 16537 -21560
rect 17161 -21594 17171 -21560
rect 17171 -21594 17195 -21560
rect 17233 -21594 17239 -21560
rect 17239 -21594 17267 -21560
rect 17305 -21594 17307 -21560
rect 17307 -21594 17339 -21560
rect 17377 -21594 17409 -21560
rect 17409 -21594 17411 -21560
rect 17449 -21594 17477 -21560
rect 17477 -21594 17483 -21560
rect 17521 -21594 17545 -21560
rect 17545 -21594 17555 -21560
rect 18179 -21594 18189 -21560
rect 18189 -21594 18213 -21560
rect 18251 -21594 18257 -21560
rect 18257 -21594 18285 -21560
rect 18323 -21594 18325 -21560
rect 18325 -21594 18357 -21560
rect 18395 -21594 18427 -21560
rect 18427 -21594 18429 -21560
rect 18467 -21594 18495 -21560
rect 18495 -21594 18501 -21560
rect 18539 -21594 18563 -21560
rect 18563 -21594 18573 -21560
rect 19197 -21594 19207 -21560
rect 19207 -21594 19231 -21560
rect 19269 -21594 19275 -21560
rect 19275 -21594 19303 -21560
rect 19341 -21594 19343 -21560
rect 19343 -21594 19375 -21560
rect 19413 -21594 19445 -21560
rect 19445 -21594 19447 -21560
rect 19485 -21594 19513 -21560
rect 19513 -21594 19519 -21560
rect 19557 -21594 19581 -21560
rect 19581 -21594 19591 -21560
rect 20215 -21594 20225 -21560
rect 20225 -21594 20249 -21560
rect 20287 -21594 20293 -21560
rect 20293 -21594 20321 -21560
rect 20359 -21594 20361 -21560
rect 20361 -21594 20393 -21560
rect 20431 -21594 20463 -21560
rect 20463 -21594 20465 -21560
rect 20503 -21594 20531 -21560
rect 20531 -21594 20537 -21560
rect 20575 -21594 20599 -21560
rect 20599 -21594 20609 -21560
rect 21233 -21594 21243 -21560
rect 21243 -21594 21267 -21560
rect 21305 -21594 21311 -21560
rect 21311 -21594 21339 -21560
rect 21377 -21594 21379 -21560
rect 21379 -21594 21411 -21560
rect 21449 -21594 21481 -21560
rect 21481 -21594 21483 -21560
rect 21521 -21594 21549 -21560
rect 21549 -21594 21555 -21560
rect 21593 -21594 21617 -21560
rect 21617 -21594 21627 -21560
rect 22251 -21594 22261 -21560
rect 22261 -21594 22285 -21560
rect 22323 -21594 22329 -21560
rect 22329 -21594 22357 -21560
rect 22395 -21594 22397 -21560
rect 22397 -21594 22429 -21560
rect 22467 -21594 22499 -21560
rect 22499 -21594 22501 -21560
rect 22539 -21594 22567 -21560
rect 22567 -21594 22573 -21560
rect 22611 -21594 22635 -21560
rect 22635 -21594 22645 -21560
rect -12289 -21699 -12255 -21667
rect -12289 -21701 -12255 -21699
rect -12289 -21767 -12255 -21739
rect -12289 -21773 -12255 -21767
rect -12289 -21835 -12255 -21811
rect -12289 -21845 -12255 -21835
rect -12289 -21903 -12255 -21883
rect -12289 -21917 -12255 -21903
rect -12289 -21971 -12255 -21955
rect -12289 -21989 -12255 -21971
rect -12289 -22039 -12255 -22027
rect -12289 -22061 -12255 -22039
rect -12289 -22107 -12255 -22099
rect -12289 -22133 -12255 -22107
rect -12289 -22175 -12255 -22171
rect -12289 -22205 -12255 -22175
rect 2580 -21677 2614 -21663
rect 2580 -21697 2614 -21677
rect 2580 -21745 2614 -21735
rect 2580 -21769 2614 -21745
rect 2580 -21813 2614 -21807
rect 2580 -21841 2614 -21813
rect 2580 -21881 2614 -21879
rect 2580 -21913 2614 -21881
rect 2580 -21983 2614 -21951
rect 2580 -21985 2614 -21983
rect 2580 -22051 2614 -22023
rect 2580 -22057 2614 -22051
rect 2580 -22119 2614 -22095
rect 2580 -22129 2614 -22119
rect 2580 -22187 2614 -22167
rect 2580 -22201 2614 -22187
rect 3598 -21677 3632 -21663
rect 3598 -21697 3632 -21677
rect 3598 -21745 3632 -21735
rect 3598 -21769 3632 -21745
rect 3598 -21813 3632 -21807
rect 3598 -21841 3632 -21813
rect 3598 -21881 3632 -21879
rect 3598 -21913 3632 -21881
rect 3598 -21983 3632 -21951
rect 3598 -21985 3632 -21983
rect 3598 -22051 3632 -22023
rect 3598 -22057 3632 -22051
rect 3598 -22119 3632 -22095
rect 3598 -22129 3632 -22119
rect 3598 -22187 3632 -22167
rect 3598 -22201 3632 -22187
rect 4616 -21677 4650 -21663
rect 4616 -21697 4650 -21677
rect 4616 -21745 4650 -21735
rect 4616 -21769 4650 -21745
rect 4616 -21813 4650 -21807
rect 4616 -21841 4650 -21813
rect 4616 -21881 4650 -21879
rect 4616 -21913 4650 -21881
rect 4616 -21983 4650 -21951
rect 4616 -21985 4650 -21983
rect 4616 -22051 4650 -22023
rect 4616 -22057 4650 -22051
rect 4616 -22119 4650 -22095
rect 4616 -22129 4650 -22119
rect 4616 -22187 4650 -22167
rect 4616 -22201 4650 -22187
rect 5634 -21677 5668 -21663
rect 5634 -21697 5668 -21677
rect 5634 -21745 5668 -21735
rect 5634 -21769 5668 -21745
rect 5634 -21813 5668 -21807
rect 5634 -21841 5668 -21813
rect 5634 -21881 5668 -21879
rect 5634 -21913 5668 -21881
rect 5634 -21983 5668 -21951
rect 5634 -21985 5668 -21983
rect 5634 -22051 5668 -22023
rect 5634 -22057 5668 -22051
rect 5634 -22119 5668 -22095
rect 5634 -22129 5668 -22119
rect 5634 -22187 5668 -22167
rect 5634 -22201 5668 -22187
rect 6652 -21677 6686 -21663
rect 6652 -21697 6686 -21677
rect 6652 -21745 6686 -21735
rect 6652 -21769 6686 -21745
rect 6652 -21813 6686 -21807
rect 6652 -21841 6686 -21813
rect 6652 -21881 6686 -21879
rect 6652 -21913 6686 -21881
rect 6652 -21983 6686 -21951
rect 6652 -21985 6686 -21983
rect 6652 -22051 6686 -22023
rect 6652 -22057 6686 -22051
rect 6652 -22119 6686 -22095
rect 6652 -22129 6686 -22119
rect 6652 -22187 6686 -22167
rect 6652 -22201 6686 -22187
rect 7670 -21677 7704 -21663
rect 7670 -21697 7704 -21677
rect 7670 -21745 7704 -21735
rect 7670 -21769 7704 -21745
rect 7670 -21813 7704 -21807
rect 7670 -21841 7704 -21813
rect 7670 -21881 7704 -21879
rect 7670 -21913 7704 -21881
rect 7670 -21983 7704 -21951
rect 7670 -21985 7704 -21983
rect 7670 -22051 7704 -22023
rect 7670 -22057 7704 -22051
rect 7670 -22119 7704 -22095
rect 7670 -22129 7704 -22119
rect 7670 -22187 7704 -22167
rect 7670 -22201 7704 -22187
rect 8688 -21677 8722 -21663
rect 8688 -21697 8722 -21677
rect 8688 -21745 8722 -21735
rect 8688 -21769 8722 -21745
rect 8688 -21813 8722 -21807
rect 8688 -21841 8722 -21813
rect 8688 -21881 8722 -21879
rect 8688 -21913 8722 -21881
rect 8688 -21983 8722 -21951
rect 8688 -21985 8722 -21983
rect 8688 -22051 8722 -22023
rect 8688 -22057 8722 -22051
rect 8688 -22119 8722 -22095
rect 8688 -22129 8722 -22119
rect 8688 -22187 8722 -22167
rect 8688 -22201 8722 -22187
rect 9706 -21677 9740 -21663
rect 9706 -21697 9740 -21677
rect 9706 -21745 9740 -21735
rect 9706 -21769 9740 -21745
rect 9706 -21813 9740 -21807
rect 9706 -21841 9740 -21813
rect 9706 -21881 9740 -21879
rect 9706 -21913 9740 -21881
rect 9706 -21983 9740 -21951
rect 9706 -21985 9740 -21983
rect 9706 -22051 9740 -22023
rect 9706 -22057 9740 -22051
rect 9706 -22119 9740 -22095
rect 9706 -22129 9740 -22119
rect 9706 -22187 9740 -22167
rect 9706 -22201 9740 -22187
rect 10724 -21677 10758 -21663
rect 10724 -21697 10758 -21677
rect 10724 -21745 10758 -21735
rect 10724 -21769 10758 -21745
rect 10724 -21813 10758 -21807
rect 10724 -21841 10758 -21813
rect 10724 -21881 10758 -21879
rect 10724 -21913 10758 -21881
rect 10724 -21983 10758 -21951
rect 10724 -21985 10758 -21983
rect 10724 -22051 10758 -22023
rect 10724 -22057 10758 -22051
rect 10724 -22119 10758 -22095
rect 10724 -22129 10758 -22119
rect 10724 -22187 10758 -22167
rect 10724 -22201 10758 -22187
rect 11742 -21677 11776 -21663
rect 11742 -21697 11776 -21677
rect 11742 -21745 11776 -21735
rect 11742 -21769 11776 -21745
rect 11742 -21813 11776 -21807
rect 11742 -21841 11776 -21813
rect 11742 -21881 11776 -21879
rect 11742 -21913 11776 -21881
rect 11742 -21983 11776 -21951
rect 11742 -21985 11776 -21983
rect 11742 -22051 11776 -22023
rect 11742 -22057 11776 -22051
rect 11742 -22119 11776 -22095
rect 11742 -22129 11776 -22119
rect 11742 -22187 11776 -22167
rect 11742 -22201 11776 -22187
rect 12760 -21677 12794 -21663
rect 12760 -21697 12794 -21677
rect 12760 -21745 12794 -21735
rect 12760 -21769 12794 -21745
rect 12760 -21813 12794 -21807
rect 12760 -21841 12794 -21813
rect 12760 -21881 12794 -21879
rect 12760 -21913 12794 -21881
rect 12760 -21983 12794 -21951
rect 12760 -21985 12794 -21983
rect 12760 -22051 12794 -22023
rect 12760 -22057 12794 -22051
rect 12760 -22119 12794 -22095
rect 12760 -22129 12794 -22119
rect 12760 -22187 12794 -22167
rect 12760 -22201 12794 -22187
rect 13778 -21677 13812 -21663
rect 13778 -21697 13812 -21677
rect 13778 -21745 13812 -21735
rect 13778 -21769 13812 -21745
rect 13778 -21813 13812 -21807
rect 13778 -21841 13812 -21813
rect 13778 -21881 13812 -21879
rect 13778 -21913 13812 -21881
rect 13778 -21983 13812 -21951
rect 13778 -21985 13812 -21983
rect 13778 -22051 13812 -22023
rect 13778 -22057 13812 -22051
rect 13778 -22119 13812 -22095
rect 13778 -22129 13812 -22119
rect 13778 -22187 13812 -22167
rect 13778 -22201 13812 -22187
rect 14796 -21677 14830 -21663
rect 14796 -21697 14830 -21677
rect 14796 -21745 14830 -21735
rect 14796 -21769 14830 -21745
rect 14796 -21813 14830 -21807
rect 14796 -21841 14830 -21813
rect 14796 -21881 14830 -21879
rect 14796 -21913 14830 -21881
rect 14796 -21983 14830 -21951
rect 14796 -21985 14830 -21983
rect 14796 -22051 14830 -22023
rect 14796 -22057 14830 -22051
rect 14796 -22119 14830 -22095
rect 14796 -22129 14830 -22119
rect 14796 -22187 14830 -22167
rect 14796 -22201 14830 -22187
rect 15814 -21677 15848 -21663
rect 15814 -21697 15848 -21677
rect 15814 -21745 15848 -21735
rect 15814 -21769 15848 -21745
rect 15814 -21813 15848 -21807
rect 15814 -21841 15848 -21813
rect 15814 -21881 15848 -21879
rect 15814 -21913 15848 -21881
rect 15814 -21983 15848 -21951
rect 15814 -21985 15848 -21983
rect 15814 -22051 15848 -22023
rect 15814 -22057 15848 -22051
rect 15814 -22119 15848 -22095
rect 15814 -22129 15848 -22119
rect 15814 -22187 15848 -22167
rect 15814 -22201 15848 -22187
rect 16832 -21677 16866 -21663
rect 16832 -21697 16866 -21677
rect 16832 -21745 16866 -21735
rect 16832 -21769 16866 -21745
rect 16832 -21813 16866 -21807
rect 16832 -21841 16866 -21813
rect 16832 -21881 16866 -21879
rect 16832 -21913 16866 -21881
rect 16832 -21983 16866 -21951
rect 16832 -21985 16866 -21983
rect 16832 -22051 16866 -22023
rect 16832 -22057 16866 -22051
rect 16832 -22119 16866 -22095
rect 16832 -22129 16866 -22119
rect 16832 -22187 16866 -22167
rect 16832 -22201 16866 -22187
rect 17850 -21677 17884 -21663
rect 17850 -21697 17884 -21677
rect 17850 -21745 17884 -21735
rect 17850 -21769 17884 -21745
rect 17850 -21813 17884 -21807
rect 17850 -21841 17884 -21813
rect 17850 -21881 17884 -21879
rect 17850 -21913 17884 -21881
rect 17850 -21983 17884 -21951
rect 17850 -21985 17884 -21983
rect 17850 -22051 17884 -22023
rect 17850 -22057 17884 -22051
rect 17850 -22119 17884 -22095
rect 17850 -22129 17884 -22119
rect 17850 -22187 17884 -22167
rect 17850 -22201 17884 -22187
rect 18868 -21677 18902 -21663
rect 18868 -21697 18902 -21677
rect 18868 -21745 18902 -21735
rect 18868 -21769 18902 -21745
rect 18868 -21813 18902 -21807
rect 18868 -21841 18902 -21813
rect 18868 -21881 18902 -21879
rect 18868 -21913 18902 -21881
rect 18868 -21983 18902 -21951
rect 18868 -21985 18902 -21983
rect 18868 -22051 18902 -22023
rect 18868 -22057 18902 -22051
rect 18868 -22119 18902 -22095
rect 18868 -22129 18902 -22119
rect 18868 -22187 18902 -22167
rect 18868 -22201 18902 -22187
rect 19886 -21677 19920 -21663
rect 19886 -21697 19920 -21677
rect 19886 -21745 19920 -21735
rect 19886 -21769 19920 -21745
rect 19886 -21813 19920 -21807
rect 19886 -21841 19920 -21813
rect 19886 -21881 19920 -21879
rect 19886 -21913 19920 -21881
rect 19886 -21983 19920 -21951
rect 19886 -21985 19920 -21983
rect 19886 -22051 19920 -22023
rect 19886 -22057 19920 -22051
rect 19886 -22119 19920 -22095
rect 19886 -22129 19920 -22119
rect 19886 -22187 19920 -22167
rect 19886 -22201 19920 -22187
rect 20904 -21677 20938 -21663
rect 20904 -21697 20938 -21677
rect 20904 -21745 20938 -21735
rect 20904 -21769 20938 -21745
rect 20904 -21813 20938 -21807
rect 20904 -21841 20938 -21813
rect 20904 -21881 20938 -21879
rect 20904 -21913 20938 -21881
rect 20904 -21983 20938 -21951
rect 20904 -21985 20938 -21983
rect 20904 -22051 20938 -22023
rect 20904 -22057 20938 -22051
rect 20904 -22119 20938 -22095
rect 20904 -22129 20938 -22119
rect 20904 -22187 20938 -22167
rect 20904 -22201 20938 -22187
rect 21922 -21677 21956 -21663
rect 21922 -21697 21956 -21677
rect 21922 -21745 21956 -21735
rect 21922 -21769 21956 -21745
rect 21922 -21813 21956 -21807
rect 21922 -21841 21956 -21813
rect 21922 -21881 21956 -21879
rect 21922 -21913 21956 -21881
rect 21922 -21983 21956 -21951
rect 21922 -21985 21956 -21983
rect 21922 -22051 21956 -22023
rect 21922 -22057 21956 -22051
rect 21922 -22119 21956 -22095
rect 21922 -22129 21956 -22119
rect 21922 -22187 21956 -22167
rect 21922 -22201 21956 -22187
rect 22940 -21677 22974 -21663
rect 22940 -21697 22974 -21677
rect 22940 -21745 22974 -21735
rect 22940 -21769 22974 -21745
rect 22940 -21813 22974 -21807
rect 22940 -21841 22974 -21813
rect 22940 -21881 22974 -21879
rect 22940 -21913 22974 -21881
rect 22940 -21983 22974 -21951
rect 22940 -21985 22974 -21983
rect 22940 -22051 22974 -22023
rect 22940 -22057 22974 -22051
rect 22940 -22119 22974 -22095
rect 22940 -22129 22974 -22119
rect 22940 -22187 22974 -22167
rect 22940 -22201 22974 -22187
rect 24855 -21597 24889 -21595
rect 24855 -21629 24889 -21597
rect 24855 -21699 24889 -21667
rect 24855 -21701 24889 -21699
rect 24855 -21767 24889 -21739
rect 24855 -21773 24889 -21767
rect 24855 -21835 24889 -21811
rect 24855 -21845 24889 -21835
rect 24855 -21903 24889 -21883
rect 24855 -21917 24889 -21903
rect 24855 -21971 24889 -21955
rect 24855 -21989 24889 -21971
rect 24855 -22039 24889 -22027
rect 24855 -22061 24889 -22039
rect 24855 -22107 24889 -22099
rect 24855 -22133 24889 -22107
rect 24855 -22175 24889 -22171
rect 24855 -22205 24889 -22175
rect -12289 -22277 -12255 -22243
rect 2909 -22304 2919 -22270
rect 2919 -22304 2943 -22270
rect 2981 -22304 2987 -22270
rect 2987 -22304 3015 -22270
rect 3053 -22304 3055 -22270
rect 3055 -22304 3087 -22270
rect 3125 -22304 3157 -22270
rect 3157 -22304 3159 -22270
rect 3197 -22304 3225 -22270
rect 3225 -22304 3231 -22270
rect 3269 -22304 3293 -22270
rect 3293 -22304 3303 -22270
rect 3927 -22304 3937 -22270
rect 3937 -22304 3961 -22270
rect 3999 -22304 4005 -22270
rect 4005 -22304 4033 -22270
rect 4071 -22304 4073 -22270
rect 4073 -22304 4105 -22270
rect 4143 -22304 4175 -22270
rect 4175 -22304 4177 -22270
rect 4215 -22304 4243 -22270
rect 4243 -22304 4249 -22270
rect 4287 -22304 4311 -22270
rect 4311 -22304 4321 -22270
rect 4945 -22304 4955 -22270
rect 4955 -22304 4979 -22270
rect 5017 -22304 5023 -22270
rect 5023 -22304 5051 -22270
rect 5089 -22304 5091 -22270
rect 5091 -22304 5123 -22270
rect 5161 -22304 5193 -22270
rect 5193 -22304 5195 -22270
rect 5233 -22304 5261 -22270
rect 5261 -22304 5267 -22270
rect 5305 -22304 5329 -22270
rect 5329 -22304 5339 -22270
rect 5963 -22304 5973 -22270
rect 5973 -22304 5997 -22270
rect 6035 -22304 6041 -22270
rect 6041 -22304 6069 -22270
rect 6107 -22304 6109 -22270
rect 6109 -22304 6141 -22270
rect 6179 -22304 6211 -22270
rect 6211 -22304 6213 -22270
rect 6251 -22304 6279 -22270
rect 6279 -22304 6285 -22270
rect 6323 -22304 6347 -22270
rect 6347 -22304 6357 -22270
rect 6981 -22304 6991 -22270
rect 6991 -22304 7015 -22270
rect 7053 -22304 7059 -22270
rect 7059 -22304 7087 -22270
rect 7125 -22304 7127 -22270
rect 7127 -22304 7159 -22270
rect 7197 -22304 7229 -22270
rect 7229 -22304 7231 -22270
rect 7269 -22304 7297 -22270
rect 7297 -22304 7303 -22270
rect 7341 -22304 7365 -22270
rect 7365 -22304 7375 -22270
rect 7999 -22304 8009 -22270
rect 8009 -22304 8033 -22270
rect 8071 -22304 8077 -22270
rect 8077 -22304 8105 -22270
rect 8143 -22304 8145 -22270
rect 8145 -22304 8177 -22270
rect 8215 -22304 8247 -22270
rect 8247 -22304 8249 -22270
rect 8287 -22304 8315 -22270
rect 8315 -22304 8321 -22270
rect 8359 -22304 8383 -22270
rect 8383 -22304 8393 -22270
rect 9017 -22304 9027 -22270
rect 9027 -22304 9051 -22270
rect 9089 -22304 9095 -22270
rect 9095 -22304 9123 -22270
rect 9161 -22304 9163 -22270
rect 9163 -22304 9195 -22270
rect 9233 -22304 9265 -22270
rect 9265 -22304 9267 -22270
rect 9305 -22304 9333 -22270
rect 9333 -22304 9339 -22270
rect 9377 -22304 9401 -22270
rect 9401 -22304 9411 -22270
rect 10035 -22304 10045 -22270
rect 10045 -22304 10069 -22270
rect 10107 -22304 10113 -22270
rect 10113 -22304 10141 -22270
rect 10179 -22304 10181 -22270
rect 10181 -22304 10213 -22270
rect 10251 -22304 10283 -22270
rect 10283 -22304 10285 -22270
rect 10323 -22304 10351 -22270
rect 10351 -22304 10357 -22270
rect 10395 -22304 10419 -22270
rect 10419 -22304 10429 -22270
rect 11053 -22304 11063 -22270
rect 11063 -22304 11087 -22270
rect 11125 -22304 11131 -22270
rect 11131 -22304 11159 -22270
rect 11197 -22304 11199 -22270
rect 11199 -22304 11231 -22270
rect 11269 -22304 11301 -22270
rect 11301 -22304 11303 -22270
rect 11341 -22304 11369 -22270
rect 11369 -22304 11375 -22270
rect 11413 -22304 11437 -22270
rect 11437 -22304 11447 -22270
rect 12071 -22304 12081 -22270
rect 12081 -22304 12105 -22270
rect 12143 -22304 12149 -22270
rect 12149 -22304 12177 -22270
rect 12215 -22304 12217 -22270
rect 12217 -22304 12249 -22270
rect 12287 -22304 12319 -22270
rect 12319 -22304 12321 -22270
rect 12359 -22304 12387 -22270
rect 12387 -22304 12393 -22270
rect 12431 -22304 12455 -22270
rect 12455 -22304 12465 -22270
rect 13089 -22304 13099 -22270
rect 13099 -22304 13123 -22270
rect 13161 -22304 13167 -22270
rect 13167 -22304 13195 -22270
rect 13233 -22304 13235 -22270
rect 13235 -22304 13267 -22270
rect 13305 -22304 13337 -22270
rect 13337 -22304 13339 -22270
rect 13377 -22304 13405 -22270
rect 13405 -22304 13411 -22270
rect 13449 -22304 13473 -22270
rect 13473 -22304 13483 -22270
rect 14107 -22304 14117 -22270
rect 14117 -22304 14141 -22270
rect 14179 -22304 14185 -22270
rect 14185 -22304 14213 -22270
rect 14251 -22304 14253 -22270
rect 14253 -22304 14285 -22270
rect 14323 -22304 14355 -22270
rect 14355 -22304 14357 -22270
rect 14395 -22304 14423 -22270
rect 14423 -22304 14429 -22270
rect 14467 -22304 14491 -22270
rect 14491 -22304 14501 -22270
rect 15125 -22304 15135 -22270
rect 15135 -22304 15159 -22270
rect 15197 -22304 15203 -22270
rect 15203 -22304 15231 -22270
rect 15269 -22304 15271 -22270
rect 15271 -22304 15303 -22270
rect 15341 -22304 15373 -22270
rect 15373 -22304 15375 -22270
rect 15413 -22304 15441 -22270
rect 15441 -22304 15447 -22270
rect 15485 -22304 15509 -22270
rect 15509 -22304 15519 -22270
rect 16143 -22304 16153 -22270
rect 16153 -22304 16177 -22270
rect 16215 -22304 16221 -22270
rect 16221 -22304 16249 -22270
rect 16287 -22304 16289 -22270
rect 16289 -22304 16321 -22270
rect 16359 -22304 16391 -22270
rect 16391 -22304 16393 -22270
rect 16431 -22304 16459 -22270
rect 16459 -22304 16465 -22270
rect 16503 -22304 16527 -22270
rect 16527 -22304 16537 -22270
rect 17161 -22304 17171 -22270
rect 17171 -22304 17195 -22270
rect 17233 -22304 17239 -22270
rect 17239 -22304 17267 -22270
rect 17305 -22304 17307 -22270
rect 17307 -22304 17339 -22270
rect 17377 -22304 17409 -22270
rect 17409 -22304 17411 -22270
rect 17449 -22304 17477 -22270
rect 17477 -22304 17483 -22270
rect 17521 -22304 17545 -22270
rect 17545 -22304 17555 -22270
rect 18179 -22304 18189 -22270
rect 18189 -22304 18213 -22270
rect 18251 -22304 18257 -22270
rect 18257 -22304 18285 -22270
rect 18323 -22304 18325 -22270
rect 18325 -22304 18357 -22270
rect 18395 -22304 18427 -22270
rect 18427 -22304 18429 -22270
rect 18467 -22304 18495 -22270
rect 18495 -22304 18501 -22270
rect 18539 -22304 18563 -22270
rect 18563 -22304 18573 -22270
rect 19197 -22304 19207 -22270
rect 19207 -22304 19231 -22270
rect 19269 -22304 19275 -22270
rect 19275 -22304 19303 -22270
rect 19341 -22304 19343 -22270
rect 19343 -22304 19375 -22270
rect 19413 -22304 19445 -22270
rect 19445 -22304 19447 -22270
rect 19485 -22304 19513 -22270
rect 19513 -22304 19519 -22270
rect 19557 -22304 19581 -22270
rect 19581 -22304 19591 -22270
rect 20215 -22304 20225 -22270
rect 20225 -22304 20249 -22270
rect 20287 -22304 20293 -22270
rect 20293 -22304 20321 -22270
rect 20359 -22304 20361 -22270
rect 20361 -22304 20393 -22270
rect 20431 -22304 20463 -22270
rect 20463 -22304 20465 -22270
rect 20503 -22304 20531 -22270
rect 20531 -22304 20537 -22270
rect 20575 -22304 20599 -22270
rect 20599 -22304 20609 -22270
rect 21233 -22304 21243 -22270
rect 21243 -22304 21267 -22270
rect 21305 -22304 21311 -22270
rect 21311 -22304 21339 -22270
rect 21377 -22304 21379 -22270
rect 21379 -22304 21411 -22270
rect 21449 -22304 21481 -22270
rect 21481 -22304 21483 -22270
rect 21521 -22304 21549 -22270
rect 21549 -22304 21555 -22270
rect 21593 -22304 21617 -22270
rect 21617 -22304 21627 -22270
rect 22251 -22304 22261 -22270
rect 22261 -22304 22285 -22270
rect 22323 -22304 22329 -22270
rect 22329 -22304 22357 -22270
rect 22395 -22304 22397 -22270
rect 22397 -22304 22429 -22270
rect 22467 -22304 22499 -22270
rect 22499 -22304 22501 -22270
rect 22539 -22304 22567 -22270
rect 22567 -22304 22573 -22270
rect 22611 -22304 22635 -22270
rect 22635 -22304 22645 -22270
rect 24855 -22277 24889 -22243
rect -12289 -22345 -12255 -22315
rect -12289 -22349 -12255 -22345
rect -12289 -22413 -12255 -22387
rect -12289 -22421 -12255 -22413
rect -12289 -22481 -12255 -22459
rect -12289 -22493 -12255 -22481
rect -12289 -22549 -12255 -22531
rect -12289 -22565 -12255 -22549
rect -12289 -22617 -12255 -22603
rect -12289 -22637 -12255 -22617
rect -12289 -22685 -12255 -22675
rect -12289 -22709 -12255 -22685
rect -12289 -22753 -12255 -22747
rect -12289 -22781 -12255 -22753
rect -12289 -22821 -12255 -22819
rect -12289 -22853 -12255 -22821
rect 24855 -22345 24889 -22315
rect 24855 -22349 24889 -22345
rect 24855 -22413 24889 -22387
rect 24855 -22421 24889 -22413
rect 24855 -22481 24889 -22459
rect 24855 -22493 24889 -22481
rect 24855 -22549 24889 -22531
rect 24855 -22565 24889 -22549
rect 24855 -22617 24889 -22603
rect 24855 -22637 24889 -22617
rect 24855 -22685 24889 -22675
rect 24855 -22709 24889 -22685
rect 24855 -22753 24889 -22747
rect 24855 -22781 24889 -22753
rect 2909 -22826 2919 -22792
rect 2919 -22826 2943 -22792
rect 2981 -22826 2987 -22792
rect 2987 -22826 3015 -22792
rect 3053 -22826 3055 -22792
rect 3055 -22826 3087 -22792
rect 3125 -22826 3157 -22792
rect 3157 -22826 3159 -22792
rect 3197 -22826 3225 -22792
rect 3225 -22826 3231 -22792
rect 3269 -22826 3293 -22792
rect 3293 -22826 3303 -22792
rect 3927 -22826 3937 -22792
rect 3937 -22826 3961 -22792
rect 3999 -22826 4005 -22792
rect 4005 -22826 4033 -22792
rect 4071 -22826 4073 -22792
rect 4073 -22826 4105 -22792
rect 4143 -22826 4175 -22792
rect 4175 -22826 4177 -22792
rect 4215 -22826 4243 -22792
rect 4243 -22826 4249 -22792
rect 4287 -22826 4311 -22792
rect 4311 -22826 4321 -22792
rect 4945 -22826 4955 -22792
rect 4955 -22826 4979 -22792
rect 5017 -22826 5023 -22792
rect 5023 -22826 5051 -22792
rect 5089 -22826 5091 -22792
rect 5091 -22826 5123 -22792
rect 5161 -22826 5193 -22792
rect 5193 -22826 5195 -22792
rect 5233 -22826 5261 -22792
rect 5261 -22826 5267 -22792
rect 5305 -22826 5329 -22792
rect 5329 -22826 5339 -22792
rect 5963 -22826 5973 -22792
rect 5973 -22826 5997 -22792
rect 6035 -22826 6041 -22792
rect 6041 -22826 6069 -22792
rect 6107 -22826 6109 -22792
rect 6109 -22826 6141 -22792
rect 6179 -22826 6211 -22792
rect 6211 -22826 6213 -22792
rect 6251 -22826 6279 -22792
rect 6279 -22826 6285 -22792
rect 6323 -22826 6347 -22792
rect 6347 -22826 6357 -22792
rect 6981 -22826 6991 -22792
rect 6991 -22826 7015 -22792
rect 7053 -22826 7059 -22792
rect 7059 -22826 7087 -22792
rect 7125 -22826 7127 -22792
rect 7127 -22826 7159 -22792
rect 7197 -22826 7229 -22792
rect 7229 -22826 7231 -22792
rect 7269 -22826 7297 -22792
rect 7297 -22826 7303 -22792
rect 7341 -22826 7365 -22792
rect 7365 -22826 7375 -22792
rect 7999 -22826 8009 -22792
rect 8009 -22826 8033 -22792
rect 8071 -22826 8077 -22792
rect 8077 -22826 8105 -22792
rect 8143 -22826 8145 -22792
rect 8145 -22826 8177 -22792
rect 8215 -22826 8247 -22792
rect 8247 -22826 8249 -22792
rect 8287 -22826 8315 -22792
rect 8315 -22826 8321 -22792
rect 8359 -22826 8383 -22792
rect 8383 -22826 8393 -22792
rect 9017 -22826 9027 -22792
rect 9027 -22826 9051 -22792
rect 9089 -22826 9095 -22792
rect 9095 -22826 9123 -22792
rect 9161 -22826 9163 -22792
rect 9163 -22826 9195 -22792
rect 9233 -22826 9265 -22792
rect 9265 -22826 9267 -22792
rect 9305 -22826 9333 -22792
rect 9333 -22826 9339 -22792
rect 9377 -22826 9401 -22792
rect 9401 -22826 9411 -22792
rect 10035 -22826 10045 -22792
rect 10045 -22826 10069 -22792
rect 10107 -22826 10113 -22792
rect 10113 -22826 10141 -22792
rect 10179 -22826 10181 -22792
rect 10181 -22826 10213 -22792
rect 10251 -22826 10283 -22792
rect 10283 -22826 10285 -22792
rect 10323 -22826 10351 -22792
rect 10351 -22826 10357 -22792
rect 10395 -22826 10419 -22792
rect 10419 -22826 10429 -22792
rect 11053 -22826 11063 -22792
rect 11063 -22826 11087 -22792
rect 11125 -22826 11131 -22792
rect 11131 -22826 11159 -22792
rect 11197 -22826 11199 -22792
rect 11199 -22826 11231 -22792
rect 11269 -22826 11301 -22792
rect 11301 -22826 11303 -22792
rect 11341 -22826 11369 -22792
rect 11369 -22826 11375 -22792
rect 11413 -22826 11437 -22792
rect 11437 -22826 11447 -22792
rect 12071 -22826 12081 -22792
rect 12081 -22826 12105 -22792
rect 12143 -22826 12149 -22792
rect 12149 -22826 12177 -22792
rect 12215 -22826 12217 -22792
rect 12217 -22826 12249 -22792
rect 12287 -22826 12319 -22792
rect 12319 -22826 12321 -22792
rect 12359 -22826 12387 -22792
rect 12387 -22826 12393 -22792
rect 12431 -22826 12455 -22792
rect 12455 -22826 12465 -22792
rect 13089 -22826 13099 -22792
rect 13099 -22826 13123 -22792
rect 13161 -22826 13167 -22792
rect 13167 -22826 13195 -22792
rect 13233 -22826 13235 -22792
rect 13235 -22826 13267 -22792
rect 13305 -22826 13337 -22792
rect 13337 -22826 13339 -22792
rect 13377 -22826 13405 -22792
rect 13405 -22826 13411 -22792
rect 13449 -22826 13473 -22792
rect 13473 -22826 13483 -22792
rect 14107 -22826 14117 -22792
rect 14117 -22826 14141 -22792
rect 14179 -22826 14185 -22792
rect 14185 -22826 14213 -22792
rect 14251 -22826 14253 -22792
rect 14253 -22826 14285 -22792
rect 14323 -22826 14355 -22792
rect 14355 -22826 14357 -22792
rect 14395 -22826 14423 -22792
rect 14423 -22826 14429 -22792
rect 14467 -22826 14491 -22792
rect 14491 -22826 14501 -22792
rect 15125 -22826 15135 -22792
rect 15135 -22826 15159 -22792
rect 15197 -22826 15203 -22792
rect 15203 -22826 15231 -22792
rect 15269 -22826 15271 -22792
rect 15271 -22826 15303 -22792
rect 15341 -22826 15373 -22792
rect 15373 -22826 15375 -22792
rect 15413 -22826 15441 -22792
rect 15441 -22826 15447 -22792
rect 15485 -22826 15509 -22792
rect 15509 -22826 15519 -22792
rect 16143 -22826 16153 -22792
rect 16153 -22826 16177 -22792
rect 16215 -22826 16221 -22792
rect 16221 -22826 16249 -22792
rect 16287 -22826 16289 -22792
rect 16289 -22826 16321 -22792
rect 16359 -22826 16391 -22792
rect 16391 -22826 16393 -22792
rect 16431 -22826 16459 -22792
rect 16459 -22826 16465 -22792
rect 16503 -22826 16527 -22792
rect 16527 -22826 16537 -22792
rect 17161 -22826 17171 -22792
rect 17171 -22826 17195 -22792
rect 17233 -22826 17239 -22792
rect 17239 -22826 17267 -22792
rect 17305 -22826 17307 -22792
rect 17307 -22826 17339 -22792
rect 17377 -22826 17409 -22792
rect 17409 -22826 17411 -22792
rect 17449 -22826 17477 -22792
rect 17477 -22826 17483 -22792
rect 17521 -22826 17545 -22792
rect 17545 -22826 17555 -22792
rect 18179 -22826 18189 -22792
rect 18189 -22826 18213 -22792
rect 18251 -22826 18257 -22792
rect 18257 -22826 18285 -22792
rect 18323 -22826 18325 -22792
rect 18325 -22826 18357 -22792
rect 18395 -22826 18427 -22792
rect 18427 -22826 18429 -22792
rect 18467 -22826 18495 -22792
rect 18495 -22826 18501 -22792
rect 18539 -22826 18563 -22792
rect 18563 -22826 18573 -22792
rect 19197 -22826 19207 -22792
rect 19207 -22826 19231 -22792
rect 19269 -22826 19275 -22792
rect 19275 -22826 19303 -22792
rect 19341 -22826 19343 -22792
rect 19343 -22826 19375 -22792
rect 19413 -22826 19445 -22792
rect 19445 -22826 19447 -22792
rect 19485 -22826 19513 -22792
rect 19513 -22826 19519 -22792
rect 19557 -22826 19581 -22792
rect 19581 -22826 19591 -22792
rect 20215 -22826 20225 -22792
rect 20225 -22826 20249 -22792
rect 20287 -22826 20293 -22792
rect 20293 -22826 20321 -22792
rect 20359 -22826 20361 -22792
rect 20361 -22826 20393 -22792
rect 20431 -22826 20463 -22792
rect 20463 -22826 20465 -22792
rect 20503 -22826 20531 -22792
rect 20531 -22826 20537 -22792
rect 20575 -22826 20599 -22792
rect 20599 -22826 20609 -22792
rect 21233 -22826 21243 -22792
rect 21243 -22826 21267 -22792
rect 21305 -22826 21311 -22792
rect 21311 -22826 21339 -22792
rect 21377 -22826 21379 -22792
rect 21379 -22826 21411 -22792
rect 21449 -22826 21481 -22792
rect 21481 -22826 21483 -22792
rect 21521 -22826 21549 -22792
rect 21549 -22826 21555 -22792
rect 21593 -22826 21617 -22792
rect 21617 -22826 21627 -22792
rect 22251 -22826 22261 -22792
rect 22261 -22826 22285 -22792
rect 22323 -22826 22329 -22792
rect 22329 -22826 22357 -22792
rect 22395 -22826 22397 -22792
rect 22397 -22826 22429 -22792
rect 22467 -22826 22499 -22792
rect 22499 -22826 22501 -22792
rect 22539 -22826 22567 -22792
rect 22567 -22826 22573 -22792
rect 22611 -22826 22635 -22792
rect 22635 -22826 22645 -22792
rect 24855 -22821 24889 -22819
rect 24855 -22853 24889 -22821
rect -12289 -22923 -12255 -22891
rect -12289 -22925 -12255 -22923
rect -12289 -22991 -12255 -22963
rect -12289 -22997 -12255 -22991
rect -12289 -23059 -12255 -23035
rect -12289 -23069 -12255 -23059
rect -12289 -23127 -12255 -23107
rect -12289 -23141 -12255 -23127
rect -12289 -23195 -12255 -23179
rect -12289 -23213 -12255 -23195
rect -12289 -23263 -12255 -23251
rect -12289 -23285 -12255 -23263
rect -12289 -23331 -12255 -23323
rect -12289 -23357 -12255 -23331
rect -12289 -23399 -12255 -23395
rect -12289 -23429 -12255 -23399
rect -12289 -23501 -12255 -23467
rect 2580 -22909 2614 -22895
rect 2580 -22929 2614 -22909
rect 2580 -22977 2614 -22967
rect 2580 -23001 2614 -22977
rect 2580 -23045 2614 -23039
rect 2580 -23073 2614 -23045
rect 2580 -23113 2614 -23111
rect 2580 -23145 2614 -23113
rect 2580 -23215 2614 -23183
rect 2580 -23217 2614 -23215
rect 2580 -23283 2614 -23255
rect 2580 -23289 2614 -23283
rect 2580 -23351 2614 -23327
rect 2580 -23361 2614 -23351
rect 2580 -23419 2614 -23399
rect 2580 -23433 2614 -23419
rect 3598 -22909 3632 -22895
rect 3598 -22929 3632 -22909
rect 3598 -22977 3632 -22967
rect 3598 -23001 3632 -22977
rect 3598 -23045 3632 -23039
rect 3598 -23073 3632 -23045
rect 3598 -23113 3632 -23111
rect 3598 -23145 3632 -23113
rect 3598 -23215 3632 -23183
rect 3598 -23217 3632 -23215
rect 3598 -23283 3632 -23255
rect 3598 -23289 3632 -23283
rect 3598 -23351 3632 -23327
rect 3598 -23361 3632 -23351
rect 3598 -23419 3632 -23399
rect 3598 -23433 3632 -23419
rect 4616 -22909 4650 -22895
rect 4616 -22929 4650 -22909
rect 4616 -22977 4650 -22967
rect 4616 -23001 4650 -22977
rect 4616 -23045 4650 -23039
rect 4616 -23073 4650 -23045
rect 4616 -23113 4650 -23111
rect 4616 -23145 4650 -23113
rect 4616 -23215 4650 -23183
rect 4616 -23217 4650 -23215
rect 4616 -23283 4650 -23255
rect 4616 -23289 4650 -23283
rect 4616 -23351 4650 -23327
rect 4616 -23361 4650 -23351
rect 4616 -23419 4650 -23399
rect 4616 -23433 4650 -23419
rect 5634 -22909 5668 -22895
rect 5634 -22929 5668 -22909
rect 5634 -22977 5668 -22967
rect 5634 -23001 5668 -22977
rect 5634 -23045 5668 -23039
rect 5634 -23073 5668 -23045
rect 5634 -23113 5668 -23111
rect 5634 -23145 5668 -23113
rect 5634 -23215 5668 -23183
rect 5634 -23217 5668 -23215
rect 5634 -23283 5668 -23255
rect 5634 -23289 5668 -23283
rect 5634 -23351 5668 -23327
rect 5634 -23361 5668 -23351
rect 5634 -23419 5668 -23399
rect 5634 -23433 5668 -23419
rect 6652 -22909 6686 -22895
rect 6652 -22929 6686 -22909
rect 6652 -22977 6686 -22967
rect 6652 -23001 6686 -22977
rect 6652 -23045 6686 -23039
rect 6652 -23073 6686 -23045
rect 6652 -23113 6686 -23111
rect 6652 -23145 6686 -23113
rect 6652 -23215 6686 -23183
rect 6652 -23217 6686 -23215
rect 6652 -23283 6686 -23255
rect 6652 -23289 6686 -23283
rect 6652 -23351 6686 -23327
rect 6652 -23361 6686 -23351
rect 6652 -23419 6686 -23399
rect 6652 -23433 6686 -23419
rect 7670 -22909 7704 -22895
rect 7670 -22929 7704 -22909
rect 7670 -22977 7704 -22967
rect 7670 -23001 7704 -22977
rect 7670 -23045 7704 -23039
rect 7670 -23073 7704 -23045
rect 7670 -23113 7704 -23111
rect 7670 -23145 7704 -23113
rect 7670 -23215 7704 -23183
rect 7670 -23217 7704 -23215
rect 7670 -23283 7704 -23255
rect 7670 -23289 7704 -23283
rect 7670 -23351 7704 -23327
rect 7670 -23361 7704 -23351
rect 7670 -23419 7704 -23399
rect 7670 -23433 7704 -23419
rect 8688 -22909 8722 -22895
rect 8688 -22929 8722 -22909
rect 8688 -22977 8722 -22967
rect 8688 -23001 8722 -22977
rect 8688 -23045 8722 -23039
rect 8688 -23073 8722 -23045
rect 8688 -23113 8722 -23111
rect 8688 -23145 8722 -23113
rect 8688 -23215 8722 -23183
rect 8688 -23217 8722 -23215
rect 8688 -23283 8722 -23255
rect 8688 -23289 8722 -23283
rect 8688 -23351 8722 -23327
rect 8688 -23361 8722 -23351
rect 8688 -23419 8722 -23399
rect 8688 -23433 8722 -23419
rect 9706 -22909 9740 -22895
rect 9706 -22929 9740 -22909
rect 9706 -22977 9740 -22967
rect 9706 -23001 9740 -22977
rect 9706 -23045 9740 -23039
rect 9706 -23073 9740 -23045
rect 9706 -23113 9740 -23111
rect 9706 -23145 9740 -23113
rect 9706 -23215 9740 -23183
rect 9706 -23217 9740 -23215
rect 9706 -23283 9740 -23255
rect 9706 -23289 9740 -23283
rect 9706 -23351 9740 -23327
rect 9706 -23361 9740 -23351
rect 9706 -23419 9740 -23399
rect 9706 -23433 9740 -23419
rect 10724 -22909 10758 -22895
rect 10724 -22929 10758 -22909
rect 10724 -22977 10758 -22967
rect 10724 -23001 10758 -22977
rect 10724 -23045 10758 -23039
rect 10724 -23073 10758 -23045
rect 10724 -23113 10758 -23111
rect 10724 -23145 10758 -23113
rect 10724 -23215 10758 -23183
rect 10724 -23217 10758 -23215
rect 10724 -23283 10758 -23255
rect 10724 -23289 10758 -23283
rect 10724 -23351 10758 -23327
rect 10724 -23361 10758 -23351
rect 10724 -23419 10758 -23399
rect 10724 -23433 10758 -23419
rect 11742 -22909 11776 -22895
rect 11742 -22929 11776 -22909
rect 11742 -22977 11776 -22967
rect 11742 -23001 11776 -22977
rect 11742 -23045 11776 -23039
rect 11742 -23073 11776 -23045
rect 11742 -23113 11776 -23111
rect 11742 -23145 11776 -23113
rect 11742 -23215 11776 -23183
rect 11742 -23217 11776 -23215
rect 11742 -23283 11776 -23255
rect 11742 -23289 11776 -23283
rect 11742 -23351 11776 -23327
rect 11742 -23361 11776 -23351
rect 11742 -23419 11776 -23399
rect 11742 -23433 11776 -23419
rect 12760 -22909 12794 -22895
rect 12760 -22929 12794 -22909
rect 12760 -22977 12794 -22967
rect 12760 -23001 12794 -22977
rect 12760 -23045 12794 -23039
rect 12760 -23073 12794 -23045
rect 12760 -23113 12794 -23111
rect 12760 -23145 12794 -23113
rect 12760 -23215 12794 -23183
rect 12760 -23217 12794 -23215
rect 12760 -23283 12794 -23255
rect 12760 -23289 12794 -23283
rect 12760 -23351 12794 -23327
rect 12760 -23361 12794 -23351
rect 12760 -23419 12794 -23399
rect 12760 -23433 12794 -23419
rect 13778 -22909 13812 -22895
rect 13778 -22929 13812 -22909
rect 13778 -22977 13812 -22967
rect 13778 -23001 13812 -22977
rect 13778 -23045 13812 -23039
rect 13778 -23073 13812 -23045
rect 13778 -23113 13812 -23111
rect 13778 -23145 13812 -23113
rect 13778 -23215 13812 -23183
rect 13778 -23217 13812 -23215
rect 13778 -23283 13812 -23255
rect 13778 -23289 13812 -23283
rect 13778 -23351 13812 -23327
rect 13778 -23361 13812 -23351
rect 13778 -23419 13812 -23399
rect 13778 -23433 13812 -23419
rect 14796 -22909 14830 -22895
rect 14796 -22929 14830 -22909
rect 14796 -22977 14830 -22967
rect 14796 -23001 14830 -22977
rect 14796 -23045 14830 -23039
rect 14796 -23073 14830 -23045
rect 14796 -23113 14830 -23111
rect 14796 -23145 14830 -23113
rect 14796 -23215 14830 -23183
rect 14796 -23217 14830 -23215
rect 14796 -23283 14830 -23255
rect 14796 -23289 14830 -23283
rect 14796 -23351 14830 -23327
rect 14796 -23361 14830 -23351
rect 14796 -23419 14830 -23399
rect 14796 -23433 14830 -23419
rect 15814 -22909 15848 -22895
rect 15814 -22929 15848 -22909
rect 15814 -22977 15848 -22967
rect 15814 -23001 15848 -22977
rect 15814 -23045 15848 -23039
rect 15814 -23073 15848 -23045
rect 15814 -23113 15848 -23111
rect 15814 -23145 15848 -23113
rect 15814 -23215 15848 -23183
rect 15814 -23217 15848 -23215
rect 15814 -23283 15848 -23255
rect 15814 -23289 15848 -23283
rect 15814 -23351 15848 -23327
rect 15814 -23361 15848 -23351
rect 15814 -23419 15848 -23399
rect 15814 -23433 15848 -23419
rect 16832 -22909 16866 -22895
rect 16832 -22929 16866 -22909
rect 16832 -22977 16866 -22967
rect 16832 -23001 16866 -22977
rect 16832 -23045 16866 -23039
rect 16832 -23073 16866 -23045
rect 16832 -23113 16866 -23111
rect 16832 -23145 16866 -23113
rect 16832 -23215 16866 -23183
rect 16832 -23217 16866 -23215
rect 16832 -23283 16866 -23255
rect 16832 -23289 16866 -23283
rect 16832 -23351 16866 -23327
rect 16832 -23361 16866 -23351
rect 16832 -23419 16866 -23399
rect 16832 -23433 16866 -23419
rect 17850 -22909 17884 -22895
rect 17850 -22929 17884 -22909
rect 17850 -22977 17884 -22967
rect 17850 -23001 17884 -22977
rect 17850 -23045 17884 -23039
rect 17850 -23073 17884 -23045
rect 17850 -23113 17884 -23111
rect 17850 -23145 17884 -23113
rect 17850 -23215 17884 -23183
rect 17850 -23217 17884 -23215
rect 17850 -23283 17884 -23255
rect 17850 -23289 17884 -23283
rect 17850 -23351 17884 -23327
rect 17850 -23361 17884 -23351
rect 17850 -23419 17884 -23399
rect 17850 -23433 17884 -23419
rect 18868 -22909 18902 -22895
rect 18868 -22929 18902 -22909
rect 18868 -22977 18902 -22967
rect 18868 -23001 18902 -22977
rect 18868 -23045 18902 -23039
rect 18868 -23073 18902 -23045
rect 18868 -23113 18902 -23111
rect 18868 -23145 18902 -23113
rect 18868 -23215 18902 -23183
rect 18868 -23217 18902 -23215
rect 18868 -23283 18902 -23255
rect 18868 -23289 18902 -23283
rect 18868 -23351 18902 -23327
rect 18868 -23361 18902 -23351
rect 18868 -23419 18902 -23399
rect 18868 -23433 18902 -23419
rect 19886 -22909 19920 -22895
rect 19886 -22929 19920 -22909
rect 19886 -22977 19920 -22967
rect 19886 -23001 19920 -22977
rect 19886 -23045 19920 -23039
rect 19886 -23073 19920 -23045
rect 19886 -23113 19920 -23111
rect 19886 -23145 19920 -23113
rect 19886 -23215 19920 -23183
rect 19886 -23217 19920 -23215
rect 19886 -23283 19920 -23255
rect 19886 -23289 19920 -23283
rect 19886 -23351 19920 -23327
rect 19886 -23361 19920 -23351
rect 19886 -23419 19920 -23399
rect 19886 -23433 19920 -23419
rect 20904 -22909 20938 -22895
rect 20904 -22929 20938 -22909
rect 20904 -22977 20938 -22967
rect 20904 -23001 20938 -22977
rect 20904 -23045 20938 -23039
rect 20904 -23073 20938 -23045
rect 20904 -23113 20938 -23111
rect 20904 -23145 20938 -23113
rect 20904 -23215 20938 -23183
rect 20904 -23217 20938 -23215
rect 20904 -23283 20938 -23255
rect 20904 -23289 20938 -23283
rect 20904 -23351 20938 -23327
rect 20904 -23361 20938 -23351
rect 20904 -23419 20938 -23399
rect 20904 -23433 20938 -23419
rect 21922 -22909 21956 -22895
rect 21922 -22929 21956 -22909
rect 21922 -22977 21956 -22967
rect 21922 -23001 21956 -22977
rect 21922 -23045 21956 -23039
rect 21922 -23073 21956 -23045
rect 21922 -23113 21956 -23111
rect 21922 -23145 21956 -23113
rect 21922 -23215 21956 -23183
rect 21922 -23217 21956 -23215
rect 21922 -23283 21956 -23255
rect 21922 -23289 21956 -23283
rect 21922 -23351 21956 -23327
rect 21922 -23361 21956 -23351
rect 21922 -23419 21956 -23399
rect 21922 -23433 21956 -23419
rect 22940 -22909 22974 -22895
rect 22940 -22929 22974 -22909
rect 22940 -22977 22974 -22967
rect 22940 -23001 22974 -22977
rect 22940 -23045 22974 -23039
rect 22940 -23073 22974 -23045
rect 22940 -23113 22974 -23111
rect 22940 -23145 22974 -23113
rect 22940 -23215 22974 -23183
rect 22940 -23217 22974 -23215
rect 22940 -23283 22974 -23255
rect 22940 -23289 22974 -23283
rect 22940 -23351 22974 -23327
rect 22940 -23361 22974 -23351
rect 22940 -23419 22974 -23399
rect 22940 -23433 22974 -23419
rect 24855 -22923 24889 -22891
rect 24855 -22925 24889 -22923
rect 24855 -22991 24889 -22963
rect 24855 -22997 24889 -22991
rect 24855 -23059 24889 -23035
rect 24855 -23069 24889 -23059
rect 24855 -23127 24889 -23107
rect 24855 -23141 24889 -23127
rect 24855 -23195 24889 -23179
rect 24855 -23213 24889 -23195
rect 24855 -23263 24889 -23251
rect 24855 -23285 24889 -23263
rect 24855 -23331 24889 -23323
rect 24855 -23357 24889 -23331
rect 24855 -23399 24889 -23395
rect 24855 -23429 24889 -23399
rect 24855 -23501 24889 -23467
rect -12289 -23569 -12255 -23539
rect -12289 -23573 -12255 -23569
rect 2909 -23536 2919 -23502
rect 2919 -23536 2943 -23502
rect 2981 -23536 2987 -23502
rect 2987 -23536 3015 -23502
rect 3053 -23536 3055 -23502
rect 3055 -23536 3087 -23502
rect 3125 -23536 3157 -23502
rect 3157 -23536 3159 -23502
rect 3197 -23536 3225 -23502
rect 3225 -23536 3231 -23502
rect 3269 -23536 3293 -23502
rect 3293 -23536 3303 -23502
rect 3927 -23536 3937 -23502
rect 3937 -23536 3961 -23502
rect 3999 -23536 4005 -23502
rect 4005 -23536 4033 -23502
rect 4071 -23536 4073 -23502
rect 4073 -23536 4105 -23502
rect 4143 -23536 4175 -23502
rect 4175 -23536 4177 -23502
rect 4215 -23536 4243 -23502
rect 4243 -23536 4249 -23502
rect 4287 -23536 4311 -23502
rect 4311 -23536 4321 -23502
rect 4945 -23536 4955 -23502
rect 4955 -23536 4979 -23502
rect 5017 -23536 5023 -23502
rect 5023 -23536 5051 -23502
rect 5089 -23536 5091 -23502
rect 5091 -23536 5123 -23502
rect 5161 -23536 5193 -23502
rect 5193 -23536 5195 -23502
rect 5233 -23536 5261 -23502
rect 5261 -23536 5267 -23502
rect 5305 -23536 5329 -23502
rect 5329 -23536 5339 -23502
rect 5963 -23536 5973 -23502
rect 5973 -23536 5997 -23502
rect 6035 -23536 6041 -23502
rect 6041 -23536 6069 -23502
rect 6107 -23536 6109 -23502
rect 6109 -23536 6141 -23502
rect 6179 -23536 6211 -23502
rect 6211 -23536 6213 -23502
rect 6251 -23536 6279 -23502
rect 6279 -23536 6285 -23502
rect 6323 -23536 6347 -23502
rect 6347 -23536 6357 -23502
rect 6981 -23536 6991 -23502
rect 6991 -23536 7015 -23502
rect 7053 -23536 7059 -23502
rect 7059 -23536 7087 -23502
rect 7125 -23536 7127 -23502
rect 7127 -23536 7159 -23502
rect 7197 -23536 7229 -23502
rect 7229 -23536 7231 -23502
rect 7269 -23536 7297 -23502
rect 7297 -23536 7303 -23502
rect 7341 -23536 7365 -23502
rect 7365 -23536 7375 -23502
rect 7999 -23536 8009 -23502
rect 8009 -23536 8033 -23502
rect 8071 -23536 8077 -23502
rect 8077 -23536 8105 -23502
rect 8143 -23536 8145 -23502
rect 8145 -23536 8177 -23502
rect 8215 -23536 8247 -23502
rect 8247 -23536 8249 -23502
rect 8287 -23536 8315 -23502
rect 8315 -23536 8321 -23502
rect 8359 -23536 8383 -23502
rect 8383 -23536 8393 -23502
rect 9017 -23536 9027 -23502
rect 9027 -23536 9051 -23502
rect 9089 -23536 9095 -23502
rect 9095 -23536 9123 -23502
rect 9161 -23536 9163 -23502
rect 9163 -23536 9195 -23502
rect 9233 -23536 9265 -23502
rect 9265 -23536 9267 -23502
rect 9305 -23536 9333 -23502
rect 9333 -23536 9339 -23502
rect 9377 -23536 9401 -23502
rect 9401 -23536 9411 -23502
rect 10035 -23536 10045 -23502
rect 10045 -23536 10069 -23502
rect 10107 -23536 10113 -23502
rect 10113 -23536 10141 -23502
rect 10179 -23536 10181 -23502
rect 10181 -23536 10213 -23502
rect 10251 -23536 10283 -23502
rect 10283 -23536 10285 -23502
rect 10323 -23536 10351 -23502
rect 10351 -23536 10357 -23502
rect 10395 -23536 10419 -23502
rect 10419 -23536 10429 -23502
rect 11053 -23536 11063 -23502
rect 11063 -23536 11087 -23502
rect 11125 -23536 11131 -23502
rect 11131 -23536 11159 -23502
rect 11197 -23536 11199 -23502
rect 11199 -23536 11231 -23502
rect 11269 -23536 11301 -23502
rect 11301 -23536 11303 -23502
rect 11341 -23536 11369 -23502
rect 11369 -23536 11375 -23502
rect 11413 -23536 11437 -23502
rect 11437 -23536 11447 -23502
rect 12071 -23536 12081 -23502
rect 12081 -23536 12105 -23502
rect 12143 -23536 12149 -23502
rect 12149 -23536 12177 -23502
rect 12215 -23536 12217 -23502
rect 12217 -23536 12249 -23502
rect 12287 -23536 12319 -23502
rect 12319 -23536 12321 -23502
rect 12359 -23536 12387 -23502
rect 12387 -23536 12393 -23502
rect 12431 -23536 12455 -23502
rect 12455 -23536 12465 -23502
rect 13089 -23536 13099 -23502
rect 13099 -23536 13123 -23502
rect 13161 -23536 13167 -23502
rect 13167 -23536 13195 -23502
rect 13233 -23536 13235 -23502
rect 13235 -23536 13267 -23502
rect 13305 -23536 13337 -23502
rect 13337 -23536 13339 -23502
rect 13377 -23536 13405 -23502
rect 13405 -23536 13411 -23502
rect 13449 -23536 13473 -23502
rect 13473 -23536 13483 -23502
rect 14107 -23536 14117 -23502
rect 14117 -23536 14141 -23502
rect 14179 -23536 14185 -23502
rect 14185 -23536 14213 -23502
rect 14251 -23536 14253 -23502
rect 14253 -23536 14285 -23502
rect 14323 -23536 14355 -23502
rect 14355 -23536 14357 -23502
rect 14395 -23536 14423 -23502
rect 14423 -23536 14429 -23502
rect 14467 -23536 14491 -23502
rect 14491 -23536 14501 -23502
rect 15125 -23536 15135 -23502
rect 15135 -23536 15159 -23502
rect 15197 -23536 15203 -23502
rect 15203 -23536 15231 -23502
rect 15269 -23536 15271 -23502
rect 15271 -23536 15303 -23502
rect 15341 -23536 15373 -23502
rect 15373 -23536 15375 -23502
rect 15413 -23536 15441 -23502
rect 15441 -23536 15447 -23502
rect 15485 -23536 15509 -23502
rect 15509 -23536 15519 -23502
rect 16143 -23536 16153 -23502
rect 16153 -23536 16177 -23502
rect 16215 -23536 16221 -23502
rect 16221 -23536 16249 -23502
rect 16287 -23536 16289 -23502
rect 16289 -23536 16321 -23502
rect 16359 -23536 16391 -23502
rect 16391 -23536 16393 -23502
rect 16431 -23536 16459 -23502
rect 16459 -23536 16465 -23502
rect 16503 -23536 16527 -23502
rect 16527 -23536 16537 -23502
rect 17161 -23536 17171 -23502
rect 17171 -23536 17195 -23502
rect 17233 -23536 17239 -23502
rect 17239 -23536 17267 -23502
rect 17305 -23536 17307 -23502
rect 17307 -23536 17339 -23502
rect 17377 -23536 17409 -23502
rect 17409 -23536 17411 -23502
rect 17449 -23536 17477 -23502
rect 17477 -23536 17483 -23502
rect 17521 -23536 17545 -23502
rect 17545 -23536 17555 -23502
rect 18179 -23536 18189 -23502
rect 18189 -23536 18213 -23502
rect 18251 -23536 18257 -23502
rect 18257 -23536 18285 -23502
rect 18323 -23536 18325 -23502
rect 18325 -23536 18357 -23502
rect 18395 -23536 18427 -23502
rect 18427 -23536 18429 -23502
rect 18467 -23536 18495 -23502
rect 18495 -23536 18501 -23502
rect 18539 -23536 18563 -23502
rect 18563 -23536 18573 -23502
rect 19197 -23536 19207 -23502
rect 19207 -23536 19231 -23502
rect 19269 -23536 19275 -23502
rect 19275 -23536 19303 -23502
rect 19341 -23536 19343 -23502
rect 19343 -23536 19375 -23502
rect 19413 -23536 19445 -23502
rect 19445 -23536 19447 -23502
rect 19485 -23536 19513 -23502
rect 19513 -23536 19519 -23502
rect 19557 -23536 19581 -23502
rect 19581 -23536 19591 -23502
rect 20215 -23536 20225 -23502
rect 20225 -23536 20249 -23502
rect 20287 -23536 20293 -23502
rect 20293 -23536 20321 -23502
rect 20359 -23536 20361 -23502
rect 20361 -23536 20393 -23502
rect 20431 -23536 20463 -23502
rect 20463 -23536 20465 -23502
rect 20503 -23536 20531 -23502
rect 20531 -23536 20537 -23502
rect 20575 -23536 20599 -23502
rect 20599 -23536 20609 -23502
rect 21233 -23536 21243 -23502
rect 21243 -23536 21267 -23502
rect 21305 -23536 21311 -23502
rect 21311 -23536 21339 -23502
rect 21377 -23536 21379 -23502
rect 21379 -23536 21411 -23502
rect 21449 -23536 21481 -23502
rect 21481 -23536 21483 -23502
rect 21521 -23536 21549 -23502
rect 21549 -23536 21555 -23502
rect 21593 -23536 21617 -23502
rect 21617 -23536 21627 -23502
rect 22251 -23536 22261 -23502
rect 22261 -23536 22285 -23502
rect 22323 -23536 22329 -23502
rect 22329 -23536 22357 -23502
rect 22395 -23536 22397 -23502
rect 22397 -23536 22429 -23502
rect 22467 -23536 22499 -23502
rect 22499 -23536 22501 -23502
rect 22539 -23536 22567 -23502
rect 22567 -23536 22573 -23502
rect 22611 -23536 22635 -23502
rect 22635 -23536 22645 -23502
rect -12289 -23637 -12255 -23611
rect -12289 -23645 -12255 -23637
rect -12289 -23705 -12255 -23683
rect -12289 -23717 -12255 -23705
rect -12289 -23773 -12255 -23755
rect -12289 -23789 -12255 -23773
rect -12289 -23841 -12255 -23827
rect -12289 -23861 -12255 -23841
rect -12289 -23909 -12255 -23899
rect -12289 -23933 -12255 -23909
rect -12289 -23977 -12255 -23971
rect -12289 -24005 -12255 -23977
rect -12289 -24045 -12255 -24043
rect -12289 -24077 -12255 -24045
rect 24855 -23569 24889 -23539
rect 24855 -23573 24889 -23569
rect 24855 -23637 24889 -23611
rect 24855 -23645 24889 -23637
rect 24855 -23705 24889 -23683
rect 24855 -23717 24889 -23705
rect 24855 -23773 24889 -23755
rect 24855 -23789 24889 -23773
rect 24855 -23841 24889 -23827
rect 24855 -23861 24889 -23841
rect 24855 -23909 24889 -23899
rect 24855 -23933 24889 -23909
rect 24855 -23977 24889 -23971
rect 24855 -24005 24889 -23977
rect 2909 -24060 2919 -24026
rect 2919 -24060 2943 -24026
rect 2981 -24060 2987 -24026
rect 2987 -24060 3015 -24026
rect 3053 -24060 3055 -24026
rect 3055 -24060 3087 -24026
rect 3125 -24060 3157 -24026
rect 3157 -24060 3159 -24026
rect 3197 -24060 3225 -24026
rect 3225 -24060 3231 -24026
rect 3269 -24060 3293 -24026
rect 3293 -24060 3303 -24026
rect 3927 -24060 3937 -24026
rect 3937 -24060 3961 -24026
rect 3999 -24060 4005 -24026
rect 4005 -24060 4033 -24026
rect 4071 -24060 4073 -24026
rect 4073 -24060 4105 -24026
rect 4143 -24060 4175 -24026
rect 4175 -24060 4177 -24026
rect 4215 -24060 4243 -24026
rect 4243 -24060 4249 -24026
rect 4287 -24060 4311 -24026
rect 4311 -24060 4321 -24026
rect 4945 -24060 4955 -24026
rect 4955 -24060 4979 -24026
rect 5017 -24060 5023 -24026
rect 5023 -24060 5051 -24026
rect 5089 -24060 5091 -24026
rect 5091 -24060 5123 -24026
rect 5161 -24060 5193 -24026
rect 5193 -24060 5195 -24026
rect 5233 -24060 5261 -24026
rect 5261 -24060 5267 -24026
rect 5305 -24060 5329 -24026
rect 5329 -24060 5339 -24026
rect 5963 -24060 5973 -24026
rect 5973 -24060 5997 -24026
rect 6035 -24060 6041 -24026
rect 6041 -24060 6069 -24026
rect 6107 -24060 6109 -24026
rect 6109 -24060 6141 -24026
rect 6179 -24060 6211 -24026
rect 6211 -24060 6213 -24026
rect 6251 -24060 6279 -24026
rect 6279 -24060 6285 -24026
rect 6323 -24060 6347 -24026
rect 6347 -24060 6357 -24026
rect 6981 -24060 6991 -24026
rect 6991 -24060 7015 -24026
rect 7053 -24060 7059 -24026
rect 7059 -24060 7087 -24026
rect 7125 -24060 7127 -24026
rect 7127 -24060 7159 -24026
rect 7197 -24060 7229 -24026
rect 7229 -24060 7231 -24026
rect 7269 -24060 7297 -24026
rect 7297 -24060 7303 -24026
rect 7341 -24060 7365 -24026
rect 7365 -24060 7375 -24026
rect 7999 -24060 8009 -24026
rect 8009 -24060 8033 -24026
rect 8071 -24060 8077 -24026
rect 8077 -24060 8105 -24026
rect 8143 -24060 8145 -24026
rect 8145 -24060 8177 -24026
rect 8215 -24060 8247 -24026
rect 8247 -24060 8249 -24026
rect 8287 -24060 8315 -24026
rect 8315 -24060 8321 -24026
rect 8359 -24060 8383 -24026
rect 8383 -24060 8393 -24026
rect 9017 -24060 9027 -24026
rect 9027 -24060 9051 -24026
rect 9089 -24060 9095 -24026
rect 9095 -24060 9123 -24026
rect 9161 -24060 9163 -24026
rect 9163 -24060 9195 -24026
rect 9233 -24060 9265 -24026
rect 9265 -24060 9267 -24026
rect 9305 -24060 9333 -24026
rect 9333 -24060 9339 -24026
rect 9377 -24060 9401 -24026
rect 9401 -24060 9411 -24026
rect 10035 -24060 10045 -24026
rect 10045 -24060 10069 -24026
rect 10107 -24060 10113 -24026
rect 10113 -24060 10141 -24026
rect 10179 -24060 10181 -24026
rect 10181 -24060 10213 -24026
rect 10251 -24060 10283 -24026
rect 10283 -24060 10285 -24026
rect 10323 -24060 10351 -24026
rect 10351 -24060 10357 -24026
rect 10395 -24060 10419 -24026
rect 10419 -24060 10429 -24026
rect 11053 -24060 11063 -24026
rect 11063 -24060 11087 -24026
rect 11125 -24060 11131 -24026
rect 11131 -24060 11159 -24026
rect 11197 -24060 11199 -24026
rect 11199 -24060 11231 -24026
rect 11269 -24060 11301 -24026
rect 11301 -24060 11303 -24026
rect 11341 -24060 11369 -24026
rect 11369 -24060 11375 -24026
rect 11413 -24060 11437 -24026
rect 11437 -24060 11447 -24026
rect 12071 -24060 12081 -24026
rect 12081 -24060 12105 -24026
rect 12143 -24060 12149 -24026
rect 12149 -24060 12177 -24026
rect 12215 -24060 12217 -24026
rect 12217 -24060 12249 -24026
rect 12287 -24060 12319 -24026
rect 12319 -24060 12321 -24026
rect 12359 -24060 12387 -24026
rect 12387 -24060 12393 -24026
rect 12431 -24060 12455 -24026
rect 12455 -24060 12465 -24026
rect 13089 -24060 13099 -24026
rect 13099 -24060 13123 -24026
rect 13161 -24060 13167 -24026
rect 13167 -24060 13195 -24026
rect 13233 -24060 13235 -24026
rect 13235 -24060 13267 -24026
rect 13305 -24060 13337 -24026
rect 13337 -24060 13339 -24026
rect 13377 -24060 13405 -24026
rect 13405 -24060 13411 -24026
rect 13449 -24060 13473 -24026
rect 13473 -24060 13483 -24026
rect 14107 -24060 14117 -24026
rect 14117 -24060 14141 -24026
rect 14179 -24060 14185 -24026
rect 14185 -24060 14213 -24026
rect 14251 -24060 14253 -24026
rect 14253 -24060 14285 -24026
rect 14323 -24060 14355 -24026
rect 14355 -24060 14357 -24026
rect 14395 -24060 14423 -24026
rect 14423 -24060 14429 -24026
rect 14467 -24060 14491 -24026
rect 14491 -24060 14501 -24026
rect 15125 -24060 15135 -24026
rect 15135 -24060 15159 -24026
rect 15197 -24060 15203 -24026
rect 15203 -24060 15231 -24026
rect 15269 -24060 15271 -24026
rect 15271 -24060 15303 -24026
rect 15341 -24060 15373 -24026
rect 15373 -24060 15375 -24026
rect 15413 -24060 15441 -24026
rect 15441 -24060 15447 -24026
rect 15485 -24060 15509 -24026
rect 15509 -24060 15519 -24026
rect 16143 -24060 16153 -24026
rect 16153 -24060 16177 -24026
rect 16215 -24060 16221 -24026
rect 16221 -24060 16249 -24026
rect 16287 -24060 16289 -24026
rect 16289 -24060 16321 -24026
rect 16359 -24060 16391 -24026
rect 16391 -24060 16393 -24026
rect 16431 -24060 16459 -24026
rect 16459 -24060 16465 -24026
rect 16503 -24060 16527 -24026
rect 16527 -24060 16537 -24026
rect 17161 -24060 17171 -24026
rect 17171 -24060 17195 -24026
rect 17233 -24060 17239 -24026
rect 17239 -24060 17267 -24026
rect 17305 -24060 17307 -24026
rect 17307 -24060 17339 -24026
rect 17377 -24060 17409 -24026
rect 17409 -24060 17411 -24026
rect 17449 -24060 17477 -24026
rect 17477 -24060 17483 -24026
rect 17521 -24060 17545 -24026
rect 17545 -24060 17555 -24026
rect 18179 -24060 18189 -24026
rect 18189 -24060 18213 -24026
rect 18251 -24060 18257 -24026
rect 18257 -24060 18285 -24026
rect 18323 -24060 18325 -24026
rect 18325 -24060 18357 -24026
rect 18395 -24060 18427 -24026
rect 18427 -24060 18429 -24026
rect 18467 -24060 18495 -24026
rect 18495 -24060 18501 -24026
rect 18539 -24060 18563 -24026
rect 18563 -24060 18573 -24026
rect 19197 -24060 19207 -24026
rect 19207 -24060 19231 -24026
rect 19269 -24060 19275 -24026
rect 19275 -24060 19303 -24026
rect 19341 -24060 19343 -24026
rect 19343 -24060 19375 -24026
rect 19413 -24060 19445 -24026
rect 19445 -24060 19447 -24026
rect 19485 -24060 19513 -24026
rect 19513 -24060 19519 -24026
rect 19557 -24060 19581 -24026
rect 19581 -24060 19591 -24026
rect 20215 -24060 20225 -24026
rect 20225 -24060 20249 -24026
rect 20287 -24060 20293 -24026
rect 20293 -24060 20321 -24026
rect 20359 -24060 20361 -24026
rect 20361 -24060 20393 -24026
rect 20431 -24060 20463 -24026
rect 20463 -24060 20465 -24026
rect 20503 -24060 20531 -24026
rect 20531 -24060 20537 -24026
rect 20575 -24060 20599 -24026
rect 20599 -24060 20609 -24026
rect 21233 -24060 21243 -24026
rect 21243 -24060 21267 -24026
rect 21305 -24060 21311 -24026
rect 21311 -24060 21339 -24026
rect 21377 -24060 21379 -24026
rect 21379 -24060 21411 -24026
rect 21449 -24060 21481 -24026
rect 21481 -24060 21483 -24026
rect 21521 -24060 21549 -24026
rect 21549 -24060 21555 -24026
rect 21593 -24060 21617 -24026
rect 21617 -24060 21627 -24026
rect 22251 -24060 22261 -24026
rect 22261 -24060 22285 -24026
rect 22323 -24060 22329 -24026
rect 22329 -24060 22357 -24026
rect 22395 -24060 22397 -24026
rect 22397 -24060 22429 -24026
rect 22467 -24060 22499 -24026
rect 22499 -24060 22501 -24026
rect 22539 -24060 22567 -24026
rect 22567 -24060 22573 -24026
rect 22611 -24060 22635 -24026
rect 22635 -24060 22645 -24026
rect 24855 -24045 24889 -24043
rect 24855 -24077 24889 -24045
rect -12289 -24147 -12255 -24115
rect -12289 -24149 -12255 -24147
rect -12289 -24215 -12255 -24187
rect -12289 -24221 -12255 -24215
rect -12289 -24283 -12255 -24259
rect -12289 -24293 -12255 -24283
rect -12289 -24351 -12255 -24331
rect -12289 -24365 -12255 -24351
rect -12289 -24419 -12255 -24403
rect -12289 -24437 -12255 -24419
rect -12289 -24487 -12255 -24475
rect -12289 -24509 -12255 -24487
rect -12289 -24555 -12255 -24547
rect -12289 -24581 -12255 -24555
rect -12289 -24623 -12255 -24619
rect -12289 -24653 -12255 -24623
rect -12289 -24725 -12255 -24691
rect 2580 -24143 2614 -24129
rect 2580 -24163 2614 -24143
rect 2580 -24211 2614 -24201
rect 2580 -24235 2614 -24211
rect 2580 -24279 2614 -24273
rect 2580 -24307 2614 -24279
rect 2580 -24347 2614 -24345
rect 2580 -24379 2614 -24347
rect 2580 -24449 2614 -24417
rect 2580 -24451 2614 -24449
rect 2580 -24517 2614 -24489
rect 2580 -24523 2614 -24517
rect 2580 -24585 2614 -24561
rect 2580 -24595 2614 -24585
rect 2580 -24653 2614 -24633
rect 2580 -24667 2614 -24653
rect 3598 -24143 3632 -24129
rect 3598 -24163 3632 -24143
rect 3598 -24211 3632 -24201
rect 3598 -24235 3632 -24211
rect 3598 -24279 3632 -24273
rect 3598 -24307 3632 -24279
rect 3598 -24347 3632 -24345
rect 3598 -24379 3632 -24347
rect 3598 -24449 3632 -24417
rect 3598 -24451 3632 -24449
rect 3598 -24517 3632 -24489
rect 3598 -24523 3632 -24517
rect 3598 -24585 3632 -24561
rect 3598 -24595 3632 -24585
rect 3598 -24653 3632 -24633
rect 3598 -24667 3632 -24653
rect 4616 -24143 4650 -24129
rect 4616 -24163 4650 -24143
rect 4616 -24211 4650 -24201
rect 4616 -24235 4650 -24211
rect 4616 -24279 4650 -24273
rect 4616 -24307 4650 -24279
rect 4616 -24347 4650 -24345
rect 4616 -24379 4650 -24347
rect 4616 -24449 4650 -24417
rect 4616 -24451 4650 -24449
rect 4616 -24517 4650 -24489
rect 4616 -24523 4650 -24517
rect 4616 -24585 4650 -24561
rect 4616 -24595 4650 -24585
rect 4616 -24653 4650 -24633
rect 4616 -24667 4650 -24653
rect 5634 -24143 5668 -24129
rect 5634 -24163 5668 -24143
rect 5634 -24211 5668 -24201
rect 5634 -24235 5668 -24211
rect 5634 -24279 5668 -24273
rect 5634 -24307 5668 -24279
rect 5634 -24347 5668 -24345
rect 5634 -24379 5668 -24347
rect 5634 -24449 5668 -24417
rect 5634 -24451 5668 -24449
rect 5634 -24517 5668 -24489
rect 5634 -24523 5668 -24517
rect 5634 -24585 5668 -24561
rect 5634 -24595 5668 -24585
rect 5634 -24653 5668 -24633
rect 5634 -24667 5668 -24653
rect 6652 -24143 6686 -24129
rect 6652 -24163 6686 -24143
rect 6652 -24211 6686 -24201
rect 6652 -24235 6686 -24211
rect 6652 -24279 6686 -24273
rect 6652 -24307 6686 -24279
rect 6652 -24347 6686 -24345
rect 6652 -24379 6686 -24347
rect 6652 -24449 6686 -24417
rect 6652 -24451 6686 -24449
rect 6652 -24517 6686 -24489
rect 6652 -24523 6686 -24517
rect 6652 -24585 6686 -24561
rect 6652 -24595 6686 -24585
rect 6652 -24653 6686 -24633
rect 6652 -24667 6686 -24653
rect 7670 -24143 7704 -24129
rect 7670 -24163 7704 -24143
rect 7670 -24211 7704 -24201
rect 7670 -24235 7704 -24211
rect 7670 -24279 7704 -24273
rect 7670 -24307 7704 -24279
rect 7670 -24347 7704 -24345
rect 7670 -24379 7704 -24347
rect 7670 -24449 7704 -24417
rect 7670 -24451 7704 -24449
rect 7670 -24517 7704 -24489
rect 7670 -24523 7704 -24517
rect 7670 -24585 7704 -24561
rect 7670 -24595 7704 -24585
rect 7670 -24653 7704 -24633
rect 7670 -24667 7704 -24653
rect 8688 -24143 8722 -24129
rect 8688 -24163 8722 -24143
rect 8688 -24211 8722 -24201
rect 8688 -24235 8722 -24211
rect 8688 -24279 8722 -24273
rect 8688 -24307 8722 -24279
rect 8688 -24347 8722 -24345
rect 8688 -24379 8722 -24347
rect 8688 -24449 8722 -24417
rect 8688 -24451 8722 -24449
rect 8688 -24517 8722 -24489
rect 8688 -24523 8722 -24517
rect 8688 -24585 8722 -24561
rect 8688 -24595 8722 -24585
rect 8688 -24653 8722 -24633
rect 8688 -24667 8722 -24653
rect 9706 -24143 9740 -24129
rect 9706 -24163 9740 -24143
rect 9706 -24211 9740 -24201
rect 9706 -24235 9740 -24211
rect 9706 -24279 9740 -24273
rect 9706 -24307 9740 -24279
rect 9706 -24347 9740 -24345
rect 9706 -24379 9740 -24347
rect 9706 -24449 9740 -24417
rect 9706 -24451 9740 -24449
rect 9706 -24517 9740 -24489
rect 9706 -24523 9740 -24517
rect 9706 -24585 9740 -24561
rect 9706 -24595 9740 -24585
rect 9706 -24653 9740 -24633
rect 9706 -24667 9740 -24653
rect 10724 -24143 10758 -24129
rect 10724 -24163 10758 -24143
rect 10724 -24211 10758 -24201
rect 10724 -24235 10758 -24211
rect 10724 -24279 10758 -24273
rect 10724 -24307 10758 -24279
rect 10724 -24347 10758 -24345
rect 10724 -24379 10758 -24347
rect 10724 -24449 10758 -24417
rect 10724 -24451 10758 -24449
rect 10724 -24517 10758 -24489
rect 10724 -24523 10758 -24517
rect 10724 -24585 10758 -24561
rect 10724 -24595 10758 -24585
rect 10724 -24653 10758 -24633
rect 10724 -24667 10758 -24653
rect 11742 -24143 11776 -24129
rect 11742 -24163 11776 -24143
rect 11742 -24211 11776 -24201
rect 11742 -24235 11776 -24211
rect 11742 -24279 11776 -24273
rect 11742 -24307 11776 -24279
rect 11742 -24347 11776 -24345
rect 11742 -24379 11776 -24347
rect 11742 -24449 11776 -24417
rect 11742 -24451 11776 -24449
rect 11742 -24517 11776 -24489
rect 11742 -24523 11776 -24517
rect 11742 -24585 11776 -24561
rect 11742 -24595 11776 -24585
rect 11742 -24653 11776 -24633
rect 11742 -24667 11776 -24653
rect 12760 -24143 12794 -24129
rect 12760 -24163 12794 -24143
rect 12760 -24211 12794 -24201
rect 12760 -24235 12794 -24211
rect 12760 -24279 12794 -24273
rect 12760 -24307 12794 -24279
rect 12760 -24347 12794 -24345
rect 12760 -24379 12794 -24347
rect 12760 -24449 12794 -24417
rect 12760 -24451 12794 -24449
rect 12760 -24517 12794 -24489
rect 12760 -24523 12794 -24517
rect 12760 -24585 12794 -24561
rect 12760 -24595 12794 -24585
rect 12760 -24653 12794 -24633
rect 12760 -24667 12794 -24653
rect 13778 -24143 13812 -24129
rect 13778 -24163 13812 -24143
rect 13778 -24211 13812 -24201
rect 13778 -24235 13812 -24211
rect 13778 -24279 13812 -24273
rect 13778 -24307 13812 -24279
rect 13778 -24347 13812 -24345
rect 13778 -24379 13812 -24347
rect 13778 -24449 13812 -24417
rect 13778 -24451 13812 -24449
rect 13778 -24517 13812 -24489
rect 13778 -24523 13812 -24517
rect 13778 -24585 13812 -24561
rect 13778 -24595 13812 -24585
rect 13778 -24653 13812 -24633
rect 13778 -24667 13812 -24653
rect 14796 -24143 14830 -24129
rect 14796 -24163 14830 -24143
rect 14796 -24211 14830 -24201
rect 14796 -24235 14830 -24211
rect 14796 -24279 14830 -24273
rect 14796 -24307 14830 -24279
rect 14796 -24347 14830 -24345
rect 14796 -24379 14830 -24347
rect 14796 -24449 14830 -24417
rect 14796 -24451 14830 -24449
rect 14796 -24517 14830 -24489
rect 14796 -24523 14830 -24517
rect 14796 -24585 14830 -24561
rect 14796 -24595 14830 -24585
rect 14796 -24653 14830 -24633
rect 14796 -24667 14830 -24653
rect 15814 -24143 15848 -24129
rect 15814 -24163 15848 -24143
rect 15814 -24211 15848 -24201
rect 15814 -24235 15848 -24211
rect 15814 -24279 15848 -24273
rect 15814 -24307 15848 -24279
rect 15814 -24347 15848 -24345
rect 15814 -24379 15848 -24347
rect 15814 -24449 15848 -24417
rect 15814 -24451 15848 -24449
rect 15814 -24517 15848 -24489
rect 15814 -24523 15848 -24517
rect 15814 -24585 15848 -24561
rect 15814 -24595 15848 -24585
rect 15814 -24653 15848 -24633
rect 15814 -24667 15848 -24653
rect 16832 -24143 16866 -24129
rect 16832 -24163 16866 -24143
rect 16832 -24211 16866 -24201
rect 16832 -24235 16866 -24211
rect 16832 -24279 16866 -24273
rect 16832 -24307 16866 -24279
rect 16832 -24347 16866 -24345
rect 16832 -24379 16866 -24347
rect 16832 -24449 16866 -24417
rect 16832 -24451 16866 -24449
rect 16832 -24517 16866 -24489
rect 16832 -24523 16866 -24517
rect 16832 -24585 16866 -24561
rect 16832 -24595 16866 -24585
rect 16832 -24653 16866 -24633
rect 16832 -24667 16866 -24653
rect 17850 -24143 17884 -24129
rect 17850 -24163 17884 -24143
rect 17850 -24211 17884 -24201
rect 17850 -24235 17884 -24211
rect 17850 -24279 17884 -24273
rect 17850 -24307 17884 -24279
rect 17850 -24347 17884 -24345
rect 17850 -24379 17884 -24347
rect 17850 -24449 17884 -24417
rect 17850 -24451 17884 -24449
rect 17850 -24517 17884 -24489
rect 17850 -24523 17884 -24517
rect 17850 -24585 17884 -24561
rect 17850 -24595 17884 -24585
rect 17850 -24653 17884 -24633
rect 17850 -24667 17884 -24653
rect 18868 -24143 18902 -24129
rect 18868 -24163 18902 -24143
rect 18868 -24211 18902 -24201
rect 18868 -24235 18902 -24211
rect 18868 -24279 18902 -24273
rect 18868 -24307 18902 -24279
rect 18868 -24347 18902 -24345
rect 18868 -24379 18902 -24347
rect 18868 -24449 18902 -24417
rect 18868 -24451 18902 -24449
rect 18868 -24517 18902 -24489
rect 18868 -24523 18902 -24517
rect 18868 -24585 18902 -24561
rect 18868 -24595 18902 -24585
rect 18868 -24653 18902 -24633
rect 18868 -24667 18902 -24653
rect 19886 -24143 19920 -24129
rect 19886 -24163 19920 -24143
rect 19886 -24211 19920 -24201
rect 19886 -24235 19920 -24211
rect 19886 -24279 19920 -24273
rect 19886 -24307 19920 -24279
rect 19886 -24347 19920 -24345
rect 19886 -24379 19920 -24347
rect 19886 -24449 19920 -24417
rect 19886 -24451 19920 -24449
rect 19886 -24517 19920 -24489
rect 19886 -24523 19920 -24517
rect 19886 -24585 19920 -24561
rect 19886 -24595 19920 -24585
rect 19886 -24653 19920 -24633
rect 19886 -24667 19920 -24653
rect 20904 -24143 20938 -24129
rect 20904 -24163 20938 -24143
rect 20904 -24211 20938 -24201
rect 20904 -24235 20938 -24211
rect 20904 -24279 20938 -24273
rect 20904 -24307 20938 -24279
rect 20904 -24347 20938 -24345
rect 20904 -24379 20938 -24347
rect 20904 -24449 20938 -24417
rect 20904 -24451 20938 -24449
rect 20904 -24517 20938 -24489
rect 20904 -24523 20938 -24517
rect 20904 -24585 20938 -24561
rect 20904 -24595 20938 -24585
rect 20904 -24653 20938 -24633
rect 20904 -24667 20938 -24653
rect 21922 -24143 21956 -24129
rect 21922 -24163 21956 -24143
rect 21922 -24211 21956 -24201
rect 21922 -24235 21956 -24211
rect 21922 -24279 21956 -24273
rect 21922 -24307 21956 -24279
rect 21922 -24347 21956 -24345
rect 21922 -24379 21956 -24347
rect 21922 -24449 21956 -24417
rect 21922 -24451 21956 -24449
rect 21922 -24517 21956 -24489
rect 21922 -24523 21956 -24517
rect 21922 -24585 21956 -24561
rect 21922 -24595 21956 -24585
rect 21922 -24653 21956 -24633
rect 21922 -24667 21956 -24653
rect 22940 -24143 22974 -24129
rect 22940 -24163 22974 -24143
rect 22940 -24211 22974 -24201
rect 22940 -24235 22974 -24211
rect 22940 -24279 22974 -24273
rect 22940 -24307 22974 -24279
rect 22940 -24347 22974 -24345
rect 22940 -24379 22974 -24347
rect 22940 -24449 22974 -24417
rect 22940 -24451 22974 -24449
rect 22940 -24517 22974 -24489
rect 22940 -24523 22974 -24517
rect 22940 -24585 22974 -24561
rect 22940 -24595 22974 -24585
rect 22940 -24653 22974 -24633
rect 22940 -24667 22974 -24653
rect 24855 -24147 24889 -24115
rect 24855 -24149 24889 -24147
rect 24855 -24215 24889 -24187
rect 24855 -24221 24889 -24215
rect 24855 -24283 24889 -24259
rect 24855 -24293 24889 -24283
rect 24855 -24351 24889 -24331
rect 24855 -24365 24889 -24351
rect 24855 -24419 24889 -24403
rect 24855 -24437 24889 -24419
rect 24855 -24487 24889 -24475
rect 24855 -24509 24889 -24487
rect 24855 -24555 24889 -24547
rect 24855 -24581 24889 -24555
rect 24855 -24623 24889 -24619
rect 24855 -24653 24889 -24623
rect 24855 -24725 24889 -24691
rect -12289 -24793 -12255 -24763
rect -12289 -24797 -12255 -24793
rect 2909 -24770 2919 -24736
rect 2919 -24770 2943 -24736
rect 2981 -24770 2987 -24736
rect 2987 -24770 3015 -24736
rect 3053 -24770 3055 -24736
rect 3055 -24770 3087 -24736
rect 3125 -24770 3157 -24736
rect 3157 -24770 3159 -24736
rect 3197 -24770 3225 -24736
rect 3225 -24770 3231 -24736
rect 3269 -24770 3293 -24736
rect 3293 -24770 3303 -24736
rect 3927 -24770 3937 -24736
rect 3937 -24770 3961 -24736
rect 3999 -24770 4005 -24736
rect 4005 -24770 4033 -24736
rect 4071 -24770 4073 -24736
rect 4073 -24770 4105 -24736
rect 4143 -24770 4175 -24736
rect 4175 -24770 4177 -24736
rect 4215 -24770 4243 -24736
rect 4243 -24770 4249 -24736
rect 4287 -24770 4311 -24736
rect 4311 -24770 4321 -24736
rect 4945 -24770 4955 -24736
rect 4955 -24770 4979 -24736
rect 5017 -24770 5023 -24736
rect 5023 -24770 5051 -24736
rect 5089 -24770 5091 -24736
rect 5091 -24770 5123 -24736
rect 5161 -24770 5193 -24736
rect 5193 -24770 5195 -24736
rect 5233 -24770 5261 -24736
rect 5261 -24770 5267 -24736
rect 5305 -24770 5329 -24736
rect 5329 -24770 5339 -24736
rect 5963 -24770 5973 -24736
rect 5973 -24770 5997 -24736
rect 6035 -24770 6041 -24736
rect 6041 -24770 6069 -24736
rect 6107 -24770 6109 -24736
rect 6109 -24770 6141 -24736
rect 6179 -24770 6211 -24736
rect 6211 -24770 6213 -24736
rect 6251 -24770 6279 -24736
rect 6279 -24770 6285 -24736
rect 6323 -24770 6347 -24736
rect 6347 -24770 6357 -24736
rect 6981 -24770 6991 -24736
rect 6991 -24770 7015 -24736
rect 7053 -24770 7059 -24736
rect 7059 -24770 7087 -24736
rect 7125 -24770 7127 -24736
rect 7127 -24770 7159 -24736
rect 7197 -24770 7229 -24736
rect 7229 -24770 7231 -24736
rect 7269 -24770 7297 -24736
rect 7297 -24770 7303 -24736
rect 7341 -24770 7365 -24736
rect 7365 -24770 7375 -24736
rect 7999 -24770 8009 -24736
rect 8009 -24770 8033 -24736
rect 8071 -24770 8077 -24736
rect 8077 -24770 8105 -24736
rect 8143 -24770 8145 -24736
rect 8145 -24770 8177 -24736
rect 8215 -24770 8247 -24736
rect 8247 -24770 8249 -24736
rect 8287 -24770 8315 -24736
rect 8315 -24770 8321 -24736
rect 8359 -24770 8383 -24736
rect 8383 -24770 8393 -24736
rect 9017 -24770 9027 -24736
rect 9027 -24770 9051 -24736
rect 9089 -24770 9095 -24736
rect 9095 -24770 9123 -24736
rect 9161 -24770 9163 -24736
rect 9163 -24770 9195 -24736
rect 9233 -24770 9265 -24736
rect 9265 -24770 9267 -24736
rect 9305 -24770 9333 -24736
rect 9333 -24770 9339 -24736
rect 9377 -24770 9401 -24736
rect 9401 -24770 9411 -24736
rect 10035 -24770 10045 -24736
rect 10045 -24770 10069 -24736
rect 10107 -24770 10113 -24736
rect 10113 -24770 10141 -24736
rect 10179 -24770 10181 -24736
rect 10181 -24770 10213 -24736
rect 10251 -24770 10283 -24736
rect 10283 -24770 10285 -24736
rect 10323 -24770 10351 -24736
rect 10351 -24770 10357 -24736
rect 10395 -24770 10419 -24736
rect 10419 -24770 10429 -24736
rect 11053 -24770 11063 -24736
rect 11063 -24770 11087 -24736
rect 11125 -24770 11131 -24736
rect 11131 -24770 11159 -24736
rect 11197 -24770 11199 -24736
rect 11199 -24770 11231 -24736
rect 11269 -24770 11301 -24736
rect 11301 -24770 11303 -24736
rect 11341 -24770 11369 -24736
rect 11369 -24770 11375 -24736
rect 11413 -24770 11437 -24736
rect 11437 -24770 11447 -24736
rect 12071 -24770 12081 -24736
rect 12081 -24770 12105 -24736
rect 12143 -24770 12149 -24736
rect 12149 -24770 12177 -24736
rect 12215 -24770 12217 -24736
rect 12217 -24770 12249 -24736
rect 12287 -24770 12319 -24736
rect 12319 -24770 12321 -24736
rect 12359 -24770 12387 -24736
rect 12387 -24770 12393 -24736
rect 12431 -24770 12455 -24736
rect 12455 -24770 12465 -24736
rect 13089 -24770 13099 -24736
rect 13099 -24770 13123 -24736
rect 13161 -24770 13167 -24736
rect 13167 -24770 13195 -24736
rect 13233 -24770 13235 -24736
rect 13235 -24770 13267 -24736
rect 13305 -24770 13337 -24736
rect 13337 -24770 13339 -24736
rect 13377 -24770 13405 -24736
rect 13405 -24770 13411 -24736
rect 13449 -24770 13473 -24736
rect 13473 -24770 13483 -24736
rect 14107 -24770 14117 -24736
rect 14117 -24770 14141 -24736
rect 14179 -24770 14185 -24736
rect 14185 -24770 14213 -24736
rect 14251 -24770 14253 -24736
rect 14253 -24770 14285 -24736
rect 14323 -24770 14355 -24736
rect 14355 -24770 14357 -24736
rect 14395 -24770 14423 -24736
rect 14423 -24770 14429 -24736
rect 14467 -24770 14491 -24736
rect 14491 -24770 14501 -24736
rect 15125 -24770 15135 -24736
rect 15135 -24770 15159 -24736
rect 15197 -24770 15203 -24736
rect 15203 -24770 15231 -24736
rect 15269 -24770 15271 -24736
rect 15271 -24770 15303 -24736
rect 15341 -24770 15373 -24736
rect 15373 -24770 15375 -24736
rect 15413 -24770 15441 -24736
rect 15441 -24770 15447 -24736
rect 15485 -24770 15509 -24736
rect 15509 -24770 15519 -24736
rect 16143 -24770 16153 -24736
rect 16153 -24770 16177 -24736
rect 16215 -24770 16221 -24736
rect 16221 -24770 16249 -24736
rect 16287 -24770 16289 -24736
rect 16289 -24770 16321 -24736
rect 16359 -24770 16391 -24736
rect 16391 -24770 16393 -24736
rect 16431 -24770 16459 -24736
rect 16459 -24770 16465 -24736
rect 16503 -24770 16527 -24736
rect 16527 -24770 16537 -24736
rect 17161 -24770 17171 -24736
rect 17171 -24770 17195 -24736
rect 17233 -24770 17239 -24736
rect 17239 -24770 17267 -24736
rect 17305 -24770 17307 -24736
rect 17307 -24770 17339 -24736
rect 17377 -24770 17409 -24736
rect 17409 -24770 17411 -24736
rect 17449 -24770 17477 -24736
rect 17477 -24770 17483 -24736
rect 17521 -24770 17545 -24736
rect 17545 -24770 17555 -24736
rect 18179 -24770 18189 -24736
rect 18189 -24770 18213 -24736
rect 18251 -24770 18257 -24736
rect 18257 -24770 18285 -24736
rect 18323 -24770 18325 -24736
rect 18325 -24770 18357 -24736
rect 18395 -24770 18427 -24736
rect 18427 -24770 18429 -24736
rect 18467 -24770 18495 -24736
rect 18495 -24770 18501 -24736
rect 18539 -24770 18563 -24736
rect 18563 -24770 18573 -24736
rect 19197 -24770 19207 -24736
rect 19207 -24770 19231 -24736
rect 19269 -24770 19275 -24736
rect 19275 -24770 19303 -24736
rect 19341 -24770 19343 -24736
rect 19343 -24770 19375 -24736
rect 19413 -24770 19445 -24736
rect 19445 -24770 19447 -24736
rect 19485 -24770 19513 -24736
rect 19513 -24770 19519 -24736
rect 19557 -24770 19581 -24736
rect 19581 -24770 19591 -24736
rect 20215 -24770 20225 -24736
rect 20225 -24770 20249 -24736
rect 20287 -24770 20293 -24736
rect 20293 -24770 20321 -24736
rect 20359 -24770 20361 -24736
rect 20361 -24770 20393 -24736
rect 20431 -24770 20463 -24736
rect 20463 -24770 20465 -24736
rect 20503 -24770 20531 -24736
rect 20531 -24770 20537 -24736
rect 20575 -24770 20599 -24736
rect 20599 -24770 20609 -24736
rect 21233 -24770 21243 -24736
rect 21243 -24770 21267 -24736
rect 21305 -24770 21311 -24736
rect 21311 -24770 21339 -24736
rect 21377 -24770 21379 -24736
rect 21379 -24770 21411 -24736
rect 21449 -24770 21481 -24736
rect 21481 -24770 21483 -24736
rect 21521 -24770 21549 -24736
rect 21549 -24770 21555 -24736
rect 21593 -24770 21617 -24736
rect 21617 -24770 21627 -24736
rect 22251 -24770 22261 -24736
rect 22261 -24770 22285 -24736
rect 22323 -24770 22329 -24736
rect 22329 -24770 22357 -24736
rect 22395 -24770 22397 -24736
rect 22397 -24770 22429 -24736
rect 22467 -24770 22499 -24736
rect 22499 -24770 22501 -24736
rect 22539 -24770 22567 -24736
rect 22567 -24770 22573 -24736
rect 22611 -24770 22635 -24736
rect 22635 -24770 22645 -24736
rect -12289 -24861 -12255 -24835
rect -12289 -24869 -12255 -24861
rect -12289 -24929 -12255 -24907
rect -12289 -24941 -12255 -24929
rect -12289 -24997 -12255 -24979
rect -12289 -25013 -12255 -24997
rect -12289 -25065 -12255 -25051
rect -12289 -25085 -12255 -25065
rect -12289 -25133 -12255 -25123
rect -12289 -25157 -12255 -25133
rect -12289 -25201 -12255 -25195
rect -12289 -25229 -12255 -25201
rect -12289 -25269 -12255 -25267
rect -12289 -25301 -12255 -25269
rect -12289 -25371 -12255 -25339
rect -12289 -25373 -12255 -25371
rect -12289 -25439 -12255 -25411
rect -12289 -25445 -12255 -25439
rect -12289 -25507 -12255 -25483
rect -12289 -25517 -12255 -25507
rect -12289 -25575 -12255 -25555
rect -12289 -25589 -12255 -25575
rect -12289 -25643 -12255 -25627
rect -12289 -25661 -12255 -25643
rect -12289 -25711 -12255 -25699
rect -12289 -25733 -12255 -25711
rect -12289 -25779 -12255 -25771
rect -12289 -25805 -12255 -25779
rect -12289 -25847 -12255 -25843
rect -12289 -25877 -12255 -25847
rect -12289 -25949 -12255 -25915
rect -12289 -26017 -12255 -25987
rect -12289 -26021 -12255 -26017
rect -12289 -26085 -12255 -26059
rect -12289 -26093 -12255 -26085
rect -12289 -26153 -12255 -26131
rect -12289 -26165 -12255 -26153
rect -12289 -26221 -12255 -26203
rect -12289 -26237 -12255 -26221
rect -12289 -26289 -12255 -26275
rect -12289 -26309 -12255 -26289
rect 24855 -24793 24889 -24763
rect 24855 -24797 24889 -24793
rect 24855 -24861 24889 -24835
rect 24855 -24869 24889 -24861
rect 24855 -24929 24889 -24907
rect 24855 -24941 24889 -24929
rect 24855 -24997 24889 -24979
rect 24855 -25013 24889 -24997
rect 24855 -25065 24889 -25051
rect 24855 -25085 24889 -25065
rect 24855 -25133 24889 -25123
rect 24855 -25157 24889 -25133
rect 24855 -25201 24889 -25195
rect 24855 -25229 24889 -25201
rect 24855 -25269 24889 -25267
rect 24855 -25301 24889 -25269
rect 24855 -25371 24889 -25339
rect 24855 -25373 24889 -25371
rect 24855 -25439 24889 -25411
rect 24855 -25445 24889 -25439
rect 24855 -25507 24889 -25483
rect 24855 -25517 24889 -25507
rect 24855 -25575 24889 -25555
rect 24855 -25589 24889 -25575
rect 24855 -25643 24889 -25627
rect 24855 -25661 24889 -25643
rect 24855 -25711 24889 -25699
rect 24855 -25733 24889 -25711
rect 24855 -25779 24889 -25771
rect 24855 -25805 24889 -25779
rect 24855 -25847 24889 -25843
rect 24855 -25877 24889 -25847
rect 24855 -25949 24889 -25915
rect 24855 -26017 24889 -25987
rect 24855 -26021 24889 -26017
rect 24855 -26085 24889 -26059
rect 24855 -26093 24889 -26085
rect 24855 -26153 24889 -26131
rect 24855 -26165 24889 -26153
rect 24855 -26221 24889 -26203
rect 24855 -26237 24889 -26221
rect 24855 -26289 24889 -26275
rect 24855 -26309 24889 -26289
rect -12221 -27189 -12187 -27155
rect -12149 -27189 -12145 -27155
rect -12145 -27189 -12115 -27155
rect -12077 -27189 -12043 -27155
rect -12005 -27189 -11975 -27155
rect -11975 -27189 -11971 -27155
rect -11933 -27189 -11907 -27155
rect -11907 -27189 -11899 -27155
rect -11861 -27189 -11839 -27155
rect -11839 -27189 -11827 -27155
rect -11789 -27189 -11771 -27155
rect -11771 -27189 -11755 -27155
rect -11717 -27189 -11703 -27155
rect -11703 -27189 -11683 -27155
rect -11645 -27189 -11635 -27155
rect -11635 -27189 -11611 -27155
rect -11573 -27189 -11567 -27155
rect -11567 -27189 -11539 -27155
rect -11501 -27189 -11499 -27155
rect -11499 -27189 -11467 -27155
rect -11429 -27189 -11397 -27155
rect -11397 -27189 -11395 -27155
rect -11357 -27189 -11329 -27155
rect -11329 -27189 -11323 -27155
rect -11285 -27189 -11261 -27155
rect -11261 -27189 -11251 -27155
rect -11213 -27189 -11193 -27155
rect -11193 -27189 -11179 -27155
rect -11141 -27189 -11125 -27155
rect -11125 -27189 -11107 -27155
rect -11069 -27189 -11057 -27155
rect -11057 -27189 -11035 -27155
rect -10997 -27189 -10989 -27155
rect -10989 -27189 -10963 -27155
rect -10925 -27189 -10921 -27155
rect -10921 -27189 -10891 -27155
rect -10853 -27189 -10819 -27155
rect -10781 -27189 -10751 -27155
rect -10751 -27189 -10747 -27155
rect -10709 -27189 -10683 -27155
rect -10683 -27189 -10675 -27155
rect -10637 -27189 -10615 -27155
rect -10615 -27189 -10603 -27155
rect -10565 -27189 -10547 -27155
rect -10547 -27189 -10531 -27155
rect -10493 -27189 -10479 -27155
rect -10479 -27189 -10459 -27155
rect -10421 -27189 -10411 -27155
rect -10411 -27189 -10387 -27155
rect -10349 -27189 -10343 -27155
rect -10343 -27189 -10315 -27155
rect -10277 -27189 -10275 -27155
rect -10275 -27189 -10243 -27155
rect -10205 -27189 -10173 -27155
rect -10173 -27189 -10171 -27155
rect -10133 -27189 -10105 -27155
rect -10105 -27189 -10099 -27155
rect -10061 -27189 -10037 -27155
rect -10037 -27189 -10027 -27155
rect -9989 -27189 -9969 -27155
rect -9969 -27189 -9955 -27155
rect -9917 -27189 -9901 -27155
rect -9901 -27189 -9883 -27155
rect -9845 -27189 -9833 -27155
rect -9833 -27189 -9811 -27155
rect -9773 -27189 -9765 -27155
rect -9765 -27189 -9739 -27155
rect -9701 -27189 -9697 -27155
rect -9697 -27189 -9667 -27155
rect -9629 -27189 -9595 -27155
rect -9557 -27189 -9527 -27155
rect -9527 -27189 -9523 -27155
rect -9485 -27189 -9459 -27155
rect -9459 -27189 -9451 -27155
rect -9413 -27189 -9391 -27155
rect -9391 -27189 -9379 -27155
rect -9341 -27189 -9323 -27155
rect -9323 -27189 -9307 -27155
rect -9269 -27189 -9255 -27155
rect -9255 -27189 -9235 -27155
rect -9197 -27189 -9187 -27155
rect -9187 -27189 -9163 -27155
rect -9125 -27189 -9119 -27155
rect -9119 -27189 -9091 -27155
rect -9053 -27189 -9051 -27155
rect -9051 -27189 -9019 -27155
rect -8981 -27189 -8949 -27155
rect -8949 -27189 -8947 -27155
rect -8909 -27189 -8881 -27155
rect -8881 -27189 -8875 -27155
rect -8837 -27189 -8813 -27155
rect -8813 -27189 -8803 -27155
rect -8765 -27189 -8745 -27155
rect -8745 -27189 -8731 -27155
rect -8693 -27189 -8677 -27155
rect -8677 -27189 -8659 -27155
rect -8621 -27189 -8609 -27155
rect -8609 -27189 -8587 -27155
rect -8549 -27189 -8541 -27155
rect -8541 -27189 -8515 -27155
rect -8477 -27189 -8473 -27155
rect -8473 -27189 -8443 -27155
rect -8405 -27189 -8371 -27155
rect -8333 -27189 -8303 -27155
rect -8303 -27189 -8299 -27155
rect -8261 -27189 -8235 -27155
rect -8235 -27189 -8227 -27155
rect -8189 -27189 -8167 -27155
rect -8167 -27189 -8155 -27155
rect -8117 -27189 -8099 -27155
rect -8099 -27189 -8083 -27155
rect -8045 -27189 -8031 -27155
rect -8031 -27189 -8011 -27155
rect -7973 -27189 -7963 -27155
rect -7963 -27189 -7939 -27155
rect -7901 -27189 -7895 -27155
rect -7895 -27189 -7867 -27155
rect -7829 -27189 -7827 -27155
rect -7827 -27189 -7795 -27155
rect -7757 -27189 -7725 -27155
rect -7725 -27189 -7723 -27155
rect -7685 -27189 -7657 -27155
rect -7657 -27189 -7651 -27155
rect -7613 -27189 -7589 -27155
rect -7589 -27189 -7579 -27155
rect -7541 -27189 -7521 -27155
rect -7521 -27189 -7507 -27155
rect -7469 -27189 -7453 -27155
rect -7453 -27189 -7435 -27155
rect -7397 -27189 -7385 -27155
rect -7385 -27189 -7363 -27155
rect -7325 -27189 -7317 -27155
rect -7317 -27189 -7291 -27155
rect -7253 -27189 -7249 -27155
rect -7249 -27189 -7219 -27155
rect -7181 -27189 -7147 -27155
rect -7109 -27189 -7079 -27155
rect -7079 -27189 -7075 -27155
rect -7037 -27189 -7011 -27155
rect -7011 -27189 -7003 -27155
rect -6965 -27189 -6943 -27155
rect -6943 -27189 -6931 -27155
rect -6893 -27189 -6875 -27155
rect -6875 -27189 -6859 -27155
rect -6821 -27189 -6807 -27155
rect -6807 -27189 -6787 -27155
rect -6749 -27189 -6739 -27155
rect -6739 -27189 -6715 -27155
rect -6677 -27189 -6671 -27155
rect -6671 -27189 -6643 -27155
rect -6605 -27189 -6603 -27155
rect -6603 -27189 -6571 -27155
rect -6533 -27189 -6501 -27155
rect -6501 -27189 -6499 -27155
rect -6461 -27189 -6433 -27155
rect -6433 -27189 -6427 -27155
rect -6389 -27189 -6365 -27155
rect -6365 -27189 -6355 -27155
rect -6317 -27189 -6297 -27155
rect -6297 -27189 -6283 -27155
rect -6245 -27189 -6229 -27155
rect -6229 -27189 -6211 -27155
rect -6173 -27189 -6161 -27155
rect -6161 -27189 -6139 -27155
rect -6101 -27189 -6093 -27155
rect -6093 -27189 -6067 -27155
rect -6029 -27189 -6025 -27155
rect -6025 -27189 -5995 -27155
rect -5957 -27189 -5923 -27155
rect -5885 -27189 -5855 -27155
rect -5855 -27189 -5851 -27155
rect -5813 -27189 -5787 -27155
rect -5787 -27189 -5779 -27155
rect -5741 -27189 -5719 -27155
rect -5719 -27189 -5707 -27155
rect -5669 -27189 -5651 -27155
rect -5651 -27189 -5635 -27155
rect -5597 -27189 -5583 -27155
rect -5583 -27189 -5563 -27155
rect -5525 -27189 -5515 -27155
rect -5515 -27189 -5491 -27155
rect -5453 -27189 -5447 -27155
rect -5447 -27189 -5419 -27155
rect -5381 -27189 -5379 -27155
rect -5379 -27189 -5347 -27155
rect -5309 -27189 -5277 -27155
rect -5277 -27189 -5275 -27155
rect -5237 -27189 -5209 -27155
rect -5209 -27189 -5203 -27155
rect -5165 -27189 -5141 -27155
rect -5141 -27189 -5131 -27155
rect -5093 -27189 -5073 -27155
rect -5073 -27189 -5059 -27155
rect -5021 -27189 -5005 -27155
rect -5005 -27189 -4987 -27155
rect -4949 -27189 -4937 -27155
rect -4937 -27189 -4915 -27155
rect -4877 -27189 -4869 -27155
rect -4869 -27189 -4843 -27155
rect -4805 -27189 -4801 -27155
rect -4801 -27189 -4771 -27155
rect -4733 -27189 -4699 -27155
rect -4661 -27189 -4631 -27155
rect -4631 -27189 -4627 -27155
rect -4589 -27189 -4563 -27155
rect -4563 -27189 -4555 -27155
rect -4517 -27189 -4495 -27155
rect -4495 -27189 -4483 -27155
rect -4445 -27189 -4427 -27155
rect -4427 -27189 -4411 -27155
rect -4373 -27189 -4359 -27155
rect -4359 -27189 -4339 -27155
rect -4301 -27189 -4291 -27155
rect -4291 -27189 -4267 -27155
rect -4229 -27189 -4223 -27155
rect -4223 -27189 -4195 -27155
rect -4157 -27189 -4155 -27155
rect -4155 -27189 -4123 -27155
rect -4085 -27189 -4053 -27155
rect -4053 -27189 -4051 -27155
rect -4013 -27189 -3985 -27155
rect -3985 -27189 -3979 -27155
rect -3941 -27189 -3917 -27155
rect -3917 -27189 -3907 -27155
rect -3869 -27189 -3849 -27155
rect -3849 -27189 -3835 -27155
rect -3797 -27189 -3781 -27155
rect -3781 -27189 -3763 -27155
rect -3725 -27189 -3713 -27155
rect -3713 -27189 -3691 -27155
rect -3653 -27189 -3645 -27155
rect -3645 -27189 -3619 -27155
rect -3581 -27189 -3577 -27155
rect -3577 -27189 -3547 -27155
rect -3509 -27189 -3475 -27155
rect -3437 -27189 -3407 -27155
rect -3407 -27189 -3403 -27155
rect -3365 -27189 -3339 -27155
rect -3339 -27189 -3331 -27155
rect -3293 -27189 -3271 -27155
rect -3271 -27189 -3259 -27155
rect -3221 -27189 -3203 -27155
rect -3203 -27189 -3187 -27155
rect -3149 -27189 -3135 -27155
rect -3135 -27189 -3115 -27155
rect -3077 -27189 -3067 -27155
rect -3067 -27189 -3043 -27155
rect -3005 -27189 -2999 -27155
rect -2999 -27189 -2971 -27155
rect -2933 -27189 -2931 -27155
rect -2931 -27189 -2899 -27155
rect -2861 -27189 -2829 -27155
rect -2829 -27189 -2827 -27155
rect -2789 -27189 -2761 -27155
rect -2761 -27189 -2755 -27155
rect -2717 -27189 -2693 -27155
rect -2693 -27189 -2683 -27155
rect -2645 -27189 -2625 -27155
rect -2625 -27189 -2611 -27155
rect -2573 -27189 -2557 -27155
rect -2557 -27189 -2539 -27155
rect -2501 -27189 -2489 -27155
rect -2489 -27189 -2467 -27155
rect -2429 -27189 -2421 -27155
rect -2421 -27189 -2395 -27155
rect -2357 -27189 -2353 -27155
rect -2353 -27189 -2323 -27155
rect -2285 -27189 -2251 -27155
rect -2213 -27189 -2183 -27155
rect -2183 -27189 -2179 -27155
rect -2141 -27189 -2115 -27155
rect -2115 -27189 -2107 -27155
rect -2069 -27189 -2047 -27155
rect -2047 -27189 -2035 -27155
rect -1997 -27189 -1979 -27155
rect -1979 -27189 -1963 -27155
rect -1925 -27189 -1911 -27155
rect -1911 -27189 -1891 -27155
rect -1853 -27189 -1843 -27155
rect -1843 -27189 -1819 -27155
rect -1781 -27189 -1775 -27155
rect -1775 -27189 -1747 -27155
rect -1709 -27189 -1707 -27155
rect -1707 -27189 -1675 -27155
rect -1637 -27189 -1605 -27155
rect -1605 -27189 -1603 -27155
rect -1565 -27189 -1537 -27155
rect -1537 -27189 -1531 -27155
rect -1493 -27189 -1469 -27155
rect -1469 -27189 -1459 -27155
rect -1421 -27189 -1401 -27155
rect -1401 -27189 -1387 -27155
rect -1349 -27189 -1333 -27155
rect -1333 -27189 -1315 -27155
rect -1277 -27189 -1265 -27155
rect -1265 -27189 -1243 -27155
rect -1205 -27189 -1197 -27155
rect -1197 -27189 -1171 -27155
rect -1133 -27189 -1129 -27155
rect -1129 -27189 -1099 -27155
rect -1061 -27189 -1027 -27155
rect -989 -27189 -959 -27155
rect -959 -27189 -955 -27155
rect -917 -27189 -891 -27155
rect -891 -27189 -883 -27155
rect -845 -27189 -823 -27155
rect -823 -27189 -811 -27155
rect -773 -27189 -755 -27155
rect -755 -27189 -739 -27155
rect -701 -27189 -687 -27155
rect -687 -27189 -667 -27155
rect -629 -27189 -619 -27155
rect -619 -27189 -595 -27155
rect -557 -27189 -551 -27155
rect -551 -27189 -523 -27155
rect -485 -27189 -483 -27155
rect -483 -27189 -451 -27155
rect -413 -27189 -381 -27155
rect -381 -27189 -379 -27155
rect -341 -27189 -313 -27155
rect -313 -27189 -307 -27155
rect -269 -27189 -245 -27155
rect -245 -27189 -235 -27155
rect -197 -27189 -177 -27155
rect -177 -27189 -163 -27155
rect -125 -27189 -109 -27155
rect -109 -27189 -91 -27155
rect -53 -27189 -41 -27155
rect -41 -27189 -19 -27155
rect 19 -27189 27 -27155
rect 27 -27189 53 -27155
rect 91 -27189 95 -27155
rect 95 -27189 125 -27155
rect 163 -27189 197 -27155
rect 235 -27189 265 -27155
rect 265 -27189 269 -27155
rect 307 -27189 333 -27155
rect 333 -27189 341 -27155
rect 379 -27189 401 -27155
rect 401 -27189 413 -27155
rect 451 -27189 469 -27155
rect 469 -27189 485 -27155
rect 523 -27189 537 -27155
rect 537 -27189 557 -27155
rect 595 -27189 605 -27155
rect 605 -27189 629 -27155
rect 667 -27189 673 -27155
rect 673 -27189 701 -27155
rect 739 -27189 741 -27155
rect 741 -27189 773 -27155
rect 811 -27189 843 -27155
rect 843 -27189 845 -27155
rect 883 -27189 911 -27155
rect 911 -27189 917 -27155
rect 955 -27189 979 -27155
rect 979 -27189 989 -27155
rect 1027 -27189 1047 -27155
rect 1047 -27189 1061 -27155
rect 1099 -27189 1115 -27155
rect 1115 -27189 1133 -27155
rect 1171 -27189 1183 -27155
rect 1183 -27189 1205 -27155
rect 1243 -27189 1251 -27155
rect 1251 -27189 1277 -27155
rect 1315 -27189 1319 -27155
rect 1319 -27189 1349 -27155
rect 1387 -27189 1421 -27155
rect 1459 -27189 1489 -27155
rect 1489 -27189 1493 -27155
rect 1531 -27189 1557 -27155
rect 1557 -27189 1565 -27155
rect 1603 -27189 1625 -27155
rect 1625 -27189 1637 -27155
rect 1675 -27189 1693 -27155
rect 1693 -27189 1709 -27155
rect 1747 -27189 1761 -27155
rect 1761 -27189 1781 -27155
rect 1819 -27189 1829 -27155
rect 1829 -27189 1853 -27155
rect 1891 -27189 1897 -27155
rect 1897 -27189 1925 -27155
rect 1963 -27189 1965 -27155
rect 1965 -27189 1997 -27155
rect 2035 -27189 2067 -27155
rect 2067 -27189 2069 -27155
rect 2107 -27189 2135 -27155
rect 2135 -27189 2141 -27155
rect 2179 -27189 2203 -27155
rect 2203 -27189 2213 -27155
rect 2251 -27189 2271 -27155
rect 2271 -27189 2285 -27155
rect 2323 -27189 2339 -27155
rect 2339 -27189 2357 -27155
rect 2395 -27189 2407 -27155
rect 2407 -27189 2429 -27155
rect 2467 -27189 2475 -27155
rect 2475 -27189 2501 -27155
rect 2539 -27189 2543 -27155
rect 2543 -27189 2573 -27155
rect 2611 -27189 2645 -27155
rect 2683 -27189 2713 -27155
rect 2713 -27189 2717 -27155
rect 2755 -27189 2781 -27155
rect 2781 -27189 2789 -27155
rect 2827 -27189 2849 -27155
rect 2849 -27189 2861 -27155
rect 2899 -27189 2917 -27155
rect 2917 -27189 2933 -27155
rect 2971 -27189 2985 -27155
rect 2985 -27189 3005 -27155
rect 3043 -27189 3053 -27155
rect 3053 -27189 3077 -27155
rect 3115 -27189 3121 -27155
rect 3121 -27189 3149 -27155
rect 3187 -27189 3189 -27155
rect 3189 -27189 3221 -27155
rect 3259 -27189 3291 -27155
rect 3291 -27189 3293 -27155
rect 3331 -27189 3359 -27155
rect 3359 -27189 3365 -27155
rect 3403 -27189 3427 -27155
rect 3427 -27189 3437 -27155
rect 3475 -27189 3495 -27155
rect 3495 -27189 3509 -27155
rect 3547 -27189 3563 -27155
rect 3563 -27189 3581 -27155
rect 3619 -27189 3631 -27155
rect 3631 -27189 3653 -27155
rect 3691 -27189 3699 -27155
rect 3699 -27189 3725 -27155
rect 3763 -27189 3767 -27155
rect 3767 -27189 3797 -27155
rect 3835 -27189 3869 -27155
rect 3907 -27189 3937 -27155
rect 3937 -27189 3941 -27155
rect 3979 -27189 4005 -27155
rect 4005 -27189 4013 -27155
rect 4051 -27189 4073 -27155
rect 4073 -27189 4085 -27155
rect 4123 -27189 4141 -27155
rect 4141 -27189 4157 -27155
rect 4195 -27189 4209 -27155
rect 4209 -27189 4229 -27155
rect 4267 -27189 4277 -27155
rect 4277 -27189 4301 -27155
rect 4339 -27189 4345 -27155
rect 4345 -27189 4373 -27155
rect 4411 -27189 4413 -27155
rect 4413 -27189 4445 -27155
rect 4483 -27189 4515 -27155
rect 4515 -27189 4517 -27155
rect 4555 -27189 4583 -27155
rect 4583 -27189 4589 -27155
rect 4627 -27189 4651 -27155
rect 4651 -27189 4661 -27155
rect 4699 -27189 4719 -27155
rect 4719 -27189 4733 -27155
rect 4771 -27189 4787 -27155
rect 4787 -27189 4805 -27155
rect 4843 -27189 4855 -27155
rect 4855 -27189 4877 -27155
rect 4915 -27189 4923 -27155
rect 4923 -27189 4949 -27155
rect 4987 -27189 4991 -27155
rect 4991 -27189 5021 -27155
rect 5059 -27189 5093 -27155
rect 5131 -27189 5161 -27155
rect 5161 -27189 5165 -27155
rect 5203 -27189 5229 -27155
rect 5229 -27189 5237 -27155
rect 5275 -27189 5297 -27155
rect 5297 -27189 5309 -27155
rect 5347 -27189 5365 -27155
rect 5365 -27189 5381 -27155
rect 5419 -27189 5433 -27155
rect 5433 -27189 5453 -27155
rect 5491 -27189 5501 -27155
rect 5501 -27189 5525 -27155
rect 5563 -27189 5569 -27155
rect 5569 -27189 5597 -27155
rect 5635 -27189 5637 -27155
rect 5637 -27189 5669 -27155
rect 5707 -27189 5739 -27155
rect 5739 -27189 5741 -27155
rect 5779 -27189 5807 -27155
rect 5807 -27189 5813 -27155
rect 5851 -27189 5875 -27155
rect 5875 -27189 5885 -27155
rect 5923 -27189 5943 -27155
rect 5943 -27189 5957 -27155
rect 5995 -27189 6011 -27155
rect 6011 -27189 6029 -27155
rect 6067 -27189 6079 -27155
rect 6079 -27189 6101 -27155
rect 6139 -27189 6147 -27155
rect 6147 -27189 6173 -27155
rect 6211 -27189 6215 -27155
rect 6215 -27189 6245 -27155
rect 6283 -27189 6317 -27155
rect 6355 -27189 6385 -27155
rect 6385 -27189 6389 -27155
rect 6427 -27189 6453 -27155
rect 6453 -27189 6461 -27155
rect 6499 -27189 6521 -27155
rect 6521 -27189 6533 -27155
rect 6571 -27189 6589 -27155
rect 6589 -27189 6605 -27155
rect 6643 -27189 6657 -27155
rect 6657 -27189 6677 -27155
rect 6715 -27189 6725 -27155
rect 6725 -27189 6749 -27155
rect 6787 -27189 6793 -27155
rect 6793 -27189 6821 -27155
rect 6859 -27189 6861 -27155
rect 6861 -27189 6893 -27155
rect 6931 -27189 6963 -27155
rect 6963 -27189 6965 -27155
rect 7003 -27189 7031 -27155
rect 7031 -27189 7037 -27155
rect 7075 -27189 7099 -27155
rect 7099 -27189 7109 -27155
rect 7147 -27189 7167 -27155
rect 7167 -27189 7181 -27155
rect 7219 -27189 7235 -27155
rect 7235 -27189 7253 -27155
rect 7291 -27189 7303 -27155
rect 7303 -27189 7325 -27155
rect 7363 -27189 7371 -27155
rect 7371 -27189 7397 -27155
rect 7435 -27189 7439 -27155
rect 7439 -27189 7469 -27155
rect 7507 -27189 7541 -27155
rect 7579 -27189 7609 -27155
rect 7609 -27189 7613 -27155
rect 7651 -27189 7677 -27155
rect 7677 -27189 7685 -27155
rect 7723 -27189 7745 -27155
rect 7745 -27189 7757 -27155
rect 7795 -27189 7813 -27155
rect 7813 -27189 7829 -27155
rect 7867 -27189 7881 -27155
rect 7881 -27189 7901 -27155
rect 7939 -27189 7949 -27155
rect 7949 -27189 7973 -27155
rect 8011 -27189 8017 -27155
rect 8017 -27189 8045 -27155
rect 8083 -27189 8085 -27155
rect 8085 -27189 8117 -27155
rect 8155 -27189 8187 -27155
rect 8187 -27189 8189 -27155
rect 8227 -27189 8255 -27155
rect 8255 -27189 8261 -27155
rect 8299 -27189 8323 -27155
rect 8323 -27189 8333 -27155
rect 8371 -27189 8391 -27155
rect 8391 -27189 8405 -27155
rect 8443 -27189 8459 -27155
rect 8459 -27189 8477 -27155
rect 8515 -27189 8527 -27155
rect 8527 -27189 8549 -27155
rect 8587 -27189 8595 -27155
rect 8595 -27189 8621 -27155
rect 8659 -27189 8663 -27155
rect 8663 -27189 8693 -27155
rect 8731 -27189 8765 -27155
rect 8803 -27189 8833 -27155
rect 8833 -27189 8837 -27155
rect 8875 -27189 8901 -27155
rect 8901 -27189 8909 -27155
rect 8947 -27189 8969 -27155
rect 8969 -27189 8981 -27155
rect 9019 -27189 9037 -27155
rect 9037 -27189 9053 -27155
rect 9091 -27189 9105 -27155
rect 9105 -27189 9125 -27155
rect 9163 -27189 9173 -27155
rect 9173 -27189 9197 -27155
rect 9235 -27189 9241 -27155
rect 9241 -27189 9269 -27155
rect 9307 -27189 9309 -27155
rect 9309 -27189 9341 -27155
rect 9379 -27189 9411 -27155
rect 9411 -27189 9413 -27155
rect 9451 -27189 9479 -27155
rect 9479 -27189 9485 -27155
rect 9523 -27189 9547 -27155
rect 9547 -27189 9557 -27155
rect 9595 -27189 9615 -27155
rect 9615 -27189 9629 -27155
rect 9667 -27189 9683 -27155
rect 9683 -27189 9701 -27155
rect 9739 -27189 9751 -27155
rect 9751 -27189 9773 -27155
rect 9811 -27189 9819 -27155
rect 9819 -27189 9845 -27155
rect 9883 -27189 9887 -27155
rect 9887 -27189 9917 -27155
rect 9955 -27189 9989 -27155
rect 10027 -27189 10057 -27155
rect 10057 -27189 10061 -27155
rect 10099 -27189 10125 -27155
rect 10125 -27189 10133 -27155
rect 10171 -27189 10193 -27155
rect 10193 -27189 10205 -27155
rect 10243 -27189 10261 -27155
rect 10261 -27189 10277 -27155
rect 10315 -27189 10329 -27155
rect 10329 -27189 10349 -27155
rect 10387 -27189 10397 -27155
rect 10397 -27189 10421 -27155
rect 10459 -27189 10465 -27155
rect 10465 -27189 10493 -27155
rect 10531 -27189 10533 -27155
rect 10533 -27189 10565 -27155
rect 10603 -27189 10635 -27155
rect 10635 -27189 10637 -27155
rect 10675 -27189 10703 -27155
rect 10703 -27189 10709 -27155
rect 10747 -27189 10771 -27155
rect 10771 -27189 10781 -27155
rect 10819 -27189 10839 -27155
rect 10839 -27189 10853 -27155
rect 10891 -27189 10907 -27155
rect 10907 -27189 10925 -27155
rect 10963 -27189 10975 -27155
rect 10975 -27189 10997 -27155
rect 11035 -27189 11043 -27155
rect 11043 -27189 11069 -27155
rect 11107 -27189 11111 -27155
rect 11111 -27189 11141 -27155
rect 11179 -27189 11213 -27155
rect 11251 -27189 11281 -27155
rect 11281 -27189 11285 -27155
rect 11323 -27189 11349 -27155
rect 11349 -27189 11357 -27155
rect 11395 -27189 11417 -27155
rect 11417 -27189 11429 -27155
rect 11467 -27189 11485 -27155
rect 11485 -27189 11501 -27155
rect 11539 -27189 11553 -27155
rect 11553 -27189 11573 -27155
rect 11611 -27189 11621 -27155
rect 11621 -27189 11645 -27155
rect 11683 -27189 11689 -27155
rect 11689 -27189 11717 -27155
rect 11755 -27189 11757 -27155
rect 11757 -27189 11789 -27155
rect 11827 -27189 11859 -27155
rect 11859 -27189 11861 -27155
rect 11899 -27189 11927 -27155
rect 11927 -27189 11933 -27155
rect 11971 -27189 11995 -27155
rect 11995 -27189 12005 -27155
rect 12043 -27189 12063 -27155
rect 12063 -27189 12077 -27155
rect 12115 -27189 12131 -27155
rect 12131 -27189 12149 -27155
rect 12187 -27189 12199 -27155
rect 12199 -27189 12221 -27155
rect 12259 -27189 12267 -27155
rect 12267 -27189 12293 -27155
rect 12331 -27189 12335 -27155
rect 12335 -27189 12365 -27155
rect 12403 -27189 12437 -27155
rect 12475 -27189 12505 -27155
rect 12505 -27189 12509 -27155
rect 12547 -27189 12573 -27155
rect 12573 -27189 12581 -27155
rect 12619 -27189 12641 -27155
rect 12641 -27189 12653 -27155
rect 12691 -27189 12709 -27155
rect 12709 -27189 12725 -27155
rect 12763 -27189 12777 -27155
rect 12777 -27189 12797 -27155
rect 12835 -27189 12845 -27155
rect 12845 -27189 12869 -27155
rect 12907 -27189 12913 -27155
rect 12913 -27189 12941 -27155
rect 12979 -27189 12981 -27155
rect 12981 -27189 13013 -27155
rect 13051 -27189 13083 -27155
rect 13083 -27189 13085 -27155
rect 13123 -27189 13151 -27155
rect 13151 -27189 13157 -27155
rect 13195 -27189 13219 -27155
rect 13219 -27189 13229 -27155
rect 13267 -27189 13287 -27155
rect 13287 -27189 13301 -27155
rect 13339 -27189 13355 -27155
rect 13355 -27189 13373 -27155
rect 13411 -27189 13423 -27155
rect 13423 -27189 13445 -27155
rect 13483 -27189 13491 -27155
rect 13491 -27189 13517 -27155
rect 13555 -27189 13559 -27155
rect 13559 -27189 13589 -27155
rect 13627 -27189 13661 -27155
rect 13699 -27189 13729 -27155
rect 13729 -27189 13733 -27155
rect 13771 -27189 13797 -27155
rect 13797 -27189 13805 -27155
rect 13843 -27189 13865 -27155
rect 13865 -27189 13877 -27155
rect 13915 -27189 13933 -27155
rect 13933 -27189 13949 -27155
rect 13987 -27189 14001 -27155
rect 14001 -27189 14021 -27155
rect 14059 -27189 14069 -27155
rect 14069 -27189 14093 -27155
rect 14131 -27189 14137 -27155
rect 14137 -27189 14165 -27155
rect 14203 -27189 14205 -27155
rect 14205 -27189 14237 -27155
rect 14275 -27189 14307 -27155
rect 14307 -27189 14309 -27155
rect 14347 -27189 14375 -27155
rect 14375 -27189 14381 -27155
rect 14419 -27189 14443 -27155
rect 14443 -27189 14453 -27155
rect 14491 -27189 14511 -27155
rect 14511 -27189 14525 -27155
rect 14563 -27189 14579 -27155
rect 14579 -27189 14597 -27155
rect 14635 -27189 14647 -27155
rect 14647 -27189 14669 -27155
rect 14707 -27189 14715 -27155
rect 14715 -27189 14741 -27155
rect 14779 -27189 14783 -27155
rect 14783 -27189 14813 -27155
rect 14851 -27189 14885 -27155
rect 14923 -27189 14953 -27155
rect 14953 -27189 14957 -27155
rect 14995 -27189 15021 -27155
rect 15021 -27189 15029 -27155
rect 15067 -27189 15089 -27155
rect 15089 -27189 15101 -27155
rect 15139 -27189 15157 -27155
rect 15157 -27189 15173 -27155
rect 15211 -27189 15225 -27155
rect 15225 -27189 15245 -27155
rect 15283 -27189 15293 -27155
rect 15293 -27189 15317 -27155
rect 15355 -27189 15361 -27155
rect 15361 -27189 15389 -27155
rect 15427 -27189 15429 -27155
rect 15429 -27189 15461 -27155
rect 15499 -27189 15531 -27155
rect 15531 -27189 15533 -27155
rect 15571 -27189 15599 -27155
rect 15599 -27189 15605 -27155
rect 15643 -27189 15667 -27155
rect 15667 -27189 15677 -27155
rect 15715 -27189 15735 -27155
rect 15735 -27189 15749 -27155
rect 15787 -27189 15803 -27155
rect 15803 -27189 15821 -27155
rect 15859 -27189 15871 -27155
rect 15871 -27189 15893 -27155
rect 15931 -27189 15939 -27155
rect 15939 -27189 15965 -27155
rect 16003 -27189 16007 -27155
rect 16007 -27189 16037 -27155
rect 16075 -27189 16109 -27155
rect 16147 -27189 16177 -27155
rect 16177 -27189 16181 -27155
rect 16219 -27189 16245 -27155
rect 16245 -27189 16253 -27155
rect 16291 -27189 16313 -27155
rect 16313 -27189 16325 -27155
rect 16363 -27189 16381 -27155
rect 16381 -27189 16397 -27155
rect 16435 -27189 16449 -27155
rect 16449 -27189 16469 -27155
rect 16507 -27189 16517 -27155
rect 16517 -27189 16541 -27155
rect 16579 -27189 16585 -27155
rect 16585 -27189 16613 -27155
rect 16651 -27189 16653 -27155
rect 16653 -27189 16685 -27155
rect 16723 -27189 16755 -27155
rect 16755 -27189 16757 -27155
rect 16795 -27189 16823 -27155
rect 16823 -27189 16829 -27155
rect 16867 -27189 16891 -27155
rect 16891 -27189 16901 -27155
rect 16939 -27189 16959 -27155
rect 16959 -27189 16973 -27155
rect 17011 -27189 17027 -27155
rect 17027 -27189 17045 -27155
rect 17083 -27189 17095 -27155
rect 17095 -27189 17117 -27155
rect 17155 -27189 17163 -27155
rect 17163 -27189 17189 -27155
rect 17227 -27189 17231 -27155
rect 17231 -27189 17261 -27155
rect 17299 -27189 17333 -27155
rect 17371 -27189 17401 -27155
rect 17401 -27189 17405 -27155
rect 17443 -27189 17469 -27155
rect 17469 -27189 17477 -27155
rect 17515 -27189 17537 -27155
rect 17537 -27189 17549 -27155
rect 17587 -27189 17605 -27155
rect 17605 -27189 17621 -27155
rect 17659 -27189 17673 -27155
rect 17673 -27189 17693 -27155
rect 17731 -27189 17741 -27155
rect 17741 -27189 17765 -27155
rect 17803 -27189 17809 -27155
rect 17809 -27189 17837 -27155
rect 17875 -27189 17877 -27155
rect 17877 -27189 17909 -27155
rect 17947 -27189 17979 -27155
rect 17979 -27189 17981 -27155
rect 18019 -27189 18047 -27155
rect 18047 -27189 18053 -27155
rect 18091 -27189 18115 -27155
rect 18115 -27189 18125 -27155
rect 18163 -27189 18183 -27155
rect 18183 -27189 18197 -27155
rect 18235 -27189 18251 -27155
rect 18251 -27189 18269 -27155
rect 18307 -27189 18319 -27155
rect 18319 -27189 18341 -27155
rect 18379 -27189 18387 -27155
rect 18387 -27189 18413 -27155
rect 18451 -27189 18455 -27155
rect 18455 -27189 18485 -27155
rect 18523 -27189 18557 -27155
rect 18595 -27189 18625 -27155
rect 18625 -27189 18629 -27155
rect 18667 -27189 18693 -27155
rect 18693 -27189 18701 -27155
rect 18739 -27189 18761 -27155
rect 18761 -27189 18773 -27155
rect 18811 -27189 18829 -27155
rect 18829 -27189 18845 -27155
rect 18883 -27189 18897 -27155
rect 18897 -27189 18917 -27155
rect 18955 -27189 18965 -27155
rect 18965 -27189 18989 -27155
rect 19027 -27189 19033 -27155
rect 19033 -27189 19061 -27155
rect 19099 -27189 19101 -27155
rect 19101 -27189 19133 -27155
rect 19171 -27189 19203 -27155
rect 19203 -27189 19205 -27155
rect 19243 -27189 19271 -27155
rect 19271 -27189 19277 -27155
rect 19315 -27189 19339 -27155
rect 19339 -27189 19349 -27155
rect 19387 -27189 19407 -27155
rect 19407 -27189 19421 -27155
rect 19459 -27189 19475 -27155
rect 19475 -27189 19493 -27155
rect 19531 -27189 19543 -27155
rect 19543 -27189 19565 -27155
rect 19603 -27189 19611 -27155
rect 19611 -27189 19637 -27155
rect 19675 -27189 19679 -27155
rect 19679 -27189 19709 -27155
rect 19747 -27189 19781 -27155
rect 19819 -27189 19849 -27155
rect 19849 -27189 19853 -27155
rect 19891 -27189 19917 -27155
rect 19917 -27189 19925 -27155
rect 19963 -27189 19985 -27155
rect 19985 -27189 19997 -27155
rect 20035 -27189 20053 -27155
rect 20053 -27189 20069 -27155
rect 20107 -27189 20121 -27155
rect 20121 -27189 20141 -27155
rect 20179 -27189 20189 -27155
rect 20189 -27189 20213 -27155
rect 20251 -27189 20257 -27155
rect 20257 -27189 20285 -27155
rect 20323 -27189 20325 -27155
rect 20325 -27189 20357 -27155
rect 20395 -27189 20427 -27155
rect 20427 -27189 20429 -27155
rect 20467 -27189 20495 -27155
rect 20495 -27189 20501 -27155
rect 20539 -27189 20563 -27155
rect 20563 -27189 20573 -27155
rect 20611 -27189 20631 -27155
rect 20631 -27189 20645 -27155
rect 20683 -27189 20699 -27155
rect 20699 -27189 20717 -27155
rect 20755 -27189 20767 -27155
rect 20767 -27189 20789 -27155
rect 20827 -27189 20835 -27155
rect 20835 -27189 20861 -27155
rect 20899 -27189 20903 -27155
rect 20903 -27189 20933 -27155
rect 20971 -27189 21005 -27155
rect 21043 -27189 21073 -27155
rect 21073 -27189 21077 -27155
rect 21115 -27189 21141 -27155
rect 21141 -27189 21149 -27155
rect 21187 -27189 21209 -27155
rect 21209 -27189 21221 -27155
rect 21259 -27189 21277 -27155
rect 21277 -27189 21293 -27155
rect 21331 -27189 21345 -27155
rect 21345 -27189 21365 -27155
rect 21403 -27189 21413 -27155
rect 21413 -27189 21437 -27155
rect 21475 -27189 21481 -27155
rect 21481 -27189 21509 -27155
rect 21547 -27189 21549 -27155
rect 21549 -27189 21581 -27155
rect 21619 -27189 21651 -27155
rect 21651 -27189 21653 -27155
rect 21691 -27189 21719 -27155
rect 21719 -27189 21725 -27155
rect 21763 -27189 21787 -27155
rect 21787 -27189 21797 -27155
rect 21835 -27189 21855 -27155
rect 21855 -27189 21869 -27155
rect 21907 -27189 21923 -27155
rect 21923 -27189 21941 -27155
rect 21979 -27189 21991 -27155
rect 21991 -27189 22013 -27155
rect 22051 -27189 22059 -27155
rect 22059 -27189 22085 -27155
rect 22123 -27189 22127 -27155
rect 22127 -27189 22157 -27155
rect 22195 -27189 22229 -27155
rect 22267 -27189 22297 -27155
rect 22297 -27189 22301 -27155
rect 22339 -27189 22365 -27155
rect 22365 -27189 22373 -27155
rect 22411 -27189 22433 -27155
rect 22433 -27189 22445 -27155
rect 22483 -27189 22501 -27155
rect 22501 -27189 22517 -27155
rect 22555 -27189 22569 -27155
rect 22569 -27189 22589 -27155
rect 22627 -27189 22637 -27155
rect 22637 -27189 22661 -27155
rect 22699 -27189 22705 -27155
rect 22705 -27189 22733 -27155
rect 22771 -27189 22773 -27155
rect 22773 -27189 22805 -27155
rect 22843 -27189 22875 -27155
rect 22875 -27189 22877 -27155
rect 22915 -27189 22943 -27155
rect 22943 -27189 22949 -27155
rect 22987 -27189 23011 -27155
rect 23011 -27189 23021 -27155
rect 23059 -27189 23079 -27155
rect 23079 -27189 23093 -27155
rect 23131 -27189 23147 -27155
rect 23147 -27189 23165 -27155
rect 23203 -27189 23215 -27155
rect 23215 -27189 23237 -27155
rect 23275 -27189 23283 -27155
rect 23283 -27189 23309 -27155
rect 23347 -27189 23351 -27155
rect 23351 -27189 23381 -27155
rect 23419 -27189 23453 -27155
rect 23491 -27189 23521 -27155
rect 23521 -27189 23525 -27155
rect 23563 -27189 23589 -27155
rect 23589 -27189 23597 -27155
rect 23635 -27189 23657 -27155
rect 23657 -27189 23669 -27155
rect 23707 -27189 23725 -27155
rect 23725 -27189 23741 -27155
rect 23779 -27189 23793 -27155
rect 23793 -27189 23813 -27155
rect 23851 -27189 23861 -27155
rect 23861 -27189 23885 -27155
rect 23923 -27189 23929 -27155
rect 23929 -27189 23957 -27155
rect 23995 -27189 23997 -27155
rect 23997 -27189 24029 -27155
rect 24067 -27189 24099 -27155
rect 24099 -27189 24101 -27155
rect 24139 -27189 24167 -27155
rect 24167 -27189 24173 -27155
rect 24211 -27189 24235 -27155
rect 24235 -27189 24245 -27155
rect 24283 -27189 24303 -27155
rect 24303 -27189 24317 -27155
rect 24355 -27189 24371 -27155
rect 24371 -27189 24389 -27155
rect 24427 -27189 24439 -27155
rect 24439 -27189 24461 -27155
rect 24499 -27189 24507 -27155
rect 24507 -27189 24533 -27155
rect 24571 -27189 24575 -27155
rect 24575 -27189 24605 -27155
rect 24643 -27189 24677 -27155
rect 24715 -27189 24745 -27155
rect 24745 -27189 24749 -27155
rect 24787 -27189 24821 -27155
<< metal1 >>
rect 372 4289 24828 4328
rect 372 4255 487 4289
rect 521 4255 559 4289
rect 593 4255 631 4289
rect 665 4255 703 4289
rect 737 4255 775 4289
rect 809 4255 847 4289
rect 881 4255 919 4289
rect 953 4255 991 4289
rect 1025 4255 1063 4289
rect 1097 4255 1135 4289
rect 1169 4255 1207 4289
rect 1241 4255 1279 4289
rect 1313 4255 1351 4289
rect 1385 4255 1423 4289
rect 1457 4255 1495 4289
rect 1529 4255 1567 4289
rect 1601 4255 1639 4289
rect 1673 4255 1711 4289
rect 1745 4255 1783 4289
rect 1817 4255 1855 4289
rect 1889 4255 1927 4289
rect 1961 4255 1999 4289
rect 2033 4255 2071 4289
rect 2105 4255 2143 4289
rect 2177 4255 2215 4289
rect 2249 4255 2287 4289
rect 2321 4255 2359 4289
rect 2393 4255 2431 4289
rect 2465 4255 2503 4289
rect 2537 4255 2575 4289
rect 2609 4255 2647 4289
rect 2681 4255 2719 4289
rect 2753 4255 2791 4289
rect 2825 4255 2863 4289
rect 2897 4255 2935 4289
rect 2969 4255 3007 4289
rect 3041 4255 3079 4289
rect 3113 4255 3151 4289
rect 3185 4255 3223 4289
rect 3257 4255 3295 4289
rect 3329 4255 3367 4289
rect 3401 4255 3439 4289
rect 3473 4255 3511 4289
rect 3545 4255 3583 4289
rect 3617 4255 3655 4289
rect 3689 4255 3727 4289
rect 3761 4255 3799 4289
rect 3833 4255 3871 4289
rect 3905 4255 3943 4289
rect 3977 4255 4015 4289
rect 4049 4255 4087 4289
rect 4121 4255 4159 4289
rect 4193 4255 4231 4289
rect 4265 4255 4303 4289
rect 4337 4255 4375 4289
rect 4409 4255 4447 4289
rect 4481 4255 4519 4289
rect 4553 4255 4591 4289
rect 4625 4255 4663 4289
rect 4697 4255 4735 4289
rect 4769 4255 4807 4289
rect 4841 4255 4879 4289
rect 4913 4255 4951 4289
rect 4985 4255 5023 4289
rect 5057 4255 5095 4289
rect 5129 4255 5167 4289
rect 5201 4255 5239 4289
rect 5273 4255 5311 4289
rect 5345 4255 5383 4289
rect 5417 4255 5455 4289
rect 5489 4255 5527 4289
rect 5561 4255 5599 4289
rect 5633 4255 5671 4289
rect 5705 4255 5743 4289
rect 5777 4255 5815 4289
rect 5849 4255 5887 4289
rect 5921 4255 5959 4289
rect 5993 4255 6031 4289
rect 6065 4255 6103 4289
rect 6137 4255 6175 4289
rect 6209 4255 6247 4289
rect 6281 4255 6319 4289
rect 6353 4255 6391 4289
rect 6425 4255 6463 4289
rect 6497 4255 6535 4289
rect 6569 4255 6607 4289
rect 6641 4255 6679 4289
rect 6713 4255 6751 4289
rect 6785 4255 6823 4289
rect 6857 4255 6895 4289
rect 6929 4255 6967 4289
rect 7001 4255 7039 4289
rect 7073 4255 7111 4289
rect 7145 4255 7183 4289
rect 7217 4255 7255 4289
rect 7289 4255 7327 4289
rect 7361 4255 7399 4289
rect 7433 4255 7471 4289
rect 7505 4255 7543 4289
rect 7577 4255 7615 4289
rect 7649 4255 7687 4289
rect 7721 4255 7759 4289
rect 7793 4255 7831 4289
rect 7865 4255 7903 4289
rect 7937 4255 7975 4289
rect 8009 4255 8047 4289
rect 8081 4255 8119 4289
rect 8153 4255 8191 4289
rect 8225 4255 8263 4289
rect 8297 4255 8335 4289
rect 8369 4255 8407 4289
rect 8441 4255 8479 4289
rect 8513 4255 8551 4289
rect 8585 4255 8623 4289
rect 8657 4255 8695 4289
rect 8729 4255 8767 4289
rect 8801 4255 8839 4289
rect 8873 4255 8911 4289
rect 8945 4255 8983 4289
rect 9017 4255 9055 4289
rect 9089 4255 9127 4289
rect 9161 4255 9199 4289
rect 9233 4255 9271 4289
rect 9305 4255 9343 4289
rect 9377 4255 9415 4289
rect 9449 4255 9487 4289
rect 9521 4255 9559 4289
rect 9593 4255 9631 4289
rect 9665 4255 9703 4289
rect 9737 4255 9775 4289
rect 9809 4255 9847 4289
rect 9881 4255 9919 4289
rect 9953 4255 9991 4289
rect 10025 4255 10063 4289
rect 10097 4255 10135 4289
rect 10169 4255 10207 4289
rect 10241 4255 10279 4289
rect 10313 4255 10351 4289
rect 10385 4255 10423 4289
rect 10457 4255 10495 4289
rect 10529 4255 10567 4289
rect 10601 4255 10639 4289
rect 10673 4255 10711 4289
rect 10745 4255 10783 4289
rect 10817 4255 10855 4289
rect 10889 4255 10927 4289
rect 10961 4255 10999 4289
rect 11033 4255 11071 4289
rect 11105 4255 11143 4289
rect 11177 4255 11215 4289
rect 11249 4255 11287 4289
rect 11321 4255 11359 4289
rect 11393 4255 11431 4289
rect 11465 4255 11503 4289
rect 11537 4255 11575 4289
rect 11609 4255 11647 4289
rect 11681 4255 11719 4289
rect 11753 4255 11791 4289
rect 11825 4255 11863 4289
rect 11897 4255 11935 4289
rect 11969 4255 12007 4289
rect 12041 4255 12079 4289
rect 12113 4255 12151 4289
rect 12185 4255 12223 4289
rect 12257 4255 12295 4289
rect 12329 4255 12367 4289
rect 12401 4255 12439 4289
rect 12473 4255 12511 4289
rect 12545 4255 12583 4289
rect 12617 4255 12655 4289
rect 12689 4255 12727 4289
rect 12761 4255 12799 4289
rect 12833 4255 12871 4289
rect 12905 4255 12943 4289
rect 12977 4255 13015 4289
rect 13049 4255 13087 4289
rect 13121 4255 13159 4289
rect 13193 4255 13231 4289
rect 13265 4255 13303 4289
rect 13337 4255 13375 4289
rect 13409 4255 13447 4289
rect 13481 4255 13519 4289
rect 13553 4255 13591 4289
rect 13625 4255 13663 4289
rect 13697 4255 13735 4289
rect 13769 4255 13807 4289
rect 13841 4255 13879 4289
rect 13913 4255 13951 4289
rect 13985 4255 14023 4289
rect 14057 4255 14095 4289
rect 14129 4255 14167 4289
rect 14201 4255 14239 4289
rect 14273 4255 14311 4289
rect 14345 4255 14383 4289
rect 14417 4255 14455 4289
rect 14489 4255 14527 4289
rect 14561 4255 14599 4289
rect 14633 4255 14671 4289
rect 14705 4255 14743 4289
rect 14777 4255 14815 4289
rect 14849 4255 14887 4289
rect 14921 4255 14959 4289
rect 14993 4255 15031 4289
rect 15065 4255 15103 4289
rect 15137 4255 15175 4289
rect 15209 4255 15247 4289
rect 15281 4255 15319 4289
rect 15353 4255 15391 4289
rect 15425 4255 15463 4289
rect 15497 4255 15535 4289
rect 15569 4255 15607 4289
rect 15641 4255 15679 4289
rect 15713 4255 15751 4289
rect 15785 4255 15823 4289
rect 15857 4255 15895 4289
rect 15929 4255 15967 4289
rect 16001 4255 16039 4289
rect 16073 4255 16111 4289
rect 16145 4255 16183 4289
rect 16217 4255 16255 4289
rect 16289 4255 16327 4289
rect 16361 4255 16399 4289
rect 16433 4255 16471 4289
rect 16505 4255 16543 4289
rect 16577 4255 16615 4289
rect 16649 4255 16687 4289
rect 16721 4255 16759 4289
rect 16793 4255 16831 4289
rect 16865 4255 16903 4289
rect 16937 4255 16975 4289
rect 17009 4255 17047 4289
rect 17081 4255 17119 4289
rect 17153 4255 17191 4289
rect 17225 4255 17263 4289
rect 17297 4255 17335 4289
rect 17369 4255 17407 4289
rect 17441 4255 17479 4289
rect 17513 4255 17551 4289
rect 17585 4255 17623 4289
rect 17657 4255 17695 4289
rect 17729 4255 17767 4289
rect 17801 4255 17839 4289
rect 17873 4255 17911 4289
rect 17945 4255 17983 4289
rect 18017 4255 18055 4289
rect 18089 4255 18127 4289
rect 18161 4255 18199 4289
rect 18233 4255 18271 4289
rect 18305 4255 18343 4289
rect 18377 4255 18415 4289
rect 18449 4255 18487 4289
rect 18521 4255 18559 4289
rect 18593 4255 18631 4289
rect 18665 4255 18703 4289
rect 18737 4255 18775 4289
rect 18809 4255 18847 4289
rect 18881 4255 18919 4289
rect 18953 4255 18991 4289
rect 19025 4255 19063 4289
rect 19097 4255 19135 4289
rect 19169 4255 19207 4289
rect 19241 4255 19279 4289
rect 19313 4255 19351 4289
rect 19385 4255 19423 4289
rect 19457 4255 19495 4289
rect 19529 4255 19567 4289
rect 19601 4255 19639 4289
rect 19673 4255 19711 4289
rect 19745 4255 19783 4289
rect 19817 4255 19855 4289
rect 19889 4255 19927 4289
rect 19961 4255 19999 4289
rect 20033 4255 20071 4289
rect 20105 4255 20143 4289
rect 20177 4255 20215 4289
rect 20249 4255 20287 4289
rect 20321 4255 20359 4289
rect 20393 4255 20431 4289
rect 20465 4255 20503 4289
rect 20537 4255 20575 4289
rect 20609 4255 20647 4289
rect 20681 4255 20719 4289
rect 20753 4255 20791 4289
rect 20825 4255 20863 4289
rect 20897 4255 20935 4289
rect 20969 4255 21007 4289
rect 21041 4255 21079 4289
rect 21113 4255 21151 4289
rect 21185 4255 21223 4289
rect 21257 4255 21295 4289
rect 21329 4255 21367 4289
rect 21401 4255 21439 4289
rect 21473 4255 21511 4289
rect 21545 4255 21583 4289
rect 21617 4255 21655 4289
rect 21689 4255 21727 4289
rect 21761 4255 21799 4289
rect 21833 4255 21871 4289
rect 21905 4255 21943 4289
rect 21977 4255 22015 4289
rect 22049 4255 22087 4289
rect 22121 4255 22159 4289
rect 22193 4255 22231 4289
rect 22265 4255 22303 4289
rect 22337 4255 22375 4289
rect 22409 4255 22447 4289
rect 22481 4255 22519 4289
rect 22553 4255 22591 4289
rect 22625 4255 22663 4289
rect 22697 4255 22735 4289
rect 22769 4255 22807 4289
rect 22841 4255 22879 4289
rect 22913 4255 22951 4289
rect 22985 4255 23023 4289
rect 23057 4255 23095 4289
rect 23129 4255 23167 4289
rect 23201 4255 23239 4289
rect 23273 4255 23311 4289
rect 23345 4255 23383 4289
rect 23417 4255 23455 4289
rect 23489 4255 23527 4289
rect 23561 4255 23599 4289
rect 23633 4255 23671 4289
rect 23705 4255 23743 4289
rect 23777 4255 23815 4289
rect 23849 4255 23887 4289
rect 23921 4255 23959 4289
rect 23993 4255 24031 4289
rect 24065 4255 24103 4289
rect 24137 4255 24175 4289
rect 24209 4255 24247 4289
rect 24281 4255 24319 4289
rect 24353 4255 24391 4289
rect 24425 4255 24463 4289
rect 24497 4255 24535 4289
rect 24569 4255 24607 4289
rect 24641 4255 24679 4289
rect 24713 4255 24828 4289
rect 372 4216 24828 4255
rect 372 4188 1094 4216
rect 372 3944 502 4188
rect 1066 3944 1094 4188
rect 372 3916 1094 3944
rect 24106 4188 24828 4216
rect 24106 3944 24134 4188
rect 24698 3944 24828 4188
rect 24106 3916 24828 3944
rect 372 3700 484 3916
rect 372 3666 411 3700
rect 445 3666 484 3700
rect 372 3628 484 3666
rect 372 3594 411 3628
rect 445 3594 484 3628
rect 3998 3817 20878 3866
rect 3998 3637 4075 3817
rect 20831 3637 20878 3817
rect 3998 3620 20878 3637
rect 3998 3598 4048 3620
rect 4108 3598 4484 3620
rect 4544 3598 4922 3620
rect 4982 3598 5356 3620
rect 5416 3600 20878 3620
rect 24716 3700 24828 3916
rect 24716 3666 24755 3700
rect 24789 3666 24828 3700
rect 24716 3628 24828 3666
rect 5416 3598 8352 3600
rect 372 3556 484 3594
rect 372 3522 411 3556
rect 445 3522 484 3556
rect 372 3484 484 3522
rect 372 3450 411 3484
rect 445 3450 484 3484
rect 372 3412 484 3450
rect 372 3378 411 3412
rect 445 3378 484 3412
rect 372 3340 484 3378
rect 372 3306 411 3340
rect 445 3306 484 3340
rect 372 3268 484 3306
rect 372 3234 411 3268
rect 445 3234 484 3268
rect 372 3196 484 3234
rect 372 3162 411 3196
rect 445 3162 484 3196
rect 372 3124 484 3162
rect 372 3090 411 3124
rect 445 3090 484 3124
rect 372 3052 484 3090
rect 372 3018 411 3052
rect 445 3018 484 3052
rect 372 2980 484 3018
rect 372 2946 411 2980
rect 445 2946 484 2980
rect 372 2908 484 2946
rect 372 2874 411 2908
rect 445 2874 484 2908
rect 372 2836 484 2874
rect 372 2802 411 2836
rect 445 2802 484 2836
rect 372 2764 484 2802
rect 372 2730 411 2764
rect 445 2730 484 2764
rect 372 2692 484 2730
rect 372 2658 411 2692
rect 445 2658 484 2692
rect 372 2620 484 2658
rect 372 2586 411 2620
rect 445 2586 484 2620
rect 372 2548 484 2586
rect 372 2514 411 2548
rect 445 2514 484 2548
rect 372 2476 484 2514
rect 372 2442 411 2476
rect 445 2442 484 2476
rect 372 2404 484 2442
rect 372 2370 411 2404
rect 445 2370 484 2404
rect 372 2332 484 2370
rect 372 2298 411 2332
rect 445 2298 484 2332
rect 372 2260 484 2298
rect 372 2226 411 2260
rect 445 2226 484 2260
rect 372 2188 484 2226
rect 372 2154 411 2188
rect 445 2154 484 2188
rect 372 2116 484 2154
rect 372 2082 411 2116
rect 445 2082 484 2116
rect 372 2044 484 2082
rect 372 2010 411 2044
rect 445 2010 484 2044
rect 372 1972 484 2010
rect 372 1938 411 1972
rect 445 1938 484 1972
rect 372 1900 484 1938
rect 8512 2124 8572 3600
rect 10548 2124 10608 3600
rect 11052 2124 11112 3600
rect 11560 2124 11620 3600
rect 12072 2124 12132 3600
rect 12586 2124 12646 3600
rect 14618 2124 14678 3600
rect 16658 2124 16718 3600
rect 17148 2124 17208 3600
rect 17668 2124 17728 3600
rect 18176 2124 18236 3600
rect 18690 2124 18750 3600
rect 20726 2124 20786 3600
rect 8512 2064 20786 2124
rect 372 1866 411 1900
rect 445 1866 484 1900
rect 372 1828 484 1866
rect 7980 1914 8052 1918
rect 7980 1862 7990 1914
rect 8042 1862 8052 1914
rect 7980 1858 8052 1862
rect 372 1794 411 1828
rect 445 1794 484 1828
rect 372 1756 484 1794
rect 372 1722 411 1756
rect 445 1722 484 1756
rect 372 1684 484 1722
rect 372 1650 411 1684
rect 445 1650 484 1684
rect 372 1612 484 1650
rect 372 1578 411 1612
rect 445 1578 484 1612
rect 372 1540 484 1578
rect 372 1506 411 1540
rect 445 1506 484 1540
rect 372 1468 484 1506
rect 372 1434 411 1468
rect 445 1434 484 1468
rect 372 1396 484 1434
rect 6474 1642 7552 1702
rect 6474 1422 6534 1642
rect 6978 1526 7038 1642
rect 7492 1436 7552 1642
rect 7986 1518 8046 1858
rect 8512 1672 8572 2064
rect 9062 1914 9134 1918
rect 9062 1862 9072 1914
rect 9124 1862 9134 1914
rect 9062 1858 9134 1862
rect 10020 1914 10092 1918
rect 10020 1862 10030 1914
rect 10082 1862 10092 1914
rect 10020 1858 10092 1862
rect 8506 1668 8578 1672
rect 8506 1616 8516 1668
rect 8568 1616 8578 1668
rect 8506 1612 8578 1616
rect 8512 1438 8572 1612
rect 9068 1516 9128 1858
rect 10026 1512 10086 1858
rect 10548 1672 10608 2064
rect 10542 1668 10614 1672
rect 10542 1616 10552 1668
rect 10604 1616 10614 1668
rect 10542 1612 10614 1616
rect 10548 1438 10608 1612
rect 11052 1518 11112 2064
rect 372 1362 411 1396
rect 445 1362 484 1396
rect 11560 1392 11620 2064
rect 12072 1518 12132 2064
rect 12586 1674 12646 2064
rect 13084 1914 13156 1918
rect 13084 1862 13094 1914
rect 13146 1862 13156 1914
rect 13084 1858 13156 1862
rect 14102 1914 14174 1918
rect 14102 1862 14112 1914
rect 14164 1862 14174 1914
rect 14102 1858 14174 1862
rect 12580 1670 12652 1674
rect 12580 1618 12590 1670
rect 12642 1618 12652 1670
rect 12580 1614 12652 1618
rect 12586 1422 12646 1614
rect 13090 1522 13150 1858
rect 14108 1516 14168 1858
rect 14618 1674 14678 2064
rect 15126 1914 15198 1918
rect 15126 1862 15136 1914
rect 15188 1862 15198 1914
rect 15126 1858 15198 1862
rect 16138 1914 16210 1918
rect 16138 1862 16148 1914
rect 16200 1862 16210 1914
rect 16138 1858 16210 1862
rect 14610 1670 14682 1674
rect 14610 1618 14620 1670
rect 14672 1618 14682 1670
rect 14610 1614 14682 1618
rect 14618 1422 14678 1614
rect 15132 1522 15192 1858
rect 16144 1522 16204 1858
rect 16658 1676 16718 2064
rect 16652 1672 16724 1676
rect 16652 1620 16662 1672
rect 16714 1620 16724 1672
rect 16652 1616 16724 1620
rect 16658 1424 16718 1616
rect 17148 1522 17208 2064
rect 17668 1676 17728 2064
rect 17662 1672 17734 1676
rect 17662 1620 17672 1672
rect 17724 1620 17734 1672
rect 17662 1616 17734 1620
rect 17668 1392 17728 1616
rect 18176 1512 18236 2064
rect 18690 1676 18750 2064
rect 19196 1914 19268 1918
rect 19196 1862 19206 1914
rect 19258 1862 19268 1914
rect 19196 1858 19268 1862
rect 20208 1914 20280 1918
rect 20208 1862 20218 1914
rect 20270 1862 20280 1914
rect 20208 1858 20280 1862
rect 18684 1672 18756 1676
rect 18684 1620 18694 1672
rect 18746 1620 18756 1672
rect 18684 1616 18756 1620
rect 18690 1434 18750 1616
rect 19202 1522 19262 1858
rect 20214 1522 20274 1858
rect 20726 1676 20786 2064
rect 24716 3594 24755 3628
rect 24789 3594 24828 3628
rect 24716 3556 24828 3594
rect 24716 3522 24755 3556
rect 24789 3522 24828 3556
rect 24716 3484 24828 3522
rect 24716 3450 24755 3484
rect 24789 3450 24828 3484
rect 24716 3412 24828 3450
rect 24716 3378 24755 3412
rect 24789 3378 24828 3412
rect 24716 3340 24828 3378
rect 24716 3306 24755 3340
rect 24789 3306 24828 3340
rect 24716 3268 24828 3306
rect 24716 3234 24755 3268
rect 24789 3234 24828 3268
rect 24716 3196 24828 3234
rect 24716 3162 24755 3196
rect 24789 3162 24828 3196
rect 24716 3124 24828 3162
rect 24716 3090 24755 3124
rect 24789 3090 24828 3124
rect 24716 3052 24828 3090
rect 24716 3018 24755 3052
rect 24789 3018 24828 3052
rect 24716 2980 24828 3018
rect 24716 2946 24755 2980
rect 24789 2946 24828 2980
rect 24716 2908 24828 2946
rect 24716 2874 24755 2908
rect 24789 2874 24828 2908
rect 24716 2836 24828 2874
rect 24716 2802 24755 2836
rect 24789 2802 24828 2836
rect 24716 2764 24828 2802
rect 24716 2730 24755 2764
rect 24789 2730 24828 2764
rect 24716 2692 24828 2730
rect 24716 2658 24755 2692
rect 24789 2658 24828 2692
rect 24716 2620 24828 2658
rect 24716 2586 24755 2620
rect 24789 2586 24828 2620
rect 24716 2548 24828 2586
rect 24716 2514 24755 2548
rect 24789 2514 24828 2548
rect 24716 2476 24828 2514
rect 24716 2442 24755 2476
rect 24789 2442 24828 2476
rect 24716 2404 24828 2442
rect 24716 2370 24755 2404
rect 24789 2370 24828 2404
rect 24716 2332 24828 2370
rect 24716 2298 24755 2332
rect 24789 2298 24828 2332
rect 24716 2260 24828 2298
rect 24716 2226 24755 2260
rect 24789 2226 24828 2260
rect 24716 2188 24828 2226
rect 24716 2154 24755 2188
rect 24789 2154 24828 2188
rect 24716 2116 24828 2154
rect 24716 2082 24755 2116
rect 24789 2082 24828 2116
rect 24716 2044 24828 2082
rect 24716 2010 24755 2044
rect 24789 2010 24828 2044
rect 24716 1972 24828 2010
rect 24716 1938 24755 1972
rect 24789 1938 24828 1972
rect 21226 1914 21298 1918
rect 21226 1862 21236 1914
rect 21288 1862 21298 1914
rect 21226 1858 21298 1862
rect 24716 1900 24828 1938
rect 24716 1866 24755 1900
rect 24789 1866 24828 1900
rect 20720 1672 20792 1676
rect 20720 1620 20730 1672
rect 20782 1620 20792 1672
rect 20720 1616 20792 1620
rect 20726 1430 20786 1616
rect 21232 1516 21292 1858
rect 24716 1828 24828 1866
rect 24716 1794 24755 1828
rect 24789 1794 24828 1828
rect 24716 1756 24828 1794
rect 24716 1722 24755 1756
rect 24789 1722 24828 1756
rect 24716 1684 24828 1722
rect 21746 1624 22826 1684
rect 21746 1432 21806 1624
rect 22248 1522 22308 1624
rect 22766 1416 22826 1624
rect 24716 1650 24755 1684
rect 24789 1650 24828 1684
rect 24716 1612 24828 1650
rect 24716 1578 24755 1612
rect 24789 1578 24828 1612
rect 24716 1540 24828 1578
rect 24716 1506 24755 1540
rect 24789 1506 24828 1540
rect 24716 1468 24828 1506
rect 24716 1434 24755 1468
rect 24789 1434 24828 1468
rect 24716 1396 24828 1434
rect 372 1324 484 1362
rect 372 1290 411 1324
rect 445 1290 484 1324
rect 372 1252 484 1290
rect 372 1218 411 1252
rect 445 1218 484 1252
rect 372 1180 484 1218
rect 372 1146 411 1180
rect 445 1146 484 1180
rect 372 1108 484 1146
rect 372 1074 411 1108
rect 445 1074 484 1108
rect 372 1036 484 1074
rect 372 1002 411 1036
rect 445 1002 484 1036
rect 372 964 484 1002
rect 372 930 411 964
rect 445 930 484 964
rect 24716 1362 24755 1396
rect 24789 1362 24828 1396
rect 24716 1324 24828 1362
rect 24716 1290 24755 1324
rect 24789 1290 24828 1324
rect 24716 1252 24828 1290
rect 24716 1218 24755 1252
rect 24789 1218 24828 1252
rect 24716 1180 24828 1218
rect 24716 1146 24755 1180
rect 24789 1146 24828 1180
rect 24716 1108 24828 1146
rect 24716 1074 24755 1108
rect 24789 1074 24828 1108
rect 24716 1036 24828 1074
rect 24716 1002 24755 1036
rect 24789 1002 24828 1036
rect 24716 964 24828 1002
rect 372 892 484 930
rect 372 858 411 892
rect 445 858 484 892
rect 372 820 484 858
rect 372 786 411 820
rect 445 786 484 820
rect 372 748 484 786
rect 372 714 411 748
rect 445 714 484 748
rect 7494 740 7554 922
rect 372 676 484 714
rect 6324 736 6396 740
rect 6324 684 6334 736
rect 6386 684 6396 736
rect 6324 680 6396 684
rect 7488 736 7560 740
rect 7488 684 7498 736
rect 7550 684 7560 736
rect 7488 680 7560 684
rect 372 642 411 676
rect 445 642 484 676
rect 372 604 484 642
rect 372 570 411 604
rect 445 570 484 604
rect 372 532 484 570
rect 372 498 411 532
rect 445 498 484 532
rect 372 460 484 498
rect 6194 532 6266 536
rect 6194 480 6204 532
rect 6256 480 6266 532
rect 6194 476 6266 480
rect 372 426 411 460
rect 445 426 484 460
rect 372 388 484 426
rect 372 354 411 388
rect 445 354 484 388
rect 372 316 484 354
rect 372 282 411 316
rect 445 282 484 316
rect 372 244 484 282
rect 372 210 411 244
rect 445 210 484 244
rect 372 172 484 210
rect 372 138 411 172
rect 445 138 484 172
rect 372 100 484 138
rect 372 66 411 100
rect 445 66 484 100
rect 372 28 484 66
rect 372 -6 411 28
rect 445 -6 484 28
rect 372 -44 484 -6
rect 372 -78 411 -44
rect 445 -78 484 -44
rect 372 -116 484 -78
rect 372 -150 411 -116
rect 445 -150 484 -116
rect 372 -188 484 -150
rect 372 -222 411 -188
rect 445 -222 484 -188
rect 372 -260 484 -222
rect 372 -294 411 -260
rect 445 -294 484 -260
rect 372 -332 484 -294
rect 372 -366 411 -332
rect 445 -366 484 -332
rect 372 -404 484 -366
rect 372 -438 411 -404
rect 445 -438 484 -404
rect 372 -476 484 -438
rect 372 -510 411 -476
rect 445 -510 484 -476
rect 372 -548 484 -510
rect 372 -582 411 -548
rect 445 -582 484 -548
rect 372 -620 484 -582
rect 372 -654 411 -620
rect 445 -654 484 -620
rect 372 -692 484 -654
rect 372 -726 411 -692
rect 445 -726 484 -692
rect 372 -764 484 -726
rect 372 -798 411 -764
rect 445 -798 484 -764
rect 372 -836 484 -798
rect 372 -870 411 -836
rect 445 -870 484 -836
rect 372 -908 484 -870
rect 372 -942 411 -908
rect 445 -942 484 -908
rect 372 -980 484 -942
rect 372 -1014 411 -980
rect 445 -1014 484 -980
rect 372 -1052 484 -1014
rect 372 -1086 411 -1052
rect 445 -1086 484 -1052
rect 372 -1124 484 -1086
rect 372 -1158 411 -1124
rect 445 -1158 484 -1124
rect 372 -1196 484 -1158
rect 372 -1230 411 -1196
rect 445 -1230 484 -1196
rect 372 -1268 484 -1230
rect 372 -1302 411 -1268
rect 445 -1302 484 -1268
rect 372 -1340 484 -1302
rect 372 -1374 411 -1340
rect 445 -1374 484 -1340
rect 372 -1412 484 -1374
rect 372 -1446 411 -1412
rect 445 -1446 484 -1412
rect 372 -1484 484 -1446
rect 372 -1518 411 -1484
rect 445 -1518 484 -1484
rect 372 -1556 484 -1518
rect 372 -1590 411 -1556
rect 445 -1590 484 -1556
rect 372 -1628 484 -1590
rect 372 -1662 411 -1628
rect 445 -1662 484 -1628
rect 372 -1700 484 -1662
rect 372 -1734 411 -1700
rect 445 -1734 484 -1700
rect 4186 -1652 4258 -1648
rect 4186 -1704 4196 -1652
rect 4248 -1704 4258 -1652
rect 4186 -1708 4258 -1704
rect 372 -1772 484 -1734
rect 372 -1806 411 -1772
rect 445 -1806 484 -1772
rect 372 -1844 484 -1806
rect 372 -1878 411 -1844
rect 445 -1878 484 -1844
rect 372 -1916 484 -1878
rect 372 -1950 411 -1916
rect 445 -1950 484 -1916
rect 372 -1988 484 -1950
rect 372 -2022 411 -1988
rect 445 -2022 484 -1988
rect 372 -2060 484 -2022
rect 372 -2094 411 -2060
rect 445 -2094 484 -2060
rect 372 -2132 484 -2094
rect 372 -2166 411 -2132
rect 445 -2166 484 -2132
rect 372 -2204 484 -2166
rect 372 -2238 411 -2204
rect 445 -2238 484 -2204
rect 372 -2276 484 -2238
rect 372 -2310 411 -2276
rect 445 -2310 484 -2276
rect 372 -2348 484 -2310
rect 372 -2382 411 -2348
rect 445 -2382 484 -2348
rect 372 -2420 484 -2382
rect 372 -2454 411 -2420
rect 445 -2454 484 -2420
rect 372 -2492 484 -2454
rect 372 -2526 411 -2492
rect 445 -2526 484 -2492
rect 372 -2564 484 -2526
rect 372 -2598 411 -2564
rect 445 -2598 484 -2564
rect 372 -2636 484 -2598
rect 372 -2670 411 -2636
rect 445 -2670 484 -2636
rect 372 -2708 484 -2670
rect 372 -2742 411 -2708
rect 445 -2742 484 -2708
rect 372 -2780 484 -2742
rect 372 -2814 411 -2780
rect 445 -2814 484 -2780
rect 372 -2852 484 -2814
rect 372 -2886 411 -2852
rect 445 -2886 484 -2852
rect 372 -2924 484 -2886
rect 372 -2958 411 -2924
rect 445 -2958 484 -2924
rect 372 -2996 484 -2958
rect 372 -3030 411 -2996
rect 445 -3030 484 -2996
rect 372 -3068 484 -3030
rect 372 -3102 411 -3068
rect 445 -3102 484 -3068
rect 372 -3140 484 -3102
rect 372 -3174 411 -3140
rect 445 -3174 484 -3140
rect 372 -3212 484 -3174
rect 372 -3246 411 -3212
rect 445 -3246 484 -3212
rect 372 -3284 484 -3246
rect 372 -3318 411 -3284
rect 445 -3318 484 -3284
rect 372 -3356 484 -3318
rect 372 -3390 411 -3356
rect 445 -3390 484 -3356
rect 372 -3428 484 -3390
rect 372 -3462 411 -3428
rect 445 -3462 484 -3428
rect 372 -3500 484 -3462
rect 372 -3534 411 -3500
rect 445 -3534 484 -3500
rect 372 -3572 484 -3534
rect 372 -3606 411 -3572
rect 445 -3606 484 -3572
rect 372 -3644 484 -3606
rect 372 -3678 411 -3644
rect 445 -3678 484 -3644
rect 372 -3716 484 -3678
rect 372 -3750 411 -3716
rect 445 -3750 484 -3716
rect 372 -3788 484 -3750
rect 372 -3822 411 -3788
rect 445 -3822 484 -3788
rect 372 -3860 484 -3822
rect 372 -3894 411 -3860
rect 445 -3894 484 -3860
rect 372 -3932 484 -3894
rect 372 -3966 411 -3932
rect 445 -3966 484 -3932
rect 372 -4004 484 -3966
rect 372 -4038 411 -4004
rect 445 -4038 484 -4004
rect 372 -4076 484 -4038
rect 372 -4110 411 -4076
rect 445 -4110 484 -4076
rect 372 -4148 484 -4110
rect 372 -4182 411 -4148
rect 445 -4182 484 -4148
rect 372 -4220 484 -4182
rect 372 -4254 411 -4220
rect 445 -4254 484 -4220
rect 372 -4292 484 -4254
rect 372 -4326 411 -4292
rect 445 -4326 484 -4292
rect 372 -4364 484 -4326
rect 372 -4398 411 -4364
rect 445 -4398 484 -4364
rect 372 -4436 484 -4398
rect 372 -4470 411 -4436
rect 445 -4470 484 -4436
rect 372 -4508 484 -4470
rect 372 -4542 411 -4508
rect 445 -4542 484 -4508
rect 372 -4580 484 -4542
rect 372 -4614 411 -4580
rect 445 -4614 484 -4580
rect 372 -4652 484 -4614
rect 372 -4686 411 -4652
rect 445 -4686 484 -4652
rect 372 -4724 484 -4686
rect 372 -4758 411 -4724
rect 445 -4758 484 -4724
rect 372 -4796 484 -4758
rect 372 -4830 411 -4796
rect 445 -4830 484 -4796
rect 372 -4868 484 -4830
rect 372 -4902 411 -4868
rect 445 -4902 484 -4868
rect 372 -4940 484 -4902
rect 372 -4974 411 -4940
rect 445 -4974 484 -4940
rect 372 -5012 484 -4974
rect 372 -5046 411 -5012
rect 445 -5046 484 -5012
rect 372 -5084 484 -5046
rect 372 -5118 411 -5084
rect 445 -5118 484 -5084
rect 372 -5156 484 -5118
rect 372 -5190 411 -5156
rect 445 -5190 484 -5156
rect 372 -5228 484 -5190
rect 372 -5262 411 -5228
rect 445 -5262 484 -5228
rect 372 -5300 484 -5262
rect 372 -5334 411 -5300
rect 445 -5334 484 -5300
rect 372 -5372 484 -5334
rect 372 -5406 411 -5372
rect 445 -5406 484 -5372
rect 372 -5444 484 -5406
rect 372 -5478 411 -5444
rect 445 -5478 484 -5444
rect 372 -5516 484 -5478
rect 372 -5550 411 -5516
rect 445 -5550 484 -5516
rect 372 -5588 484 -5550
rect 372 -5622 411 -5588
rect 445 -5622 484 -5588
rect 372 -5660 484 -5622
rect 372 -5694 411 -5660
rect 445 -5694 484 -5660
rect 372 -5732 484 -5694
rect 372 -5766 411 -5732
rect 445 -5766 484 -5732
rect 372 -5804 484 -5766
rect 372 -5838 411 -5804
rect 445 -5838 484 -5804
rect 372 -5876 484 -5838
rect 372 -5910 411 -5876
rect 445 -5910 484 -5876
rect 372 -5948 484 -5910
rect 372 -5982 411 -5948
rect 445 -5982 484 -5948
rect 372 -6020 484 -5982
rect 372 -6054 411 -6020
rect 445 -6054 484 -6020
rect 372 -6092 484 -6054
rect 372 -6126 411 -6092
rect 445 -6126 484 -6092
rect 372 -6164 484 -6126
rect 372 -6198 411 -6164
rect 445 -6198 484 -6164
rect 372 -6236 484 -6198
rect 372 -6270 411 -6236
rect 445 -6270 484 -6236
rect 372 -6308 484 -6270
rect 372 -6342 411 -6308
rect 445 -6342 484 -6308
rect 372 -6380 484 -6342
rect 372 -6414 411 -6380
rect 445 -6414 484 -6380
rect 372 -6452 484 -6414
rect 372 -6486 411 -6452
rect 445 -6486 484 -6452
rect 372 -6524 484 -6486
rect 372 -6558 411 -6524
rect 445 -6558 484 -6524
rect 372 -6596 484 -6558
rect 372 -6630 411 -6596
rect 445 -6630 484 -6596
rect 372 -6668 484 -6630
rect 372 -6702 411 -6668
rect 445 -6702 484 -6668
rect 372 -6740 484 -6702
rect 372 -6774 411 -6740
rect 445 -6774 484 -6740
rect 372 -6812 484 -6774
rect 372 -6846 411 -6812
rect 445 -6846 484 -6812
rect 372 -6884 484 -6846
rect 372 -6918 411 -6884
rect 445 -6918 484 -6884
rect 372 -6956 484 -6918
rect 2014 -5024 3236 -4964
rect 2014 -6940 2074 -5024
rect 2156 -5238 2216 -5024
rect 2668 -5128 2728 -5024
rect 3176 -5240 3236 -5024
rect 3676 -5906 3736 -5824
rect 3670 -5910 3742 -5906
rect 3670 -5962 3680 -5910
rect 3732 -5962 3742 -5910
rect 3670 -5966 3742 -5962
rect 3778 -6022 3850 -6018
rect 3778 -6074 3788 -6022
rect 3840 -6074 3850 -6022
rect 3778 -6078 3850 -6074
rect 3784 -6158 3844 -6078
rect 372 -6990 411 -6956
rect 445 -6990 484 -6956
rect 372 -7028 484 -6990
rect 2008 -6944 2080 -6940
rect 2008 -6996 2018 -6944
rect 2070 -6996 2080 -6944
rect 2008 -7000 2080 -6996
rect 372 -7062 411 -7028
rect 445 -7062 484 -7028
rect 372 -7100 484 -7062
rect 372 -7134 411 -7100
rect 445 -7134 484 -7100
rect 372 -7172 484 -7134
rect 372 -7206 411 -7172
rect 445 -7206 484 -7172
rect 372 -7244 484 -7206
rect 372 -7278 411 -7244
rect 445 -7278 484 -7244
rect 372 -7316 484 -7278
rect 372 -7350 411 -7316
rect 445 -7350 484 -7316
rect 372 -7388 484 -7350
rect 372 -7422 411 -7388
rect 445 -7422 484 -7388
rect 372 -7460 484 -7422
rect 372 -7494 411 -7460
rect 445 -7494 484 -7460
rect 372 -7532 484 -7494
rect 372 -7566 411 -7532
rect 445 -7566 484 -7532
rect 372 -7604 484 -7566
rect 372 -7638 411 -7604
rect 445 -7638 484 -7604
rect 372 -7676 484 -7638
rect 372 -7710 411 -7676
rect 445 -7710 484 -7676
rect 372 -7748 484 -7710
rect 372 -7782 411 -7748
rect 445 -7782 484 -7748
rect 372 -7820 484 -7782
rect 372 -7854 411 -7820
rect 445 -7854 484 -7820
rect 372 -7892 484 -7854
rect 372 -7926 411 -7892
rect 445 -7926 484 -7892
rect 372 -7964 484 -7926
rect 372 -7998 411 -7964
rect 445 -7998 484 -7964
rect 372 -8036 484 -7998
rect 372 -8070 411 -8036
rect 445 -8070 484 -8036
rect 372 -8108 484 -8070
rect 1888 -8028 1948 -8022
rect 2014 -8028 2074 -7000
rect 2154 -7050 2214 -6738
rect 2656 -7050 2716 -6856
rect 3174 -7050 3234 -6746
rect 2154 -7054 3240 -7050
rect 2154 -7106 3178 -7054
rect 3230 -7106 3240 -7054
rect 2154 -7110 3240 -7106
rect 2154 -7312 2214 -7110
rect 2656 -7188 2716 -7110
rect 3174 -7316 3234 -7110
rect 3684 -7194 3744 -6860
rect 3690 -7974 3750 -7888
rect 3684 -7978 3756 -7974
rect 1888 -8032 3238 -8028
rect 1888 -8084 1892 -8032
rect 1944 -8084 3238 -8032
rect 3684 -8030 3694 -7978
rect 3746 -8030 3756 -7978
rect 3684 -8034 3756 -8030
rect 1888 -8088 3238 -8084
rect 1888 -8094 1948 -8088
rect 372 -8142 411 -8108
rect 445 -8142 484 -8108
rect 372 -8180 484 -8142
rect 372 -8214 411 -8180
rect 445 -8214 484 -8180
rect 372 -8252 484 -8214
rect 372 -8286 411 -8252
rect 445 -8286 484 -8252
rect 372 -8324 484 -8286
rect 372 -8358 411 -8324
rect 445 -8358 484 -8324
rect 2152 -8336 2212 -8088
rect 2660 -8226 2720 -8088
rect 3178 -8332 3238 -8088
rect 3790 -8078 3862 -8074
rect 3790 -8130 3800 -8078
rect 3852 -8130 3862 -8078
rect 3790 -8134 3862 -8130
rect 3796 -8222 3856 -8134
rect 4192 -8358 4252 -1708
rect 6200 -2080 6260 476
rect 6330 -1934 6390 680
rect 7488 532 7560 536
rect 7488 480 7498 532
rect 7550 480 7560 532
rect 7488 476 7560 480
rect 7494 288 7554 476
rect 7998 376 8058 834
rect 8514 286 8574 926
rect 9530 636 9590 914
rect 9524 632 9596 636
rect 9524 580 9534 632
rect 9586 580 9596 632
rect 9524 576 9596 580
rect 10538 296 10602 944
rect 11560 632 11632 636
rect 11560 580 11570 632
rect 11622 580 11632 632
rect 11560 576 11632 580
rect 11566 288 11626 576
rect 12574 292 12638 940
rect 13092 378 13152 836
rect 13604 740 13664 926
rect 13598 736 13670 740
rect 13598 684 13608 736
rect 13660 684 13670 736
rect 13598 680 13670 684
rect 13594 532 13666 536
rect 13594 480 13604 532
rect 13656 480 13666 532
rect 13594 476 13666 480
rect 13600 300 13660 476
rect 14110 384 14170 842
rect 14616 294 14680 942
rect 15126 376 15186 839
rect 15638 740 15698 924
rect 15632 736 15704 740
rect 15632 684 15642 736
rect 15694 684 15704 736
rect 15632 680 15704 684
rect 16138 536 16198 839
rect 15630 532 15702 536
rect 15630 480 15640 532
rect 15692 480 15702 532
rect 15630 476 15702 480
rect 16132 532 16204 536
rect 16132 480 16142 532
rect 16194 480 16204 532
rect 16132 476 16204 480
rect 15636 294 15696 476
rect 16138 376 16198 476
rect 16654 278 16718 926
rect 17666 632 17738 636
rect 17666 580 17676 632
rect 17728 580 17738 632
rect 17666 576 17738 580
rect 17152 532 17224 536
rect 17152 480 17162 532
rect 17214 480 17224 532
rect 17152 476 17224 480
rect 17158 382 17218 476
rect 17672 302 17732 576
rect 18178 532 18250 536
rect 18690 532 18750 934
rect 24716 930 24755 964
rect 24789 930 24828 964
rect 19706 636 19766 918
rect 19700 632 19772 636
rect 19700 580 19710 632
rect 19762 580 19772 632
rect 19700 576 19772 580
rect 20730 538 20790 924
rect 18178 480 18188 532
rect 18240 480 18250 532
rect 18178 476 18250 480
rect 18684 528 18756 532
rect 18684 476 18694 528
rect 18746 476 18756 528
rect 18184 382 18244 476
rect 18684 472 18756 476
rect 19198 528 19270 532
rect 19198 476 19208 528
rect 19260 476 19270 528
rect 19198 472 19270 476
rect 19702 528 19774 532
rect 19702 476 19712 528
rect 19764 476 19774 528
rect 19702 472 19774 476
rect 20208 528 20280 532
rect 20208 476 20218 528
rect 20270 476 20280 528
rect 20208 472 20280 476
rect 20730 528 20794 538
rect 20730 476 20738 528
rect 20790 476 20794 528
rect 18690 282 18750 472
rect 19204 380 19264 472
rect 19708 298 19768 472
rect 20214 380 20274 472
rect 20730 466 20794 476
rect 20730 290 20790 466
rect 21210 382 21270 845
rect 21746 740 21806 926
rect 24716 892 24828 930
rect 24716 858 24755 892
rect 24789 858 24828 892
rect 24716 820 24828 858
rect 24716 786 24755 820
rect 24789 786 24828 820
rect 24716 748 24828 786
rect 21740 736 21812 740
rect 21740 684 21750 736
rect 21802 684 21812 736
rect 21740 680 21812 684
rect 22990 736 23062 740
rect 22990 684 23000 736
rect 23052 684 23062 736
rect 22990 680 23062 684
rect 24716 714 24755 748
rect 24789 714 24828 748
rect 21750 464 22820 524
rect 21750 298 21810 464
rect 22256 390 22316 464
rect 22760 292 22820 464
rect 14618 -204 14678 -202
rect 6476 -400 6536 -214
rect 6988 -400 7048 -312
rect 7494 -400 7554 -220
rect 10546 -224 10606 -222
rect 6476 -460 7554 -400
rect 7488 -604 7548 -602
rect 6478 -664 7548 -604
rect 6478 -842 6538 -664
rect 6988 -744 7048 -664
rect 7488 -842 7548 -664
rect 7980 -618 8040 -296
rect 7980 -670 7984 -618
rect 8036 -670 8040 -618
rect 7980 -754 8040 -670
rect 8510 -396 8570 -224
rect 9008 -396 9068 -302
rect 9528 -396 9588 -230
rect 10036 -396 10096 -298
rect 8510 -402 10096 -396
rect 10546 -398 10610 -224
rect 8510 -454 10040 -402
rect 10092 -454 10096 -402
rect 8510 -456 10096 -454
rect 8510 -862 8570 -456
rect 10036 -464 10096 -456
rect 10540 -402 10612 -398
rect 10540 -454 10550 -402
rect 10602 -454 10612 -402
rect 10540 -458 10612 -454
rect 9522 -502 9598 -496
rect 9522 -554 9534 -502
rect 9586 -554 9598 -502
rect 9522 -560 9598 -554
rect 9012 -618 9084 -614
rect 9012 -670 9022 -618
rect 9074 -670 9084 -618
rect 9012 -674 9084 -670
rect 9528 -654 9592 -560
rect 10024 -618 10096 -614
rect 9018 -754 9078 -674
rect 9528 -856 9594 -654
rect 10024 -670 10034 -618
rect 10086 -670 10096 -618
rect 10024 -674 10096 -670
rect 10030 -758 10090 -674
rect 9528 -860 9592 -856
rect 10546 -858 10610 -458
rect 11040 -606 11100 -310
rect 11564 -496 11628 -214
rect 12580 -216 12640 -214
rect 11398 -502 11628 -496
rect 11398 -554 11410 -502
rect 11462 -554 11628 -502
rect 11398 -560 11628 -554
rect 12064 -606 12124 -310
rect 12580 -398 12644 -216
rect 12574 -402 12646 -398
rect 12574 -454 12584 -402
rect 12636 -454 12646 -402
rect 12574 -458 12646 -454
rect 11034 -610 11106 -606
rect 11034 -662 11044 -610
rect 11096 -662 11106 -610
rect 11034 -666 11106 -662
rect 12058 -610 12130 -606
rect 12058 -662 12068 -610
rect 12120 -662 12130 -610
rect 12058 -666 12130 -662
rect 12580 -870 12644 -458
rect 13092 -606 13152 -296
rect 13086 -610 13158 -606
rect 13086 -662 13096 -610
rect 13148 -662 13158 -610
rect 13086 -666 13158 -662
rect 13092 -754 13152 -666
rect 14120 -764 14180 -306
rect 14618 -400 14682 -204
rect 16654 -208 16714 -206
rect 14612 -404 14684 -400
rect 14612 -456 14622 -404
rect 14674 -456 14684 -404
rect 14612 -460 14684 -456
rect 14618 -850 14682 -460
rect 15138 -754 15198 -291
rect 15638 -498 15698 -220
rect 15632 -502 15704 -498
rect 15632 -554 15642 -502
rect 15694 -554 15704 -502
rect 15632 -558 15704 -554
rect 16138 -758 16198 -295
rect 16654 -400 16718 -208
rect 18690 -400 18750 -214
rect 19192 -400 19252 -308
rect 16648 -404 16720 -400
rect 16648 -456 16658 -404
rect 16710 -456 16720 -404
rect 16648 -460 16720 -456
rect 17148 -404 17220 -400
rect 17148 -456 17158 -404
rect 17210 -456 17220 -404
rect 17148 -460 17220 -456
rect 17662 -404 17734 -400
rect 17662 -456 17672 -404
rect 17724 -456 17734 -404
rect 17662 -460 17734 -456
rect 18186 -404 18258 -400
rect 18186 -456 18196 -404
rect 18248 -456 18258 -404
rect 18186 -460 18258 -456
rect 18684 -404 18756 -400
rect 18684 -456 18694 -404
rect 18746 -456 18756 -404
rect 18684 -460 18756 -456
rect 19186 -404 19258 -400
rect 19706 -402 19766 -180
rect 20724 -220 20784 -218
rect 20214 -402 20274 -296
rect 20724 -402 20788 -220
rect 19186 -456 19196 -404
rect 19248 -456 19258 -404
rect 19186 -460 19258 -456
rect 19700 -406 19772 -402
rect 19700 -458 19710 -406
rect 19762 -458 19772 -406
rect 16654 -862 16718 -460
rect 17154 -754 17214 -460
rect 17668 -864 17728 -460
rect 18192 -754 18252 -460
rect 18690 -864 18750 -460
rect 19700 -462 19772 -458
rect 20208 -406 20280 -402
rect 20208 -458 20218 -406
rect 20270 -458 20280 -406
rect 20208 -462 20280 -458
rect 20718 -406 20790 -402
rect 20718 -458 20728 -406
rect 20780 -458 20790 -406
rect 20718 -462 20790 -458
rect 19190 -618 19262 -614
rect 19190 -670 19200 -618
rect 19252 -670 19262 -618
rect 19190 -674 19262 -670
rect 20202 -618 20274 -614
rect 20202 -670 20212 -618
rect 20264 -670 20274 -618
rect 20202 -674 20274 -670
rect 19196 -756 19256 -674
rect 20208 -750 20268 -674
rect 20724 -856 20788 -462
rect 21210 -614 21270 -297
rect 21746 -498 21806 -220
rect 21740 -502 21812 -498
rect 21740 -554 21750 -502
rect 21802 -554 21812 -502
rect 21740 -558 21812 -554
rect 21748 -612 21808 -610
rect 21204 -618 21276 -614
rect 21204 -670 21214 -618
rect 21266 -670 21276 -618
rect 21204 -674 21276 -670
rect 21748 -672 22820 -612
rect 21210 -760 21270 -674
rect 21748 -836 21808 -672
rect 22252 -748 22312 -672
rect 22760 -860 22820 -672
rect 7488 -1594 7552 -1344
rect 7044 -1654 7552 -1594
rect 6324 -1938 6396 -1934
rect 6324 -1990 6334 -1938
rect 6386 -1990 6396 -1938
rect 6324 -1994 6396 -1990
rect 6200 -2140 6620 -2080
rect 6560 -4952 6620 -2140
rect 6680 -4346 6752 -4342
rect 6680 -4398 6690 -4346
rect 6742 -4398 6752 -4346
rect 6680 -4402 6752 -4398
rect 6554 -4956 6626 -4952
rect 5210 -5020 6420 -4960
rect 6554 -5008 6564 -4956
rect 6616 -5008 6626 -4956
rect 6554 -5012 6626 -5008
rect 5210 -5236 5270 -5020
rect 5722 -5124 5782 -5020
rect 6228 -5234 6288 -5020
rect 4568 -6018 4628 -5822
rect 4692 -5910 4764 -5906
rect 4692 -5962 4702 -5910
rect 4754 -5962 4764 -5910
rect 4692 -5966 4764 -5962
rect 4562 -6022 4634 -6018
rect 4562 -6074 4572 -6022
rect 4624 -6074 4634 -6022
rect 4562 -6078 4634 -6074
rect 4698 -6154 4758 -5966
rect 4702 -7190 4762 -6856
rect 5208 -6940 5268 -6710
rect 5722 -6940 5782 -6856
rect 6228 -6940 6288 -6750
rect 5202 -6944 6288 -6940
rect 5202 -6996 5212 -6944
rect 5264 -6996 6288 -6944
rect 5202 -7000 6288 -6996
rect 5208 -7308 5268 -7000
rect 5722 -7194 5782 -7000
rect 6228 -7288 6288 -7000
rect 6360 -7050 6420 -5020
rect 6354 -7054 6426 -7050
rect 6354 -7106 6364 -7054
rect 6416 -7106 6426 -7054
rect 6354 -7110 6426 -7106
rect 4582 -8074 4642 -7888
rect 4694 -7978 4766 -7974
rect 4694 -8030 4704 -7978
rect 4756 -8030 4766 -7978
rect 6360 -8028 6420 -7110
rect 6546 -7182 6618 -7178
rect 6546 -7234 6556 -7182
rect 6608 -7234 6618 -7182
rect 6546 -7238 6618 -7234
rect 4694 -8034 4766 -8030
rect 4576 -8078 4648 -8074
rect 4576 -8130 4586 -8078
rect 4638 -8130 4648 -8078
rect 4576 -8134 4648 -8130
rect 4700 -8224 4760 -8034
rect 5208 -8088 6420 -8028
rect 5208 -8314 5268 -8088
rect 5710 -8226 5770 -8088
rect 6228 -8352 6288 -8088
rect 372 -8396 484 -8358
rect 372 -8430 411 -8396
rect 445 -8430 484 -8396
rect 372 -8468 484 -8430
rect 372 -8502 411 -8468
rect 445 -8502 484 -8468
rect 372 -8540 484 -8502
rect 372 -8574 411 -8540
rect 445 -8574 484 -8540
rect 372 -8612 484 -8574
rect 372 -8646 411 -8612
rect 445 -8646 484 -8612
rect 372 -8684 484 -8646
rect 372 -8718 411 -8684
rect 445 -8718 484 -8684
rect 372 -8756 484 -8718
rect 372 -8790 411 -8756
rect 445 -8790 484 -8756
rect 372 -8828 484 -8790
rect 372 -8862 411 -8828
rect 445 -8862 484 -8828
rect 372 -8900 484 -8862
rect 372 -8934 411 -8900
rect 445 -8934 484 -8900
rect 372 -8972 484 -8934
rect 372 -9006 411 -8972
rect 445 -9006 484 -8972
rect 372 -9044 484 -9006
rect 372 -9078 411 -9044
rect 445 -9078 484 -9044
rect 372 -9116 484 -9078
rect 372 -9150 411 -9116
rect 445 -9150 484 -9116
rect 1402 -9084 1462 -9078
rect 3682 -9084 3742 -8916
rect 1402 -9088 3742 -9084
rect 1402 -9140 1406 -9088
rect 1458 -9140 3742 -9088
rect 1402 -9144 3742 -9140
rect 1402 -9150 1462 -9144
rect 372 -9188 484 -9150
rect 372 -9222 411 -9188
rect 445 -9222 484 -9188
rect 372 -9260 484 -9222
rect 372 -9294 411 -9260
rect 445 -9294 484 -9260
rect 372 -9332 484 -9294
rect 1542 -9260 1602 -9254
rect 4688 -9260 4748 -8909
rect 1542 -9264 4748 -9260
rect 1542 -9316 1546 -9264
rect 1598 -9316 4748 -9264
rect 1542 -9320 4748 -9316
rect 1542 -9326 1602 -9320
rect 372 -9366 411 -9332
rect 445 -9366 484 -9332
rect 372 -9404 484 -9366
rect 372 -9438 411 -9404
rect 445 -9438 484 -9404
rect 372 -9476 484 -9438
rect 372 -9510 411 -9476
rect 445 -9510 484 -9476
rect 2442 -9434 2502 -9428
rect 5210 -9434 5270 -8778
rect 2442 -9438 5270 -9434
rect 2442 -9490 2446 -9438
rect 2498 -9490 5270 -9438
rect 2442 -9494 5270 -9490
rect 2442 -9500 2502 -9494
rect 372 -9548 484 -9510
rect 372 -9582 411 -9548
rect 445 -9582 484 -9548
rect 372 -9620 484 -9582
rect 372 -9654 411 -9620
rect 445 -9654 484 -9620
rect 1282 -9584 1342 -9578
rect 6552 -9584 6612 -7238
rect 6686 -8330 6746 -4402
rect 6796 -4956 6868 -4952
rect 6796 -5008 6806 -4956
rect 6858 -5008 6868 -4956
rect 6796 -5012 6868 -5008
rect 6802 -7074 6862 -5012
rect 7044 -5916 7104 -1654
rect 7488 -1784 7552 -1654
rect 7482 -1790 7558 -1784
rect 7482 -1842 7494 -1790
rect 7546 -1842 7558 -1790
rect 7482 -1848 7558 -1842
rect 7312 -1938 7372 -1928
rect 7312 -1990 7316 -1938
rect 7368 -1990 7372 -1938
rect 7312 -4870 7372 -1990
rect 7990 -2040 8050 -1446
rect 8510 -1536 8570 -1350
rect 10546 -1362 10606 -1360
rect 8504 -1540 8576 -1536
rect 8504 -1592 8514 -1540
rect 8566 -1592 8576 -1540
rect 8504 -1596 8576 -1592
rect 9032 -2040 9092 -1440
rect 9526 -1646 9590 -1362
rect 9520 -1652 9596 -1646
rect 9520 -1704 9532 -1652
rect 9584 -1704 9596 -1652
rect 9520 -1710 9596 -1704
rect 10032 -2040 10092 -1446
rect 10546 -1536 10610 -1362
rect 11068 -1536 11128 -1436
rect 11566 -1536 11626 -1330
rect 12580 -1354 12640 -1352
rect 10540 -1540 10612 -1536
rect 10540 -1592 10550 -1540
rect 10602 -1592 10612 -1540
rect 10540 -1596 10612 -1592
rect 11062 -1540 11134 -1536
rect 11062 -1592 11072 -1540
rect 11124 -1592 11134 -1540
rect 11062 -1596 11134 -1592
rect 11560 -1540 11632 -1536
rect 11560 -1592 11570 -1540
rect 11622 -1592 11632 -1540
rect 11560 -1596 11632 -1592
rect 12040 -1544 12100 -1444
rect 12580 -1532 12644 -1354
rect 12040 -1596 12044 -1544
rect 12096 -1596 12100 -1544
rect 7422 -2044 7494 -2040
rect 7422 -2096 7432 -2044
rect 7484 -2096 7494 -2044
rect 7422 -2100 7494 -2096
rect 7984 -2044 8056 -2040
rect 7984 -2096 7994 -2044
rect 8046 -2096 8056 -2044
rect 7984 -2100 8056 -2096
rect 9026 -2044 9098 -2040
rect 9026 -2096 9036 -2044
rect 9088 -2096 9098 -2044
rect 9026 -2100 9098 -2096
rect 10026 -2044 10098 -2040
rect 10026 -2096 10036 -2044
rect 10088 -2096 10098 -2044
rect 10026 -2100 10098 -2096
rect 7428 -4682 7488 -2100
rect 12040 -2138 12100 -1596
rect 12548 -1536 12644 -1532
rect 12548 -1541 12646 -1536
rect 12548 -1593 12568 -1541
rect 12620 -1593 12646 -1541
rect 12548 -1596 12646 -1593
rect 13034 -1540 13106 -1536
rect 13034 -1592 13044 -1540
rect 13096 -1592 13106 -1540
rect 13034 -1596 13106 -1592
rect 12548 -2138 12608 -1596
rect 13040 -2138 13100 -1596
rect 13194 -2040 13254 -1444
rect 13598 -1794 13662 -1354
rect 13598 -1846 13604 -1794
rect 13656 -1846 13662 -1794
rect 13598 -1858 13662 -1846
rect 14084 -1538 14144 -1528
rect 14084 -1590 14088 -1538
rect 14140 -1590 14144 -1538
rect 13188 -2044 13260 -2040
rect 13188 -2096 13198 -2044
rect 13250 -2096 13260 -2044
rect 13188 -2100 13260 -2096
rect 14084 -2138 14144 -1590
rect 14204 -2040 14264 -1444
rect 14616 -1536 14676 -1326
rect 16654 -1346 16714 -1344
rect 14610 -1540 14682 -1536
rect 14610 -1592 14620 -1540
rect 14672 -1592 14682 -1540
rect 14610 -1596 14682 -1592
rect 15146 -2040 15206 -1444
rect 15634 -1930 15698 -1350
rect 16128 -1538 16188 -1528
rect 16654 -1534 16718 -1346
rect 16128 -1590 16132 -1538
rect 16184 -1590 16188 -1538
rect 15628 -1936 15704 -1930
rect 15628 -1988 15640 -1936
rect 15692 -1988 15704 -1936
rect 15628 -1994 15704 -1988
rect 14198 -2044 14270 -2040
rect 14198 -2096 14208 -2044
rect 14260 -2096 14270 -2044
rect 14198 -2100 14270 -2096
rect 15140 -2044 15212 -2040
rect 15140 -2096 15150 -2044
rect 15202 -2096 15212 -2044
rect 15140 -2100 15212 -2096
rect 16128 -2138 16188 -1590
rect 16622 -1538 16718 -1534
rect 16622 -1543 16720 -1538
rect 16622 -1595 16642 -1543
rect 16694 -1595 16720 -1543
rect 16622 -1598 16720 -1595
rect 17150 -1548 17210 -1430
rect 17672 -1534 17732 -940
rect 18690 -1358 18750 -1356
rect 16622 -2138 16682 -1598
rect 17150 -1600 17154 -1548
rect 17206 -1600 17210 -1548
rect 17150 -2138 17210 -1600
rect 17638 -1545 17732 -1534
rect 17638 -1597 17659 -1545
rect 17711 -1597 17732 -1545
rect 17638 -1608 17732 -1597
rect 18150 -1548 18210 -1436
rect 18690 -1540 18754 -1358
rect 18150 -1600 18154 -1548
rect 18206 -1600 18210 -1548
rect 18684 -1544 18756 -1540
rect 18684 -1596 18694 -1544
rect 18746 -1596 18756 -1544
rect 18684 -1600 18756 -1596
rect 17638 -2138 17698 -1608
rect 18150 -2138 18210 -1600
rect 19706 -1646 19770 -1352
rect 20724 -1358 20784 -1356
rect 20724 -1540 20788 -1358
rect 20718 -1544 20790 -1540
rect 20718 -1596 20728 -1544
rect 20780 -1596 20790 -1544
rect 20718 -1600 20790 -1596
rect 19700 -1652 19776 -1646
rect 19700 -1704 19712 -1652
rect 19764 -1704 19776 -1652
rect 19700 -1710 19776 -1704
rect 21740 -1934 21800 -1298
rect 22996 -1778 23056 680
rect 22992 -1790 23056 -1778
rect 22992 -1842 22998 -1790
rect 23050 -1842 23056 -1790
rect 22992 -1854 23056 -1842
rect 21734 -1938 21806 -1934
rect 21734 -1990 21744 -1938
rect 21796 -1990 21806 -1938
rect 21734 -1994 21806 -1990
rect 9704 -2198 19944 -2138
rect 7536 -2246 7608 -2242
rect 7536 -2298 7546 -2246
rect 7598 -2298 7608 -2246
rect 7536 -2302 7608 -2298
rect 7542 -4216 7602 -2302
rect 7668 -3176 7728 -2994
rect 8180 -3176 8240 -3086
rect 8686 -3176 8746 -3000
rect 7668 -3178 8746 -3176
rect 7668 -3182 8752 -3178
rect 7668 -3234 8690 -3182
rect 8742 -3234 8752 -3182
rect 7668 -3236 8752 -3234
rect 8680 -3238 8752 -3236
rect 9190 -3286 9250 -3084
rect 9184 -3290 9256 -3286
rect 9184 -3342 9194 -3290
rect 9246 -3342 9256 -3290
rect 9184 -3346 9256 -3342
rect 9190 -3424 9250 -3346
rect 7668 -4216 7728 -4000
rect 8170 -4216 8230 -4110
rect 8682 -4210 8742 -4026
rect 8676 -4214 8748 -4210
rect 8676 -4216 8686 -4214
rect 7542 -4266 8686 -4216
rect 8738 -4266 8748 -4214
rect 7542 -4276 8748 -4266
rect 9188 -4348 9248 -4122
rect 9188 -4400 9192 -4348
rect 9244 -4400 9248 -4348
rect 9188 -4410 9248 -4400
rect 9704 -4552 9764 -2198
rect 10714 -2246 10786 -2242
rect 10714 -2298 10724 -2246
rect 10776 -2298 10786 -2246
rect 10714 -2302 10786 -2298
rect 10720 -2512 10780 -2302
rect 10210 -3280 10270 -3071
rect 10714 -3182 10786 -3178
rect 10714 -3234 10724 -3182
rect 10776 -3234 10786 -3182
rect 10714 -3238 10786 -3234
rect 10210 -3290 10272 -3280
rect 10210 -3342 10216 -3290
rect 10268 -3342 10272 -3290
rect 10210 -3352 10272 -3342
rect 10210 -3414 10270 -3352
rect 10720 -3526 10780 -3238
rect 11232 -3280 11292 -3091
rect 11230 -3290 11292 -3280
rect 11230 -3342 11234 -3290
rect 11286 -3342 11292 -3290
rect 11230 -3352 11292 -3342
rect 11232 -3434 11292 -3352
rect 10202 -4352 10262 -4106
rect 10202 -4404 10206 -4352
rect 10258 -4404 10262 -4352
rect 10202 -4414 10262 -4404
rect 11234 -4344 11294 -4118
rect 11234 -4396 11238 -4344
rect 11290 -4396 11294 -4344
rect 11234 -4406 11294 -4396
rect 11742 -4552 11802 -2198
rect 12252 -3280 12312 -3081
rect 12762 -3178 12822 -2960
rect 12756 -3182 12828 -3178
rect 12756 -3234 12766 -3182
rect 12818 -3234 12828 -3182
rect 12756 -3238 12828 -3234
rect 12252 -3290 12314 -3280
rect 12252 -3342 12258 -3290
rect 12310 -3342 12314 -3290
rect 12252 -3352 12314 -3342
rect 13268 -3290 13328 -3075
rect 13268 -3342 13272 -3290
rect 13324 -3342 13328 -3290
rect 12252 -3424 12312 -3352
rect 13268 -3418 13328 -3342
rect 12232 -4344 12292 -4112
rect 12762 -4210 12822 -3990
rect 12756 -4214 12828 -4210
rect 12756 -4266 12766 -4214
rect 12818 -4266 12828 -4214
rect 12756 -4270 12828 -4266
rect 12232 -4396 12236 -4344
rect 12288 -4396 12292 -4344
rect 12232 -4406 12292 -4396
rect 13276 -4344 13336 -4096
rect 13276 -4396 13280 -4344
rect 13332 -4396 13336 -4344
rect 13276 -4406 13336 -4396
rect 13780 -4552 13840 -2198
rect 14782 -2246 14854 -2242
rect 14782 -2298 14792 -2246
rect 14844 -2298 14854 -2246
rect 14782 -2302 14854 -2298
rect 14788 -2522 14848 -2302
rect 14284 -3280 14344 -3081
rect 14782 -3182 14854 -3178
rect 14782 -3234 14792 -3182
rect 14844 -3234 14854 -3182
rect 14782 -3238 14854 -3234
rect 14284 -3290 14346 -3280
rect 14284 -3342 14290 -3290
rect 14342 -3342 14346 -3290
rect 14284 -3352 14346 -3342
rect 14284 -3424 14344 -3352
rect 14788 -3542 14848 -3238
rect 15294 -3280 15354 -3081
rect 15294 -3290 15356 -3280
rect 15294 -3342 15300 -3290
rect 15352 -3342 15356 -3290
rect 15294 -3352 15356 -3342
rect 15294 -3424 15354 -3352
rect 14280 -4348 14340 -4106
rect 14280 -4400 14284 -4348
rect 14336 -4400 14340 -4348
rect 14280 -4410 14340 -4400
rect 14798 -4460 14858 -3964
rect 15296 -4348 15356 -4102
rect 15296 -4400 15300 -4348
rect 15352 -4400 15356 -4348
rect 15296 -4410 15356 -4400
rect 14588 -4520 14858 -4460
rect 9704 -4556 14146 -4552
rect 9704 -4608 14084 -4556
rect 14136 -4608 14146 -4556
rect 9704 -4612 14146 -4608
rect 7428 -4742 11596 -4682
rect 7306 -4874 7378 -4870
rect 7306 -4926 7316 -4874
rect 7368 -4926 7378 -4874
rect 7306 -4930 7378 -4926
rect 8472 -4874 8544 -4870
rect 8472 -4926 8482 -4874
rect 8534 -4926 8544 -4874
rect 8472 -4930 8544 -4926
rect 7038 -5920 7110 -5916
rect 7038 -5972 7048 -5920
rect 7100 -5972 7110 -5920
rect 7038 -5976 7110 -5972
rect 6796 -7078 6868 -7074
rect 6796 -7130 6806 -7078
rect 6858 -7130 6868 -7078
rect 6796 -7134 6868 -7130
rect 6792 -7292 6864 -7288
rect 6792 -7344 6802 -7292
rect 6854 -7344 6864 -7292
rect 6792 -7348 6864 -7344
rect 6680 -8334 6752 -8330
rect 6680 -8386 6690 -8334
rect 6742 -8386 6752 -8334
rect 6680 -8390 6752 -8386
rect 1282 -9588 6612 -9584
rect 1282 -9640 1286 -9588
rect 1338 -9640 6612 -9588
rect 1282 -9644 6612 -9640
rect 1282 -9650 1342 -9644
rect 372 -9692 484 -9654
rect 372 -9726 411 -9692
rect 445 -9726 484 -9692
rect -13992 -10402 -2722 -10122
rect 372 -10242 484 -9726
rect 2336 -9846 2396 -9840
rect 6798 -9846 6858 -7348
rect 7044 -9588 7104 -5976
rect 7174 -6018 7246 -6014
rect 7174 -6070 7184 -6018
rect 7236 -6070 7246 -6018
rect 7174 -6074 7246 -6070
rect 7038 -9592 7110 -9588
rect 7038 -9644 7048 -9592
rect 7100 -9644 7110 -9592
rect 7038 -9648 7110 -9644
rect 7180 -9718 7240 -6074
rect 7312 -8538 7372 -4930
rect 8478 -5110 8538 -4930
rect 9494 -5130 9554 -4742
rect 10508 -4874 10580 -4870
rect 10508 -4926 10518 -4874
rect 10570 -4926 10580 -4874
rect 10508 -4930 10580 -4926
rect 11016 -4876 11092 -4870
rect 11016 -4928 11028 -4876
rect 11080 -4928 11092 -4876
rect 10514 -5108 10574 -4930
rect 11016 -4934 11092 -4928
rect 11022 -5028 11086 -4934
rect 11536 -5138 11596 -4742
rect 12040 -5028 12100 -4612
rect 7460 -5818 7520 -5624
rect 7974 -5818 8034 -5722
rect 8476 -5818 8536 -5636
rect 7460 -5878 8536 -5818
rect 8966 -6120 9026 -5714
rect 9496 -5818 9556 -5636
rect 9490 -5822 9562 -5818
rect 9490 -5874 9500 -5822
rect 9552 -5874 9562 -5822
rect 9490 -5878 9562 -5874
rect 10004 -5872 10064 -5713
rect 11010 -5872 11070 -5713
rect 11532 -5818 11592 -5632
rect 12042 -5814 12102 -5718
rect 12548 -5814 12608 -4612
rect 13040 -5024 13100 -4612
rect 14078 -5022 14138 -4612
rect 13062 -5814 13122 -5722
rect 13568 -5814 13628 -5636
rect 14072 -5814 14132 -5720
rect 9496 -6014 9556 -5878
rect 10004 -5932 11070 -5872
rect 11526 -5822 11598 -5818
rect 11526 -5874 11536 -5822
rect 11588 -5874 11598 -5822
rect 11526 -5878 11598 -5874
rect 11868 -5820 11940 -5816
rect 11868 -5872 11878 -5820
rect 11930 -5872 11940 -5820
rect 11868 -5876 11940 -5872
rect 12042 -5874 14132 -5814
rect 14588 -5816 14648 -4520
rect 15816 -4556 15876 -2198
rect 17846 -2858 17906 -2198
rect 18858 -2246 18930 -2242
rect 18858 -2298 18868 -2246
rect 18920 -2298 18930 -2246
rect 18858 -2302 18930 -2298
rect 18864 -2512 18924 -2302
rect 16316 -3280 16376 -3075
rect 16830 -3178 16890 -2960
rect 16824 -3182 16896 -3178
rect 16824 -3234 16834 -3182
rect 16886 -3234 16896 -3182
rect 16824 -3238 16896 -3234
rect 17330 -3280 17390 -3075
rect 16316 -3290 16378 -3280
rect 16316 -3342 16322 -3290
rect 16374 -3342 16378 -3290
rect 16316 -3352 16378 -3342
rect 17330 -3290 17392 -3280
rect 17330 -3342 17336 -3290
rect 17388 -3342 17392 -3290
rect 17330 -3352 17392 -3342
rect 16316 -3418 16376 -3352
rect 17330 -3418 17390 -3352
rect 16300 -4348 16360 -4112
rect 16830 -4210 16890 -3974
rect 16824 -4214 16896 -4210
rect 16824 -4266 16834 -4214
rect 16886 -4266 16896 -4214
rect 16824 -4270 16896 -4266
rect 16300 -4400 16304 -4348
rect 16356 -4400 16360 -4348
rect 16300 -4410 16360 -4400
rect 17332 -4344 17392 -4118
rect 17332 -4396 17336 -4344
rect 17388 -4396 17392 -4344
rect 17332 -4406 17392 -4396
rect 15816 -4608 15820 -4556
rect 15872 -4608 15876 -4556
rect 15090 -4754 15166 -4748
rect 15090 -4806 15102 -4754
rect 15154 -4806 15166 -4754
rect 15090 -4812 15166 -4806
rect 15096 -4870 15160 -4812
rect 15816 -4842 15876 -4608
rect 17846 -4452 17906 -2952
rect 18362 -3280 18422 -3075
rect 18860 -3182 18932 -3178
rect 18860 -3234 18870 -3182
rect 18922 -3234 18932 -3182
rect 18860 -3238 18932 -3234
rect 18362 -3290 18424 -3280
rect 18362 -3342 18368 -3290
rect 18420 -3342 18424 -3290
rect 18362 -3352 18424 -3342
rect 18362 -3418 18422 -3352
rect 18866 -3548 18926 -3238
rect 19372 -3280 19432 -3075
rect 19372 -3290 19434 -3280
rect 19372 -3342 19378 -3290
rect 19430 -3342 19434 -3290
rect 19372 -3352 19434 -3342
rect 19372 -3418 19432 -3352
rect 18348 -4348 18408 -4106
rect 18348 -4400 18352 -4348
rect 18404 -4400 18408 -4348
rect 18348 -4410 18408 -4400
rect 19376 -4348 19436 -4112
rect 19376 -4400 19380 -4348
rect 19432 -4400 19436 -4348
rect 19376 -4410 19436 -4400
rect 19884 -4452 19944 -2198
rect 22054 -2246 22126 -2242
rect 22054 -2298 22064 -2246
rect 22116 -2298 22126 -2246
rect 22054 -2302 22126 -2298
rect 20394 -3280 20454 -3081
rect 20902 -3176 20962 -2948
rect 21424 -3176 21484 -3088
rect 21918 -3176 21978 -2998
rect 20902 -3178 21978 -3176
rect 20896 -3182 21978 -3178
rect 20896 -3234 20906 -3182
rect 20958 -3234 21978 -3182
rect 20896 -3236 21978 -3234
rect 20896 -3238 20968 -3236
rect 20394 -3290 20456 -3280
rect 20394 -3342 20400 -3290
rect 20452 -3342 20456 -3290
rect 20394 -3352 20456 -3342
rect 20394 -3424 20454 -3352
rect 20396 -4348 20456 -4106
rect 20898 -4206 20958 -3980
rect 21386 -4206 21446 -4112
rect 21918 -4206 21978 -3984
rect 22060 -4206 22120 -2302
rect 20896 -4210 22120 -4206
rect 20892 -4214 22120 -4210
rect 20892 -4266 20902 -4214
rect 20954 -4266 22120 -4214
rect 20892 -4270 20964 -4266
rect 20396 -4400 20400 -4348
rect 20452 -4400 20456 -4348
rect 20396 -4410 20456 -4400
rect 22848 -4346 22920 -4342
rect 22848 -4398 22858 -4346
rect 22910 -4398 22920 -4346
rect 22848 -4402 22920 -4398
rect 17846 -4512 19944 -4452
rect 17846 -4842 17906 -4512
rect 21708 -4572 21780 -4568
rect 21708 -4624 21718 -4572
rect 21770 -4624 21780 -4572
rect 21708 -4628 21780 -4624
rect 19154 -4754 19230 -4748
rect 19154 -4806 19166 -4754
rect 19218 -4806 19230 -4754
rect 19154 -4812 19230 -4806
rect 20178 -4754 20254 -4748
rect 20178 -4806 20190 -4754
rect 20242 -4806 20254 -4754
rect 20178 -4812 20254 -4806
rect 21190 -4754 21266 -4748
rect 21190 -4806 21202 -4754
rect 21254 -4806 21266 -4754
rect 21190 -4812 21266 -4806
rect 15092 -4876 15168 -4870
rect 15092 -4928 15104 -4876
rect 15156 -4928 15168 -4876
rect 15816 -4902 18210 -4842
rect 19160 -4866 19224 -4812
rect 15092 -4934 15168 -4928
rect 15096 -5022 15160 -4934
rect 16128 -5028 16188 -4902
rect 14582 -5820 14654 -5816
rect 14582 -5872 14592 -5820
rect 14644 -5872 14654 -5820
rect 9490 -6018 9562 -6014
rect 9490 -6070 9500 -6018
rect 9552 -6070 9562 -6018
rect 9490 -6074 9562 -6070
rect 10004 -6120 10064 -5932
rect 10510 -6016 10582 -6012
rect 10510 -6068 10520 -6016
rect 10572 -6068 10582 -6016
rect 10510 -6072 10582 -6068
rect 8476 -6128 8548 -6124
rect 8476 -6180 8486 -6128
rect 8538 -6180 8548 -6128
rect 8476 -6184 8548 -6180
rect 8966 -6180 10064 -6120
rect 10516 -6124 10576 -6072
rect 8482 -6366 8542 -6184
rect 8966 -6282 9026 -6180
rect 10004 -6287 10064 -6180
rect 10510 -6128 10582 -6124
rect 10510 -6180 10520 -6128
rect 10572 -6180 10582 -6128
rect 10510 -6184 10582 -6180
rect 10516 -6362 10576 -6184
rect 11010 -6287 11070 -5932
rect 11874 -6130 11934 -5876
rect 11532 -6190 11934 -6130
rect 11532 -6398 11592 -6190
rect 12548 -6384 12608 -5874
rect 14582 -5876 14654 -5872
rect 15606 -6012 15666 -5582
rect 16116 -5814 16176 -5722
rect 16622 -5814 16682 -4902
rect 17150 -5032 17210 -4902
rect 17142 -5814 17202 -5721
rect 17638 -5814 17698 -4902
rect 18150 -5038 18210 -4902
rect 18654 -4874 18726 -4870
rect 18654 -4926 18664 -4874
rect 18716 -4926 18726 -4874
rect 18654 -4930 18726 -4926
rect 18660 -5112 18720 -4930
rect 19160 -5028 19224 -4930
rect 20184 -5022 20248 -4812
rect 20688 -4874 20760 -4870
rect 20688 -4926 20698 -4874
rect 20750 -4926 20760 -4874
rect 20688 -4930 20760 -4926
rect 20694 -5108 20754 -4930
rect 21196 -5018 21260 -4812
rect 21714 -4866 21774 -4628
rect 21714 -4926 22790 -4866
rect 21714 -5120 21774 -4926
rect 22228 -5022 22288 -4926
rect 22730 -5108 22790 -4926
rect 18154 -5814 18214 -5724
rect 16116 -5874 18214 -5814
rect 15600 -6016 15672 -6012
rect 15600 -6068 15610 -6016
rect 15662 -6068 15672 -6016
rect 15600 -6072 15672 -6068
rect 13566 -6130 13638 -6126
rect 13566 -6182 13576 -6130
rect 13628 -6182 13638 -6130
rect 13566 -6186 13638 -6182
rect 15600 -6130 15672 -6126
rect 15600 -6182 15610 -6130
rect 15662 -6182 15672 -6130
rect 15600 -6186 15672 -6182
rect 13572 -6368 13632 -6186
rect 15606 -6370 15666 -6186
rect 17638 -6360 17698 -5874
rect 18656 -6130 18728 -6126
rect 18656 -6182 18666 -6130
rect 18718 -6182 18728 -6130
rect 18656 -6186 18728 -6182
rect 18662 -6368 18722 -6186
rect 19162 -6287 19222 -5713
rect 19676 -5818 19736 -5636
rect 19670 -5822 19742 -5818
rect 19670 -5874 19680 -5822
rect 19732 -5874 19742 -5822
rect 19670 -5878 19742 -5874
rect 20186 -6287 20246 -5713
rect 20690 -6130 20762 -6126
rect 20690 -6182 20700 -6130
rect 20752 -6182 20762 -6130
rect 20690 -6186 20762 -6182
rect 20696 -6364 20756 -6186
rect 21192 -6281 21252 -5707
rect 21712 -5818 21772 -5632
rect 21706 -5822 21778 -5818
rect 21706 -5874 21716 -5822
rect 21768 -5874 21778 -5822
rect 21706 -5878 21778 -5874
rect 21714 -6180 22790 -6120
rect 21714 -6374 21774 -6180
rect 22228 -6276 22288 -6180
rect 22730 -6362 22790 -6180
rect 7464 -7074 7524 -6880
rect 7978 -7074 8038 -6978
rect 8480 -7074 8540 -6892
rect 7464 -7134 8540 -7074
rect 7464 -7288 7524 -7134
rect 7458 -7292 7530 -7288
rect 7458 -7344 7468 -7292
rect 7520 -7344 7530 -7292
rect 7458 -7348 7530 -7344
rect 7462 -7458 8538 -7398
rect 7462 -7630 7522 -7458
rect 7976 -7532 8036 -7458
rect 8478 -7618 8538 -7458
rect 8960 -7542 9020 -6968
rect 9498 -7182 9558 -6890
rect 9498 -7234 9502 -7182
rect 9554 -7234 9558 -7182
rect 9498 -7244 9558 -7234
rect 9492 -7386 9564 -7382
rect 9492 -7438 9502 -7386
rect 9554 -7438 9564 -7386
rect 9492 -7442 9564 -7438
rect 9498 -7620 9558 -7442
rect 9998 -7543 10058 -6968
rect 11004 -7543 11064 -6968
rect 11534 -7178 11594 -6886
rect 12054 -7070 12114 -6977
rect 12550 -7070 12610 -6886
rect 13066 -7070 13126 -6980
rect 12054 -7130 13126 -7070
rect 13562 -7078 13634 -7074
rect 13562 -7130 13572 -7078
rect 13624 -7130 13634 -7078
rect 11528 -7182 11600 -7178
rect 11528 -7234 11538 -7182
rect 11590 -7234 11600 -7182
rect 11528 -7238 11600 -7234
rect 11526 -7284 11598 -7280
rect 11526 -7336 11536 -7284
rect 11588 -7336 11598 -7284
rect 11526 -7340 11598 -7336
rect 11532 -7382 11592 -7340
rect 11526 -7386 11598 -7382
rect 11526 -7438 11536 -7386
rect 11588 -7438 11598 -7386
rect 11526 -7442 11598 -7438
rect 11532 -7624 11592 -7442
rect 12550 -7634 12610 -7130
rect 13562 -7134 13634 -7130
rect 13568 -7620 13628 -7134
rect 14070 -7236 14130 -6974
rect 14588 -7074 14648 -6892
rect 14582 -7078 14654 -7074
rect 14582 -7130 14592 -7078
rect 14644 -7130 14654 -7078
rect 14582 -7134 14654 -7130
rect 15100 -7236 15160 -6962
rect 14070 -7296 15160 -7236
rect 14070 -7548 14130 -7296
rect 14582 -7384 14654 -7380
rect 14582 -7436 14592 -7384
rect 14644 -7436 14654 -7384
rect 14582 -7440 14654 -7436
rect 14588 -7618 14648 -7440
rect 15100 -7536 15160 -7296
rect 15606 -7380 15666 -6888
rect 15600 -7384 15672 -7380
rect 15600 -7436 15610 -7384
rect 15662 -7436 15672 -7384
rect 15600 -7440 15672 -7436
rect 16112 -7536 16172 -6962
rect 16624 -7074 16684 -6888
rect 17142 -7072 17202 -6979
rect 17638 -7072 17698 -6888
rect 18154 -7072 18214 -6982
rect 16618 -7078 16690 -7074
rect 16618 -7130 16628 -7078
rect 16680 -7130 16690 -7078
rect 16618 -7134 16690 -7130
rect 17142 -7132 18214 -7072
rect 16616 -7384 16688 -7380
rect 16616 -7436 16626 -7384
rect 16678 -7436 16688 -7384
rect 16616 -7440 16688 -7436
rect 16622 -7622 16682 -7440
rect 17638 -7626 17698 -7132
rect 18652 -7182 18724 -7178
rect 18652 -7234 18662 -7182
rect 18714 -7234 18724 -7182
rect 18652 -7238 18724 -7234
rect 18658 -7628 18718 -7238
rect 19156 -7543 19216 -6968
rect 19520 -7064 19592 -7060
rect 19520 -7116 19530 -7064
rect 19582 -7116 19592 -7064
rect 19520 -7120 19592 -7116
rect 19526 -7380 19586 -7120
rect 19674 -7170 19734 -6880
rect 19668 -7174 19740 -7170
rect 19668 -7226 19678 -7174
rect 19730 -7226 19740 -7174
rect 19668 -7230 19740 -7226
rect 19520 -7384 19592 -7380
rect 19520 -7436 19530 -7384
rect 19582 -7436 19592 -7384
rect 19520 -7440 19592 -7436
rect 19672 -7382 19744 -7378
rect 19672 -7434 19682 -7382
rect 19734 -7434 19744 -7382
rect 19672 -7438 19744 -7434
rect 19678 -7616 19738 -7438
rect 20180 -7543 20240 -6968
rect 20694 -7280 20754 -6888
rect 20688 -7284 20760 -7280
rect 20688 -7336 20698 -7284
rect 20750 -7336 20760 -7284
rect 20688 -7340 20760 -7336
rect 21186 -7537 21246 -6962
rect 21714 -7170 21774 -6876
rect 22854 -7170 22914 -4402
rect 22996 -4574 23056 -1854
rect 24716 676 24828 714
rect 24716 642 24755 676
rect 24789 642 24828 676
rect 24716 604 24828 642
rect 24716 570 24755 604
rect 24789 570 24828 604
rect 24716 532 24828 570
rect 24716 498 24755 532
rect 24789 498 24828 532
rect 24716 460 24828 498
rect 24716 426 24755 460
rect 24789 426 24828 460
rect 24716 388 24828 426
rect 24716 354 24755 388
rect 24789 354 24828 388
rect 24716 316 24828 354
rect 24716 282 24755 316
rect 24789 282 24828 316
rect 24716 244 24828 282
rect 24716 210 24755 244
rect 24789 210 24828 244
rect 24716 172 24828 210
rect 24716 138 24755 172
rect 24789 138 24828 172
rect 24716 100 24828 138
rect 24716 66 24755 100
rect 24789 66 24828 100
rect 24716 28 24828 66
rect 24716 -6 24755 28
rect 24789 -6 24828 28
rect 24716 -44 24828 -6
rect 24716 -78 24755 -44
rect 24789 -78 24828 -44
rect 24716 -116 24828 -78
rect 24716 -150 24755 -116
rect 24789 -150 24828 -116
rect 24716 -188 24828 -150
rect 24716 -222 24755 -188
rect 24789 -222 24828 -188
rect 24716 -260 24828 -222
rect 24716 -294 24755 -260
rect 24789 -294 24828 -260
rect 24716 -332 24828 -294
rect 24716 -366 24755 -332
rect 24789 -366 24828 -332
rect 24716 -404 24828 -366
rect 24716 -438 24755 -404
rect 24789 -438 24828 -404
rect 24716 -476 24828 -438
rect 24716 -510 24755 -476
rect 24789 -510 24828 -476
rect 24716 -548 24828 -510
rect 24716 -582 24755 -548
rect 24789 -582 24828 -548
rect 24716 -620 24828 -582
rect 24716 -654 24755 -620
rect 24789 -654 24828 -620
rect 24716 -692 24828 -654
rect 24716 -726 24755 -692
rect 24789 -726 24828 -692
rect 24716 -764 24828 -726
rect 24716 -798 24755 -764
rect 24789 -798 24828 -764
rect 24716 -836 24828 -798
rect 24716 -870 24755 -836
rect 24789 -870 24828 -836
rect 24716 -908 24828 -870
rect 24716 -942 24755 -908
rect 24789 -942 24828 -908
rect 24716 -980 24828 -942
rect 24716 -1014 24755 -980
rect 24789 -1014 24828 -980
rect 24716 -1052 24828 -1014
rect 24716 -1086 24755 -1052
rect 24789 -1086 24828 -1052
rect 24716 -1124 24828 -1086
rect 24716 -1158 24755 -1124
rect 24789 -1158 24828 -1124
rect 24716 -1196 24828 -1158
rect 24716 -1230 24755 -1196
rect 24789 -1230 24828 -1196
rect 24716 -1268 24828 -1230
rect 24716 -1302 24755 -1268
rect 24789 -1302 24828 -1268
rect 24716 -1340 24828 -1302
rect 24716 -1374 24755 -1340
rect 24789 -1374 24828 -1340
rect 24716 -1412 24828 -1374
rect 24716 -1446 24755 -1412
rect 24789 -1446 24828 -1412
rect 24716 -1484 24828 -1446
rect 24716 -1518 24755 -1484
rect 24789 -1518 24828 -1484
rect 24716 -1556 24828 -1518
rect 24716 -1590 24755 -1556
rect 24789 -1590 24828 -1556
rect 24716 -1628 24828 -1590
rect 24716 -1662 24755 -1628
rect 24789 -1662 24828 -1628
rect 24716 -1700 24828 -1662
rect 24716 -1734 24755 -1700
rect 24789 -1734 24828 -1700
rect 24716 -1772 24828 -1734
rect 24716 -1806 24755 -1772
rect 24789 -1806 24828 -1772
rect 24716 -1844 24828 -1806
rect 24716 -1878 24755 -1844
rect 24789 -1878 24828 -1844
rect 24716 -1916 24828 -1878
rect 24716 -1950 24755 -1916
rect 24789 -1950 24828 -1916
rect 24716 -1988 24828 -1950
rect 24716 -2022 24755 -1988
rect 24789 -2022 24828 -1988
rect 24716 -2060 24828 -2022
rect 24716 -2094 24755 -2060
rect 24789 -2094 24828 -2060
rect 24716 -2132 24828 -2094
rect 24716 -2166 24755 -2132
rect 24789 -2166 24828 -2132
rect 24716 -2204 24828 -2166
rect 24716 -2238 24755 -2204
rect 24789 -2238 24828 -2204
rect 24716 -2276 24828 -2238
rect 24716 -2310 24755 -2276
rect 24789 -2310 24828 -2276
rect 24716 -2348 24828 -2310
rect 24716 -2382 24755 -2348
rect 24789 -2382 24828 -2348
rect 24716 -2420 24828 -2382
rect 24716 -2454 24755 -2420
rect 24789 -2454 24828 -2420
rect 24716 -2492 24828 -2454
rect 24716 -2526 24755 -2492
rect 24789 -2526 24828 -2492
rect 24716 -2564 24828 -2526
rect 24716 -2598 24755 -2564
rect 24789 -2598 24828 -2564
rect 24716 -2636 24828 -2598
rect 24716 -2670 24755 -2636
rect 24789 -2670 24828 -2636
rect 24716 -2708 24828 -2670
rect 24716 -2742 24755 -2708
rect 24789 -2742 24828 -2708
rect 24716 -2780 24828 -2742
rect 24716 -2814 24755 -2780
rect 24789 -2814 24828 -2780
rect 24716 -2852 24828 -2814
rect 24716 -2886 24755 -2852
rect 24789 -2886 24828 -2852
rect 24716 -2924 24828 -2886
rect 24716 -2958 24755 -2924
rect 24789 -2958 24828 -2924
rect 24716 -2996 24828 -2958
rect 24716 -3030 24755 -2996
rect 24789 -3030 24828 -2996
rect 24716 -3068 24828 -3030
rect 24716 -3102 24755 -3068
rect 24789 -3102 24828 -3068
rect 24716 -3140 24828 -3102
rect 24716 -3174 24755 -3140
rect 24789 -3174 24828 -3140
rect 24716 -3212 24828 -3174
rect 24716 -3246 24755 -3212
rect 24789 -3246 24828 -3212
rect 24716 -3284 24828 -3246
rect 24716 -3318 24755 -3284
rect 24789 -3318 24828 -3284
rect 24716 -3356 24828 -3318
rect 24716 -3390 24755 -3356
rect 24789 -3390 24828 -3356
rect 24716 -3428 24828 -3390
rect 24716 -3462 24755 -3428
rect 24789 -3462 24828 -3428
rect 24716 -3500 24828 -3462
rect 24716 -3534 24755 -3500
rect 24789 -3534 24828 -3500
rect 24716 -3572 24828 -3534
rect 24716 -3606 24755 -3572
rect 24789 -3606 24828 -3572
rect 24716 -3644 24828 -3606
rect 24716 -3678 24755 -3644
rect 24789 -3678 24828 -3644
rect 24716 -3716 24828 -3678
rect 24716 -3750 24755 -3716
rect 24789 -3750 24828 -3716
rect 24716 -3788 24828 -3750
rect 24716 -3822 24755 -3788
rect 24789 -3822 24828 -3788
rect 24716 -3860 24828 -3822
rect 24716 -3894 24755 -3860
rect 24789 -3894 24828 -3860
rect 24716 -3932 24828 -3894
rect 24716 -3966 24755 -3932
rect 24789 -3966 24828 -3932
rect 24716 -4004 24828 -3966
rect 24716 -4038 24755 -4004
rect 24789 -4038 24828 -4004
rect 24716 -4076 24828 -4038
rect 24716 -4110 24755 -4076
rect 24789 -4110 24828 -4076
rect 24716 -4148 24828 -4110
rect 24716 -4182 24755 -4148
rect 24789 -4182 24828 -4148
rect 23284 -4214 23356 -4210
rect 23284 -4266 23294 -4214
rect 23346 -4266 23356 -4214
rect 23284 -4270 23356 -4266
rect 24716 -4220 24828 -4182
rect 24716 -4254 24755 -4220
rect 24789 -4254 24828 -4220
rect 22996 -4626 23000 -4574
rect 23052 -4626 23056 -4574
rect 22996 -4636 23056 -4626
rect 23132 -4874 23204 -4870
rect 23132 -4926 23142 -4874
rect 23194 -4926 23204 -4874
rect 23132 -4930 23204 -4926
rect 22972 -6016 23044 -6012
rect 22972 -6068 22982 -6016
rect 23034 -6068 23044 -6016
rect 22972 -6072 23044 -6068
rect 21708 -7174 21780 -7170
rect 21708 -7226 21718 -7174
rect 21770 -7226 21780 -7174
rect 21708 -7230 21780 -7226
rect 22848 -7174 22920 -7170
rect 22848 -7226 22858 -7174
rect 22910 -7226 22920 -7174
rect 22848 -7230 22920 -7226
rect 21706 -7382 21778 -7378
rect 21706 -7434 21716 -7382
rect 21768 -7434 21778 -7382
rect 21706 -7438 21778 -7434
rect 21712 -7620 21772 -7438
rect 8480 -8330 8540 -8144
rect 8474 -8334 8546 -8330
rect 8474 -8386 8484 -8334
rect 8536 -8386 8546 -8334
rect 8474 -8390 8546 -8386
rect 7306 -8542 7378 -8538
rect 7306 -8594 7316 -8542
rect 7368 -8594 7378 -8542
rect 7306 -8598 7378 -8594
rect 7462 -8696 8538 -8636
rect 7462 -8890 7522 -8696
rect 7976 -8792 8036 -8696
rect 8478 -8878 8538 -8696
rect 8972 -8792 9032 -8218
rect 9488 -8644 9560 -8640
rect 9488 -8696 9498 -8644
rect 9550 -8696 9560 -8644
rect 9488 -8700 9560 -8696
rect 9494 -8878 9554 -8700
rect 10010 -8792 10070 -8218
rect 10516 -8330 10576 -8148
rect 10510 -8334 10582 -8330
rect 10510 -8386 10520 -8334
rect 10572 -8386 10582 -8334
rect 10510 -8390 10582 -8386
rect 10516 -8438 10576 -8390
rect 10510 -8442 10582 -8438
rect 10510 -8494 10520 -8442
rect 10572 -8494 10582 -8442
rect 10510 -8498 10582 -8494
rect 11016 -8488 11076 -8218
rect 11534 -8322 11594 -8153
rect 12052 -8322 12112 -8229
rect 12548 -8322 12608 -8138
rect 13064 -8322 13124 -8232
rect 11528 -8326 11600 -8322
rect 11528 -8378 11538 -8326
rect 11590 -8378 11600 -8326
rect 11528 -8382 11600 -8378
rect 12052 -8382 13124 -8322
rect 13330 -8326 13402 -8322
rect 13330 -8378 13340 -8326
rect 13392 -8378 13402 -8326
rect 13570 -8328 13630 -8142
rect 13330 -8382 13402 -8378
rect 13564 -8332 13636 -8328
rect 11016 -8548 11792 -8488
rect 11016 -8792 11076 -8548
rect 11522 -8644 11594 -8640
rect 11522 -8696 11532 -8644
rect 11584 -8696 11594 -8644
rect 11732 -8652 11792 -8548
rect 11522 -8700 11594 -8696
rect 11726 -8656 11798 -8652
rect 11528 -8882 11588 -8700
rect 11726 -8708 11736 -8656
rect 11788 -8708 11798 -8656
rect 11726 -8712 11798 -8708
rect 12548 -8910 12608 -8382
rect 13336 -8592 13396 -8382
rect 13564 -8384 13574 -8332
rect 13626 -8384 13636 -8332
rect 13564 -8388 13636 -8384
rect 14066 -8450 14126 -8228
rect 15094 -8450 15154 -8234
rect 15606 -8328 15666 -8146
rect 15600 -8332 15672 -8328
rect 15600 -8384 15610 -8332
rect 15662 -8384 15672 -8332
rect 15600 -8388 15672 -8384
rect 14066 -8510 15154 -8450
rect 15598 -8442 15670 -8438
rect 15598 -8494 15608 -8442
rect 15660 -8494 15670 -8442
rect 15598 -8498 15670 -8494
rect 13336 -8652 14644 -8592
rect 14584 -8904 14644 -8652
rect 15094 -8656 15154 -8510
rect 15094 -8708 15098 -8656
rect 15150 -8708 15154 -8656
rect 15094 -8790 15154 -8708
rect 15604 -8916 15664 -8498
rect 16110 -8656 16170 -8226
rect 17140 -8324 17200 -8231
rect 17636 -8324 17696 -8140
rect 18152 -8324 18212 -8234
rect 17140 -8384 18212 -8324
rect 18660 -8326 18720 -8140
rect 18654 -8330 18726 -8326
rect 18654 -8382 18664 -8330
rect 18716 -8382 18726 -8330
rect 16110 -8708 16114 -8656
rect 16166 -8708 16170 -8656
rect 16110 -8718 16170 -8708
rect 17636 -8890 17696 -8384
rect 18654 -8386 18726 -8382
rect 19168 -8646 19228 -8218
rect 19676 -8644 19748 -8640
rect 19168 -8656 19230 -8646
rect 19168 -8708 19174 -8656
rect 19226 -8708 19230 -8656
rect 19676 -8696 19686 -8644
rect 19738 -8696 19748 -8644
rect 19676 -8700 19748 -8696
rect 19168 -8718 19230 -8708
rect 19168 -8792 19228 -8718
rect 19682 -8878 19742 -8700
rect 20192 -8792 20252 -8218
rect 20696 -8326 20756 -8144
rect 20690 -8330 20762 -8326
rect 20690 -8382 20700 -8330
rect 20752 -8382 20762 -8330
rect 20690 -8386 20762 -8382
rect 21198 -8786 21258 -8212
rect 21712 -8330 21772 -8136
rect 22226 -8330 22286 -8234
rect 22728 -8330 22788 -8148
rect 21712 -8390 22788 -8330
rect 22854 -8438 22914 -7230
rect 22978 -7378 23038 -6072
rect 22972 -7382 23044 -7378
rect 22972 -7434 22982 -7382
rect 23034 -7434 23044 -7382
rect 22972 -7438 23044 -7434
rect 22848 -8442 22920 -8438
rect 22848 -8494 22858 -8442
rect 22910 -8494 22920 -8442
rect 22848 -8498 22920 -8494
rect 21710 -8644 21782 -8640
rect 21710 -8696 21720 -8644
rect 21772 -8696 21782 -8644
rect 21710 -8700 21782 -8696
rect 21716 -8882 21776 -8700
rect 8476 -9588 8536 -9402
rect 8470 -9592 8542 -9588
rect 8470 -9644 8480 -9592
rect 8532 -9644 8542 -9592
rect 8470 -9648 8542 -9644
rect 8984 -9702 9044 -9490
rect 10008 -9702 10068 -9482
rect 10512 -9588 10572 -9406
rect 10506 -9592 10578 -9588
rect 10506 -9644 10516 -9592
rect 10568 -9644 10578 -9592
rect 10506 -9648 10578 -9644
rect 11014 -9702 11074 -9482
rect 7174 -9722 7246 -9718
rect 7174 -9774 7184 -9722
rect 7236 -9774 7246 -9722
rect 7174 -9778 7246 -9774
rect 8984 -9762 11074 -9702
rect 2332 -9850 6858 -9846
rect 2332 -9902 2340 -9850
rect 2392 -9902 6858 -9850
rect 2332 -9906 6858 -9902
rect 2336 -9912 2396 -9906
rect 2216 -9964 2276 -9958
rect 7180 -9964 7240 -9778
rect 2216 -9968 7240 -9964
rect 2216 -10020 2220 -9968
rect 2272 -10020 7240 -9968
rect 2216 -10024 7240 -10020
rect 2216 -10030 2276 -10024
rect 1770 -10082 1830 -10076
rect 8984 -10082 9044 -9762
rect 11014 -9972 11074 -9762
rect 11534 -9858 11594 -9392
rect 12052 -9582 12112 -9487
rect 12548 -9582 12608 -9396
rect 13064 -9582 13124 -9490
rect 13570 -9582 13630 -9384
rect 14080 -9582 14140 -9490
rect 16106 -9582 16166 -9490
rect 16622 -9582 16682 -9400
rect 17140 -9582 17200 -9489
rect 17636 -9582 17696 -9398
rect 18152 -9582 18212 -9492
rect 12052 -9642 18212 -9582
rect 18664 -9588 18724 -9402
rect 18658 -9592 18730 -9588
rect 18658 -9644 18668 -9592
rect 18720 -9644 18730 -9592
rect 18658 -9648 18730 -9644
rect 19172 -9700 19232 -9474
rect 20192 -9700 20252 -9482
rect 20700 -9588 20760 -9406
rect 20694 -9592 20766 -9588
rect 20694 -9644 20704 -9592
rect 20756 -9644 20766 -9592
rect 20694 -9648 20766 -9644
rect 21194 -9700 21254 -9482
rect 21714 -9584 21774 -9390
rect 22228 -9584 22288 -9488
rect 22730 -9584 22790 -9402
rect 21714 -9644 22790 -9584
rect 19172 -9760 21254 -9700
rect 11528 -9862 11600 -9858
rect 11528 -9914 11538 -9862
rect 11590 -9914 11600 -9862
rect 11528 -9918 11600 -9914
rect 19172 -9972 19232 -9760
rect 23138 -9858 23198 -4930
rect 23290 -6126 23350 -4270
rect 24716 -4292 24828 -4254
rect 24716 -4326 24755 -4292
rect 24789 -4326 24828 -4292
rect 24716 -4364 24828 -4326
rect 24716 -4398 24755 -4364
rect 24789 -4398 24828 -4364
rect 24716 -4436 24828 -4398
rect 24716 -4470 24755 -4436
rect 24789 -4470 24828 -4436
rect 24716 -4508 24828 -4470
rect 24716 -4542 24755 -4508
rect 24789 -4542 24828 -4508
rect 24716 -4580 24828 -4542
rect 24716 -4614 24755 -4580
rect 24789 -4614 24828 -4580
rect 24716 -4652 24828 -4614
rect 24716 -4686 24755 -4652
rect 24789 -4686 24828 -4652
rect 24716 -4724 24828 -4686
rect 24716 -4758 24755 -4724
rect 24789 -4758 24828 -4724
rect 24716 -4796 24828 -4758
rect 24716 -4830 24755 -4796
rect 24789 -4830 24828 -4796
rect 24716 -4868 24828 -4830
rect 24716 -4902 24755 -4868
rect 24789 -4902 24828 -4868
rect 24716 -4940 24828 -4902
rect 24716 -4974 24755 -4940
rect 24789 -4974 24828 -4940
rect 24716 -5012 24828 -4974
rect 24716 -5046 24755 -5012
rect 24789 -5046 24828 -5012
rect 24716 -5084 24828 -5046
rect 24716 -5118 24755 -5084
rect 24789 -5118 24828 -5084
rect 24716 -5156 24828 -5118
rect 24716 -5190 24755 -5156
rect 24789 -5190 24828 -5156
rect 24716 -5228 24828 -5190
rect 24716 -5262 24755 -5228
rect 24789 -5262 24828 -5228
rect 24716 -5300 24828 -5262
rect 24716 -5334 24755 -5300
rect 24789 -5334 24828 -5300
rect 24716 -5372 24828 -5334
rect 24716 -5406 24755 -5372
rect 24789 -5406 24828 -5372
rect 24716 -5444 24828 -5406
rect 24716 -5478 24755 -5444
rect 24789 -5478 24828 -5444
rect 24716 -5516 24828 -5478
rect 24716 -5550 24755 -5516
rect 24789 -5550 24828 -5516
rect 24716 -5588 24828 -5550
rect 24716 -5622 24755 -5588
rect 24789 -5622 24828 -5588
rect 24716 -5660 24828 -5622
rect 24716 -5694 24755 -5660
rect 24789 -5694 24828 -5660
rect 24716 -5732 24828 -5694
rect 24716 -5766 24755 -5732
rect 24789 -5766 24828 -5732
rect 24716 -5804 24828 -5766
rect 24716 -5838 24755 -5804
rect 24789 -5838 24828 -5804
rect 24716 -5876 24828 -5838
rect 24716 -5910 24755 -5876
rect 24789 -5910 24828 -5876
rect 24716 -5948 24828 -5910
rect 24716 -5982 24755 -5948
rect 24789 -5982 24828 -5948
rect 24716 -6020 24828 -5982
rect 24716 -6054 24755 -6020
rect 24789 -6054 24828 -6020
rect 24716 -6092 24828 -6054
rect 24716 -6126 24755 -6092
rect 24789 -6126 24828 -6092
rect 23284 -6130 23356 -6126
rect 23284 -6182 23294 -6130
rect 23346 -6182 23356 -6130
rect 23284 -6186 23356 -6182
rect 24716 -6164 24828 -6126
rect 24716 -6198 24755 -6164
rect 24789 -6198 24828 -6164
rect 24716 -6236 24828 -6198
rect 24716 -6270 24755 -6236
rect 24789 -6270 24828 -6236
rect 24716 -6308 24828 -6270
rect 24716 -6342 24755 -6308
rect 24789 -6342 24828 -6308
rect 24716 -6380 24828 -6342
rect 24716 -6414 24755 -6380
rect 24789 -6414 24828 -6380
rect 24716 -6452 24828 -6414
rect 24716 -6486 24755 -6452
rect 24789 -6486 24828 -6452
rect 24716 -6524 24828 -6486
rect 24716 -6558 24755 -6524
rect 24789 -6558 24828 -6524
rect 24716 -6596 24828 -6558
rect 24716 -6630 24755 -6596
rect 24789 -6630 24828 -6596
rect 24716 -6668 24828 -6630
rect 24716 -6702 24755 -6668
rect 24789 -6702 24828 -6668
rect 24716 -6740 24828 -6702
rect 24716 -6774 24755 -6740
rect 24789 -6774 24828 -6740
rect 24716 -6812 24828 -6774
rect 24716 -6846 24755 -6812
rect 24789 -6846 24828 -6812
rect 24716 -6884 24828 -6846
rect 24716 -6918 24755 -6884
rect 24789 -6918 24828 -6884
rect 24716 -6956 24828 -6918
rect 24716 -6990 24755 -6956
rect 24789 -6990 24828 -6956
rect 24716 -7028 24828 -6990
rect 24716 -7062 24755 -7028
rect 24789 -7062 24828 -7028
rect 24716 -7100 24828 -7062
rect 24716 -7134 24755 -7100
rect 24789 -7134 24828 -7100
rect 24716 -7172 24828 -7134
rect 24716 -7206 24755 -7172
rect 24789 -7206 24828 -7172
rect 24716 -7244 24828 -7206
rect 24716 -7278 24755 -7244
rect 24789 -7278 24828 -7244
rect 24716 -7316 24828 -7278
rect 24716 -7350 24755 -7316
rect 24789 -7350 24828 -7316
rect 24716 -7388 24828 -7350
rect 24716 -7422 24755 -7388
rect 24789 -7422 24828 -7388
rect 24716 -7460 24828 -7422
rect 24716 -7494 24755 -7460
rect 24789 -7494 24828 -7460
rect 24716 -7532 24828 -7494
rect 24716 -7566 24755 -7532
rect 24789 -7566 24828 -7532
rect 24716 -7604 24828 -7566
rect 24716 -7638 24755 -7604
rect 24789 -7638 24828 -7604
rect 24716 -7676 24828 -7638
rect 24716 -7710 24755 -7676
rect 24789 -7710 24828 -7676
rect 24716 -7748 24828 -7710
rect 24716 -7782 24755 -7748
rect 24789 -7782 24828 -7748
rect 24716 -7820 24828 -7782
rect 24716 -7854 24755 -7820
rect 24789 -7854 24828 -7820
rect 24716 -7892 24828 -7854
rect 24716 -7926 24755 -7892
rect 24789 -7926 24828 -7892
rect 24716 -7964 24828 -7926
rect 24716 -7998 24755 -7964
rect 24789 -7998 24828 -7964
rect 24716 -8036 24828 -7998
rect 24716 -8070 24755 -8036
rect 24789 -8070 24828 -8036
rect 24716 -8108 24828 -8070
rect 24716 -8142 24755 -8108
rect 24789 -8142 24828 -8108
rect 24716 -8180 24828 -8142
rect 24716 -8214 24755 -8180
rect 24789 -8214 24828 -8180
rect 24716 -8252 24828 -8214
rect 24716 -8286 24755 -8252
rect 24789 -8286 24828 -8252
rect 24716 -8324 24828 -8286
rect 24716 -8358 24755 -8324
rect 24789 -8358 24828 -8324
rect 24716 -8396 24828 -8358
rect 24716 -8430 24755 -8396
rect 24789 -8430 24828 -8396
rect 24716 -8468 24828 -8430
rect 24716 -8502 24755 -8468
rect 24789 -8502 24828 -8468
rect 24716 -8540 24828 -8502
rect 24716 -8574 24755 -8540
rect 24789 -8574 24828 -8540
rect 24716 -8612 24828 -8574
rect 24716 -8646 24755 -8612
rect 24789 -8646 24828 -8612
rect 24716 -8684 24828 -8646
rect 24716 -8718 24755 -8684
rect 24789 -8718 24828 -8684
rect 24716 -8756 24828 -8718
rect 24716 -8790 24755 -8756
rect 24789 -8790 24828 -8756
rect 24716 -8828 24828 -8790
rect 24716 -8862 24755 -8828
rect 24789 -8862 24828 -8828
rect 24716 -8900 24828 -8862
rect 24716 -8934 24755 -8900
rect 24789 -8934 24828 -8900
rect 24716 -8972 24828 -8934
rect 24716 -9006 24755 -8972
rect 24789 -9006 24828 -8972
rect 24716 -9044 24828 -9006
rect 24716 -9078 24755 -9044
rect 24789 -9078 24828 -9044
rect 24716 -9116 24828 -9078
rect 24716 -9150 24755 -9116
rect 24789 -9150 24828 -9116
rect 24716 -9188 24828 -9150
rect 24716 -9222 24755 -9188
rect 24789 -9222 24828 -9188
rect 24716 -9260 24828 -9222
rect 24716 -9294 24755 -9260
rect 24789 -9294 24828 -9260
rect 24716 -9332 24828 -9294
rect 24716 -9366 24755 -9332
rect 24789 -9366 24828 -9332
rect 24716 -9404 24828 -9366
rect 24716 -9438 24755 -9404
rect 24789 -9438 24828 -9404
rect 24716 -9476 24828 -9438
rect 24716 -9510 24755 -9476
rect 24789 -9510 24828 -9476
rect 24716 -9548 24828 -9510
rect 24716 -9582 24755 -9548
rect 24789 -9582 24828 -9548
rect 24716 -9620 24828 -9582
rect 24716 -9654 24755 -9620
rect 24789 -9654 24828 -9620
rect 24716 -9692 24828 -9654
rect 24716 -9726 24755 -9692
rect 24789 -9726 24828 -9692
rect 23132 -9862 23204 -9858
rect 23132 -9914 23142 -9862
rect 23194 -9914 23204 -9862
rect 23132 -9918 23204 -9914
rect 11014 -10032 19232 -9972
rect 1770 -10086 9044 -10082
rect 1770 -10138 1774 -10086
rect 1826 -10138 9044 -10086
rect 1770 -10142 9044 -10138
rect 1770 -10148 1830 -10142
rect 24716 -10242 24828 -9726
rect 372 -10281 24828 -10242
rect 372 -10315 487 -10281
rect 521 -10315 559 -10281
rect 593 -10315 631 -10281
rect 665 -10315 703 -10281
rect 737 -10315 775 -10281
rect 809 -10315 847 -10281
rect 881 -10315 919 -10281
rect 953 -10315 991 -10281
rect 1025 -10315 1063 -10281
rect 1097 -10315 1135 -10281
rect 1169 -10315 1207 -10281
rect 1241 -10315 1279 -10281
rect 1313 -10315 1351 -10281
rect 1385 -10315 1423 -10281
rect 1457 -10315 1495 -10281
rect 1529 -10315 1567 -10281
rect 1601 -10315 1639 -10281
rect 1673 -10315 1711 -10281
rect 1745 -10315 1783 -10281
rect 1817 -10315 1855 -10281
rect 1889 -10315 1927 -10281
rect 1961 -10315 1999 -10281
rect 2033 -10315 2071 -10281
rect 2105 -10315 2143 -10281
rect 2177 -10315 2215 -10281
rect 2249 -10315 2287 -10281
rect 2321 -10315 2359 -10281
rect 2393 -10315 2431 -10281
rect 2465 -10315 2503 -10281
rect 2537 -10315 2575 -10281
rect 2609 -10315 2647 -10281
rect 2681 -10315 2719 -10281
rect 2753 -10315 2791 -10281
rect 2825 -10315 2863 -10281
rect 2897 -10315 2935 -10281
rect 2969 -10315 3007 -10281
rect 3041 -10315 3079 -10281
rect 3113 -10315 3151 -10281
rect 3185 -10315 3223 -10281
rect 3257 -10315 3295 -10281
rect 3329 -10315 3367 -10281
rect 3401 -10315 3439 -10281
rect 3473 -10315 3511 -10281
rect 3545 -10315 3583 -10281
rect 3617 -10315 3655 -10281
rect 3689 -10315 3727 -10281
rect 3761 -10315 3799 -10281
rect 3833 -10315 3871 -10281
rect 3905 -10315 3943 -10281
rect 3977 -10315 4015 -10281
rect 4049 -10315 4087 -10281
rect 4121 -10315 4159 -10281
rect 4193 -10315 4231 -10281
rect 4265 -10315 4303 -10281
rect 4337 -10315 4375 -10281
rect 4409 -10315 4447 -10281
rect 4481 -10315 4519 -10281
rect 4553 -10315 4591 -10281
rect 4625 -10315 4663 -10281
rect 4697 -10315 4735 -10281
rect 4769 -10315 4807 -10281
rect 4841 -10315 4879 -10281
rect 4913 -10315 4951 -10281
rect 4985 -10315 5023 -10281
rect 5057 -10315 5095 -10281
rect 5129 -10315 5167 -10281
rect 5201 -10315 5239 -10281
rect 5273 -10315 5311 -10281
rect 5345 -10315 5383 -10281
rect 5417 -10315 5455 -10281
rect 5489 -10315 5527 -10281
rect 5561 -10315 5599 -10281
rect 5633 -10315 5671 -10281
rect 5705 -10315 5743 -10281
rect 5777 -10315 5815 -10281
rect 5849 -10315 5887 -10281
rect 5921 -10315 5959 -10281
rect 5993 -10315 6031 -10281
rect 6065 -10315 6103 -10281
rect 6137 -10315 6175 -10281
rect 6209 -10315 6247 -10281
rect 6281 -10315 6319 -10281
rect 6353 -10315 6391 -10281
rect 6425 -10315 6463 -10281
rect 6497 -10315 6535 -10281
rect 6569 -10315 6607 -10281
rect 6641 -10315 6679 -10281
rect 6713 -10315 6751 -10281
rect 6785 -10315 6823 -10281
rect 6857 -10315 6895 -10281
rect 6929 -10315 6967 -10281
rect 7001 -10315 7039 -10281
rect 7073 -10315 7111 -10281
rect 7145 -10315 7183 -10281
rect 7217 -10315 7255 -10281
rect 7289 -10315 7327 -10281
rect 7361 -10315 7399 -10281
rect 7433 -10315 7471 -10281
rect 7505 -10315 7543 -10281
rect 7577 -10315 7615 -10281
rect 7649 -10315 7687 -10281
rect 7721 -10315 7759 -10281
rect 7793 -10315 7831 -10281
rect 7865 -10315 7903 -10281
rect 7937 -10315 7975 -10281
rect 8009 -10315 8047 -10281
rect 8081 -10315 8119 -10281
rect 8153 -10315 8191 -10281
rect 8225 -10315 8263 -10281
rect 8297 -10315 8335 -10281
rect 8369 -10315 8407 -10281
rect 8441 -10315 8479 -10281
rect 8513 -10315 8551 -10281
rect 8585 -10315 8623 -10281
rect 8657 -10315 8695 -10281
rect 8729 -10315 8767 -10281
rect 8801 -10315 8839 -10281
rect 8873 -10315 8911 -10281
rect 8945 -10315 8983 -10281
rect 9017 -10315 9055 -10281
rect 9089 -10315 9127 -10281
rect 9161 -10315 9199 -10281
rect 9233 -10315 9271 -10281
rect 9305 -10315 9343 -10281
rect 9377 -10315 9415 -10281
rect 9449 -10315 9487 -10281
rect 9521 -10315 9559 -10281
rect 9593 -10315 9631 -10281
rect 9665 -10315 9703 -10281
rect 9737 -10315 9775 -10281
rect 9809 -10315 9847 -10281
rect 9881 -10315 9919 -10281
rect 9953 -10315 9991 -10281
rect 10025 -10315 10063 -10281
rect 10097 -10315 10135 -10281
rect 10169 -10315 10207 -10281
rect 10241 -10315 10279 -10281
rect 10313 -10315 10351 -10281
rect 10385 -10315 10423 -10281
rect 10457 -10315 10495 -10281
rect 10529 -10315 10567 -10281
rect 10601 -10315 10639 -10281
rect 10673 -10315 10711 -10281
rect 10745 -10315 10783 -10281
rect 10817 -10315 10855 -10281
rect 10889 -10315 10927 -10281
rect 10961 -10315 10999 -10281
rect 11033 -10315 11071 -10281
rect 11105 -10315 11143 -10281
rect 11177 -10315 11215 -10281
rect 11249 -10315 11287 -10281
rect 11321 -10315 11359 -10281
rect 11393 -10315 11431 -10281
rect 11465 -10315 11503 -10281
rect 11537 -10315 11575 -10281
rect 11609 -10315 11647 -10281
rect 11681 -10315 11719 -10281
rect 11753 -10315 11791 -10281
rect 11825 -10315 11863 -10281
rect 11897 -10315 11935 -10281
rect 11969 -10315 12007 -10281
rect 12041 -10315 12079 -10281
rect 12113 -10315 12151 -10281
rect 12185 -10315 12223 -10281
rect 12257 -10315 12295 -10281
rect 12329 -10315 12367 -10281
rect 12401 -10315 12439 -10281
rect 12473 -10315 12511 -10281
rect 12545 -10315 12583 -10281
rect 12617 -10315 12655 -10281
rect 12689 -10315 12727 -10281
rect 12761 -10315 12799 -10281
rect 12833 -10315 12871 -10281
rect 12905 -10315 12943 -10281
rect 12977 -10315 13015 -10281
rect 13049 -10315 13087 -10281
rect 13121 -10315 13159 -10281
rect 13193 -10315 13231 -10281
rect 13265 -10315 13303 -10281
rect 13337 -10315 13375 -10281
rect 13409 -10315 13447 -10281
rect 13481 -10315 13519 -10281
rect 13553 -10315 13591 -10281
rect 13625 -10315 13663 -10281
rect 13697 -10315 13735 -10281
rect 13769 -10315 13807 -10281
rect 13841 -10315 13879 -10281
rect 13913 -10315 13951 -10281
rect 13985 -10315 14023 -10281
rect 14057 -10315 14095 -10281
rect 14129 -10315 14167 -10281
rect 14201 -10315 14239 -10281
rect 14273 -10315 14311 -10281
rect 14345 -10315 14383 -10281
rect 14417 -10315 14455 -10281
rect 14489 -10315 14527 -10281
rect 14561 -10315 14599 -10281
rect 14633 -10315 14671 -10281
rect 14705 -10315 14743 -10281
rect 14777 -10315 14815 -10281
rect 14849 -10315 14887 -10281
rect 14921 -10315 14959 -10281
rect 14993 -10315 15031 -10281
rect 15065 -10315 15103 -10281
rect 15137 -10315 15175 -10281
rect 15209 -10315 15247 -10281
rect 15281 -10315 15319 -10281
rect 15353 -10315 15391 -10281
rect 15425 -10315 15463 -10281
rect 15497 -10315 15535 -10281
rect 15569 -10315 15607 -10281
rect 15641 -10315 15679 -10281
rect 15713 -10315 15751 -10281
rect 15785 -10315 15823 -10281
rect 15857 -10315 15895 -10281
rect 15929 -10315 15967 -10281
rect 16001 -10315 16039 -10281
rect 16073 -10315 16111 -10281
rect 16145 -10315 16183 -10281
rect 16217 -10315 16255 -10281
rect 16289 -10315 16327 -10281
rect 16361 -10315 16399 -10281
rect 16433 -10315 16471 -10281
rect 16505 -10315 16543 -10281
rect 16577 -10315 16615 -10281
rect 16649 -10315 16687 -10281
rect 16721 -10315 16759 -10281
rect 16793 -10315 16831 -10281
rect 16865 -10315 16903 -10281
rect 16937 -10315 16975 -10281
rect 17009 -10315 17047 -10281
rect 17081 -10315 17119 -10281
rect 17153 -10315 17191 -10281
rect 17225 -10315 17263 -10281
rect 17297 -10315 17335 -10281
rect 17369 -10315 17407 -10281
rect 17441 -10315 17479 -10281
rect 17513 -10315 17551 -10281
rect 17585 -10315 17623 -10281
rect 17657 -10315 17695 -10281
rect 17729 -10315 17767 -10281
rect 17801 -10315 17839 -10281
rect 17873 -10315 17911 -10281
rect 17945 -10315 17983 -10281
rect 18017 -10315 18055 -10281
rect 18089 -10315 18127 -10281
rect 18161 -10315 18199 -10281
rect 18233 -10315 18271 -10281
rect 18305 -10315 18343 -10281
rect 18377 -10315 18415 -10281
rect 18449 -10315 18487 -10281
rect 18521 -10315 18559 -10281
rect 18593 -10315 18631 -10281
rect 18665 -10315 18703 -10281
rect 18737 -10315 18775 -10281
rect 18809 -10315 18847 -10281
rect 18881 -10315 18919 -10281
rect 18953 -10315 18991 -10281
rect 19025 -10315 19063 -10281
rect 19097 -10315 19135 -10281
rect 19169 -10315 19207 -10281
rect 19241 -10315 19279 -10281
rect 19313 -10315 19351 -10281
rect 19385 -10315 19423 -10281
rect 19457 -10315 19495 -10281
rect 19529 -10315 19567 -10281
rect 19601 -10315 19639 -10281
rect 19673 -10315 19711 -10281
rect 19745 -10315 19783 -10281
rect 19817 -10315 19855 -10281
rect 19889 -10315 19927 -10281
rect 19961 -10315 19999 -10281
rect 20033 -10315 20071 -10281
rect 20105 -10315 20143 -10281
rect 20177 -10315 20215 -10281
rect 20249 -10315 20287 -10281
rect 20321 -10315 20359 -10281
rect 20393 -10315 20431 -10281
rect 20465 -10315 20503 -10281
rect 20537 -10315 20575 -10281
rect 20609 -10315 20647 -10281
rect 20681 -10315 20719 -10281
rect 20753 -10315 20791 -10281
rect 20825 -10315 20863 -10281
rect 20897 -10315 20935 -10281
rect 20969 -10315 21007 -10281
rect 21041 -10315 21079 -10281
rect 21113 -10315 21151 -10281
rect 21185 -10315 21223 -10281
rect 21257 -10315 21295 -10281
rect 21329 -10315 21367 -10281
rect 21401 -10315 21439 -10281
rect 21473 -10315 21511 -10281
rect 21545 -10315 21583 -10281
rect 21617 -10315 21655 -10281
rect 21689 -10315 21727 -10281
rect 21761 -10315 21799 -10281
rect 21833 -10315 21871 -10281
rect 21905 -10315 21943 -10281
rect 21977 -10315 22015 -10281
rect 22049 -10315 22087 -10281
rect 22121 -10315 22159 -10281
rect 22193 -10315 22231 -10281
rect 22265 -10315 22303 -10281
rect 22337 -10315 22375 -10281
rect 22409 -10315 22447 -10281
rect 22481 -10315 22519 -10281
rect 22553 -10315 22591 -10281
rect 22625 -10315 22663 -10281
rect 22697 -10315 22735 -10281
rect 22769 -10315 22807 -10281
rect 22841 -10315 22879 -10281
rect 22913 -10315 22951 -10281
rect 22985 -10315 23023 -10281
rect 23057 -10315 23095 -10281
rect 23129 -10315 23167 -10281
rect 23201 -10315 23239 -10281
rect 23273 -10315 23311 -10281
rect 23345 -10315 23383 -10281
rect 23417 -10315 23455 -10281
rect 23489 -10315 23527 -10281
rect 23561 -10315 23599 -10281
rect 23633 -10315 23671 -10281
rect 23705 -10315 23743 -10281
rect 23777 -10315 23815 -10281
rect 23849 -10315 23887 -10281
rect 23921 -10315 23959 -10281
rect 23993 -10315 24031 -10281
rect 24065 -10315 24103 -10281
rect 24137 -10315 24175 -10281
rect 24209 -10315 24247 -10281
rect 24281 -10315 24319 -10281
rect 24353 -10315 24391 -10281
rect 24425 -10315 24463 -10281
rect 24497 -10315 24535 -10281
rect 24569 -10315 24607 -10281
rect 24641 -10315 24679 -10281
rect 24713 -10315 24828 -10281
rect 372 -10354 24828 -10315
rect -13992 -10646 -13618 -10402
rect -2878 -10646 -2722 -10402
rect -13992 -10978 -2722 -10646
rect -13992 -11172 -1640 -10978
rect -13992 -11211 24928 -11172
rect -13992 -11245 -12221 -11211
rect -12187 -11245 -12149 -11211
rect -12115 -11245 -12077 -11211
rect -12043 -11245 -12005 -11211
rect -11971 -11245 -11933 -11211
rect -11899 -11245 -11861 -11211
rect -11827 -11245 -11789 -11211
rect -11755 -11245 -11717 -11211
rect -11683 -11245 -11645 -11211
rect -11611 -11245 -11573 -11211
rect -11539 -11245 -11501 -11211
rect -11467 -11245 -11429 -11211
rect -11395 -11245 -11357 -11211
rect -11323 -11245 -11285 -11211
rect -11251 -11245 -11213 -11211
rect -11179 -11245 -11141 -11211
rect -11107 -11245 -11069 -11211
rect -11035 -11245 -10997 -11211
rect -10963 -11245 -10925 -11211
rect -10891 -11245 -10853 -11211
rect -10819 -11245 -10781 -11211
rect -10747 -11245 -10709 -11211
rect -10675 -11245 -10637 -11211
rect -10603 -11245 -10565 -11211
rect -10531 -11245 -10493 -11211
rect -10459 -11245 -10421 -11211
rect -10387 -11245 -10349 -11211
rect -10315 -11245 -10277 -11211
rect -10243 -11245 -10205 -11211
rect -10171 -11245 -10133 -11211
rect -10099 -11245 -10061 -11211
rect -10027 -11245 -9989 -11211
rect -9955 -11245 -9917 -11211
rect -9883 -11245 -9845 -11211
rect -9811 -11245 -9773 -11211
rect -9739 -11245 -9701 -11211
rect -9667 -11245 -9629 -11211
rect -9595 -11245 -9557 -11211
rect -9523 -11245 -9485 -11211
rect -9451 -11245 -9413 -11211
rect -9379 -11245 -9341 -11211
rect -9307 -11245 -9269 -11211
rect -9235 -11245 -9197 -11211
rect -9163 -11245 -9125 -11211
rect -9091 -11245 -9053 -11211
rect -9019 -11245 -8981 -11211
rect -8947 -11245 -8909 -11211
rect -8875 -11245 -8837 -11211
rect -8803 -11245 -8765 -11211
rect -8731 -11245 -8693 -11211
rect -8659 -11245 -8621 -11211
rect -8587 -11245 -8549 -11211
rect -8515 -11245 -8477 -11211
rect -8443 -11245 -8405 -11211
rect -8371 -11245 -8333 -11211
rect -8299 -11245 -8261 -11211
rect -8227 -11245 -8189 -11211
rect -8155 -11245 -8117 -11211
rect -8083 -11245 -8045 -11211
rect -8011 -11245 -7973 -11211
rect -7939 -11245 -7901 -11211
rect -7867 -11245 -7829 -11211
rect -7795 -11245 -7757 -11211
rect -7723 -11245 -7685 -11211
rect -7651 -11245 -7613 -11211
rect -7579 -11245 -7541 -11211
rect -7507 -11245 -7469 -11211
rect -7435 -11245 -7397 -11211
rect -7363 -11245 -7325 -11211
rect -7291 -11245 -7253 -11211
rect -7219 -11245 -7181 -11211
rect -7147 -11245 -7109 -11211
rect -7075 -11245 -7037 -11211
rect -7003 -11245 -6965 -11211
rect -6931 -11245 -6893 -11211
rect -6859 -11245 -6821 -11211
rect -6787 -11245 -6749 -11211
rect -6715 -11245 -6677 -11211
rect -6643 -11245 -6605 -11211
rect -6571 -11245 -6533 -11211
rect -6499 -11245 -6461 -11211
rect -6427 -11245 -6389 -11211
rect -6355 -11245 -6317 -11211
rect -6283 -11245 -6245 -11211
rect -6211 -11245 -6173 -11211
rect -6139 -11245 -6101 -11211
rect -6067 -11245 -6029 -11211
rect -5995 -11245 -5957 -11211
rect -5923 -11245 -5885 -11211
rect -5851 -11245 -5813 -11211
rect -5779 -11245 -5741 -11211
rect -5707 -11245 -5669 -11211
rect -5635 -11245 -5597 -11211
rect -5563 -11245 -5525 -11211
rect -5491 -11245 -5453 -11211
rect -5419 -11245 -5381 -11211
rect -5347 -11245 -5309 -11211
rect -5275 -11245 -5237 -11211
rect -5203 -11245 -5165 -11211
rect -5131 -11245 -5093 -11211
rect -5059 -11245 -5021 -11211
rect -4987 -11245 -4949 -11211
rect -4915 -11245 -4877 -11211
rect -4843 -11245 -4805 -11211
rect -4771 -11245 -4733 -11211
rect -4699 -11245 -4661 -11211
rect -4627 -11245 -4589 -11211
rect -4555 -11245 -4517 -11211
rect -4483 -11245 -4445 -11211
rect -4411 -11245 -4373 -11211
rect -4339 -11245 -4301 -11211
rect -4267 -11245 -4229 -11211
rect -4195 -11245 -4157 -11211
rect -4123 -11245 -4085 -11211
rect -4051 -11245 -4013 -11211
rect -3979 -11245 -3941 -11211
rect -3907 -11245 -3869 -11211
rect -3835 -11245 -3797 -11211
rect -3763 -11245 -3725 -11211
rect -3691 -11245 -3653 -11211
rect -3619 -11245 -3581 -11211
rect -3547 -11245 -3509 -11211
rect -3475 -11245 -3437 -11211
rect -3403 -11245 -3365 -11211
rect -3331 -11245 -3293 -11211
rect -3259 -11245 -3221 -11211
rect -3187 -11245 -3149 -11211
rect -3115 -11245 -3077 -11211
rect -3043 -11245 -3005 -11211
rect -2971 -11245 -2933 -11211
rect -2899 -11245 -2861 -11211
rect -2827 -11245 -2789 -11211
rect -2755 -11245 -2717 -11211
rect -2683 -11245 -2645 -11211
rect -2611 -11245 -2573 -11211
rect -2539 -11245 -2501 -11211
rect -2467 -11245 -2429 -11211
rect -2395 -11245 -2357 -11211
rect -2323 -11245 -2285 -11211
rect -2251 -11245 -2213 -11211
rect -2179 -11245 -2141 -11211
rect -2107 -11245 -2069 -11211
rect -2035 -11245 -1997 -11211
rect -1963 -11245 -1925 -11211
rect -1891 -11245 -1853 -11211
rect -1819 -11245 -1781 -11211
rect -1747 -11245 -1709 -11211
rect -1675 -11245 -1637 -11211
rect -1603 -11245 -1565 -11211
rect -1531 -11245 -1493 -11211
rect -1459 -11245 -1421 -11211
rect -1387 -11245 -1349 -11211
rect -1315 -11245 -1277 -11211
rect -1243 -11245 -1205 -11211
rect -1171 -11245 -1133 -11211
rect -1099 -11245 -1061 -11211
rect -1027 -11245 -989 -11211
rect -955 -11245 -917 -11211
rect -883 -11245 -845 -11211
rect -811 -11245 -773 -11211
rect -739 -11245 -701 -11211
rect -667 -11245 -629 -11211
rect -595 -11245 -557 -11211
rect -523 -11245 -485 -11211
rect -451 -11245 -413 -11211
rect -379 -11245 -341 -11211
rect -307 -11245 -269 -11211
rect -235 -11245 -197 -11211
rect -163 -11245 -125 -11211
rect -91 -11245 -53 -11211
rect -19 -11245 19 -11211
rect 53 -11245 91 -11211
rect 125 -11245 163 -11211
rect 197 -11245 235 -11211
rect 269 -11245 307 -11211
rect 341 -11245 379 -11211
rect 413 -11245 451 -11211
rect 485 -11245 523 -11211
rect 557 -11245 595 -11211
rect 629 -11245 667 -11211
rect 701 -11245 739 -11211
rect 773 -11245 811 -11211
rect 845 -11245 883 -11211
rect 917 -11245 955 -11211
rect 989 -11245 1027 -11211
rect 1061 -11245 1099 -11211
rect 1133 -11245 1171 -11211
rect 1205 -11245 1243 -11211
rect 1277 -11245 1315 -11211
rect 1349 -11245 1387 -11211
rect 1421 -11245 1459 -11211
rect 1493 -11245 1531 -11211
rect 1565 -11245 1603 -11211
rect 1637 -11245 1675 -11211
rect 1709 -11245 1747 -11211
rect 1781 -11245 1819 -11211
rect 1853 -11245 1891 -11211
rect 1925 -11245 1963 -11211
rect 1997 -11245 2035 -11211
rect 2069 -11245 2107 -11211
rect 2141 -11245 2179 -11211
rect 2213 -11245 2251 -11211
rect 2285 -11245 2323 -11211
rect 2357 -11245 2395 -11211
rect 2429 -11245 2467 -11211
rect 2501 -11245 2539 -11211
rect 2573 -11245 2611 -11211
rect 2645 -11245 2683 -11211
rect 2717 -11245 2755 -11211
rect 2789 -11245 2827 -11211
rect 2861 -11245 2899 -11211
rect 2933 -11245 2971 -11211
rect 3005 -11245 3043 -11211
rect 3077 -11245 3115 -11211
rect 3149 -11245 3187 -11211
rect 3221 -11245 3259 -11211
rect 3293 -11245 3331 -11211
rect 3365 -11245 3403 -11211
rect 3437 -11245 3475 -11211
rect 3509 -11245 3547 -11211
rect 3581 -11245 3619 -11211
rect 3653 -11245 3691 -11211
rect 3725 -11245 3763 -11211
rect 3797 -11245 3835 -11211
rect 3869 -11245 3907 -11211
rect 3941 -11245 3979 -11211
rect 4013 -11245 4051 -11211
rect 4085 -11245 4123 -11211
rect 4157 -11245 4195 -11211
rect 4229 -11245 4267 -11211
rect 4301 -11245 4339 -11211
rect 4373 -11245 4411 -11211
rect 4445 -11245 4483 -11211
rect 4517 -11245 4555 -11211
rect 4589 -11245 4627 -11211
rect 4661 -11245 4699 -11211
rect 4733 -11245 4771 -11211
rect 4805 -11245 4843 -11211
rect 4877 -11245 4915 -11211
rect 4949 -11245 4987 -11211
rect 5021 -11245 5059 -11211
rect 5093 -11245 5131 -11211
rect 5165 -11245 5203 -11211
rect 5237 -11245 5275 -11211
rect 5309 -11245 5347 -11211
rect 5381 -11245 5419 -11211
rect 5453 -11245 5491 -11211
rect 5525 -11245 5563 -11211
rect 5597 -11245 5635 -11211
rect 5669 -11245 5707 -11211
rect 5741 -11245 5779 -11211
rect 5813 -11245 5851 -11211
rect 5885 -11245 5923 -11211
rect 5957 -11245 5995 -11211
rect 6029 -11245 6067 -11211
rect 6101 -11245 6139 -11211
rect 6173 -11245 6211 -11211
rect 6245 -11245 6283 -11211
rect 6317 -11245 6355 -11211
rect 6389 -11245 6427 -11211
rect 6461 -11245 6499 -11211
rect 6533 -11245 6571 -11211
rect 6605 -11245 6643 -11211
rect 6677 -11245 6715 -11211
rect 6749 -11245 6787 -11211
rect 6821 -11245 6859 -11211
rect 6893 -11245 6931 -11211
rect 6965 -11245 7003 -11211
rect 7037 -11245 7075 -11211
rect 7109 -11245 7147 -11211
rect 7181 -11245 7219 -11211
rect 7253 -11245 7291 -11211
rect 7325 -11245 7363 -11211
rect 7397 -11245 7435 -11211
rect 7469 -11245 7507 -11211
rect 7541 -11245 7579 -11211
rect 7613 -11245 7651 -11211
rect 7685 -11245 7723 -11211
rect 7757 -11245 7795 -11211
rect 7829 -11245 7867 -11211
rect 7901 -11245 7939 -11211
rect 7973 -11245 8011 -11211
rect 8045 -11245 8083 -11211
rect 8117 -11245 8155 -11211
rect 8189 -11245 8227 -11211
rect 8261 -11245 8299 -11211
rect 8333 -11245 8371 -11211
rect 8405 -11245 8443 -11211
rect 8477 -11245 8515 -11211
rect 8549 -11245 8587 -11211
rect 8621 -11245 8659 -11211
rect 8693 -11245 8731 -11211
rect 8765 -11245 8803 -11211
rect 8837 -11245 8875 -11211
rect 8909 -11245 8947 -11211
rect 8981 -11245 9019 -11211
rect 9053 -11245 9091 -11211
rect 9125 -11245 9163 -11211
rect 9197 -11245 9235 -11211
rect 9269 -11245 9307 -11211
rect 9341 -11245 9379 -11211
rect 9413 -11245 9451 -11211
rect 9485 -11245 9523 -11211
rect 9557 -11245 9595 -11211
rect 9629 -11245 9667 -11211
rect 9701 -11245 9739 -11211
rect 9773 -11245 9811 -11211
rect 9845 -11245 9883 -11211
rect 9917 -11245 9955 -11211
rect 9989 -11245 10027 -11211
rect 10061 -11245 10099 -11211
rect 10133 -11245 10171 -11211
rect 10205 -11245 10243 -11211
rect 10277 -11245 10315 -11211
rect 10349 -11245 10387 -11211
rect 10421 -11245 10459 -11211
rect 10493 -11245 10531 -11211
rect 10565 -11245 10603 -11211
rect 10637 -11245 10675 -11211
rect 10709 -11245 10747 -11211
rect 10781 -11245 10819 -11211
rect 10853 -11245 10891 -11211
rect 10925 -11245 10963 -11211
rect 10997 -11245 11035 -11211
rect 11069 -11245 11107 -11211
rect 11141 -11245 11179 -11211
rect 11213 -11245 11251 -11211
rect 11285 -11245 11323 -11211
rect 11357 -11245 11395 -11211
rect 11429 -11245 11467 -11211
rect 11501 -11245 11539 -11211
rect 11573 -11245 11611 -11211
rect 11645 -11245 11683 -11211
rect 11717 -11245 11755 -11211
rect 11789 -11245 11827 -11211
rect 11861 -11245 11899 -11211
rect 11933 -11245 11971 -11211
rect 12005 -11245 12043 -11211
rect 12077 -11245 12115 -11211
rect 12149 -11245 12187 -11211
rect 12221 -11245 12259 -11211
rect 12293 -11245 12331 -11211
rect 12365 -11245 12403 -11211
rect 12437 -11245 12475 -11211
rect 12509 -11245 12547 -11211
rect 12581 -11245 12619 -11211
rect 12653 -11245 12691 -11211
rect 12725 -11245 12763 -11211
rect 12797 -11245 12835 -11211
rect 12869 -11245 12907 -11211
rect 12941 -11245 12979 -11211
rect 13013 -11245 13051 -11211
rect 13085 -11245 13123 -11211
rect 13157 -11245 13195 -11211
rect 13229 -11245 13267 -11211
rect 13301 -11245 13339 -11211
rect 13373 -11245 13411 -11211
rect 13445 -11245 13483 -11211
rect 13517 -11245 13555 -11211
rect 13589 -11245 13627 -11211
rect 13661 -11245 13699 -11211
rect 13733 -11245 13771 -11211
rect 13805 -11245 13843 -11211
rect 13877 -11245 13915 -11211
rect 13949 -11245 13987 -11211
rect 14021 -11245 14059 -11211
rect 14093 -11245 14131 -11211
rect 14165 -11245 14203 -11211
rect 14237 -11245 14275 -11211
rect 14309 -11245 14347 -11211
rect 14381 -11245 14419 -11211
rect 14453 -11245 14491 -11211
rect 14525 -11245 14563 -11211
rect 14597 -11245 14635 -11211
rect 14669 -11245 14707 -11211
rect 14741 -11245 14779 -11211
rect 14813 -11245 14851 -11211
rect 14885 -11245 14923 -11211
rect 14957 -11245 14995 -11211
rect 15029 -11245 15067 -11211
rect 15101 -11245 15139 -11211
rect 15173 -11245 15211 -11211
rect 15245 -11245 15283 -11211
rect 15317 -11245 15355 -11211
rect 15389 -11245 15427 -11211
rect 15461 -11245 15499 -11211
rect 15533 -11245 15571 -11211
rect 15605 -11245 15643 -11211
rect 15677 -11245 15715 -11211
rect 15749 -11245 15787 -11211
rect 15821 -11245 15859 -11211
rect 15893 -11245 15931 -11211
rect 15965 -11245 16003 -11211
rect 16037 -11245 16075 -11211
rect 16109 -11245 16147 -11211
rect 16181 -11245 16219 -11211
rect 16253 -11245 16291 -11211
rect 16325 -11245 16363 -11211
rect 16397 -11245 16435 -11211
rect 16469 -11245 16507 -11211
rect 16541 -11245 16579 -11211
rect 16613 -11245 16651 -11211
rect 16685 -11245 16723 -11211
rect 16757 -11245 16795 -11211
rect 16829 -11245 16867 -11211
rect 16901 -11245 16939 -11211
rect 16973 -11245 17011 -11211
rect 17045 -11245 17083 -11211
rect 17117 -11245 17155 -11211
rect 17189 -11245 17227 -11211
rect 17261 -11245 17299 -11211
rect 17333 -11245 17371 -11211
rect 17405 -11245 17443 -11211
rect 17477 -11245 17515 -11211
rect 17549 -11245 17587 -11211
rect 17621 -11245 17659 -11211
rect 17693 -11245 17731 -11211
rect 17765 -11245 17803 -11211
rect 17837 -11245 17875 -11211
rect 17909 -11245 17947 -11211
rect 17981 -11245 18019 -11211
rect 18053 -11245 18091 -11211
rect 18125 -11245 18163 -11211
rect 18197 -11245 18235 -11211
rect 18269 -11245 18307 -11211
rect 18341 -11245 18379 -11211
rect 18413 -11245 18451 -11211
rect 18485 -11245 18523 -11211
rect 18557 -11245 18595 -11211
rect 18629 -11245 18667 -11211
rect 18701 -11245 18739 -11211
rect 18773 -11245 18811 -11211
rect 18845 -11245 18883 -11211
rect 18917 -11245 18955 -11211
rect 18989 -11245 19027 -11211
rect 19061 -11245 19099 -11211
rect 19133 -11245 19171 -11211
rect 19205 -11245 19243 -11211
rect 19277 -11245 19315 -11211
rect 19349 -11245 19387 -11211
rect 19421 -11245 19459 -11211
rect 19493 -11245 19531 -11211
rect 19565 -11245 19603 -11211
rect 19637 -11245 19675 -11211
rect 19709 -11245 19747 -11211
rect 19781 -11245 19819 -11211
rect 19853 -11245 19891 -11211
rect 19925 -11245 19963 -11211
rect 19997 -11245 20035 -11211
rect 20069 -11245 20107 -11211
rect 20141 -11245 20179 -11211
rect 20213 -11245 20251 -11211
rect 20285 -11245 20323 -11211
rect 20357 -11245 20395 -11211
rect 20429 -11245 20467 -11211
rect 20501 -11245 20539 -11211
rect 20573 -11245 20611 -11211
rect 20645 -11245 20683 -11211
rect 20717 -11245 20755 -11211
rect 20789 -11245 20827 -11211
rect 20861 -11245 20899 -11211
rect 20933 -11245 20971 -11211
rect 21005 -11245 21043 -11211
rect 21077 -11245 21115 -11211
rect 21149 -11245 21187 -11211
rect 21221 -11245 21259 -11211
rect 21293 -11245 21331 -11211
rect 21365 -11245 21403 -11211
rect 21437 -11245 21475 -11211
rect 21509 -11245 21547 -11211
rect 21581 -11245 21619 -11211
rect 21653 -11245 21691 -11211
rect 21725 -11245 21763 -11211
rect 21797 -11245 21835 -11211
rect 21869 -11245 21907 -11211
rect 21941 -11245 21979 -11211
rect 22013 -11245 22051 -11211
rect 22085 -11245 22123 -11211
rect 22157 -11245 22195 -11211
rect 22229 -11245 22267 -11211
rect 22301 -11245 22339 -11211
rect 22373 -11245 22411 -11211
rect 22445 -11245 22483 -11211
rect 22517 -11245 22555 -11211
rect 22589 -11245 22627 -11211
rect 22661 -11245 22699 -11211
rect 22733 -11245 22771 -11211
rect 22805 -11245 22843 -11211
rect 22877 -11245 22915 -11211
rect 22949 -11245 22987 -11211
rect 23021 -11245 23059 -11211
rect 23093 -11245 23131 -11211
rect 23165 -11245 23203 -11211
rect 23237 -11245 23275 -11211
rect 23309 -11245 23347 -11211
rect 23381 -11245 23419 -11211
rect 23453 -11245 23491 -11211
rect 23525 -11245 23563 -11211
rect 23597 -11245 23635 -11211
rect 23669 -11245 23707 -11211
rect 23741 -11245 23779 -11211
rect 23813 -11245 23851 -11211
rect 23885 -11245 23923 -11211
rect 23957 -11245 23995 -11211
rect 24029 -11245 24067 -11211
rect 24101 -11245 24139 -11211
rect 24173 -11245 24211 -11211
rect 24245 -11245 24283 -11211
rect 24317 -11245 24355 -11211
rect 24389 -11245 24427 -11211
rect 24461 -11245 24499 -11211
rect 24533 -11245 24571 -11211
rect 24605 -11245 24643 -11211
rect 24677 -11245 24715 -11211
rect 24749 -11245 24787 -11211
rect 24821 -11245 24928 -11211
rect -13992 -11284 24928 -11245
rect -13992 -11300 -1642 -11284
rect -12328 -12091 -12216 -11300
rect 2210 -11352 2282 -11348
rect 1888 -11362 1948 -11352
rect 1888 -11414 1892 -11362
rect 1944 -11414 1948 -11362
rect 2210 -11404 2220 -11352
rect 2272 -11404 2282 -11352
rect 2210 -11408 2282 -11404
rect 2336 -11360 2396 -11350
rect 1764 -11462 1836 -11458
rect 1536 -11478 1608 -11474
rect 1276 -11498 1348 -11494
rect 1276 -11550 1286 -11498
rect 1338 -11550 1348 -11498
rect 1276 -11554 1348 -11550
rect 1396 -11496 1468 -11492
rect 1396 -11548 1406 -11496
rect 1458 -11548 1468 -11496
rect 1536 -11530 1546 -11478
rect 1598 -11530 1608 -11478
rect 1764 -11514 1774 -11462
rect 1826 -11514 1836 -11462
rect 1764 -11518 1836 -11514
rect 1536 -11534 1608 -11530
rect 1396 -11552 1468 -11548
rect 1144 -11626 1216 -11622
rect 1144 -11678 1154 -11626
rect 1206 -11678 1216 -11626
rect 1144 -11682 1216 -11678
rect -12328 -12125 -12289 -12091
rect -12255 -12125 -12216 -12091
rect -12328 -12163 -12216 -12125
rect -12328 -12197 -12289 -12163
rect -12255 -12197 -12216 -12163
rect -12328 -12235 -12216 -12197
rect -12328 -12269 -12289 -12235
rect -12255 -12269 -12216 -12235
rect -12328 -12307 -12216 -12269
rect -1568 -12224 -1496 -12220
rect -1568 -12276 -1558 -12224
rect -1506 -12276 -1496 -12224
rect -1568 -12280 -1496 -12276
rect -12328 -12341 -12289 -12307
rect -12255 -12341 -12216 -12307
rect -1562 -12324 -1502 -12280
rect -12328 -12379 -12216 -12341
rect -12328 -12413 -12289 -12379
rect -12255 -12413 -12216 -12379
rect -12328 -12451 -12216 -12413
rect -12328 -12485 -12289 -12451
rect -12255 -12485 -12216 -12451
rect -12328 -12523 -12216 -12485
rect -12328 -12557 -12289 -12523
rect -12255 -12557 -12216 -12523
rect -9196 -12384 -1502 -12324
rect -9196 -12543 -9136 -12384
rect -8686 -12434 -8626 -12384
rect -8902 -12440 -8414 -12434
rect -8902 -12474 -8855 -12440
rect -8821 -12474 -8783 -12440
rect -8749 -12474 -8711 -12440
rect -8677 -12474 -8639 -12440
rect -8605 -12474 -8567 -12440
rect -8533 -12474 -8495 -12440
rect -8461 -12474 -8414 -12440
rect -8902 -12480 -8414 -12474
rect -9196 -12554 -9184 -12543
rect -12328 -12595 -12216 -12557
rect -12328 -12629 -12289 -12595
rect -12255 -12629 -12216 -12595
rect -12328 -12667 -12216 -12629
rect -12328 -12701 -12289 -12667
rect -12255 -12701 -12216 -12667
rect -12328 -12739 -12216 -12701
rect -12328 -12773 -12289 -12739
rect -12255 -12773 -12216 -12739
rect -12328 -12811 -12216 -12773
rect -12328 -12845 -12289 -12811
rect -12255 -12845 -12216 -12811
rect -12328 -12883 -12216 -12845
rect -12328 -12917 -12289 -12883
rect -12255 -12917 -12216 -12883
rect -12328 -12955 -12216 -12917
rect -12328 -12989 -12289 -12955
rect -12255 -12989 -12216 -12955
rect -12328 -13027 -12216 -12989
rect -12328 -13061 -12289 -13027
rect -12255 -13061 -12216 -13027
rect -12328 -13099 -12216 -13061
rect -9190 -12577 -9184 -12554
rect -9150 -12554 -9136 -12543
rect -8180 -12543 -8120 -12384
rect -7678 -12434 -7618 -12384
rect -6650 -12434 -6590 -12384
rect -7884 -12440 -7396 -12434
rect -7884 -12474 -7837 -12440
rect -7803 -12474 -7765 -12440
rect -7731 -12474 -7693 -12440
rect -7659 -12474 -7621 -12440
rect -7587 -12474 -7549 -12440
rect -7515 -12474 -7477 -12440
rect -7443 -12474 -7396 -12440
rect -7884 -12480 -7396 -12474
rect -6866 -12440 -6378 -12434
rect -6866 -12474 -6819 -12440
rect -6785 -12474 -6747 -12440
rect -6713 -12474 -6675 -12440
rect -6641 -12474 -6603 -12440
rect -6569 -12474 -6531 -12440
rect -6497 -12474 -6459 -12440
rect -6425 -12474 -6378 -12440
rect -6866 -12480 -6378 -12474
rect -8180 -12548 -8166 -12543
rect -9150 -12577 -9144 -12554
rect -9190 -12615 -9144 -12577
rect -9190 -12649 -9184 -12615
rect -9150 -12649 -9144 -12615
rect -9190 -12687 -9144 -12649
rect -9190 -12721 -9184 -12687
rect -9150 -12721 -9144 -12687
rect -9190 -12759 -9144 -12721
rect -9190 -12793 -9184 -12759
rect -9150 -12793 -9144 -12759
rect -9190 -12831 -9144 -12793
rect -9190 -12865 -9184 -12831
rect -9150 -12865 -9144 -12831
rect -9190 -12903 -9144 -12865
rect -9190 -12937 -9184 -12903
rect -9150 -12937 -9144 -12903
rect -9190 -12975 -9144 -12937
rect -9190 -13009 -9184 -12975
rect -9150 -13009 -9144 -12975
rect -9190 -13047 -9144 -13009
rect -9190 -13081 -9184 -13047
rect -9150 -13081 -9144 -13047
rect -8172 -12577 -8166 -12548
rect -8132 -12548 -8120 -12543
rect -7154 -12543 -7108 -12512
rect -8132 -12577 -8126 -12548
rect -8172 -12615 -8126 -12577
rect -8172 -12649 -8166 -12615
rect -8132 -12649 -8126 -12615
rect -8172 -12687 -8126 -12649
rect -8172 -12721 -8166 -12687
rect -8132 -12721 -8126 -12687
rect -8172 -12759 -8126 -12721
rect -8172 -12793 -8166 -12759
rect -8132 -12793 -8126 -12759
rect -8172 -12831 -8126 -12793
rect -8172 -12865 -8166 -12831
rect -8132 -12865 -8126 -12831
rect -8172 -12903 -8126 -12865
rect -8172 -12937 -8166 -12903
rect -8132 -12937 -8126 -12903
rect -8172 -12975 -8126 -12937
rect -8172 -13009 -8166 -12975
rect -8132 -13009 -8126 -12975
rect -8172 -13047 -8126 -13009
rect -8172 -13078 -8166 -13047
rect -9190 -13082 -9144 -13081
rect -8180 -13081 -8166 -13078
rect -8132 -13078 -8126 -13047
rect -7154 -12577 -7148 -12543
rect -7114 -12577 -7108 -12543
rect -6142 -12543 -6082 -12384
rect -5636 -12434 -5576 -12384
rect -4622 -12434 -4562 -12384
rect -5848 -12440 -5360 -12434
rect -5848 -12474 -5801 -12440
rect -5767 -12474 -5729 -12440
rect -5695 -12474 -5657 -12440
rect -5623 -12474 -5585 -12440
rect -5551 -12474 -5513 -12440
rect -5479 -12474 -5441 -12440
rect -5407 -12474 -5360 -12440
rect -5848 -12480 -5360 -12474
rect -4830 -12440 -4342 -12434
rect -4830 -12474 -4783 -12440
rect -4749 -12474 -4711 -12440
rect -4677 -12474 -4639 -12440
rect -4605 -12474 -4567 -12440
rect -4533 -12474 -4495 -12440
rect -4461 -12474 -4423 -12440
rect -4389 -12474 -4342 -12440
rect -4830 -12480 -4342 -12474
rect -6142 -12562 -6130 -12543
rect -7154 -12615 -7108 -12577
rect -7154 -12649 -7148 -12615
rect -7114 -12649 -7108 -12615
rect -7154 -12687 -7108 -12649
rect -7154 -12721 -7148 -12687
rect -7114 -12721 -7108 -12687
rect -7154 -12759 -7108 -12721
rect -7154 -12793 -7148 -12759
rect -7114 -12793 -7108 -12759
rect -7154 -12831 -7108 -12793
rect -7154 -12865 -7148 -12831
rect -7114 -12865 -7108 -12831
rect -7154 -12903 -7108 -12865
rect -7154 -12937 -7148 -12903
rect -7114 -12937 -7108 -12903
rect -7154 -12975 -7108 -12937
rect -7154 -13009 -7148 -12975
rect -7114 -13009 -7108 -12975
rect -7154 -13047 -7108 -13009
rect -7154 -13076 -7148 -13047
rect -8132 -13081 -8120 -13078
rect -12328 -13133 -12289 -13099
rect -12255 -13133 -12216 -13099
rect -12328 -13171 -12216 -13133
rect -12328 -13205 -12289 -13171
rect -12255 -13205 -12216 -13171
rect -12328 -13243 -12216 -13205
rect -12328 -13277 -12289 -13243
rect -12255 -13277 -12216 -13243
rect -12328 -13315 -12216 -13277
rect -12328 -13349 -12289 -13315
rect -12255 -13349 -12216 -13315
rect -12328 -13387 -12216 -13349
rect -9200 -13361 -9140 -13082
rect -8902 -13150 -8414 -13144
rect -8902 -13184 -8855 -13150
rect -8821 -13184 -8783 -13150
rect -8749 -13184 -8711 -13150
rect -8677 -13184 -8639 -13150
rect -8605 -13184 -8567 -13150
rect -8533 -13184 -8495 -13150
rect -8461 -13184 -8414 -13150
rect -8902 -13190 -8414 -13184
rect -8686 -13252 -8626 -13190
rect -8902 -13258 -8414 -13252
rect -8902 -13292 -8855 -13258
rect -8821 -13292 -8783 -13258
rect -8749 -13292 -8711 -13258
rect -8677 -13292 -8639 -13258
rect -8605 -13292 -8567 -13258
rect -8533 -13292 -8495 -13258
rect -8461 -13292 -8414 -13258
rect -8902 -13298 -8414 -13292
rect -9200 -13372 -9184 -13361
rect -12328 -13421 -12289 -13387
rect -12255 -13421 -12216 -13387
rect -12328 -13459 -12216 -13421
rect -12328 -13493 -12289 -13459
rect -12255 -13493 -12216 -13459
rect -12328 -13531 -12216 -13493
rect -12328 -13565 -12289 -13531
rect -12255 -13565 -12216 -13531
rect -12328 -13603 -12216 -13565
rect -12328 -13637 -12289 -13603
rect -12255 -13637 -12216 -13603
rect -12328 -13675 -12216 -13637
rect -12328 -13709 -12289 -13675
rect -12255 -13709 -12216 -13675
rect -12328 -13747 -12216 -13709
rect -12328 -13781 -12289 -13747
rect -12255 -13781 -12216 -13747
rect -12328 -13819 -12216 -13781
rect -12328 -13853 -12289 -13819
rect -12255 -13853 -12216 -13819
rect -12328 -13891 -12216 -13853
rect -12328 -13925 -12289 -13891
rect -12255 -13925 -12216 -13891
rect -9190 -13395 -9184 -13372
rect -9150 -13372 -9140 -13361
rect -8180 -13361 -8120 -13081
rect -7160 -13081 -7148 -13076
rect -7114 -13076 -7108 -13047
rect -6136 -12577 -6130 -12562
rect -6096 -12562 -6082 -12543
rect -5118 -12543 -5072 -12512
rect -4106 -12524 -4046 -12384
rect -3590 -12434 -3530 -12384
rect -2584 -12434 -2524 -12384
rect -3812 -12440 -3324 -12434
rect -3812 -12474 -3765 -12440
rect -3731 -12474 -3693 -12440
rect -3659 -12474 -3621 -12440
rect -3587 -12474 -3549 -12440
rect -3515 -12474 -3477 -12440
rect -3443 -12474 -3405 -12440
rect -3371 -12474 -3324 -12440
rect -3812 -12480 -3324 -12474
rect -2794 -12440 -2306 -12434
rect -2794 -12474 -2747 -12440
rect -2713 -12474 -2675 -12440
rect -2641 -12474 -2603 -12440
rect -2569 -12474 -2531 -12440
rect -2497 -12474 -2459 -12440
rect -2425 -12474 -2387 -12440
rect -2353 -12474 -2306 -12440
rect -2794 -12480 -2306 -12474
rect -6096 -12577 -6090 -12562
rect -6136 -12615 -6090 -12577
rect -6136 -12649 -6130 -12615
rect -6096 -12649 -6090 -12615
rect -6136 -12687 -6090 -12649
rect -6136 -12721 -6130 -12687
rect -6096 -12721 -6090 -12687
rect -6136 -12759 -6090 -12721
rect -6136 -12793 -6130 -12759
rect -6096 -12793 -6090 -12759
rect -6136 -12831 -6090 -12793
rect -6136 -12865 -6130 -12831
rect -6096 -12865 -6090 -12831
rect -6136 -12903 -6090 -12865
rect -6136 -12937 -6130 -12903
rect -6096 -12937 -6090 -12903
rect -6136 -12975 -6090 -12937
rect -6136 -13009 -6130 -12975
rect -6096 -13009 -6090 -12975
rect -6136 -13047 -6090 -13009
rect -7114 -13081 -7100 -13076
rect -6136 -13080 -6130 -13047
rect -7884 -13150 -7396 -13144
rect -7884 -13184 -7837 -13150
rect -7803 -13184 -7765 -13150
rect -7731 -13184 -7693 -13150
rect -7659 -13184 -7621 -13150
rect -7587 -13184 -7549 -13150
rect -7515 -13184 -7477 -13150
rect -7443 -13184 -7396 -13150
rect -7884 -13190 -7396 -13184
rect -7682 -13252 -7622 -13190
rect -7884 -13258 -7396 -13252
rect -7884 -13292 -7837 -13258
rect -7803 -13292 -7765 -13258
rect -7731 -13292 -7693 -13258
rect -7659 -13292 -7621 -13258
rect -7587 -13292 -7549 -13258
rect -7515 -13292 -7477 -13258
rect -7443 -13292 -7396 -13258
rect -7884 -13298 -7396 -13292
rect -8180 -13368 -8166 -13361
rect -9150 -13395 -9144 -13372
rect -9190 -13433 -9144 -13395
rect -9190 -13467 -9184 -13433
rect -9150 -13467 -9144 -13433
rect -9190 -13505 -9144 -13467
rect -9190 -13539 -9184 -13505
rect -9150 -13539 -9144 -13505
rect -9190 -13577 -9144 -13539
rect -9190 -13611 -9184 -13577
rect -9150 -13611 -9144 -13577
rect -9190 -13649 -9144 -13611
rect -9190 -13683 -9184 -13649
rect -9150 -13683 -9144 -13649
rect -9190 -13721 -9144 -13683
rect -9190 -13755 -9184 -13721
rect -9150 -13755 -9144 -13721
rect -9190 -13793 -9144 -13755
rect -9190 -13827 -9184 -13793
rect -9150 -13827 -9144 -13793
rect -9190 -13865 -9144 -13827
rect -9190 -13896 -9184 -13865
rect -12328 -13963 -12216 -13925
rect -12328 -13997 -12289 -13963
rect -12255 -13997 -12216 -13963
rect -12328 -14035 -12216 -13997
rect -12328 -14069 -12289 -14035
rect -12255 -14069 -12216 -14035
rect -12328 -14107 -12216 -14069
rect -12328 -14141 -12289 -14107
rect -12255 -14141 -12216 -14107
rect -12328 -14179 -12216 -14141
rect -12328 -14213 -12289 -14179
rect -12255 -14213 -12216 -14179
rect -9198 -13899 -9184 -13896
rect -9150 -13896 -9144 -13865
rect -8172 -13395 -8166 -13368
rect -8132 -13368 -8120 -13361
rect -7160 -13361 -7100 -13081
rect -6142 -13081 -6130 -13080
rect -6096 -13080 -6090 -13047
rect -5118 -12577 -5112 -12543
rect -5078 -12577 -5072 -12543
rect -4108 -12543 -4046 -12524
rect -4108 -12558 -4094 -12543
rect -4106 -12570 -4094 -12558
rect -5118 -12615 -5072 -12577
rect -5118 -12649 -5112 -12615
rect -5078 -12649 -5072 -12615
rect -5118 -12687 -5072 -12649
rect -5118 -12721 -5112 -12687
rect -5078 -12721 -5072 -12687
rect -5118 -12759 -5072 -12721
rect -5118 -12793 -5112 -12759
rect -5078 -12793 -5072 -12759
rect -5118 -12831 -5072 -12793
rect -5118 -12865 -5112 -12831
rect -5078 -12865 -5072 -12831
rect -5118 -12903 -5072 -12865
rect -5118 -12937 -5112 -12903
rect -5078 -12937 -5072 -12903
rect -5118 -12975 -5072 -12937
rect -5118 -13009 -5112 -12975
rect -5078 -13009 -5072 -12975
rect -5118 -13047 -5072 -13009
rect -5118 -13072 -5112 -13047
rect -6096 -13081 -6082 -13080
rect -6866 -13150 -6378 -13144
rect -6866 -13184 -6819 -13150
rect -6785 -13184 -6747 -13150
rect -6713 -13184 -6675 -13150
rect -6641 -13184 -6603 -13150
rect -6569 -13184 -6531 -13150
rect -6497 -13184 -6459 -13150
rect -6425 -13184 -6378 -13150
rect -6866 -13190 -6378 -13184
rect -6652 -13252 -6592 -13190
rect -6866 -13258 -6378 -13252
rect -6866 -13292 -6819 -13258
rect -6785 -13292 -6747 -13258
rect -6713 -13292 -6675 -13258
rect -6641 -13292 -6603 -13258
rect -6569 -13292 -6531 -13258
rect -6497 -13292 -6459 -13258
rect -6425 -13292 -6378 -13258
rect -6866 -13298 -6378 -13292
rect -7160 -13366 -7148 -13361
rect -8132 -13395 -8126 -13368
rect -8172 -13433 -8126 -13395
rect -8172 -13467 -8166 -13433
rect -8132 -13467 -8126 -13433
rect -8172 -13505 -8126 -13467
rect -8172 -13539 -8166 -13505
rect -8132 -13539 -8126 -13505
rect -8172 -13577 -8126 -13539
rect -8172 -13611 -8166 -13577
rect -8132 -13611 -8126 -13577
rect -8172 -13649 -8126 -13611
rect -8172 -13683 -8166 -13649
rect -8132 -13683 -8126 -13649
rect -8172 -13721 -8126 -13683
rect -8172 -13755 -8166 -13721
rect -8132 -13755 -8126 -13721
rect -8172 -13793 -8126 -13755
rect -8172 -13827 -8166 -13793
rect -8132 -13827 -8126 -13793
rect -8172 -13865 -8126 -13827
rect -8172 -13892 -8166 -13865
rect -9150 -13899 -9138 -13896
rect -9198 -14179 -9138 -13899
rect -8178 -13899 -8166 -13892
rect -8132 -13892 -8126 -13865
rect -7154 -13395 -7148 -13366
rect -7114 -13366 -7100 -13361
rect -6142 -13361 -6082 -13081
rect -5122 -13081 -5112 -13072
rect -5078 -13072 -5072 -13047
rect -4100 -12577 -4094 -12570
rect -4060 -12570 -4046 -12543
rect -3082 -12543 -3036 -12512
rect -4060 -12577 -4054 -12570
rect -4100 -12615 -4054 -12577
rect -4100 -12649 -4094 -12615
rect -4060 -12649 -4054 -12615
rect -4100 -12687 -4054 -12649
rect -4100 -12721 -4094 -12687
rect -4060 -12721 -4054 -12687
rect -4100 -12759 -4054 -12721
rect -4100 -12793 -4094 -12759
rect -4060 -12793 -4054 -12759
rect -4100 -12831 -4054 -12793
rect -4100 -12865 -4094 -12831
rect -4060 -12865 -4054 -12831
rect -4100 -12903 -4054 -12865
rect -4100 -12937 -4094 -12903
rect -4060 -12937 -4054 -12903
rect -4100 -12975 -4054 -12937
rect -4100 -13009 -4094 -12975
rect -4060 -13009 -4054 -12975
rect -4100 -13047 -4054 -13009
rect -5078 -13081 -5062 -13072
rect -4100 -13080 -4094 -13047
rect -5848 -13150 -5360 -13144
rect -5848 -13184 -5801 -13150
rect -5767 -13184 -5729 -13150
rect -5695 -13184 -5657 -13150
rect -5623 -13184 -5585 -13150
rect -5551 -13184 -5513 -13150
rect -5479 -13184 -5441 -13150
rect -5407 -13184 -5360 -13150
rect -5848 -13190 -5360 -13184
rect -5650 -13252 -5590 -13190
rect -5848 -13258 -5360 -13252
rect -5848 -13292 -5801 -13258
rect -5767 -13292 -5729 -13258
rect -5695 -13292 -5657 -13258
rect -5623 -13292 -5585 -13258
rect -5551 -13292 -5513 -13258
rect -5479 -13292 -5441 -13258
rect -5407 -13292 -5360 -13258
rect -5848 -13298 -5360 -13292
rect -7114 -13395 -7108 -13366
rect -6142 -13370 -6130 -13361
rect -7154 -13433 -7108 -13395
rect -7154 -13467 -7148 -13433
rect -7114 -13467 -7108 -13433
rect -7154 -13505 -7108 -13467
rect -7154 -13539 -7148 -13505
rect -7114 -13539 -7108 -13505
rect -7154 -13577 -7108 -13539
rect -7154 -13611 -7148 -13577
rect -7114 -13611 -7108 -13577
rect -7154 -13649 -7108 -13611
rect -7154 -13683 -7148 -13649
rect -7114 -13683 -7108 -13649
rect -7154 -13721 -7108 -13683
rect -7154 -13755 -7148 -13721
rect -7114 -13755 -7108 -13721
rect -7154 -13793 -7108 -13755
rect -7154 -13827 -7148 -13793
rect -7114 -13827 -7108 -13793
rect -7154 -13865 -7108 -13827
rect -7154 -13890 -7148 -13865
rect -8132 -13899 -8118 -13892
rect -8902 -13968 -8414 -13962
rect -8902 -14002 -8855 -13968
rect -8821 -14002 -8783 -13968
rect -8749 -14002 -8711 -13968
rect -8677 -14002 -8639 -13968
rect -8605 -14002 -8567 -13968
rect -8533 -14002 -8495 -13968
rect -8461 -14002 -8414 -13968
rect -8902 -14008 -8414 -14002
rect -8686 -14070 -8626 -14008
rect -8902 -14076 -8414 -14070
rect -8902 -14110 -8855 -14076
rect -8821 -14110 -8783 -14076
rect -8749 -14110 -8711 -14076
rect -8677 -14110 -8639 -14076
rect -8605 -14110 -8567 -14076
rect -8533 -14110 -8495 -14076
rect -8461 -14110 -8414 -14076
rect -8902 -14116 -8414 -14110
rect -9198 -14186 -9184 -14179
rect -12328 -14251 -12216 -14213
rect -12328 -14285 -12289 -14251
rect -12255 -14285 -12216 -14251
rect -12328 -14323 -12216 -14285
rect -12328 -14357 -12289 -14323
rect -12255 -14357 -12216 -14323
rect -12328 -14395 -12216 -14357
rect -12328 -14429 -12289 -14395
rect -12255 -14429 -12216 -14395
rect -12328 -14467 -12216 -14429
rect -12328 -14501 -12289 -14467
rect -12255 -14501 -12216 -14467
rect -12328 -14539 -12216 -14501
rect -12328 -14573 -12289 -14539
rect -12255 -14573 -12216 -14539
rect -12328 -14611 -12216 -14573
rect -12328 -14645 -12289 -14611
rect -12255 -14645 -12216 -14611
rect -12328 -14683 -12216 -14645
rect -12328 -14717 -12289 -14683
rect -12255 -14717 -12216 -14683
rect -12328 -14755 -12216 -14717
rect -9190 -14213 -9184 -14186
rect -9150 -14186 -9138 -14179
rect -8178 -14179 -8118 -13899
rect -7158 -13899 -7148 -13890
rect -7114 -13890 -7108 -13865
rect -6136 -13395 -6130 -13370
rect -6096 -13370 -6082 -13361
rect -5122 -13361 -5062 -13081
rect -4110 -13081 -4094 -13080
rect -4060 -13080 -4054 -13047
rect -3082 -12577 -3076 -12543
rect -3042 -12577 -3036 -12543
rect -2072 -12543 -2012 -12384
rect -1562 -12434 -1502 -12384
rect -42 -12358 30 -12354
rect -42 -12410 -32 -12358
rect 20 -12410 30 -12358
rect -42 -12414 30 -12410
rect -1776 -12440 -1288 -12434
rect -1776 -12474 -1729 -12440
rect -1695 -12474 -1657 -12440
rect -1623 -12474 -1585 -12440
rect -1551 -12474 -1513 -12440
rect -1479 -12474 -1441 -12440
rect -1407 -12474 -1369 -12440
rect -1335 -12474 -1288 -12440
rect -1776 -12480 -1288 -12474
rect -758 -12440 -270 -12434
rect -758 -12474 -711 -12440
rect -677 -12474 -639 -12440
rect -605 -12474 -567 -12440
rect -533 -12474 -495 -12440
rect -461 -12474 -423 -12440
rect -389 -12474 -351 -12440
rect -317 -12474 -270 -12440
rect -758 -12480 -270 -12474
rect -2072 -12560 -2058 -12543
rect -3082 -12615 -3036 -12577
rect -3082 -12649 -3076 -12615
rect -3042 -12649 -3036 -12615
rect -3082 -12687 -3036 -12649
rect -3082 -12721 -3076 -12687
rect -3042 -12721 -3036 -12687
rect -3082 -12759 -3036 -12721
rect -3082 -12793 -3076 -12759
rect -3042 -12793 -3036 -12759
rect -3082 -12831 -3036 -12793
rect -3082 -12865 -3076 -12831
rect -3042 -12865 -3036 -12831
rect -3082 -12903 -3036 -12865
rect -3082 -12937 -3076 -12903
rect -3042 -12937 -3036 -12903
rect -3082 -12975 -3036 -12937
rect -3082 -13009 -3076 -12975
rect -3042 -13009 -3036 -12975
rect -3082 -13047 -3036 -13009
rect -3082 -13080 -3076 -13047
rect -4060 -13081 -4050 -13080
rect -4830 -13150 -4342 -13144
rect -4830 -13184 -4783 -13150
rect -4749 -13184 -4711 -13150
rect -4677 -13184 -4639 -13150
rect -4605 -13184 -4567 -13150
rect -4533 -13184 -4495 -13150
rect -4461 -13184 -4423 -13150
rect -4389 -13184 -4342 -13150
rect -4830 -13190 -4342 -13184
rect -4620 -13252 -4560 -13190
rect -4830 -13258 -4342 -13252
rect -4830 -13292 -4783 -13258
rect -4749 -13292 -4711 -13258
rect -4677 -13292 -4639 -13258
rect -4605 -13292 -4567 -13258
rect -4533 -13292 -4495 -13258
rect -4461 -13292 -4423 -13258
rect -4389 -13292 -4342 -13258
rect -4830 -13298 -4342 -13292
rect -5122 -13362 -5112 -13361
rect -6096 -13395 -6090 -13370
rect -6136 -13433 -6090 -13395
rect -6136 -13467 -6130 -13433
rect -6096 -13467 -6090 -13433
rect -6136 -13505 -6090 -13467
rect -6136 -13539 -6130 -13505
rect -6096 -13539 -6090 -13505
rect -6136 -13577 -6090 -13539
rect -6136 -13611 -6130 -13577
rect -6096 -13611 -6090 -13577
rect -6136 -13649 -6090 -13611
rect -6136 -13683 -6130 -13649
rect -6096 -13683 -6090 -13649
rect -6136 -13721 -6090 -13683
rect -6136 -13755 -6130 -13721
rect -6096 -13755 -6090 -13721
rect -6136 -13793 -6090 -13755
rect -6136 -13827 -6130 -13793
rect -6096 -13827 -6090 -13793
rect -6136 -13865 -6090 -13827
rect -7114 -13899 -7098 -13890
rect -6136 -13894 -6130 -13865
rect -7884 -13968 -7396 -13962
rect -7884 -14002 -7837 -13968
rect -7803 -14002 -7765 -13968
rect -7731 -14002 -7693 -13968
rect -7659 -14002 -7621 -13968
rect -7587 -14002 -7549 -13968
rect -7515 -14002 -7477 -13968
rect -7443 -14002 -7396 -13968
rect -7884 -14008 -7396 -14002
rect -7670 -14070 -7610 -14008
rect -7884 -14076 -7396 -14070
rect -7884 -14110 -7837 -14076
rect -7803 -14110 -7765 -14076
rect -7731 -14110 -7693 -14076
rect -7659 -14110 -7621 -14076
rect -7587 -14110 -7549 -14076
rect -7515 -14110 -7477 -14076
rect -7443 -14110 -7396 -14076
rect -7884 -14116 -7396 -14110
rect -8178 -14182 -8166 -14179
rect -9150 -14213 -9144 -14186
rect -9190 -14251 -9144 -14213
rect -9190 -14285 -9184 -14251
rect -9150 -14285 -9144 -14251
rect -9190 -14323 -9144 -14285
rect -9190 -14357 -9184 -14323
rect -9150 -14357 -9144 -14323
rect -9190 -14395 -9144 -14357
rect -9190 -14429 -9184 -14395
rect -9150 -14429 -9144 -14395
rect -9190 -14467 -9144 -14429
rect -9190 -14501 -9184 -14467
rect -9150 -14501 -9144 -14467
rect -9190 -14539 -9144 -14501
rect -9190 -14573 -9184 -14539
rect -9150 -14573 -9144 -14539
rect -9190 -14611 -9144 -14573
rect -9190 -14645 -9184 -14611
rect -9150 -14645 -9144 -14611
rect -9190 -14683 -9144 -14645
rect -9190 -14717 -9184 -14683
rect -9150 -14717 -9144 -14683
rect -9190 -14724 -9144 -14717
rect -8172 -14213 -8166 -14182
rect -8132 -14182 -8118 -14179
rect -7158 -14179 -7098 -13899
rect -6140 -13899 -6130 -13894
rect -6096 -13894 -6090 -13865
rect -5118 -13395 -5112 -13362
rect -5078 -13362 -5062 -13361
rect -4110 -13361 -4050 -13081
rect -3088 -13081 -3076 -13080
rect -3042 -13080 -3036 -13047
rect -2064 -12577 -2058 -12560
rect -2024 -12560 -2012 -12543
rect -1046 -12543 -1000 -12512
rect -2024 -12577 -2018 -12560
rect -2064 -12615 -2018 -12577
rect -2064 -12649 -2058 -12615
rect -2024 -12649 -2018 -12615
rect -2064 -12687 -2018 -12649
rect -2064 -12721 -2058 -12687
rect -2024 -12721 -2018 -12687
rect -2064 -12759 -2018 -12721
rect -2064 -12793 -2058 -12759
rect -2024 -12793 -2018 -12759
rect -2064 -12831 -2018 -12793
rect -2064 -12865 -2058 -12831
rect -2024 -12865 -2018 -12831
rect -2064 -12903 -2018 -12865
rect -2064 -12937 -2058 -12903
rect -2024 -12937 -2018 -12903
rect -2064 -12975 -2018 -12937
rect -2064 -13009 -2058 -12975
rect -2024 -13009 -2018 -12975
rect -2064 -13047 -2018 -13009
rect -2064 -13080 -2058 -13047
rect -3042 -13081 -3028 -13080
rect -3812 -13150 -3324 -13144
rect -3812 -13184 -3765 -13150
rect -3731 -13184 -3693 -13150
rect -3659 -13184 -3621 -13150
rect -3587 -13184 -3549 -13150
rect -3515 -13184 -3477 -13150
rect -3443 -13184 -3405 -13150
rect -3371 -13184 -3324 -13150
rect -3812 -13190 -3324 -13184
rect -3604 -13252 -3544 -13190
rect -3812 -13258 -3324 -13252
rect -3812 -13292 -3765 -13258
rect -3731 -13292 -3693 -13258
rect -3659 -13292 -3621 -13258
rect -3587 -13292 -3549 -13258
rect -3515 -13292 -3477 -13258
rect -3443 -13292 -3405 -13258
rect -3371 -13292 -3324 -13258
rect -3812 -13298 -3324 -13292
rect -5078 -13395 -5072 -13362
rect -4110 -13370 -4094 -13361
rect -5118 -13433 -5072 -13395
rect -5118 -13467 -5112 -13433
rect -5078 -13467 -5072 -13433
rect -5118 -13505 -5072 -13467
rect -5118 -13539 -5112 -13505
rect -5078 -13539 -5072 -13505
rect -5118 -13577 -5072 -13539
rect -5118 -13611 -5112 -13577
rect -5078 -13611 -5072 -13577
rect -5118 -13649 -5072 -13611
rect -5118 -13683 -5112 -13649
rect -5078 -13683 -5072 -13649
rect -5118 -13721 -5072 -13683
rect -5118 -13755 -5112 -13721
rect -5078 -13755 -5072 -13721
rect -5118 -13793 -5072 -13755
rect -5118 -13827 -5112 -13793
rect -5078 -13827 -5072 -13793
rect -5118 -13865 -5072 -13827
rect -5118 -13886 -5112 -13865
rect -6096 -13899 -6080 -13894
rect -6866 -13968 -6378 -13962
rect -6866 -14002 -6819 -13968
rect -6785 -14002 -6747 -13968
rect -6713 -14002 -6675 -13968
rect -6641 -14002 -6603 -13968
rect -6569 -14002 -6531 -13968
rect -6497 -14002 -6459 -13968
rect -6425 -14002 -6378 -13968
rect -6866 -14008 -6378 -14002
rect -6652 -14070 -6592 -14008
rect -6866 -14076 -6378 -14070
rect -6866 -14110 -6819 -14076
rect -6785 -14110 -6747 -14076
rect -6713 -14110 -6675 -14076
rect -6641 -14110 -6603 -14076
rect -6569 -14110 -6531 -14076
rect -6497 -14110 -6459 -14076
rect -6425 -14110 -6378 -14076
rect -6866 -14116 -6378 -14110
rect -7158 -14180 -7148 -14179
rect -8132 -14213 -8126 -14182
rect -8172 -14251 -8126 -14213
rect -8172 -14285 -8166 -14251
rect -8132 -14285 -8126 -14251
rect -8172 -14323 -8126 -14285
rect -8172 -14357 -8166 -14323
rect -8132 -14357 -8126 -14323
rect -8172 -14395 -8126 -14357
rect -8172 -14429 -8166 -14395
rect -8132 -14429 -8126 -14395
rect -8172 -14467 -8126 -14429
rect -8172 -14501 -8166 -14467
rect -8132 -14501 -8126 -14467
rect -8172 -14539 -8126 -14501
rect -8172 -14573 -8166 -14539
rect -8132 -14573 -8126 -14539
rect -8172 -14611 -8126 -14573
rect -8172 -14645 -8166 -14611
rect -8132 -14645 -8126 -14611
rect -8172 -14683 -8126 -14645
rect -8172 -14717 -8166 -14683
rect -8132 -14717 -8126 -14683
rect -8172 -14720 -8126 -14717
rect -7154 -14213 -7148 -14180
rect -7114 -14180 -7098 -14179
rect -6140 -14179 -6080 -13899
rect -5120 -13899 -5112 -13886
rect -5078 -13886 -5072 -13865
rect -4100 -13395 -4094 -13370
rect -4060 -13370 -4050 -13361
rect -3088 -13361 -3028 -13081
rect -2068 -13081 -2058 -13080
rect -2024 -13080 -2018 -13047
rect -1046 -12577 -1040 -12543
rect -1006 -12577 -1000 -12543
rect -36 -12543 24 -12414
rect -36 -12560 -22 -12543
rect -1046 -12615 -1000 -12577
rect -1046 -12649 -1040 -12615
rect -1006 -12649 -1000 -12615
rect -1046 -12687 -1000 -12649
rect -1046 -12721 -1040 -12687
rect -1006 -12721 -1000 -12687
rect -1046 -12759 -1000 -12721
rect -1046 -12793 -1040 -12759
rect -1006 -12793 -1000 -12759
rect -1046 -12831 -1000 -12793
rect -1046 -12865 -1040 -12831
rect -1006 -12865 -1000 -12831
rect -1046 -12903 -1000 -12865
rect -1046 -12937 -1040 -12903
rect -1006 -12937 -1000 -12903
rect -1046 -12975 -1000 -12937
rect -1046 -13009 -1040 -12975
rect -1006 -13009 -1000 -12975
rect -1046 -13047 -1000 -13009
rect -1046 -13076 -1040 -13047
rect -2024 -13081 -2008 -13080
rect -2794 -13150 -2306 -13144
rect -2794 -13184 -2747 -13150
rect -2713 -13184 -2675 -13150
rect -2641 -13184 -2603 -13150
rect -2569 -13184 -2531 -13150
rect -2497 -13184 -2459 -13150
rect -2425 -13184 -2387 -13150
rect -2353 -13184 -2306 -13150
rect -2794 -13190 -2306 -13184
rect -2582 -13252 -2522 -13190
rect -2794 -13258 -2306 -13252
rect -2794 -13292 -2747 -13258
rect -2713 -13292 -2675 -13258
rect -2641 -13292 -2603 -13258
rect -2569 -13292 -2531 -13258
rect -2497 -13292 -2459 -13258
rect -2425 -13292 -2387 -13258
rect -2353 -13292 -2306 -13258
rect -2794 -13298 -2306 -13292
rect -3088 -13370 -3076 -13361
rect -4060 -13395 -4054 -13370
rect -4100 -13433 -4054 -13395
rect -4100 -13467 -4094 -13433
rect -4060 -13467 -4054 -13433
rect -4100 -13505 -4054 -13467
rect -4100 -13539 -4094 -13505
rect -4060 -13539 -4054 -13505
rect -4100 -13577 -4054 -13539
rect -4100 -13611 -4094 -13577
rect -4060 -13611 -4054 -13577
rect -4100 -13649 -4054 -13611
rect -4100 -13683 -4094 -13649
rect -4060 -13683 -4054 -13649
rect -4100 -13721 -4054 -13683
rect -4100 -13755 -4094 -13721
rect -4060 -13755 -4054 -13721
rect -4100 -13793 -4054 -13755
rect -4100 -13827 -4094 -13793
rect -4060 -13827 -4054 -13793
rect -4100 -13865 -4054 -13827
rect -5078 -13899 -5060 -13886
rect -4100 -13894 -4094 -13865
rect -5848 -13968 -5360 -13962
rect -5848 -14002 -5801 -13968
rect -5767 -14002 -5729 -13968
rect -5695 -14002 -5657 -13968
rect -5623 -14002 -5585 -13968
rect -5551 -14002 -5513 -13968
rect -5479 -14002 -5441 -13968
rect -5407 -14002 -5360 -13968
rect -5848 -14008 -5360 -14002
rect -5650 -14070 -5590 -14008
rect -5848 -14076 -5360 -14070
rect -5848 -14110 -5801 -14076
rect -5767 -14110 -5729 -14076
rect -5695 -14110 -5657 -14076
rect -5623 -14110 -5585 -14076
rect -5551 -14110 -5513 -14076
rect -5479 -14110 -5441 -14076
rect -5407 -14110 -5360 -14076
rect -5848 -14116 -5360 -14110
rect -5120 -14176 -5060 -13899
rect -4108 -13899 -4094 -13894
rect -4060 -13894 -4054 -13865
rect -3082 -13395 -3076 -13370
rect -3042 -13370 -3028 -13361
rect -2068 -13361 -2008 -13081
rect -1052 -13081 -1040 -13076
rect -1006 -13076 -1000 -13047
rect -28 -12577 -22 -12560
rect 12 -12560 24 -12543
rect 12 -12577 18 -12560
rect -28 -12615 18 -12577
rect -28 -12649 -22 -12615
rect 12 -12649 18 -12615
rect -28 -12687 18 -12649
rect -28 -12721 -22 -12687
rect 12 -12721 18 -12687
rect -28 -12759 18 -12721
rect -28 -12793 -22 -12759
rect 12 -12793 18 -12759
rect -28 -12831 18 -12793
rect -28 -12865 -22 -12831
rect 12 -12865 18 -12831
rect -28 -12903 18 -12865
rect -28 -12937 -22 -12903
rect 12 -12937 18 -12903
rect -28 -12975 18 -12937
rect -28 -13009 -22 -12975
rect 12 -13009 18 -12975
rect -28 -13047 18 -13009
rect -1006 -13081 -992 -13076
rect -28 -13080 -22 -13047
rect -1776 -13150 -1288 -13144
rect -1776 -13184 -1729 -13150
rect -1695 -13184 -1657 -13150
rect -1623 -13184 -1585 -13150
rect -1551 -13184 -1513 -13150
rect -1479 -13184 -1441 -13150
rect -1407 -13184 -1369 -13150
rect -1335 -13184 -1288 -13150
rect -1776 -13190 -1288 -13184
rect -1570 -13252 -1510 -13190
rect -1776 -13258 -1288 -13252
rect -1776 -13292 -1729 -13258
rect -1695 -13292 -1657 -13258
rect -1623 -13292 -1585 -13258
rect -1551 -13292 -1513 -13258
rect -1479 -13292 -1441 -13258
rect -1407 -13292 -1369 -13258
rect -1335 -13292 -1288 -13258
rect -1776 -13298 -1288 -13292
rect -2068 -13370 -2058 -13361
rect -3042 -13395 -3036 -13370
rect -3082 -13433 -3036 -13395
rect -3082 -13467 -3076 -13433
rect -3042 -13467 -3036 -13433
rect -3082 -13505 -3036 -13467
rect -3082 -13539 -3076 -13505
rect -3042 -13539 -3036 -13505
rect -3082 -13577 -3036 -13539
rect -3082 -13611 -3076 -13577
rect -3042 -13611 -3036 -13577
rect -3082 -13649 -3036 -13611
rect -3082 -13683 -3076 -13649
rect -3042 -13683 -3036 -13649
rect -3082 -13721 -3036 -13683
rect -3082 -13755 -3076 -13721
rect -3042 -13755 -3036 -13721
rect -3082 -13793 -3036 -13755
rect -3082 -13827 -3076 -13793
rect -3042 -13827 -3036 -13793
rect -3082 -13865 -3036 -13827
rect -3082 -13894 -3076 -13865
rect -4060 -13899 -4048 -13894
rect -4830 -13968 -4342 -13962
rect -4830 -14002 -4783 -13968
rect -4749 -14002 -4711 -13968
rect -4677 -14002 -4639 -13968
rect -4605 -14002 -4567 -13968
rect -4533 -14002 -4495 -13968
rect -4461 -14002 -4423 -13968
rect -4389 -14002 -4342 -13968
rect -4830 -14008 -4342 -14002
rect -4620 -14070 -4560 -14008
rect -4830 -14076 -4342 -14070
rect -4830 -14110 -4783 -14076
rect -4749 -14110 -4711 -14076
rect -4677 -14110 -4639 -14076
rect -4605 -14110 -4567 -14076
rect -4533 -14110 -4495 -14076
rect -4461 -14110 -4423 -14076
rect -4389 -14110 -4342 -14076
rect -4830 -14116 -4342 -14110
rect -7114 -14213 -7108 -14180
rect -6140 -14184 -6130 -14179
rect -7154 -14251 -7108 -14213
rect -7154 -14285 -7148 -14251
rect -7114 -14285 -7108 -14251
rect -7154 -14323 -7108 -14285
rect -7154 -14357 -7148 -14323
rect -7114 -14357 -7108 -14323
rect -7154 -14395 -7108 -14357
rect -7154 -14429 -7148 -14395
rect -7114 -14429 -7108 -14395
rect -7154 -14467 -7108 -14429
rect -7154 -14501 -7148 -14467
rect -7114 -14501 -7108 -14467
rect -7154 -14539 -7108 -14501
rect -7154 -14573 -7148 -14539
rect -7114 -14573 -7108 -14539
rect -7154 -14611 -7108 -14573
rect -7154 -14645 -7148 -14611
rect -7114 -14645 -7108 -14611
rect -7154 -14683 -7108 -14645
rect -7154 -14717 -7148 -14683
rect -7114 -14717 -7108 -14683
rect -7154 -14718 -7108 -14717
rect -6136 -14213 -6130 -14184
rect -6096 -14184 -6080 -14179
rect -5118 -14179 -5072 -14176
rect -6096 -14213 -6090 -14184
rect -6136 -14251 -6090 -14213
rect -6136 -14285 -6130 -14251
rect -6096 -14285 -6090 -14251
rect -6136 -14323 -6090 -14285
rect -6136 -14357 -6130 -14323
rect -6096 -14357 -6090 -14323
rect -6136 -14395 -6090 -14357
rect -6136 -14429 -6130 -14395
rect -6096 -14429 -6090 -14395
rect -6136 -14467 -6090 -14429
rect -6136 -14501 -6130 -14467
rect -6096 -14501 -6090 -14467
rect -6136 -14539 -6090 -14501
rect -6136 -14573 -6130 -14539
rect -6096 -14573 -6090 -14539
rect -6136 -14611 -6090 -14573
rect -6136 -14645 -6130 -14611
rect -6096 -14645 -6090 -14611
rect -6136 -14683 -6090 -14645
rect -6136 -14717 -6130 -14683
rect -6096 -14717 -6090 -14683
rect -5118 -14213 -5112 -14179
rect -5078 -14213 -5072 -14179
rect -4108 -14179 -4048 -13899
rect -3086 -13899 -3076 -13894
rect -3042 -13894 -3036 -13865
rect -2064 -13395 -2058 -13370
rect -2024 -13370 -2008 -13361
rect -1052 -13361 -992 -13081
rect -30 -13081 -22 -13080
rect 12 -13080 18 -13047
rect 12 -13081 30 -13080
rect -758 -13150 -270 -13144
rect -758 -13184 -711 -13150
rect -677 -13184 -639 -13150
rect -605 -13184 -567 -13150
rect -533 -13184 -495 -13150
rect -461 -13184 -423 -13150
rect -389 -13184 -351 -13150
rect -317 -13184 -270 -13150
rect -758 -13190 -270 -13184
rect -550 -13252 -490 -13190
rect -758 -13258 -270 -13252
rect -758 -13292 -711 -13258
rect -677 -13292 -639 -13258
rect -605 -13292 -567 -13258
rect -533 -13292 -495 -13258
rect -461 -13292 -423 -13258
rect -389 -13292 -351 -13258
rect -317 -13292 -270 -13258
rect -758 -13298 -270 -13292
rect -1052 -13366 -1040 -13361
rect -2024 -13395 -2018 -13370
rect -2064 -13433 -2018 -13395
rect -2064 -13467 -2058 -13433
rect -2024 -13467 -2018 -13433
rect -2064 -13505 -2018 -13467
rect -2064 -13539 -2058 -13505
rect -2024 -13539 -2018 -13505
rect -2064 -13577 -2018 -13539
rect -2064 -13611 -2058 -13577
rect -2024 -13611 -2018 -13577
rect -2064 -13649 -2018 -13611
rect -2064 -13683 -2058 -13649
rect -2024 -13683 -2018 -13649
rect -2064 -13721 -2018 -13683
rect -2064 -13755 -2058 -13721
rect -2024 -13755 -2018 -13721
rect -2064 -13793 -2018 -13755
rect -2064 -13827 -2058 -13793
rect -2024 -13827 -2018 -13793
rect -2064 -13865 -2018 -13827
rect -2064 -13894 -2058 -13865
rect -3042 -13899 -3026 -13894
rect -3812 -13968 -3324 -13962
rect -3812 -14002 -3765 -13968
rect -3731 -14002 -3693 -13968
rect -3659 -14002 -3621 -13968
rect -3587 -14002 -3549 -13968
rect -3515 -14002 -3477 -13968
rect -3443 -14002 -3405 -13968
rect -3371 -14002 -3324 -13968
rect -3812 -14008 -3324 -14002
rect -3604 -14070 -3544 -14008
rect -3812 -14076 -3324 -14070
rect -3812 -14110 -3765 -14076
rect -3731 -14110 -3693 -14076
rect -3659 -14110 -3621 -14076
rect -3587 -14110 -3549 -14076
rect -3515 -14110 -3477 -14076
rect -3443 -14110 -3405 -14076
rect -3371 -14110 -3324 -14076
rect -3812 -14116 -3324 -14110
rect -4108 -14184 -4094 -14179
rect -5118 -14251 -5072 -14213
rect -5118 -14285 -5112 -14251
rect -5078 -14285 -5072 -14251
rect -5118 -14323 -5072 -14285
rect -5118 -14357 -5112 -14323
rect -5078 -14357 -5072 -14323
rect -5118 -14395 -5072 -14357
rect -5118 -14429 -5112 -14395
rect -5078 -14429 -5072 -14395
rect -5118 -14467 -5072 -14429
rect -5118 -14501 -5112 -14467
rect -5078 -14501 -5072 -14467
rect -5118 -14539 -5072 -14501
rect -5118 -14573 -5112 -14539
rect -5078 -14573 -5072 -14539
rect -5118 -14611 -5072 -14573
rect -5118 -14645 -5112 -14611
rect -5078 -14645 -5072 -14611
rect -5118 -14683 -5072 -14645
rect -5118 -14714 -5112 -14683
rect -12328 -14789 -12289 -14755
rect -12255 -14789 -12216 -14755
rect -12328 -14827 -12216 -14789
rect -12328 -14861 -12289 -14827
rect -12255 -14861 -12216 -14827
rect -12328 -14899 -12216 -14861
rect -12328 -14933 -12289 -14899
rect -12255 -14933 -12216 -14899
rect -12328 -14971 -12216 -14933
rect -12328 -15005 -12289 -14971
rect -12255 -15005 -12216 -14971
rect -12328 -15043 -12216 -15005
rect -9198 -14997 -9138 -14724
rect -8902 -14786 -8414 -14780
rect -8902 -14820 -8855 -14786
rect -8821 -14820 -8783 -14786
rect -8749 -14820 -8711 -14786
rect -8677 -14820 -8639 -14786
rect -8605 -14820 -8567 -14786
rect -8533 -14820 -8495 -14786
rect -8461 -14820 -8414 -14786
rect -8902 -14826 -8414 -14820
rect -8692 -14888 -8632 -14826
rect -8902 -14894 -8414 -14888
rect -8902 -14928 -8855 -14894
rect -8821 -14928 -8783 -14894
rect -8749 -14928 -8711 -14894
rect -8677 -14928 -8639 -14894
rect -8605 -14928 -8567 -14894
rect -8533 -14928 -8495 -14894
rect -8461 -14928 -8414 -14894
rect -8902 -14934 -8414 -14928
rect -9198 -15014 -9184 -14997
rect -12328 -15077 -12289 -15043
rect -12255 -15077 -12216 -15043
rect -12328 -15115 -12216 -15077
rect -12328 -15149 -12289 -15115
rect -12255 -15149 -12216 -15115
rect -12328 -15187 -12216 -15149
rect -12328 -15221 -12289 -15187
rect -12255 -15221 -12216 -15187
rect -12328 -15259 -12216 -15221
rect -12328 -15293 -12289 -15259
rect -12255 -15293 -12216 -15259
rect -12328 -15331 -12216 -15293
rect -12328 -15365 -12289 -15331
rect -12255 -15365 -12216 -15331
rect -12328 -15403 -12216 -15365
rect -12328 -15437 -12289 -15403
rect -12255 -15437 -12216 -15403
rect -12328 -15475 -12216 -15437
rect -12328 -15509 -12289 -15475
rect -12255 -15509 -12216 -15475
rect -12328 -15547 -12216 -15509
rect -9190 -15031 -9184 -15014
rect -9150 -15014 -9138 -14997
rect -8178 -14997 -8118 -14720
rect -7884 -14786 -7396 -14780
rect -7884 -14820 -7837 -14786
rect -7803 -14820 -7765 -14786
rect -7731 -14820 -7693 -14786
rect -7659 -14820 -7621 -14786
rect -7587 -14820 -7549 -14786
rect -7515 -14820 -7477 -14786
rect -7443 -14820 -7396 -14786
rect -7884 -14826 -7396 -14820
rect -7670 -14888 -7610 -14826
rect -7884 -14894 -7396 -14888
rect -7884 -14928 -7837 -14894
rect -7803 -14928 -7765 -14894
rect -7731 -14928 -7693 -14894
rect -7659 -14928 -7621 -14894
rect -7587 -14928 -7549 -14894
rect -7515 -14928 -7477 -14894
rect -7443 -14928 -7396 -14894
rect -7884 -14934 -7396 -14928
rect -8178 -15010 -8166 -14997
rect -9150 -15031 -9144 -15014
rect -9190 -15069 -9144 -15031
rect -9190 -15103 -9184 -15069
rect -9150 -15103 -9144 -15069
rect -9190 -15141 -9144 -15103
rect -9190 -15175 -9184 -15141
rect -9150 -15175 -9144 -15141
rect -9190 -15213 -9144 -15175
rect -9190 -15247 -9184 -15213
rect -9150 -15247 -9144 -15213
rect -9190 -15285 -9144 -15247
rect -9190 -15319 -9184 -15285
rect -9150 -15319 -9144 -15285
rect -9190 -15357 -9144 -15319
rect -9190 -15391 -9184 -15357
rect -9150 -15391 -9144 -15357
rect -9190 -15429 -9144 -15391
rect -9190 -15463 -9184 -15429
rect -9150 -15463 -9144 -15429
rect -9190 -15501 -9144 -15463
rect -9190 -15535 -9184 -15501
rect -9150 -15535 -9144 -15501
rect -8172 -15031 -8166 -15010
rect -8132 -15010 -8118 -14997
rect -7158 -14997 -7098 -14718
rect -6136 -14722 -6090 -14717
rect -5120 -14717 -5112 -14714
rect -5078 -14714 -5072 -14683
rect -4100 -14213 -4094 -14184
rect -4060 -14184 -4048 -14179
rect -3086 -14179 -3026 -13899
rect -2066 -13899 -2058 -13894
rect -2024 -13894 -2018 -13865
rect -1046 -13395 -1040 -13366
rect -1006 -13366 -992 -13361
rect -30 -13361 30 -13081
rect -1006 -13395 -1000 -13366
rect -30 -13370 -22 -13361
rect -1046 -13433 -1000 -13395
rect -1046 -13467 -1040 -13433
rect -1006 -13467 -1000 -13433
rect -1046 -13505 -1000 -13467
rect -1046 -13539 -1040 -13505
rect -1006 -13539 -1000 -13505
rect -1046 -13577 -1000 -13539
rect -1046 -13611 -1040 -13577
rect -1006 -13611 -1000 -13577
rect -1046 -13649 -1000 -13611
rect -1046 -13683 -1040 -13649
rect -1006 -13683 -1000 -13649
rect -1046 -13721 -1000 -13683
rect -1046 -13755 -1040 -13721
rect -1006 -13755 -1000 -13721
rect -1046 -13793 -1000 -13755
rect -1046 -13827 -1040 -13793
rect -1006 -13827 -1000 -13793
rect -1046 -13865 -1000 -13827
rect -1046 -13890 -1040 -13865
rect -2024 -13899 -2006 -13894
rect -2794 -13968 -2306 -13962
rect -2794 -14002 -2747 -13968
rect -2713 -14002 -2675 -13968
rect -2641 -14002 -2603 -13968
rect -2569 -14002 -2531 -13968
rect -2497 -14002 -2459 -13968
rect -2425 -14002 -2387 -13968
rect -2353 -14002 -2306 -13968
rect -2794 -14008 -2306 -14002
rect -2582 -14070 -2522 -14008
rect -2794 -14076 -2306 -14070
rect -2794 -14110 -2747 -14076
rect -2713 -14110 -2675 -14076
rect -2641 -14110 -2603 -14076
rect -2569 -14110 -2531 -14076
rect -2497 -14110 -2459 -14076
rect -2425 -14110 -2387 -14076
rect -2353 -14110 -2306 -14076
rect -2794 -14116 -2306 -14110
rect -3086 -14184 -3076 -14179
rect -4060 -14213 -4054 -14184
rect -4100 -14251 -4054 -14213
rect -4100 -14285 -4094 -14251
rect -4060 -14285 -4054 -14251
rect -4100 -14323 -4054 -14285
rect -4100 -14357 -4094 -14323
rect -4060 -14357 -4054 -14323
rect -4100 -14395 -4054 -14357
rect -4100 -14429 -4094 -14395
rect -4060 -14429 -4054 -14395
rect -4100 -14467 -4054 -14429
rect -4100 -14501 -4094 -14467
rect -4060 -14501 -4054 -14467
rect -4100 -14539 -4054 -14501
rect -4100 -14573 -4094 -14539
rect -4060 -14573 -4054 -14539
rect -4100 -14611 -4054 -14573
rect -4100 -14645 -4094 -14611
rect -4060 -14645 -4054 -14611
rect -4100 -14683 -4054 -14645
rect -5078 -14717 -5060 -14714
rect -6866 -14786 -6378 -14780
rect -6866 -14820 -6819 -14786
rect -6785 -14820 -6747 -14786
rect -6713 -14820 -6675 -14786
rect -6641 -14820 -6603 -14786
rect -6569 -14820 -6531 -14786
rect -6497 -14820 -6459 -14786
rect -6425 -14820 -6378 -14786
rect -6866 -14826 -6378 -14820
rect -6658 -14888 -6598 -14826
rect -6866 -14894 -6378 -14888
rect -6866 -14928 -6819 -14894
rect -6785 -14928 -6747 -14894
rect -6713 -14928 -6675 -14894
rect -6641 -14928 -6603 -14894
rect -6569 -14928 -6531 -14894
rect -6497 -14928 -6459 -14894
rect -6425 -14928 -6378 -14894
rect -6866 -14934 -6378 -14928
rect -7158 -15008 -7148 -14997
rect -8132 -15031 -8126 -15010
rect -8172 -15069 -8126 -15031
rect -8172 -15103 -8166 -15069
rect -8132 -15103 -8126 -15069
rect -8172 -15141 -8126 -15103
rect -8172 -15175 -8166 -15141
rect -8132 -15175 -8126 -15141
rect -8172 -15213 -8126 -15175
rect -8172 -15247 -8166 -15213
rect -8132 -15247 -8126 -15213
rect -8172 -15285 -8126 -15247
rect -8172 -15319 -8166 -15285
rect -8132 -15319 -8126 -15285
rect -8172 -15357 -8126 -15319
rect -8172 -15391 -8166 -15357
rect -8132 -15391 -8126 -15357
rect -8172 -15429 -8126 -15391
rect -8172 -15463 -8166 -15429
rect -8132 -15463 -8126 -15429
rect -8172 -15501 -8126 -15463
rect -8172 -15532 -8166 -15501
rect -9190 -15536 -9144 -15535
rect -8178 -15535 -8166 -15532
rect -8132 -15532 -8126 -15501
rect -7154 -15031 -7148 -15008
rect -7114 -15008 -7098 -14997
rect -6140 -14997 -6080 -14722
rect -5848 -14786 -5360 -14780
rect -5848 -14820 -5801 -14786
rect -5767 -14820 -5729 -14786
rect -5695 -14820 -5657 -14786
rect -5623 -14820 -5585 -14786
rect -5551 -14820 -5513 -14786
rect -5479 -14820 -5441 -14786
rect -5407 -14820 -5360 -14786
rect -5848 -14826 -5360 -14820
rect -5656 -14888 -5596 -14826
rect -5848 -14894 -5360 -14888
rect -5848 -14928 -5801 -14894
rect -5767 -14928 -5729 -14894
rect -5695 -14928 -5657 -14894
rect -5623 -14928 -5585 -14894
rect -5551 -14928 -5513 -14894
rect -5479 -14928 -5441 -14894
rect -5407 -14928 -5360 -14894
rect -5848 -14934 -5360 -14928
rect -7114 -15031 -7108 -15008
rect -6140 -15012 -6130 -14997
rect -7154 -15069 -7108 -15031
rect -7154 -15103 -7148 -15069
rect -7114 -15103 -7108 -15069
rect -7154 -15141 -7108 -15103
rect -7154 -15175 -7148 -15141
rect -7114 -15175 -7108 -15141
rect -7154 -15213 -7108 -15175
rect -7154 -15247 -7148 -15213
rect -7114 -15247 -7108 -15213
rect -7154 -15285 -7108 -15247
rect -7154 -15319 -7148 -15285
rect -7114 -15319 -7108 -15285
rect -7154 -15357 -7108 -15319
rect -7154 -15391 -7148 -15357
rect -7114 -15391 -7108 -15357
rect -7154 -15429 -7108 -15391
rect -7154 -15463 -7148 -15429
rect -7114 -15463 -7108 -15429
rect -7154 -15501 -7108 -15463
rect -7154 -15530 -7148 -15501
rect -8132 -15535 -8118 -15532
rect -12328 -15581 -12289 -15547
rect -12255 -15581 -12216 -15547
rect -12328 -15619 -12216 -15581
rect -12328 -15653 -12289 -15619
rect -12255 -15653 -12216 -15619
rect -12328 -15691 -12216 -15653
rect -12328 -15725 -12289 -15691
rect -12255 -15725 -12216 -15691
rect -12328 -15763 -12216 -15725
rect -12328 -15797 -12289 -15763
rect -12255 -15797 -12216 -15763
rect -12328 -15835 -12216 -15797
rect -9198 -15815 -9138 -15536
rect -8902 -15604 -8414 -15598
rect -8902 -15638 -8855 -15604
rect -8821 -15638 -8783 -15604
rect -8749 -15638 -8711 -15604
rect -8677 -15638 -8639 -15604
rect -8605 -15638 -8567 -15604
rect -8533 -15638 -8495 -15604
rect -8461 -15638 -8414 -15604
rect -8902 -15644 -8414 -15638
rect -8694 -15706 -8634 -15644
rect -8902 -15712 -8414 -15706
rect -8902 -15746 -8855 -15712
rect -8821 -15746 -8783 -15712
rect -8749 -15746 -8711 -15712
rect -8677 -15746 -8639 -15712
rect -8605 -15746 -8567 -15712
rect -8533 -15746 -8495 -15712
rect -8461 -15746 -8414 -15712
rect -8902 -15752 -8414 -15746
rect -9198 -15826 -9184 -15815
rect -12328 -15869 -12289 -15835
rect -12255 -15869 -12216 -15835
rect -12328 -15907 -12216 -15869
rect -12328 -15941 -12289 -15907
rect -12255 -15941 -12216 -15907
rect -12328 -15979 -12216 -15941
rect -12328 -16013 -12289 -15979
rect -12255 -16013 -12216 -15979
rect -12328 -16051 -12216 -16013
rect -12328 -16085 -12289 -16051
rect -12255 -16085 -12216 -16051
rect -12328 -16123 -12216 -16085
rect -12328 -16157 -12289 -16123
rect -12255 -16157 -12216 -16123
rect -12328 -16195 -12216 -16157
rect -12328 -16229 -12289 -16195
rect -12255 -16229 -12216 -16195
rect -12328 -16267 -12216 -16229
rect -12328 -16301 -12289 -16267
rect -12255 -16301 -12216 -16267
rect -12328 -16339 -12216 -16301
rect -12328 -16373 -12289 -16339
rect -12255 -16373 -12216 -16339
rect -9190 -15849 -9184 -15826
rect -9150 -15826 -9138 -15815
rect -8178 -15815 -8118 -15535
rect -7158 -15535 -7148 -15530
rect -7114 -15530 -7108 -15501
rect -6136 -15031 -6130 -15012
rect -6096 -15012 -6080 -14997
rect -5120 -14997 -5060 -14717
rect -4100 -14717 -4094 -14683
rect -4060 -14717 -4054 -14683
rect -4100 -14722 -4054 -14717
rect -3082 -14213 -3076 -14184
rect -3042 -14184 -3026 -14179
rect -2066 -14179 -2006 -13899
rect -1050 -13899 -1040 -13890
rect -1006 -13890 -1000 -13865
rect -28 -13395 -22 -13370
rect 12 -13370 30 -13361
rect 12 -13395 18 -13370
rect -28 -13433 18 -13395
rect -28 -13467 -22 -13433
rect 12 -13467 18 -13433
rect -28 -13505 18 -13467
rect -28 -13539 -22 -13505
rect 12 -13539 18 -13505
rect -28 -13577 18 -13539
rect -28 -13611 -22 -13577
rect 12 -13611 18 -13577
rect -28 -13649 18 -13611
rect -28 -13683 -22 -13649
rect 12 -13683 18 -13649
rect -28 -13721 18 -13683
rect -28 -13755 -22 -13721
rect 12 -13755 18 -13721
rect -28 -13793 18 -13755
rect -28 -13827 -22 -13793
rect 12 -13827 18 -13793
rect -28 -13865 18 -13827
rect -1006 -13899 -990 -13890
rect -1776 -13968 -1288 -13962
rect -1776 -14002 -1729 -13968
rect -1695 -14002 -1657 -13968
rect -1623 -14002 -1585 -13968
rect -1551 -14002 -1513 -13968
rect -1479 -14002 -1441 -13968
rect -1407 -14002 -1369 -13968
rect -1335 -14002 -1288 -13968
rect -1776 -14008 -1288 -14002
rect -1570 -14070 -1510 -14008
rect -1776 -14076 -1288 -14070
rect -1776 -14110 -1729 -14076
rect -1695 -14110 -1657 -14076
rect -1623 -14110 -1585 -14076
rect -1551 -14110 -1513 -14076
rect -1479 -14110 -1441 -14076
rect -1407 -14110 -1369 -14076
rect -1335 -14110 -1288 -14076
rect -1776 -14116 -1288 -14110
rect -2066 -14184 -2058 -14179
rect -3042 -14213 -3036 -14184
rect -3082 -14251 -3036 -14213
rect -3082 -14285 -3076 -14251
rect -3042 -14285 -3036 -14251
rect -3082 -14323 -3036 -14285
rect -3082 -14357 -3076 -14323
rect -3042 -14357 -3036 -14323
rect -3082 -14395 -3036 -14357
rect -3082 -14429 -3076 -14395
rect -3042 -14429 -3036 -14395
rect -3082 -14467 -3036 -14429
rect -3082 -14501 -3076 -14467
rect -3042 -14501 -3036 -14467
rect -3082 -14539 -3036 -14501
rect -3082 -14573 -3076 -14539
rect -3042 -14573 -3036 -14539
rect -3082 -14611 -3036 -14573
rect -3082 -14645 -3076 -14611
rect -3042 -14645 -3036 -14611
rect -3082 -14683 -3036 -14645
rect -3082 -14717 -3076 -14683
rect -3042 -14717 -3036 -14683
rect -3082 -14722 -3036 -14717
rect -2064 -14213 -2058 -14184
rect -2024 -14184 -2006 -14179
rect -1050 -14179 -990 -13899
rect -28 -13899 -22 -13865
rect 12 -13894 18 -13865
rect 12 -13899 32 -13894
rect -758 -13968 -270 -13962
rect -758 -14002 -711 -13968
rect -677 -14002 -639 -13968
rect -605 -14002 -567 -13968
rect -533 -14002 -495 -13968
rect -461 -14002 -423 -13968
rect -389 -14002 -351 -13968
rect -317 -14002 -270 -13968
rect -758 -14008 -270 -14002
rect -550 -14070 -490 -14008
rect -758 -14076 -270 -14070
rect -758 -14110 -711 -14076
rect -677 -14110 -639 -14076
rect -605 -14110 -567 -14076
rect -533 -14110 -495 -14076
rect -461 -14110 -423 -14076
rect -389 -14110 -351 -14076
rect -317 -14110 -270 -14076
rect -758 -14116 -270 -14110
rect -1050 -14180 -1040 -14179
rect -2024 -14213 -2018 -14184
rect -2064 -14251 -2018 -14213
rect -2064 -14285 -2058 -14251
rect -2024 -14285 -2018 -14251
rect -2064 -14323 -2018 -14285
rect -2064 -14357 -2058 -14323
rect -2024 -14357 -2018 -14323
rect -2064 -14395 -2018 -14357
rect -2064 -14429 -2058 -14395
rect -2024 -14429 -2018 -14395
rect -2064 -14467 -2018 -14429
rect -2064 -14501 -2058 -14467
rect -2024 -14501 -2018 -14467
rect -2064 -14539 -2018 -14501
rect -2064 -14573 -2058 -14539
rect -2024 -14573 -2018 -14539
rect -2064 -14611 -2018 -14573
rect -2064 -14645 -2058 -14611
rect -2024 -14645 -2018 -14611
rect -2064 -14683 -2018 -14645
rect -2064 -14717 -2058 -14683
rect -2024 -14717 -2018 -14683
rect -2064 -14722 -2018 -14717
rect -1046 -14213 -1040 -14180
rect -1006 -14180 -990 -14179
rect -28 -14179 32 -13899
rect -1006 -14213 -1000 -14180
rect -1046 -14251 -1000 -14213
rect -1046 -14285 -1040 -14251
rect -1006 -14285 -1000 -14251
rect -1046 -14323 -1000 -14285
rect -1046 -14357 -1040 -14323
rect -1006 -14357 -1000 -14323
rect -1046 -14395 -1000 -14357
rect -1046 -14429 -1040 -14395
rect -1006 -14429 -1000 -14395
rect -1046 -14467 -1000 -14429
rect -1046 -14501 -1040 -14467
rect -1006 -14501 -1000 -14467
rect -1046 -14539 -1000 -14501
rect -1046 -14573 -1040 -14539
rect -1006 -14573 -1000 -14539
rect -1046 -14611 -1000 -14573
rect -1046 -14645 -1040 -14611
rect -1006 -14645 -1000 -14611
rect -1046 -14683 -1000 -14645
rect -1046 -14717 -1040 -14683
rect -1006 -14717 -1000 -14683
rect -1046 -14718 -1000 -14717
rect -28 -14213 -22 -14179
rect 12 -14184 32 -14179
rect 12 -14213 18 -14184
rect -28 -14251 18 -14213
rect -28 -14285 -22 -14251
rect 12 -14285 18 -14251
rect -28 -14323 18 -14285
rect -28 -14357 -22 -14323
rect 12 -14357 18 -14323
rect -28 -14395 18 -14357
rect -28 -14429 -22 -14395
rect 12 -14429 18 -14395
rect -28 -14467 18 -14429
rect -28 -14501 -22 -14467
rect 12 -14501 18 -14467
rect -28 -14539 18 -14501
rect -28 -14573 -22 -14539
rect 12 -14573 18 -14539
rect -28 -14611 18 -14573
rect -28 -14645 -22 -14611
rect 12 -14645 18 -14611
rect -28 -14683 18 -14645
rect -28 -14717 -22 -14683
rect 12 -14717 18 -14683
rect -4830 -14786 -4342 -14780
rect -4830 -14820 -4783 -14786
rect -4749 -14820 -4711 -14786
rect -4677 -14820 -4639 -14786
rect -4605 -14820 -4567 -14786
rect -4533 -14820 -4495 -14786
rect -4461 -14820 -4423 -14786
rect -4389 -14820 -4342 -14786
rect -4830 -14826 -4342 -14820
rect -4626 -14888 -4566 -14826
rect -4830 -14894 -4342 -14888
rect -4830 -14928 -4783 -14894
rect -4749 -14928 -4711 -14894
rect -4677 -14928 -4639 -14894
rect -4605 -14928 -4567 -14894
rect -4533 -14928 -4495 -14894
rect -4461 -14928 -4423 -14894
rect -4389 -14928 -4342 -14894
rect -4830 -14934 -4342 -14928
rect -5120 -15004 -5112 -14997
rect -6096 -15031 -6090 -15012
rect -6136 -15069 -6090 -15031
rect -6136 -15103 -6130 -15069
rect -6096 -15103 -6090 -15069
rect -6136 -15141 -6090 -15103
rect -6136 -15175 -6130 -15141
rect -6096 -15175 -6090 -15141
rect -6136 -15213 -6090 -15175
rect -6136 -15247 -6130 -15213
rect -6096 -15247 -6090 -15213
rect -6136 -15285 -6090 -15247
rect -6136 -15319 -6130 -15285
rect -6096 -15319 -6090 -15285
rect -6136 -15357 -6090 -15319
rect -6136 -15391 -6130 -15357
rect -6096 -15391 -6090 -15357
rect -6136 -15429 -6090 -15391
rect -6136 -15463 -6130 -15429
rect -6096 -15463 -6090 -15429
rect -6136 -15501 -6090 -15463
rect -7114 -15535 -7098 -15530
rect -6136 -15534 -6130 -15501
rect -7884 -15604 -7396 -15598
rect -7884 -15638 -7837 -15604
rect -7803 -15638 -7765 -15604
rect -7731 -15638 -7693 -15604
rect -7659 -15638 -7621 -15604
rect -7587 -15638 -7549 -15604
rect -7515 -15638 -7477 -15604
rect -7443 -15638 -7396 -15604
rect -7884 -15644 -7396 -15638
rect -7676 -15706 -7616 -15644
rect -7884 -15712 -7396 -15706
rect -7884 -15746 -7837 -15712
rect -7803 -15746 -7765 -15712
rect -7731 -15746 -7693 -15712
rect -7659 -15746 -7621 -15712
rect -7587 -15746 -7549 -15712
rect -7515 -15746 -7477 -15712
rect -7443 -15746 -7396 -15712
rect -7884 -15752 -7396 -15746
rect -8178 -15822 -8166 -15815
rect -9150 -15849 -9144 -15826
rect -9190 -15887 -9144 -15849
rect -9190 -15921 -9184 -15887
rect -9150 -15921 -9144 -15887
rect -9190 -15959 -9144 -15921
rect -9190 -15993 -9184 -15959
rect -9150 -15993 -9144 -15959
rect -9190 -16031 -9144 -15993
rect -9190 -16065 -9184 -16031
rect -9150 -16065 -9144 -16031
rect -9190 -16103 -9144 -16065
rect -9190 -16137 -9184 -16103
rect -9150 -16137 -9144 -16103
rect -9190 -16175 -9144 -16137
rect -9190 -16209 -9184 -16175
rect -9150 -16209 -9144 -16175
rect -9190 -16247 -9144 -16209
rect -9190 -16281 -9184 -16247
rect -9150 -16281 -9144 -16247
rect -9190 -16319 -9144 -16281
rect -9190 -16353 -9184 -16319
rect -9150 -16353 -9144 -16319
rect -8172 -15849 -8166 -15822
rect -8132 -15822 -8118 -15815
rect -7158 -15815 -7098 -15535
rect -6140 -15535 -6130 -15534
rect -6096 -15534 -6090 -15501
rect -5118 -15031 -5112 -15004
rect -5078 -15004 -5060 -14997
rect -4108 -14997 -4048 -14722
rect -3812 -14786 -3324 -14780
rect -3812 -14820 -3765 -14786
rect -3731 -14820 -3693 -14786
rect -3659 -14820 -3621 -14786
rect -3587 -14820 -3549 -14786
rect -3515 -14820 -3477 -14786
rect -3443 -14820 -3405 -14786
rect -3371 -14820 -3324 -14786
rect -3812 -14826 -3324 -14820
rect -3610 -14888 -3550 -14826
rect -3812 -14894 -3324 -14888
rect -3812 -14928 -3765 -14894
rect -3731 -14928 -3693 -14894
rect -3659 -14928 -3621 -14894
rect -3587 -14928 -3549 -14894
rect -3515 -14928 -3477 -14894
rect -3443 -14928 -3405 -14894
rect -3371 -14928 -3324 -14894
rect -3812 -14934 -3324 -14928
rect -5078 -15031 -5072 -15004
rect -4108 -15012 -4094 -14997
rect -5118 -15069 -5072 -15031
rect -5118 -15103 -5112 -15069
rect -5078 -15103 -5072 -15069
rect -5118 -15141 -5072 -15103
rect -5118 -15175 -5112 -15141
rect -5078 -15175 -5072 -15141
rect -5118 -15213 -5072 -15175
rect -5118 -15247 -5112 -15213
rect -5078 -15247 -5072 -15213
rect -5118 -15285 -5072 -15247
rect -5118 -15319 -5112 -15285
rect -5078 -15319 -5072 -15285
rect -5118 -15357 -5072 -15319
rect -5118 -15391 -5112 -15357
rect -5078 -15391 -5072 -15357
rect -5118 -15429 -5072 -15391
rect -5118 -15463 -5112 -15429
rect -5078 -15463 -5072 -15429
rect -5118 -15501 -5072 -15463
rect -5118 -15526 -5112 -15501
rect -6096 -15535 -6080 -15534
rect -6866 -15604 -6378 -15598
rect -6866 -15638 -6819 -15604
rect -6785 -15638 -6747 -15604
rect -6713 -15638 -6675 -15604
rect -6641 -15638 -6603 -15604
rect -6569 -15638 -6531 -15604
rect -6497 -15638 -6459 -15604
rect -6425 -15638 -6378 -15604
rect -6866 -15644 -6378 -15638
rect -6660 -15706 -6600 -15644
rect -6866 -15712 -6378 -15706
rect -6866 -15746 -6819 -15712
rect -6785 -15746 -6747 -15712
rect -6713 -15746 -6675 -15712
rect -6641 -15746 -6603 -15712
rect -6569 -15746 -6531 -15712
rect -6497 -15746 -6459 -15712
rect -6425 -15746 -6378 -15712
rect -6866 -15752 -6378 -15746
rect -7158 -15820 -7148 -15815
rect -8132 -15849 -8126 -15822
rect -8172 -15887 -8126 -15849
rect -8172 -15921 -8166 -15887
rect -8132 -15921 -8126 -15887
rect -8172 -15959 -8126 -15921
rect -8172 -15993 -8166 -15959
rect -8132 -15993 -8126 -15959
rect -8172 -16031 -8126 -15993
rect -8172 -16065 -8166 -16031
rect -8132 -16065 -8126 -16031
rect -8172 -16103 -8126 -16065
rect -8172 -16137 -8166 -16103
rect -8132 -16137 -8126 -16103
rect -8172 -16175 -8126 -16137
rect -8172 -16209 -8166 -16175
rect -8132 -16209 -8126 -16175
rect -8172 -16247 -8126 -16209
rect -8172 -16281 -8166 -16247
rect -8132 -16281 -8126 -16247
rect -8172 -16319 -8126 -16281
rect -8172 -16352 -8166 -16319
rect -9190 -16356 -9144 -16353
rect -8178 -16353 -8166 -16352
rect -8132 -16352 -8126 -16319
rect -7154 -15849 -7148 -15820
rect -7114 -15820 -7098 -15815
rect -6140 -15815 -6080 -15535
rect -5120 -15535 -5112 -15526
rect -5078 -15526 -5072 -15501
rect -4100 -15031 -4094 -15012
rect -4060 -15012 -4048 -14997
rect -3086 -14997 -3026 -14722
rect -2794 -14786 -2306 -14780
rect -2794 -14820 -2747 -14786
rect -2713 -14820 -2675 -14786
rect -2641 -14820 -2603 -14786
rect -2569 -14820 -2531 -14786
rect -2497 -14820 -2459 -14786
rect -2425 -14820 -2387 -14786
rect -2353 -14820 -2306 -14786
rect -2794 -14826 -2306 -14820
rect -2588 -14888 -2528 -14826
rect -2794 -14894 -2306 -14888
rect -2794 -14928 -2747 -14894
rect -2713 -14928 -2675 -14894
rect -2641 -14928 -2603 -14894
rect -2569 -14928 -2531 -14894
rect -2497 -14928 -2459 -14894
rect -2425 -14928 -2387 -14894
rect -2353 -14928 -2306 -14894
rect -2794 -14934 -2306 -14928
rect -3086 -15012 -3076 -14997
rect -4060 -15031 -4054 -15012
rect -4100 -15069 -4054 -15031
rect -4100 -15103 -4094 -15069
rect -4060 -15103 -4054 -15069
rect -4100 -15141 -4054 -15103
rect -4100 -15175 -4094 -15141
rect -4060 -15175 -4054 -15141
rect -4100 -15213 -4054 -15175
rect -4100 -15247 -4094 -15213
rect -4060 -15247 -4054 -15213
rect -4100 -15285 -4054 -15247
rect -4100 -15319 -4094 -15285
rect -4060 -15319 -4054 -15285
rect -4100 -15357 -4054 -15319
rect -4100 -15391 -4094 -15357
rect -4060 -15391 -4054 -15357
rect -4100 -15429 -4054 -15391
rect -4100 -15463 -4094 -15429
rect -4060 -15463 -4054 -15429
rect -4100 -15501 -4054 -15463
rect -5078 -15535 -5060 -15526
rect -4100 -15534 -4094 -15501
rect -5848 -15604 -5360 -15598
rect -5848 -15638 -5801 -15604
rect -5767 -15638 -5729 -15604
rect -5695 -15638 -5657 -15604
rect -5623 -15638 -5585 -15604
rect -5551 -15638 -5513 -15604
rect -5479 -15638 -5441 -15604
rect -5407 -15638 -5360 -15604
rect -5848 -15644 -5360 -15638
rect -5658 -15706 -5598 -15644
rect -5848 -15712 -5360 -15706
rect -5848 -15746 -5801 -15712
rect -5767 -15746 -5729 -15712
rect -5695 -15746 -5657 -15712
rect -5623 -15746 -5585 -15712
rect -5551 -15746 -5513 -15712
rect -5479 -15746 -5441 -15712
rect -5407 -15746 -5360 -15712
rect -5848 -15752 -5360 -15746
rect -7114 -15849 -7108 -15820
rect -6140 -15824 -6130 -15815
rect -7154 -15887 -7108 -15849
rect -7154 -15921 -7148 -15887
rect -7114 -15921 -7108 -15887
rect -7154 -15959 -7108 -15921
rect -7154 -15993 -7148 -15959
rect -7114 -15993 -7108 -15959
rect -7154 -16031 -7108 -15993
rect -7154 -16065 -7148 -16031
rect -7114 -16065 -7108 -16031
rect -7154 -16103 -7108 -16065
rect -7154 -16137 -7148 -16103
rect -7114 -16137 -7108 -16103
rect -7154 -16175 -7108 -16137
rect -7154 -16209 -7148 -16175
rect -7114 -16209 -7108 -16175
rect -7154 -16247 -7108 -16209
rect -7154 -16281 -7148 -16247
rect -7114 -16281 -7108 -16247
rect -7154 -16319 -7108 -16281
rect -7154 -16350 -7148 -16319
rect -8132 -16353 -8118 -16352
rect -12328 -16411 -12216 -16373
rect -12328 -16445 -12289 -16411
rect -12255 -16445 -12216 -16411
rect -12328 -16483 -12216 -16445
rect -12328 -16517 -12289 -16483
rect -12255 -16517 -12216 -16483
rect -12328 -16555 -12216 -16517
rect -12328 -16589 -12289 -16555
rect -12255 -16589 -12216 -16555
rect -12328 -16627 -12216 -16589
rect -12328 -16661 -12289 -16627
rect -12255 -16661 -12216 -16627
rect -9198 -16633 -9138 -16356
rect -8902 -16422 -8414 -16416
rect -8902 -16456 -8855 -16422
rect -8821 -16456 -8783 -16422
rect -8749 -16456 -8711 -16422
rect -8677 -16456 -8639 -16422
rect -8605 -16456 -8567 -16422
rect -8533 -16456 -8495 -16422
rect -8461 -16456 -8414 -16422
rect -8902 -16462 -8414 -16456
rect -8692 -16524 -8632 -16462
rect -8902 -16530 -8414 -16524
rect -8902 -16564 -8855 -16530
rect -8821 -16564 -8783 -16530
rect -8749 -16564 -8711 -16530
rect -8677 -16564 -8639 -16530
rect -8605 -16564 -8567 -16530
rect -8533 -16564 -8495 -16530
rect -8461 -16564 -8414 -16530
rect -8902 -16570 -8414 -16564
rect -9198 -16646 -9184 -16633
rect -12328 -16699 -12216 -16661
rect -12328 -16733 -12289 -16699
rect -12255 -16733 -12216 -16699
rect -12328 -16771 -12216 -16733
rect -12328 -16805 -12289 -16771
rect -12255 -16805 -12216 -16771
rect -12328 -16843 -12216 -16805
rect -12328 -16877 -12289 -16843
rect -12255 -16877 -12216 -16843
rect -12328 -16915 -12216 -16877
rect -12328 -16949 -12289 -16915
rect -12255 -16949 -12216 -16915
rect -12328 -16987 -12216 -16949
rect -12328 -17021 -12289 -16987
rect -12255 -17021 -12216 -16987
rect -12328 -17059 -12216 -17021
rect -12328 -17093 -12289 -17059
rect -12255 -17093 -12216 -17059
rect -12328 -17131 -12216 -17093
rect -12328 -17165 -12289 -17131
rect -12255 -17165 -12216 -17131
rect -12328 -17203 -12216 -17165
rect -9190 -16667 -9184 -16646
rect -9150 -16646 -9138 -16633
rect -8178 -16633 -8118 -16353
rect -7158 -16353 -7148 -16350
rect -7114 -16350 -7108 -16319
rect -6136 -15849 -6130 -15824
rect -6096 -15824 -6080 -15815
rect -5120 -15815 -5060 -15535
rect -4108 -15535 -4094 -15534
rect -4060 -15534 -4054 -15501
rect -3082 -15031 -3076 -15012
rect -3042 -15012 -3026 -14997
rect -2066 -14997 -2006 -14722
rect -1776 -14786 -1288 -14780
rect -1776 -14820 -1729 -14786
rect -1695 -14820 -1657 -14786
rect -1623 -14820 -1585 -14786
rect -1551 -14820 -1513 -14786
rect -1479 -14820 -1441 -14786
rect -1407 -14820 -1369 -14786
rect -1335 -14820 -1288 -14786
rect -1776 -14826 -1288 -14820
rect -1576 -14888 -1516 -14826
rect -1776 -14894 -1288 -14888
rect -1776 -14928 -1729 -14894
rect -1695 -14928 -1657 -14894
rect -1623 -14928 -1585 -14894
rect -1551 -14928 -1513 -14894
rect -1479 -14928 -1441 -14894
rect -1407 -14928 -1369 -14894
rect -1335 -14928 -1288 -14894
rect -1776 -14934 -1288 -14928
rect -2066 -15012 -2058 -14997
rect -3042 -15031 -3036 -15012
rect -3082 -15069 -3036 -15031
rect -3082 -15103 -3076 -15069
rect -3042 -15103 -3036 -15069
rect -3082 -15141 -3036 -15103
rect -3082 -15175 -3076 -15141
rect -3042 -15175 -3036 -15141
rect -3082 -15213 -3036 -15175
rect -3082 -15247 -3076 -15213
rect -3042 -15247 -3036 -15213
rect -3082 -15285 -3036 -15247
rect -3082 -15319 -3076 -15285
rect -3042 -15319 -3036 -15285
rect -3082 -15357 -3036 -15319
rect -3082 -15391 -3076 -15357
rect -3042 -15391 -3036 -15357
rect -3082 -15429 -3036 -15391
rect -3082 -15463 -3076 -15429
rect -3042 -15463 -3036 -15429
rect -3082 -15501 -3036 -15463
rect -3082 -15534 -3076 -15501
rect -4060 -15535 -4048 -15534
rect -4830 -15604 -4342 -15598
rect -4830 -15638 -4783 -15604
rect -4749 -15638 -4711 -15604
rect -4677 -15638 -4639 -15604
rect -4605 -15638 -4567 -15604
rect -4533 -15638 -4495 -15604
rect -4461 -15638 -4423 -15604
rect -4389 -15638 -4342 -15604
rect -4830 -15644 -4342 -15638
rect -4628 -15706 -4568 -15644
rect -4830 -15712 -4342 -15706
rect -4830 -15746 -4783 -15712
rect -4749 -15746 -4711 -15712
rect -4677 -15746 -4639 -15712
rect -4605 -15746 -4567 -15712
rect -4533 -15746 -4495 -15712
rect -4461 -15746 -4423 -15712
rect -4389 -15746 -4342 -15712
rect -4830 -15752 -4342 -15746
rect -5120 -15816 -5112 -15815
rect -6096 -15849 -6090 -15824
rect -6136 -15887 -6090 -15849
rect -6136 -15921 -6130 -15887
rect -6096 -15921 -6090 -15887
rect -6136 -15959 -6090 -15921
rect -6136 -15993 -6130 -15959
rect -6096 -15993 -6090 -15959
rect -6136 -16031 -6090 -15993
rect -6136 -16065 -6130 -16031
rect -6096 -16065 -6090 -16031
rect -6136 -16103 -6090 -16065
rect -6136 -16137 -6130 -16103
rect -6096 -16137 -6090 -16103
rect -6136 -16175 -6090 -16137
rect -6136 -16209 -6130 -16175
rect -6096 -16209 -6090 -16175
rect -6136 -16247 -6090 -16209
rect -6136 -16281 -6130 -16247
rect -6096 -16281 -6090 -16247
rect -6136 -16319 -6090 -16281
rect -7114 -16353 -7098 -16350
rect -7884 -16422 -7396 -16416
rect -7884 -16456 -7837 -16422
rect -7803 -16456 -7765 -16422
rect -7731 -16456 -7693 -16422
rect -7659 -16456 -7621 -16422
rect -7587 -16456 -7549 -16422
rect -7515 -16456 -7477 -16422
rect -7443 -16456 -7396 -16422
rect -7884 -16462 -7396 -16456
rect -7678 -16524 -7618 -16462
rect -7884 -16530 -7396 -16524
rect -7884 -16564 -7837 -16530
rect -7803 -16564 -7765 -16530
rect -7731 -16564 -7693 -16530
rect -7659 -16564 -7621 -16530
rect -7587 -16564 -7549 -16530
rect -7515 -16564 -7477 -16530
rect -7443 -16564 -7396 -16530
rect -7884 -16570 -7396 -16564
rect -8178 -16642 -8166 -16633
rect -9150 -16667 -9144 -16646
rect -9190 -16705 -9144 -16667
rect -9190 -16739 -9184 -16705
rect -9150 -16739 -9144 -16705
rect -9190 -16777 -9144 -16739
rect -9190 -16811 -9184 -16777
rect -9150 -16811 -9144 -16777
rect -9190 -16849 -9144 -16811
rect -9190 -16883 -9184 -16849
rect -9150 -16883 -9144 -16849
rect -9190 -16921 -9144 -16883
rect -9190 -16955 -9184 -16921
rect -9150 -16955 -9144 -16921
rect -9190 -16993 -9144 -16955
rect -9190 -17027 -9184 -16993
rect -9150 -17027 -9144 -16993
rect -9190 -17065 -9144 -17027
rect -9190 -17099 -9184 -17065
rect -9150 -17099 -9144 -17065
rect -9190 -17137 -9144 -17099
rect -9190 -17168 -9184 -17137
rect -12328 -17237 -12289 -17203
rect -12255 -17237 -12216 -17203
rect -12328 -17275 -12216 -17237
rect -12328 -17309 -12289 -17275
rect -12255 -17309 -12216 -17275
rect -12328 -17347 -12216 -17309
rect -12328 -17381 -12289 -17347
rect -12255 -17381 -12216 -17347
rect -12328 -17419 -12216 -17381
rect -12328 -17453 -12289 -17419
rect -12255 -17453 -12216 -17419
rect -12328 -17491 -12216 -17453
rect -9198 -17171 -9184 -17168
rect -9150 -17168 -9144 -17137
rect -8172 -16667 -8166 -16642
rect -8132 -16642 -8118 -16633
rect -7158 -16633 -7098 -16353
rect -6136 -16353 -6130 -16319
rect -6096 -16353 -6090 -16319
rect -5118 -15849 -5112 -15816
rect -5078 -15816 -5060 -15815
rect -4108 -15815 -4048 -15535
rect -3086 -15535 -3076 -15534
rect -3042 -15534 -3036 -15501
rect -2064 -15031 -2058 -15012
rect -2024 -15012 -2006 -14997
rect -1050 -14997 -990 -14718
rect -28 -14722 18 -14717
rect -758 -14786 -270 -14780
rect -758 -14820 -711 -14786
rect -677 -14820 -639 -14786
rect -605 -14820 -567 -14786
rect -533 -14820 -495 -14786
rect -461 -14820 -423 -14786
rect -389 -14820 -351 -14786
rect -317 -14820 -270 -14786
rect -758 -14826 -270 -14820
rect -556 -14888 -496 -14826
rect -758 -14894 -270 -14888
rect -758 -14928 -711 -14894
rect -677 -14928 -639 -14894
rect -605 -14928 -567 -14894
rect -533 -14928 -495 -14894
rect -461 -14928 -423 -14894
rect -389 -14928 -351 -14894
rect -317 -14928 -270 -14894
rect -758 -14934 -270 -14928
rect -1050 -15008 -1040 -14997
rect -2024 -15031 -2018 -15012
rect -2064 -15069 -2018 -15031
rect -2064 -15103 -2058 -15069
rect -2024 -15103 -2018 -15069
rect -2064 -15141 -2018 -15103
rect -2064 -15175 -2058 -15141
rect -2024 -15175 -2018 -15141
rect -2064 -15213 -2018 -15175
rect -2064 -15247 -2058 -15213
rect -2024 -15247 -2018 -15213
rect -2064 -15285 -2018 -15247
rect -2064 -15319 -2058 -15285
rect -2024 -15319 -2018 -15285
rect -2064 -15357 -2018 -15319
rect -2064 -15391 -2058 -15357
rect -2024 -15391 -2018 -15357
rect -2064 -15429 -2018 -15391
rect -2064 -15463 -2058 -15429
rect -2024 -15463 -2018 -15429
rect -2064 -15501 -2018 -15463
rect -2064 -15534 -2058 -15501
rect -3042 -15535 -3026 -15534
rect -3812 -15604 -3324 -15598
rect -3812 -15638 -3765 -15604
rect -3731 -15638 -3693 -15604
rect -3659 -15638 -3621 -15604
rect -3587 -15638 -3549 -15604
rect -3515 -15638 -3477 -15604
rect -3443 -15638 -3405 -15604
rect -3371 -15638 -3324 -15604
rect -3812 -15644 -3324 -15638
rect -3612 -15706 -3552 -15644
rect -3812 -15712 -3324 -15706
rect -3812 -15746 -3765 -15712
rect -3731 -15746 -3693 -15712
rect -3659 -15746 -3621 -15712
rect -3587 -15746 -3549 -15712
rect -3515 -15746 -3477 -15712
rect -3443 -15746 -3405 -15712
rect -3371 -15746 -3324 -15712
rect -3812 -15752 -3324 -15746
rect -5078 -15849 -5072 -15816
rect -4108 -15824 -4094 -15815
rect -5118 -15887 -5072 -15849
rect -5118 -15921 -5112 -15887
rect -5078 -15921 -5072 -15887
rect -5118 -15959 -5072 -15921
rect -5118 -15993 -5112 -15959
rect -5078 -15993 -5072 -15959
rect -5118 -16031 -5072 -15993
rect -5118 -16065 -5112 -16031
rect -5078 -16065 -5072 -16031
rect -5118 -16103 -5072 -16065
rect -5118 -16137 -5112 -16103
rect -5078 -16137 -5072 -16103
rect -5118 -16175 -5072 -16137
rect -5118 -16209 -5112 -16175
rect -5078 -16209 -5072 -16175
rect -5118 -16247 -5072 -16209
rect -5118 -16281 -5112 -16247
rect -5078 -16281 -5072 -16247
rect -5118 -16319 -5072 -16281
rect -5118 -16346 -5112 -16319
rect -6136 -16354 -6090 -16353
rect -5120 -16353 -5112 -16346
rect -5078 -16346 -5072 -16319
rect -4100 -15849 -4094 -15824
rect -4060 -15824 -4048 -15815
rect -3086 -15815 -3026 -15535
rect -2066 -15535 -2058 -15534
rect -2024 -15534 -2018 -15501
rect -1046 -15031 -1040 -15008
rect -1006 -15008 -990 -14997
rect -28 -14997 32 -14722
rect -1006 -15031 -1000 -15008
rect -1046 -15069 -1000 -15031
rect -1046 -15103 -1040 -15069
rect -1006 -15103 -1000 -15069
rect -1046 -15141 -1000 -15103
rect -1046 -15175 -1040 -15141
rect -1006 -15175 -1000 -15141
rect -1046 -15213 -1000 -15175
rect -1046 -15247 -1040 -15213
rect -1006 -15247 -1000 -15213
rect -1046 -15285 -1000 -15247
rect -1046 -15319 -1040 -15285
rect -1006 -15319 -1000 -15285
rect -1046 -15357 -1000 -15319
rect -1046 -15391 -1040 -15357
rect -1006 -15391 -1000 -15357
rect -1046 -15429 -1000 -15391
rect -1046 -15463 -1040 -15429
rect -1006 -15463 -1000 -15429
rect -1046 -15501 -1000 -15463
rect -1046 -15530 -1040 -15501
rect -2024 -15535 -2006 -15534
rect -2794 -15604 -2306 -15598
rect -2794 -15638 -2747 -15604
rect -2713 -15638 -2675 -15604
rect -2641 -15638 -2603 -15604
rect -2569 -15638 -2531 -15604
rect -2497 -15638 -2459 -15604
rect -2425 -15638 -2387 -15604
rect -2353 -15638 -2306 -15604
rect -2794 -15644 -2306 -15638
rect -2590 -15706 -2530 -15644
rect -2794 -15712 -2306 -15706
rect -2794 -15746 -2747 -15712
rect -2713 -15746 -2675 -15712
rect -2641 -15746 -2603 -15712
rect -2569 -15746 -2531 -15712
rect -2497 -15746 -2459 -15712
rect -2425 -15746 -2387 -15712
rect -2353 -15746 -2306 -15712
rect -2794 -15752 -2306 -15746
rect -3086 -15824 -3076 -15815
rect -4060 -15849 -4054 -15824
rect -4100 -15887 -4054 -15849
rect -4100 -15921 -4094 -15887
rect -4060 -15921 -4054 -15887
rect -4100 -15959 -4054 -15921
rect -4100 -15993 -4094 -15959
rect -4060 -15993 -4054 -15959
rect -4100 -16031 -4054 -15993
rect -4100 -16065 -4094 -16031
rect -4060 -16065 -4054 -16031
rect -4100 -16103 -4054 -16065
rect -4100 -16137 -4094 -16103
rect -4060 -16137 -4054 -16103
rect -4100 -16175 -4054 -16137
rect -4100 -16209 -4094 -16175
rect -4060 -16209 -4054 -16175
rect -4100 -16247 -4054 -16209
rect -4100 -16281 -4094 -16247
rect -4060 -16281 -4054 -16247
rect -4100 -16319 -4054 -16281
rect -5078 -16353 -5060 -16346
rect -6866 -16422 -6378 -16416
rect -6866 -16456 -6819 -16422
rect -6785 -16456 -6747 -16422
rect -6713 -16456 -6675 -16422
rect -6641 -16456 -6603 -16422
rect -6569 -16456 -6531 -16422
rect -6497 -16456 -6459 -16422
rect -6425 -16456 -6378 -16422
rect -6866 -16462 -6378 -16456
rect -6658 -16524 -6598 -16462
rect -6866 -16530 -6378 -16524
rect -6866 -16564 -6819 -16530
rect -6785 -16564 -6747 -16530
rect -6713 -16564 -6675 -16530
rect -6641 -16564 -6603 -16530
rect -6569 -16564 -6531 -16530
rect -6497 -16564 -6459 -16530
rect -6425 -16564 -6378 -16530
rect -6866 -16570 -6378 -16564
rect -7158 -16640 -7148 -16633
rect -8132 -16667 -8126 -16642
rect -8172 -16705 -8126 -16667
rect -8172 -16739 -8166 -16705
rect -8132 -16739 -8126 -16705
rect -8172 -16777 -8126 -16739
rect -8172 -16811 -8166 -16777
rect -8132 -16811 -8126 -16777
rect -8172 -16849 -8126 -16811
rect -8172 -16883 -8166 -16849
rect -8132 -16883 -8126 -16849
rect -8172 -16921 -8126 -16883
rect -8172 -16955 -8166 -16921
rect -8132 -16955 -8126 -16921
rect -8172 -16993 -8126 -16955
rect -8172 -17027 -8166 -16993
rect -8132 -17027 -8126 -16993
rect -8172 -17065 -8126 -17027
rect -8172 -17099 -8166 -17065
rect -8132 -17099 -8126 -17065
rect -8172 -17137 -8126 -17099
rect -8172 -17164 -8166 -17137
rect -9150 -17171 -9138 -17168
rect -9198 -17451 -9138 -17171
rect -8178 -17171 -8166 -17164
rect -8132 -17164 -8126 -17137
rect -7154 -16667 -7148 -16640
rect -7114 -16640 -7098 -16633
rect -6140 -16633 -6080 -16354
rect -5848 -16422 -5360 -16416
rect -5848 -16456 -5801 -16422
rect -5767 -16456 -5729 -16422
rect -5695 -16456 -5657 -16422
rect -5623 -16456 -5585 -16422
rect -5551 -16456 -5513 -16422
rect -5479 -16456 -5441 -16422
rect -5407 -16456 -5360 -16422
rect -5848 -16462 -5360 -16456
rect -5656 -16524 -5596 -16462
rect -5848 -16530 -5360 -16524
rect -5848 -16564 -5801 -16530
rect -5767 -16564 -5729 -16530
rect -5695 -16564 -5657 -16530
rect -5623 -16564 -5585 -16530
rect -5551 -16564 -5513 -16530
rect -5479 -16564 -5441 -16530
rect -5407 -16564 -5360 -16530
rect -5848 -16570 -5360 -16564
rect -7114 -16667 -7108 -16640
rect -6140 -16644 -6130 -16633
rect -7154 -16705 -7108 -16667
rect -7154 -16739 -7148 -16705
rect -7114 -16739 -7108 -16705
rect -7154 -16777 -7108 -16739
rect -7154 -16811 -7148 -16777
rect -7114 -16811 -7108 -16777
rect -7154 -16849 -7108 -16811
rect -7154 -16883 -7148 -16849
rect -7114 -16883 -7108 -16849
rect -7154 -16921 -7108 -16883
rect -7154 -16955 -7148 -16921
rect -7114 -16955 -7108 -16921
rect -7154 -16993 -7108 -16955
rect -7154 -17027 -7148 -16993
rect -7114 -17027 -7108 -16993
rect -7154 -17065 -7108 -17027
rect -7154 -17099 -7148 -17065
rect -7114 -17099 -7108 -17065
rect -7154 -17137 -7108 -17099
rect -7154 -17162 -7148 -17137
rect -8132 -17171 -8118 -17164
rect -8902 -17240 -8414 -17234
rect -8902 -17274 -8855 -17240
rect -8821 -17274 -8783 -17240
rect -8749 -17274 -8711 -17240
rect -8677 -17274 -8639 -17240
rect -8605 -17274 -8567 -17240
rect -8533 -17274 -8495 -17240
rect -8461 -17274 -8414 -17240
rect -8902 -17280 -8414 -17274
rect -8690 -17342 -8630 -17280
rect -8902 -17348 -8414 -17342
rect -8902 -17382 -8855 -17348
rect -8821 -17382 -8783 -17348
rect -8749 -17382 -8711 -17348
rect -8677 -17382 -8639 -17348
rect -8605 -17382 -8567 -17348
rect -8533 -17382 -8495 -17348
rect -8461 -17382 -8414 -17348
rect -8902 -17388 -8414 -17382
rect -9198 -17458 -9184 -17451
rect -12328 -17525 -12289 -17491
rect -12255 -17525 -12216 -17491
rect -12328 -17563 -12216 -17525
rect -12328 -17597 -12289 -17563
rect -12255 -17597 -12216 -17563
rect -12328 -17635 -12216 -17597
rect -12328 -17669 -12289 -17635
rect -12255 -17669 -12216 -17635
rect -12328 -17707 -12216 -17669
rect -12328 -17741 -12289 -17707
rect -12255 -17741 -12216 -17707
rect -12328 -17779 -12216 -17741
rect -12328 -17813 -12289 -17779
rect -12255 -17813 -12216 -17779
rect -12328 -17851 -12216 -17813
rect -12328 -17885 -12289 -17851
rect -12255 -17885 -12216 -17851
rect -12328 -17923 -12216 -17885
rect -12328 -17957 -12289 -17923
rect -12255 -17957 -12216 -17923
rect -12328 -17995 -12216 -17957
rect -9190 -17485 -9184 -17458
rect -9150 -17458 -9138 -17451
rect -8178 -17451 -8118 -17171
rect -7158 -17171 -7148 -17162
rect -7114 -17162 -7108 -17137
rect -6136 -16667 -6130 -16644
rect -6096 -16644 -6080 -16633
rect -5120 -16633 -5060 -16353
rect -4100 -16353 -4094 -16319
rect -4060 -16353 -4054 -16319
rect -4100 -16354 -4054 -16353
rect -3082 -15849 -3076 -15824
rect -3042 -15824 -3026 -15815
rect -2066 -15815 -2006 -15535
rect -1050 -15535 -1040 -15530
rect -1006 -15530 -1000 -15501
rect -28 -15031 -22 -14997
rect 12 -15012 32 -14997
rect 12 -15031 18 -15012
rect -28 -15069 18 -15031
rect -28 -15103 -22 -15069
rect 12 -15103 18 -15069
rect -28 -15141 18 -15103
rect -28 -15175 -22 -15141
rect 12 -15175 18 -15141
rect -28 -15213 18 -15175
rect -28 -15247 -22 -15213
rect 12 -15247 18 -15213
rect -28 -15285 18 -15247
rect -28 -15319 -22 -15285
rect 12 -15319 18 -15285
rect -28 -15357 18 -15319
rect -28 -15391 -22 -15357
rect 12 -15391 18 -15357
rect -28 -15429 18 -15391
rect -28 -15463 -22 -15429
rect 12 -15463 18 -15429
rect -28 -15501 18 -15463
rect -1006 -15535 -990 -15530
rect -1776 -15604 -1288 -15598
rect -1776 -15638 -1729 -15604
rect -1695 -15638 -1657 -15604
rect -1623 -15638 -1585 -15604
rect -1551 -15638 -1513 -15604
rect -1479 -15638 -1441 -15604
rect -1407 -15638 -1369 -15604
rect -1335 -15638 -1288 -15604
rect -1776 -15644 -1288 -15638
rect -1578 -15706 -1518 -15644
rect -1776 -15712 -1288 -15706
rect -1776 -15746 -1729 -15712
rect -1695 -15746 -1657 -15712
rect -1623 -15746 -1585 -15712
rect -1551 -15746 -1513 -15712
rect -1479 -15746 -1441 -15712
rect -1407 -15746 -1369 -15712
rect -1335 -15746 -1288 -15712
rect -1776 -15752 -1288 -15746
rect -2066 -15824 -2058 -15815
rect -3042 -15849 -3036 -15824
rect -3082 -15887 -3036 -15849
rect -3082 -15921 -3076 -15887
rect -3042 -15921 -3036 -15887
rect -3082 -15959 -3036 -15921
rect -3082 -15993 -3076 -15959
rect -3042 -15993 -3036 -15959
rect -3082 -16031 -3036 -15993
rect -3082 -16065 -3076 -16031
rect -3042 -16065 -3036 -16031
rect -3082 -16103 -3036 -16065
rect -3082 -16137 -3076 -16103
rect -3042 -16137 -3036 -16103
rect -3082 -16175 -3036 -16137
rect -3082 -16209 -3076 -16175
rect -3042 -16209 -3036 -16175
rect -3082 -16247 -3036 -16209
rect -3082 -16281 -3076 -16247
rect -3042 -16281 -3036 -16247
rect -3082 -16319 -3036 -16281
rect -3082 -16353 -3076 -16319
rect -3042 -16353 -3036 -16319
rect -3082 -16354 -3036 -16353
rect -2064 -15849 -2058 -15824
rect -2024 -15824 -2006 -15815
rect -1050 -15815 -990 -15535
rect -28 -15535 -22 -15501
rect 12 -15534 18 -15501
rect 12 -15535 32 -15534
rect -758 -15604 -270 -15598
rect -758 -15638 -711 -15604
rect -677 -15638 -639 -15604
rect -605 -15638 -567 -15604
rect -533 -15638 -495 -15604
rect -461 -15638 -423 -15604
rect -389 -15638 -351 -15604
rect -317 -15638 -270 -15604
rect -758 -15644 -270 -15638
rect -558 -15706 -498 -15644
rect -758 -15712 -270 -15706
rect -758 -15746 -711 -15712
rect -677 -15746 -639 -15712
rect -605 -15746 -567 -15712
rect -533 -15746 -495 -15712
rect -461 -15746 -423 -15712
rect -389 -15746 -351 -15712
rect -317 -15746 -270 -15712
rect -758 -15752 -270 -15746
rect -1050 -15820 -1040 -15815
rect -2024 -15849 -2018 -15824
rect -2064 -15887 -2018 -15849
rect -2064 -15921 -2058 -15887
rect -2024 -15921 -2018 -15887
rect -2064 -15959 -2018 -15921
rect -2064 -15993 -2058 -15959
rect -2024 -15993 -2018 -15959
rect -2064 -16031 -2018 -15993
rect -2064 -16065 -2058 -16031
rect -2024 -16065 -2018 -16031
rect -2064 -16103 -2018 -16065
rect -2064 -16137 -2058 -16103
rect -2024 -16137 -2018 -16103
rect -2064 -16175 -2018 -16137
rect -2064 -16209 -2058 -16175
rect -2024 -16209 -2018 -16175
rect -2064 -16247 -2018 -16209
rect -2064 -16281 -2058 -16247
rect -2024 -16281 -2018 -16247
rect -2064 -16319 -2018 -16281
rect -2064 -16353 -2058 -16319
rect -2024 -16353 -2018 -16319
rect -1046 -15849 -1040 -15820
rect -1006 -15820 -990 -15815
rect -28 -15815 32 -15535
rect -1006 -15849 -1000 -15820
rect -1046 -15887 -1000 -15849
rect -1046 -15921 -1040 -15887
rect -1006 -15921 -1000 -15887
rect -1046 -15959 -1000 -15921
rect -1046 -15993 -1040 -15959
rect -1006 -15993 -1000 -15959
rect -1046 -16031 -1000 -15993
rect -1046 -16065 -1040 -16031
rect -1006 -16065 -1000 -16031
rect -1046 -16103 -1000 -16065
rect -1046 -16137 -1040 -16103
rect -1006 -16137 -1000 -16103
rect -1046 -16175 -1000 -16137
rect -1046 -16209 -1040 -16175
rect -1006 -16209 -1000 -16175
rect -1046 -16247 -1000 -16209
rect -1046 -16281 -1040 -16247
rect -1006 -16281 -1000 -16247
rect -1046 -16319 -1000 -16281
rect -1046 -16350 -1040 -16319
rect -2064 -16354 -2018 -16353
rect -1050 -16353 -1040 -16350
rect -1006 -16350 -1000 -16319
rect -28 -15849 -22 -15815
rect 12 -15824 32 -15815
rect 12 -15849 18 -15824
rect -28 -15887 18 -15849
rect -28 -15921 -22 -15887
rect 12 -15921 18 -15887
rect -28 -15959 18 -15921
rect -28 -15993 -22 -15959
rect 12 -15993 18 -15959
rect -28 -16031 18 -15993
rect -28 -16065 -22 -16031
rect 12 -16065 18 -16031
rect -28 -16103 18 -16065
rect -28 -16137 -22 -16103
rect 12 -16137 18 -16103
rect -28 -16175 18 -16137
rect -28 -16209 -22 -16175
rect 12 -16209 18 -16175
rect -28 -16247 18 -16209
rect -28 -16281 -22 -16247
rect 12 -16281 18 -16247
rect -28 -16319 18 -16281
rect -1006 -16353 -990 -16350
rect -4830 -16422 -4342 -16416
rect -4830 -16456 -4783 -16422
rect -4749 -16456 -4711 -16422
rect -4677 -16456 -4639 -16422
rect -4605 -16456 -4567 -16422
rect -4533 -16456 -4495 -16422
rect -4461 -16456 -4423 -16422
rect -4389 -16456 -4342 -16422
rect -4830 -16462 -4342 -16456
rect -4626 -16524 -4566 -16462
rect -4830 -16530 -4342 -16524
rect -4830 -16564 -4783 -16530
rect -4749 -16564 -4711 -16530
rect -4677 -16564 -4639 -16530
rect -4605 -16564 -4567 -16530
rect -4533 -16564 -4495 -16530
rect -4461 -16564 -4423 -16530
rect -4389 -16564 -4342 -16530
rect -4830 -16570 -4342 -16564
rect -5120 -16636 -5112 -16633
rect -6096 -16667 -6090 -16644
rect -6136 -16705 -6090 -16667
rect -6136 -16739 -6130 -16705
rect -6096 -16739 -6090 -16705
rect -6136 -16777 -6090 -16739
rect -6136 -16811 -6130 -16777
rect -6096 -16811 -6090 -16777
rect -6136 -16849 -6090 -16811
rect -6136 -16883 -6130 -16849
rect -6096 -16883 -6090 -16849
rect -6136 -16921 -6090 -16883
rect -6136 -16955 -6130 -16921
rect -6096 -16955 -6090 -16921
rect -6136 -16993 -6090 -16955
rect -6136 -17027 -6130 -16993
rect -6096 -17027 -6090 -16993
rect -6136 -17065 -6090 -17027
rect -6136 -17099 -6130 -17065
rect -6096 -17099 -6090 -17065
rect -6136 -17137 -6090 -17099
rect -7114 -17171 -7098 -17162
rect -6136 -17166 -6130 -17137
rect -7884 -17240 -7396 -17234
rect -7884 -17274 -7837 -17240
rect -7803 -17274 -7765 -17240
rect -7731 -17274 -7693 -17240
rect -7659 -17274 -7621 -17240
rect -7587 -17274 -7549 -17240
rect -7515 -17274 -7477 -17240
rect -7443 -17274 -7396 -17240
rect -7884 -17280 -7396 -17274
rect -7676 -17342 -7616 -17280
rect -7884 -17348 -7396 -17342
rect -7884 -17382 -7837 -17348
rect -7803 -17382 -7765 -17348
rect -7731 -17382 -7693 -17348
rect -7659 -17382 -7621 -17348
rect -7587 -17382 -7549 -17348
rect -7515 -17382 -7477 -17348
rect -7443 -17382 -7396 -17348
rect -7884 -17388 -7396 -17382
rect -8178 -17454 -8166 -17451
rect -9150 -17485 -9144 -17458
rect -9190 -17523 -9144 -17485
rect -9190 -17557 -9184 -17523
rect -9150 -17557 -9144 -17523
rect -9190 -17595 -9144 -17557
rect -9190 -17629 -9184 -17595
rect -9150 -17629 -9144 -17595
rect -9190 -17667 -9144 -17629
rect -9190 -17701 -9184 -17667
rect -9150 -17701 -9144 -17667
rect -9190 -17739 -9144 -17701
rect -9190 -17773 -9184 -17739
rect -9150 -17773 -9144 -17739
rect -9190 -17811 -9144 -17773
rect -9190 -17845 -9184 -17811
rect -9150 -17845 -9144 -17811
rect -9190 -17883 -9144 -17845
rect -9190 -17917 -9184 -17883
rect -9150 -17917 -9144 -17883
rect -9190 -17955 -9144 -17917
rect -9190 -17986 -9184 -17955
rect -12328 -18029 -12289 -17995
rect -12255 -18029 -12216 -17995
rect -12328 -18067 -12216 -18029
rect -12328 -18101 -12289 -18067
rect -12255 -18101 -12216 -18067
rect -12328 -18139 -12216 -18101
rect -12328 -18173 -12289 -18139
rect -12255 -18173 -12216 -18139
rect -12328 -18211 -12216 -18173
rect -12328 -18245 -12289 -18211
rect -12255 -18245 -12216 -18211
rect -12328 -18283 -12216 -18245
rect -9198 -17989 -9184 -17986
rect -9150 -17986 -9144 -17955
rect -8172 -17485 -8166 -17454
rect -8132 -17454 -8118 -17451
rect -7158 -17451 -7098 -17171
rect -6140 -17171 -6130 -17166
rect -6096 -17166 -6090 -17137
rect -5118 -16667 -5112 -16636
rect -5078 -16636 -5060 -16633
rect -4108 -16633 -4048 -16354
rect -3812 -16422 -3324 -16416
rect -3812 -16456 -3765 -16422
rect -3731 -16456 -3693 -16422
rect -3659 -16456 -3621 -16422
rect -3587 -16456 -3549 -16422
rect -3515 -16456 -3477 -16422
rect -3443 -16456 -3405 -16422
rect -3371 -16456 -3324 -16422
rect -3812 -16462 -3324 -16456
rect -3610 -16524 -3550 -16462
rect -3812 -16530 -3324 -16524
rect -3812 -16564 -3765 -16530
rect -3731 -16564 -3693 -16530
rect -3659 -16564 -3621 -16530
rect -3587 -16564 -3549 -16530
rect -3515 -16564 -3477 -16530
rect -3443 -16564 -3405 -16530
rect -3371 -16564 -3324 -16530
rect -3812 -16570 -3324 -16564
rect -5078 -16667 -5072 -16636
rect -4108 -16644 -4094 -16633
rect -5118 -16705 -5072 -16667
rect -5118 -16739 -5112 -16705
rect -5078 -16739 -5072 -16705
rect -5118 -16777 -5072 -16739
rect -5118 -16811 -5112 -16777
rect -5078 -16811 -5072 -16777
rect -5118 -16849 -5072 -16811
rect -5118 -16883 -5112 -16849
rect -5078 -16883 -5072 -16849
rect -5118 -16921 -5072 -16883
rect -5118 -16955 -5112 -16921
rect -5078 -16955 -5072 -16921
rect -5118 -16993 -5072 -16955
rect -5118 -17027 -5112 -16993
rect -5078 -17027 -5072 -16993
rect -5118 -17065 -5072 -17027
rect -5118 -17099 -5112 -17065
rect -5078 -17099 -5072 -17065
rect -5118 -17137 -5072 -17099
rect -5118 -17158 -5112 -17137
rect -6096 -17171 -6080 -17166
rect -6866 -17240 -6378 -17234
rect -6866 -17274 -6819 -17240
rect -6785 -17274 -6747 -17240
rect -6713 -17274 -6675 -17240
rect -6641 -17274 -6603 -17240
rect -6569 -17274 -6531 -17240
rect -6497 -17274 -6459 -17240
rect -6425 -17274 -6378 -17240
rect -6866 -17280 -6378 -17274
rect -6656 -17342 -6596 -17280
rect -6866 -17348 -6378 -17342
rect -6866 -17382 -6819 -17348
rect -6785 -17382 -6747 -17348
rect -6713 -17382 -6675 -17348
rect -6641 -17382 -6603 -17348
rect -6569 -17382 -6531 -17348
rect -6497 -17382 -6459 -17348
rect -6425 -17382 -6378 -17348
rect -6866 -17388 -6378 -17382
rect -7158 -17452 -7148 -17451
rect -8132 -17485 -8126 -17454
rect -8172 -17523 -8126 -17485
rect -8172 -17557 -8166 -17523
rect -8132 -17557 -8126 -17523
rect -8172 -17595 -8126 -17557
rect -8172 -17629 -8166 -17595
rect -8132 -17629 -8126 -17595
rect -8172 -17667 -8126 -17629
rect -8172 -17701 -8166 -17667
rect -8132 -17701 -8126 -17667
rect -8172 -17739 -8126 -17701
rect -8172 -17773 -8166 -17739
rect -8132 -17773 -8126 -17739
rect -8172 -17811 -8126 -17773
rect -8172 -17845 -8166 -17811
rect -8132 -17845 -8126 -17811
rect -8172 -17883 -8126 -17845
rect -8172 -17917 -8166 -17883
rect -8132 -17917 -8126 -17883
rect -8172 -17955 -8126 -17917
rect -8172 -17982 -8166 -17955
rect -9150 -17989 -9138 -17986
rect -9198 -18269 -9138 -17989
rect -8178 -17989 -8166 -17982
rect -8132 -17982 -8126 -17955
rect -7154 -17485 -7148 -17452
rect -7114 -17452 -7098 -17451
rect -6140 -17451 -6080 -17171
rect -5120 -17171 -5112 -17158
rect -5078 -17158 -5072 -17137
rect -4100 -16667 -4094 -16644
rect -4060 -16644 -4048 -16633
rect -3086 -16633 -3026 -16354
rect -2794 -16422 -2306 -16416
rect -2794 -16456 -2747 -16422
rect -2713 -16456 -2675 -16422
rect -2641 -16456 -2603 -16422
rect -2569 -16456 -2531 -16422
rect -2497 -16456 -2459 -16422
rect -2425 -16456 -2387 -16422
rect -2353 -16456 -2306 -16422
rect -2794 -16462 -2306 -16456
rect -2588 -16524 -2528 -16462
rect -2794 -16530 -2306 -16524
rect -2794 -16564 -2747 -16530
rect -2713 -16564 -2675 -16530
rect -2641 -16564 -2603 -16530
rect -2569 -16564 -2531 -16530
rect -2497 -16564 -2459 -16530
rect -2425 -16564 -2387 -16530
rect -2353 -16564 -2306 -16530
rect -2794 -16570 -2306 -16564
rect -3086 -16644 -3076 -16633
rect -4060 -16667 -4054 -16644
rect -4100 -16705 -4054 -16667
rect -4100 -16739 -4094 -16705
rect -4060 -16739 -4054 -16705
rect -4100 -16777 -4054 -16739
rect -4100 -16811 -4094 -16777
rect -4060 -16811 -4054 -16777
rect -4100 -16849 -4054 -16811
rect -4100 -16883 -4094 -16849
rect -4060 -16883 -4054 -16849
rect -4100 -16921 -4054 -16883
rect -4100 -16955 -4094 -16921
rect -4060 -16955 -4054 -16921
rect -4100 -16993 -4054 -16955
rect -4100 -17027 -4094 -16993
rect -4060 -17027 -4054 -16993
rect -4100 -17065 -4054 -17027
rect -4100 -17099 -4094 -17065
rect -4060 -17099 -4054 -17065
rect -4100 -17137 -4054 -17099
rect -5078 -17171 -5060 -17158
rect -4100 -17166 -4094 -17137
rect -5848 -17240 -5360 -17234
rect -5848 -17274 -5801 -17240
rect -5767 -17274 -5729 -17240
rect -5695 -17274 -5657 -17240
rect -5623 -17274 -5585 -17240
rect -5551 -17274 -5513 -17240
rect -5479 -17274 -5441 -17240
rect -5407 -17274 -5360 -17240
rect -5848 -17280 -5360 -17274
rect -5654 -17342 -5594 -17280
rect -5848 -17348 -5360 -17342
rect -5848 -17382 -5801 -17348
rect -5767 -17382 -5729 -17348
rect -5695 -17382 -5657 -17348
rect -5623 -17382 -5585 -17348
rect -5551 -17382 -5513 -17348
rect -5479 -17382 -5441 -17348
rect -5407 -17382 -5360 -17348
rect -5848 -17388 -5360 -17382
rect -5120 -17448 -5060 -17171
rect -4108 -17171 -4094 -17166
rect -4060 -17166 -4054 -17137
rect -3082 -16667 -3076 -16644
rect -3042 -16644 -3026 -16633
rect -2066 -16633 -2006 -16354
rect -1776 -16422 -1288 -16416
rect -1776 -16456 -1729 -16422
rect -1695 -16456 -1657 -16422
rect -1623 -16456 -1585 -16422
rect -1551 -16456 -1513 -16422
rect -1479 -16456 -1441 -16422
rect -1407 -16456 -1369 -16422
rect -1335 -16456 -1288 -16422
rect -1776 -16462 -1288 -16456
rect -1576 -16524 -1516 -16462
rect -1776 -16530 -1288 -16524
rect -1776 -16564 -1729 -16530
rect -1695 -16564 -1657 -16530
rect -1623 -16564 -1585 -16530
rect -1551 -16564 -1513 -16530
rect -1479 -16564 -1441 -16530
rect -1407 -16564 -1369 -16530
rect -1335 -16564 -1288 -16530
rect -1776 -16570 -1288 -16564
rect -2066 -16644 -2058 -16633
rect -3042 -16667 -3036 -16644
rect -3082 -16705 -3036 -16667
rect -3082 -16739 -3076 -16705
rect -3042 -16739 -3036 -16705
rect -3082 -16777 -3036 -16739
rect -3082 -16811 -3076 -16777
rect -3042 -16811 -3036 -16777
rect -3082 -16849 -3036 -16811
rect -3082 -16883 -3076 -16849
rect -3042 -16883 -3036 -16849
rect -3082 -16921 -3036 -16883
rect -3082 -16955 -3076 -16921
rect -3042 -16955 -3036 -16921
rect -3082 -16993 -3036 -16955
rect -3082 -17027 -3076 -16993
rect -3042 -17027 -3036 -16993
rect -3082 -17065 -3036 -17027
rect -3082 -17099 -3076 -17065
rect -3042 -17099 -3036 -17065
rect -3082 -17137 -3036 -17099
rect -3082 -17166 -3076 -17137
rect -4060 -17171 -4048 -17166
rect -4830 -17240 -4342 -17234
rect -4830 -17274 -4783 -17240
rect -4749 -17274 -4711 -17240
rect -4677 -17274 -4639 -17240
rect -4605 -17274 -4567 -17240
rect -4533 -17274 -4495 -17240
rect -4461 -17274 -4423 -17240
rect -4389 -17274 -4342 -17240
rect -4830 -17280 -4342 -17274
rect -4624 -17342 -4564 -17280
rect -4830 -17348 -4342 -17342
rect -4830 -17382 -4783 -17348
rect -4749 -17382 -4711 -17348
rect -4677 -17382 -4639 -17348
rect -4605 -17382 -4567 -17348
rect -4533 -17382 -4495 -17348
rect -4461 -17382 -4423 -17348
rect -4389 -17382 -4342 -17348
rect -4830 -17388 -4342 -17382
rect -7114 -17485 -7108 -17452
rect -6140 -17456 -6130 -17451
rect -7154 -17523 -7108 -17485
rect -7154 -17557 -7148 -17523
rect -7114 -17557 -7108 -17523
rect -7154 -17595 -7108 -17557
rect -7154 -17629 -7148 -17595
rect -7114 -17629 -7108 -17595
rect -7154 -17667 -7108 -17629
rect -7154 -17701 -7148 -17667
rect -7114 -17701 -7108 -17667
rect -7154 -17739 -7108 -17701
rect -7154 -17773 -7148 -17739
rect -7114 -17773 -7108 -17739
rect -7154 -17811 -7108 -17773
rect -7154 -17845 -7148 -17811
rect -7114 -17845 -7108 -17811
rect -7154 -17883 -7108 -17845
rect -7154 -17917 -7148 -17883
rect -7114 -17917 -7108 -17883
rect -7154 -17955 -7108 -17917
rect -7154 -17980 -7148 -17955
rect -8132 -17989 -8118 -17982
rect -8902 -18058 -8414 -18052
rect -8902 -18092 -8855 -18058
rect -8821 -18092 -8783 -18058
rect -8749 -18092 -8711 -18058
rect -8677 -18092 -8639 -18058
rect -8605 -18092 -8567 -18058
rect -8533 -18092 -8495 -18058
rect -8461 -18092 -8414 -18058
rect -8902 -18098 -8414 -18092
rect -8688 -18160 -8628 -18098
rect -8902 -18166 -8414 -18160
rect -8902 -18200 -8855 -18166
rect -8821 -18200 -8783 -18166
rect -8749 -18200 -8711 -18166
rect -8677 -18200 -8639 -18166
rect -8605 -18200 -8567 -18166
rect -8533 -18200 -8495 -18166
rect -8461 -18200 -8414 -18166
rect -8902 -18206 -8414 -18200
rect -9198 -18276 -9184 -18269
rect -12328 -18317 -12289 -18283
rect -12255 -18317 -12216 -18283
rect -12328 -18355 -12216 -18317
rect -12328 -18389 -12289 -18355
rect -12255 -18389 -12216 -18355
rect -12328 -18427 -12216 -18389
rect -12328 -18461 -12289 -18427
rect -12255 -18461 -12216 -18427
rect -12328 -18499 -12216 -18461
rect -12328 -18533 -12289 -18499
rect -12255 -18533 -12216 -18499
rect -12328 -18571 -12216 -18533
rect -12328 -18605 -12289 -18571
rect -12255 -18605 -12216 -18571
rect -12328 -18643 -12216 -18605
rect -12328 -18677 -12289 -18643
rect -12255 -18677 -12216 -18643
rect -12328 -18715 -12216 -18677
rect -12328 -18749 -12289 -18715
rect -12255 -18749 -12216 -18715
rect -12328 -18787 -12216 -18749
rect -12328 -18821 -12289 -18787
rect -12255 -18821 -12216 -18787
rect -12328 -18859 -12216 -18821
rect -9190 -18303 -9184 -18276
rect -9150 -18276 -9138 -18269
rect -8178 -18269 -8118 -17989
rect -7158 -17989 -7148 -17980
rect -7114 -17980 -7108 -17955
rect -6136 -17485 -6130 -17456
rect -6096 -17456 -6080 -17451
rect -5118 -17451 -5072 -17448
rect -6096 -17485 -6090 -17456
rect -6136 -17523 -6090 -17485
rect -6136 -17557 -6130 -17523
rect -6096 -17557 -6090 -17523
rect -6136 -17595 -6090 -17557
rect -6136 -17629 -6130 -17595
rect -6096 -17629 -6090 -17595
rect -6136 -17667 -6090 -17629
rect -6136 -17701 -6130 -17667
rect -6096 -17701 -6090 -17667
rect -6136 -17739 -6090 -17701
rect -6136 -17773 -6130 -17739
rect -6096 -17773 -6090 -17739
rect -6136 -17811 -6090 -17773
rect -6136 -17845 -6130 -17811
rect -6096 -17845 -6090 -17811
rect -6136 -17883 -6090 -17845
rect -6136 -17917 -6130 -17883
rect -6096 -17917 -6090 -17883
rect -6136 -17955 -6090 -17917
rect -7114 -17989 -7098 -17980
rect -6136 -17984 -6130 -17955
rect -7884 -18058 -7396 -18052
rect -7884 -18092 -7837 -18058
rect -7803 -18092 -7765 -18058
rect -7731 -18092 -7693 -18058
rect -7659 -18092 -7621 -18058
rect -7587 -18092 -7549 -18058
rect -7515 -18092 -7477 -18058
rect -7443 -18092 -7396 -18058
rect -7884 -18098 -7396 -18092
rect -7674 -18160 -7614 -18098
rect -7884 -18166 -7396 -18160
rect -7884 -18200 -7837 -18166
rect -7803 -18200 -7765 -18166
rect -7731 -18200 -7693 -18166
rect -7659 -18200 -7621 -18166
rect -7587 -18200 -7549 -18166
rect -7515 -18200 -7477 -18166
rect -7443 -18200 -7396 -18166
rect -7884 -18206 -7396 -18200
rect -8178 -18272 -8166 -18269
rect -9150 -18303 -9144 -18276
rect -9190 -18341 -9144 -18303
rect -9190 -18375 -9184 -18341
rect -9150 -18375 -9144 -18341
rect -9190 -18413 -9144 -18375
rect -9190 -18447 -9184 -18413
rect -9150 -18447 -9144 -18413
rect -9190 -18485 -9144 -18447
rect -9190 -18519 -9184 -18485
rect -9150 -18519 -9144 -18485
rect -9190 -18557 -9144 -18519
rect -9190 -18591 -9184 -18557
rect -9150 -18591 -9144 -18557
rect -9190 -18629 -9144 -18591
rect -9190 -18663 -9184 -18629
rect -9150 -18663 -9144 -18629
rect -9190 -18701 -9144 -18663
rect -9190 -18735 -9184 -18701
rect -9150 -18735 -9144 -18701
rect -9190 -18773 -9144 -18735
rect -9190 -18807 -9184 -18773
rect -9150 -18807 -9144 -18773
rect -9190 -18838 -9144 -18807
rect -8172 -18303 -8166 -18272
rect -8132 -18272 -8118 -18269
rect -7158 -18269 -7098 -17989
rect -6140 -17989 -6130 -17984
rect -6096 -17984 -6090 -17955
rect -5118 -17485 -5112 -17451
rect -5078 -17485 -5072 -17451
rect -4108 -17451 -4048 -17171
rect -3086 -17171 -3076 -17166
rect -3042 -17166 -3036 -17137
rect -2064 -16667 -2058 -16644
rect -2024 -16644 -2006 -16633
rect -1050 -16633 -990 -16353
rect -28 -16353 -22 -16319
rect 12 -16353 18 -16319
rect -28 -16354 18 -16353
rect -758 -16422 -270 -16416
rect -758 -16456 -711 -16422
rect -677 -16456 -639 -16422
rect -605 -16456 -567 -16422
rect -533 -16456 -495 -16422
rect -461 -16456 -423 -16422
rect -389 -16456 -351 -16422
rect -317 -16456 -270 -16422
rect -758 -16462 -270 -16456
rect -556 -16524 -496 -16462
rect -758 -16530 -270 -16524
rect -758 -16564 -711 -16530
rect -677 -16564 -639 -16530
rect -605 -16564 -567 -16530
rect -533 -16564 -495 -16530
rect -461 -16564 -423 -16530
rect -389 -16564 -351 -16530
rect -317 -16564 -270 -16530
rect -758 -16570 -270 -16564
rect -1050 -16640 -1040 -16633
rect -2024 -16667 -2018 -16644
rect -2064 -16705 -2018 -16667
rect -2064 -16739 -2058 -16705
rect -2024 -16739 -2018 -16705
rect -2064 -16777 -2018 -16739
rect -2064 -16811 -2058 -16777
rect -2024 -16811 -2018 -16777
rect -2064 -16849 -2018 -16811
rect -2064 -16883 -2058 -16849
rect -2024 -16883 -2018 -16849
rect -2064 -16921 -2018 -16883
rect -2064 -16955 -2058 -16921
rect -2024 -16955 -2018 -16921
rect -2064 -16993 -2018 -16955
rect -2064 -17027 -2058 -16993
rect -2024 -17027 -2018 -16993
rect -2064 -17065 -2018 -17027
rect -2064 -17099 -2058 -17065
rect -2024 -17099 -2018 -17065
rect -2064 -17137 -2018 -17099
rect -2064 -17166 -2058 -17137
rect -3042 -17171 -3026 -17166
rect -3812 -17240 -3324 -17234
rect -3812 -17274 -3765 -17240
rect -3731 -17274 -3693 -17240
rect -3659 -17274 -3621 -17240
rect -3587 -17274 -3549 -17240
rect -3515 -17274 -3477 -17240
rect -3443 -17274 -3405 -17240
rect -3371 -17274 -3324 -17240
rect -3812 -17280 -3324 -17274
rect -3608 -17342 -3548 -17280
rect -3812 -17348 -3324 -17342
rect -3812 -17382 -3765 -17348
rect -3731 -17382 -3693 -17348
rect -3659 -17382 -3621 -17348
rect -3587 -17382 -3549 -17348
rect -3515 -17382 -3477 -17348
rect -3443 -17382 -3405 -17348
rect -3371 -17382 -3324 -17348
rect -3812 -17388 -3324 -17382
rect -4108 -17456 -4094 -17451
rect -5118 -17523 -5072 -17485
rect -5118 -17557 -5112 -17523
rect -5078 -17557 -5072 -17523
rect -5118 -17595 -5072 -17557
rect -5118 -17629 -5112 -17595
rect -5078 -17629 -5072 -17595
rect -5118 -17667 -5072 -17629
rect -5118 -17701 -5112 -17667
rect -5078 -17701 -5072 -17667
rect -5118 -17739 -5072 -17701
rect -5118 -17773 -5112 -17739
rect -5078 -17773 -5072 -17739
rect -5118 -17811 -5072 -17773
rect -5118 -17845 -5112 -17811
rect -5078 -17845 -5072 -17811
rect -5118 -17883 -5072 -17845
rect -5118 -17917 -5112 -17883
rect -5078 -17917 -5072 -17883
rect -5118 -17955 -5072 -17917
rect -5118 -17976 -5112 -17955
rect -6096 -17989 -6080 -17984
rect -6866 -18058 -6378 -18052
rect -6866 -18092 -6819 -18058
rect -6785 -18092 -6747 -18058
rect -6713 -18092 -6675 -18058
rect -6641 -18092 -6603 -18058
rect -6569 -18092 -6531 -18058
rect -6497 -18092 -6459 -18058
rect -6425 -18092 -6378 -18058
rect -6866 -18098 -6378 -18092
rect -6654 -18160 -6594 -18098
rect -6866 -18166 -6378 -18160
rect -6866 -18200 -6819 -18166
rect -6785 -18200 -6747 -18166
rect -6713 -18200 -6675 -18166
rect -6641 -18200 -6603 -18166
rect -6569 -18200 -6531 -18166
rect -6497 -18200 -6459 -18166
rect -6425 -18200 -6378 -18166
rect -6866 -18206 -6378 -18200
rect -7158 -18270 -7148 -18269
rect -8132 -18303 -8126 -18272
rect -8172 -18341 -8126 -18303
rect -8172 -18375 -8166 -18341
rect -8132 -18375 -8126 -18341
rect -8172 -18413 -8126 -18375
rect -8172 -18447 -8166 -18413
rect -8132 -18447 -8126 -18413
rect -8172 -18485 -8126 -18447
rect -8172 -18519 -8166 -18485
rect -8132 -18519 -8126 -18485
rect -8172 -18557 -8126 -18519
rect -8172 -18591 -8166 -18557
rect -8132 -18591 -8126 -18557
rect -8172 -18629 -8126 -18591
rect -8172 -18663 -8166 -18629
rect -8132 -18663 -8126 -18629
rect -8172 -18701 -8126 -18663
rect -8172 -18735 -8166 -18701
rect -8132 -18735 -8126 -18701
rect -8172 -18773 -8126 -18735
rect -8172 -18807 -8166 -18773
rect -8132 -18807 -8126 -18773
rect -7154 -18303 -7148 -18270
rect -7114 -18270 -7098 -18269
rect -6140 -18269 -6080 -17989
rect -5120 -17989 -5112 -17976
rect -5078 -17976 -5072 -17955
rect -4100 -17485 -4094 -17456
rect -4060 -17456 -4048 -17451
rect -3086 -17451 -3026 -17171
rect -2066 -17171 -2058 -17166
rect -2024 -17166 -2018 -17137
rect -1046 -16667 -1040 -16640
rect -1006 -16640 -990 -16633
rect -28 -16633 32 -16354
rect -1006 -16667 -1000 -16640
rect -1046 -16705 -1000 -16667
rect -1046 -16739 -1040 -16705
rect -1006 -16739 -1000 -16705
rect -1046 -16777 -1000 -16739
rect -1046 -16811 -1040 -16777
rect -1006 -16811 -1000 -16777
rect -1046 -16849 -1000 -16811
rect -1046 -16883 -1040 -16849
rect -1006 -16883 -1000 -16849
rect -1046 -16921 -1000 -16883
rect -1046 -16955 -1040 -16921
rect -1006 -16955 -1000 -16921
rect -1046 -16993 -1000 -16955
rect -1046 -17027 -1040 -16993
rect -1006 -17027 -1000 -16993
rect -1046 -17065 -1000 -17027
rect -1046 -17099 -1040 -17065
rect -1006 -17099 -1000 -17065
rect -1046 -17137 -1000 -17099
rect -1046 -17162 -1040 -17137
rect -2024 -17171 -2006 -17166
rect -2794 -17240 -2306 -17234
rect -2794 -17274 -2747 -17240
rect -2713 -17274 -2675 -17240
rect -2641 -17274 -2603 -17240
rect -2569 -17274 -2531 -17240
rect -2497 -17274 -2459 -17240
rect -2425 -17274 -2387 -17240
rect -2353 -17274 -2306 -17240
rect -2794 -17280 -2306 -17274
rect -2586 -17342 -2526 -17280
rect -2794 -17348 -2306 -17342
rect -2794 -17382 -2747 -17348
rect -2713 -17382 -2675 -17348
rect -2641 -17382 -2603 -17348
rect -2569 -17382 -2531 -17348
rect -2497 -17382 -2459 -17348
rect -2425 -17382 -2387 -17348
rect -2353 -17382 -2306 -17348
rect -2794 -17388 -2306 -17382
rect -3086 -17456 -3076 -17451
rect -4060 -17485 -4054 -17456
rect -4100 -17523 -4054 -17485
rect -4100 -17557 -4094 -17523
rect -4060 -17557 -4054 -17523
rect -4100 -17595 -4054 -17557
rect -4100 -17629 -4094 -17595
rect -4060 -17629 -4054 -17595
rect -4100 -17667 -4054 -17629
rect -4100 -17701 -4094 -17667
rect -4060 -17701 -4054 -17667
rect -4100 -17739 -4054 -17701
rect -4100 -17773 -4094 -17739
rect -4060 -17773 -4054 -17739
rect -4100 -17811 -4054 -17773
rect -4100 -17845 -4094 -17811
rect -4060 -17845 -4054 -17811
rect -4100 -17883 -4054 -17845
rect -4100 -17917 -4094 -17883
rect -4060 -17917 -4054 -17883
rect -4100 -17955 -4054 -17917
rect -5078 -17989 -5060 -17976
rect -4100 -17984 -4094 -17955
rect -5848 -18058 -5360 -18052
rect -5848 -18092 -5801 -18058
rect -5767 -18092 -5729 -18058
rect -5695 -18092 -5657 -18058
rect -5623 -18092 -5585 -18058
rect -5551 -18092 -5513 -18058
rect -5479 -18092 -5441 -18058
rect -5407 -18092 -5360 -18058
rect -5848 -18098 -5360 -18092
rect -5652 -18160 -5592 -18098
rect -5848 -18166 -5360 -18160
rect -5848 -18200 -5801 -18166
rect -5767 -18200 -5729 -18166
rect -5695 -18200 -5657 -18166
rect -5623 -18200 -5585 -18166
rect -5551 -18200 -5513 -18166
rect -5479 -18200 -5441 -18166
rect -5407 -18200 -5360 -18166
rect -5848 -18206 -5360 -18200
rect -5120 -18266 -5060 -17989
rect -4108 -17989 -4094 -17984
rect -4060 -17984 -4054 -17955
rect -3082 -17485 -3076 -17456
rect -3042 -17456 -3026 -17451
rect -2066 -17451 -2006 -17171
rect -1050 -17171 -1040 -17162
rect -1006 -17162 -1000 -17137
rect -28 -16667 -22 -16633
rect 12 -16644 32 -16633
rect 12 -16667 18 -16644
rect -28 -16705 18 -16667
rect -28 -16739 -22 -16705
rect 12 -16739 18 -16705
rect -28 -16777 18 -16739
rect -28 -16811 -22 -16777
rect 12 -16811 18 -16777
rect -28 -16849 18 -16811
rect -28 -16883 -22 -16849
rect 12 -16883 18 -16849
rect -28 -16921 18 -16883
rect -28 -16955 -22 -16921
rect 12 -16955 18 -16921
rect -28 -16993 18 -16955
rect -28 -17027 -22 -16993
rect 12 -17027 18 -16993
rect -28 -17065 18 -17027
rect -28 -17099 -22 -17065
rect 12 -17099 18 -17065
rect -28 -17137 18 -17099
rect -1006 -17171 -990 -17162
rect -1776 -17240 -1288 -17234
rect -1776 -17274 -1729 -17240
rect -1695 -17274 -1657 -17240
rect -1623 -17274 -1585 -17240
rect -1551 -17274 -1513 -17240
rect -1479 -17274 -1441 -17240
rect -1407 -17274 -1369 -17240
rect -1335 -17274 -1288 -17240
rect -1776 -17280 -1288 -17274
rect -1574 -17342 -1514 -17280
rect -1776 -17348 -1288 -17342
rect -1776 -17382 -1729 -17348
rect -1695 -17382 -1657 -17348
rect -1623 -17382 -1585 -17348
rect -1551 -17382 -1513 -17348
rect -1479 -17382 -1441 -17348
rect -1407 -17382 -1369 -17348
rect -1335 -17382 -1288 -17348
rect -1776 -17388 -1288 -17382
rect -2066 -17456 -2058 -17451
rect -3042 -17485 -3036 -17456
rect -3082 -17523 -3036 -17485
rect -3082 -17557 -3076 -17523
rect -3042 -17557 -3036 -17523
rect -3082 -17595 -3036 -17557
rect -3082 -17629 -3076 -17595
rect -3042 -17629 -3036 -17595
rect -3082 -17667 -3036 -17629
rect -3082 -17701 -3076 -17667
rect -3042 -17701 -3036 -17667
rect -3082 -17739 -3036 -17701
rect -3082 -17773 -3076 -17739
rect -3042 -17773 -3036 -17739
rect -3082 -17811 -3036 -17773
rect -3082 -17845 -3076 -17811
rect -3042 -17845 -3036 -17811
rect -3082 -17883 -3036 -17845
rect -3082 -17917 -3076 -17883
rect -3042 -17917 -3036 -17883
rect -3082 -17955 -3036 -17917
rect -3082 -17984 -3076 -17955
rect -4060 -17989 -4048 -17984
rect -4830 -18058 -4342 -18052
rect -4830 -18092 -4783 -18058
rect -4749 -18092 -4711 -18058
rect -4677 -18092 -4639 -18058
rect -4605 -18092 -4567 -18058
rect -4533 -18092 -4495 -18058
rect -4461 -18092 -4423 -18058
rect -4389 -18092 -4342 -18058
rect -4830 -18098 -4342 -18092
rect -4622 -18160 -4562 -18098
rect -4830 -18166 -4342 -18160
rect -4830 -18200 -4783 -18166
rect -4749 -18200 -4711 -18166
rect -4677 -18200 -4639 -18166
rect -4605 -18200 -4567 -18166
rect -4533 -18200 -4495 -18166
rect -4461 -18200 -4423 -18166
rect -4389 -18200 -4342 -18166
rect -4830 -18206 -4342 -18200
rect -7114 -18303 -7108 -18270
rect -6140 -18274 -6130 -18269
rect -7154 -18341 -7108 -18303
rect -7154 -18375 -7148 -18341
rect -7114 -18375 -7108 -18341
rect -7154 -18413 -7108 -18375
rect -7154 -18447 -7148 -18413
rect -7114 -18447 -7108 -18413
rect -7154 -18485 -7108 -18447
rect -7154 -18519 -7148 -18485
rect -7114 -18519 -7108 -18485
rect -7154 -18557 -7108 -18519
rect -7154 -18591 -7148 -18557
rect -7114 -18591 -7108 -18557
rect -7154 -18629 -7108 -18591
rect -7154 -18663 -7148 -18629
rect -7114 -18663 -7108 -18629
rect -7154 -18701 -7108 -18663
rect -7154 -18735 -7148 -18701
rect -7114 -18735 -7108 -18701
rect -7154 -18773 -7108 -18735
rect -7154 -18780 -7148 -18773
rect -8172 -18838 -8126 -18807
rect -7164 -18807 -7148 -18780
rect -7114 -18780 -7108 -18773
rect -6136 -18303 -6130 -18274
rect -6096 -18274 -6080 -18269
rect -5118 -18269 -5072 -18266
rect -6096 -18303 -6090 -18274
rect -6136 -18341 -6090 -18303
rect -6136 -18375 -6130 -18341
rect -6096 -18375 -6090 -18341
rect -6136 -18413 -6090 -18375
rect -6136 -18447 -6130 -18413
rect -6096 -18447 -6090 -18413
rect -6136 -18485 -6090 -18447
rect -6136 -18519 -6130 -18485
rect -6096 -18519 -6090 -18485
rect -6136 -18557 -6090 -18519
rect -6136 -18591 -6130 -18557
rect -6096 -18591 -6090 -18557
rect -6136 -18629 -6090 -18591
rect -6136 -18663 -6130 -18629
rect -6096 -18663 -6090 -18629
rect -6136 -18701 -6090 -18663
rect -6136 -18735 -6130 -18701
rect -6096 -18735 -6090 -18701
rect -6136 -18773 -6090 -18735
rect -7114 -18807 -7104 -18780
rect -12328 -18893 -12289 -18859
rect -12255 -18893 -12216 -18859
rect -12328 -18931 -12216 -18893
rect -8902 -18876 -8414 -18870
rect -8902 -18910 -8855 -18876
rect -8821 -18910 -8783 -18876
rect -8749 -18910 -8711 -18876
rect -8677 -18910 -8639 -18876
rect -8605 -18910 -8567 -18876
rect -8533 -18910 -8495 -18876
rect -8461 -18910 -8414 -18876
rect -8902 -18916 -8414 -18910
rect -7884 -18876 -7396 -18870
rect -7884 -18910 -7837 -18876
rect -7803 -18910 -7765 -18876
rect -7731 -18910 -7693 -18876
rect -7659 -18910 -7621 -18876
rect -7587 -18910 -7549 -18876
rect -7515 -18910 -7477 -18876
rect -7443 -18910 -7396 -18876
rect -7884 -18916 -7672 -18910
rect -7612 -18916 -7396 -18910
rect -12328 -18965 -12289 -18931
rect -12255 -18965 -12216 -18931
rect -12328 -19003 -12216 -18965
rect -12328 -19037 -12289 -19003
rect -12255 -19037 -12216 -19003
rect -12328 -19075 -12216 -19037
rect -7164 -19000 -7104 -18807
rect -6136 -18807 -6130 -18773
rect -6096 -18807 -6090 -18773
rect -5118 -18303 -5112 -18269
rect -5078 -18303 -5072 -18269
rect -4108 -18269 -4048 -17989
rect -3086 -17989 -3076 -17984
rect -3042 -17984 -3036 -17955
rect -2064 -17485 -2058 -17456
rect -2024 -17456 -2006 -17451
rect -1050 -17451 -990 -17171
rect -28 -17171 -22 -17137
rect 12 -17166 18 -17137
rect 12 -17171 32 -17166
rect -758 -17240 -270 -17234
rect -758 -17274 -711 -17240
rect -677 -17274 -639 -17240
rect -605 -17274 -567 -17240
rect -533 -17274 -495 -17240
rect -461 -17274 -423 -17240
rect -389 -17274 -351 -17240
rect -317 -17274 -270 -17240
rect -758 -17280 -270 -17274
rect -554 -17342 -494 -17280
rect -758 -17348 -270 -17342
rect -758 -17382 -711 -17348
rect -677 -17382 -639 -17348
rect -605 -17382 -567 -17348
rect -533 -17382 -495 -17348
rect -461 -17382 -423 -17348
rect -389 -17382 -351 -17348
rect -317 -17382 -270 -17348
rect -758 -17388 -270 -17382
rect -1050 -17452 -1040 -17451
rect -2024 -17485 -2018 -17456
rect -2064 -17523 -2018 -17485
rect -2064 -17557 -2058 -17523
rect -2024 -17557 -2018 -17523
rect -2064 -17595 -2018 -17557
rect -2064 -17629 -2058 -17595
rect -2024 -17629 -2018 -17595
rect -2064 -17667 -2018 -17629
rect -2064 -17701 -2058 -17667
rect -2024 -17701 -2018 -17667
rect -2064 -17739 -2018 -17701
rect -2064 -17773 -2058 -17739
rect -2024 -17773 -2018 -17739
rect -2064 -17811 -2018 -17773
rect -2064 -17845 -2058 -17811
rect -2024 -17845 -2018 -17811
rect -2064 -17883 -2018 -17845
rect -2064 -17917 -2058 -17883
rect -2024 -17917 -2018 -17883
rect -2064 -17955 -2018 -17917
rect -2064 -17984 -2058 -17955
rect -3042 -17989 -3026 -17984
rect -3812 -18058 -3324 -18052
rect -3812 -18092 -3765 -18058
rect -3731 -18092 -3693 -18058
rect -3659 -18092 -3621 -18058
rect -3587 -18092 -3549 -18058
rect -3515 -18092 -3477 -18058
rect -3443 -18092 -3405 -18058
rect -3371 -18092 -3324 -18058
rect -3812 -18098 -3324 -18092
rect -3606 -18160 -3546 -18098
rect -3812 -18166 -3324 -18160
rect -3812 -18200 -3765 -18166
rect -3731 -18200 -3693 -18166
rect -3659 -18200 -3621 -18166
rect -3587 -18200 -3549 -18166
rect -3515 -18200 -3477 -18166
rect -3443 -18200 -3405 -18166
rect -3371 -18200 -3324 -18166
rect -3812 -18206 -3324 -18200
rect -4108 -18274 -4094 -18269
rect -5118 -18341 -5072 -18303
rect -5118 -18375 -5112 -18341
rect -5078 -18375 -5072 -18341
rect -5118 -18413 -5072 -18375
rect -5118 -18447 -5112 -18413
rect -5078 -18447 -5072 -18413
rect -5118 -18485 -5072 -18447
rect -5118 -18519 -5112 -18485
rect -5078 -18519 -5072 -18485
rect -5118 -18557 -5072 -18519
rect -5118 -18591 -5112 -18557
rect -5078 -18591 -5072 -18557
rect -5118 -18629 -5072 -18591
rect -5118 -18663 -5112 -18629
rect -5078 -18663 -5072 -18629
rect -5118 -18701 -5072 -18663
rect -5118 -18735 -5112 -18701
rect -5078 -18735 -5072 -18701
rect -5118 -18773 -5072 -18735
rect -5118 -18778 -5112 -18773
rect -6136 -18838 -6090 -18807
rect -5126 -18807 -5112 -18778
rect -5078 -18778 -5072 -18773
rect -4100 -18303 -4094 -18274
rect -4060 -18274 -4048 -18269
rect -3086 -18269 -3026 -17989
rect -2066 -17989 -2058 -17984
rect -2024 -17984 -2018 -17955
rect -1046 -17485 -1040 -17452
rect -1006 -17452 -990 -17451
rect -28 -17451 32 -17171
rect -1006 -17485 -1000 -17452
rect -1046 -17523 -1000 -17485
rect -1046 -17557 -1040 -17523
rect -1006 -17557 -1000 -17523
rect -1046 -17595 -1000 -17557
rect -1046 -17629 -1040 -17595
rect -1006 -17629 -1000 -17595
rect -1046 -17667 -1000 -17629
rect -1046 -17701 -1040 -17667
rect -1006 -17701 -1000 -17667
rect -1046 -17739 -1000 -17701
rect -1046 -17773 -1040 -17739
rect -1006 -17773 -1000 -17739
rect -1046 -17811 -1000 -17773
rect -1046 -17845 -1040 -17811
rect -1006 -17845 -1000 -17811
rect -1046 -17883 -1000 -17845
rect -1046 -17917 -1040 -17883
rect -1006 -17917 -1000 -17883
rect -1046 -17955 -1000 -17917
rect -1046 -17980 -1040 -17955
rect -2024 -17989 -2006 -17984
rect -2794 -18058 -2306 -18052
rect -2794 -18092 -2747 -18058
rect -2713 -18092 -2675 -18058
rect -2641 -18092 -2603 -18058
rect -2569 -18092 -2531 -18058
rect -2497 -18092 -2459 -18058
rect -2425 -18092 -2387 -18058
rect -2353 -18092 -2306 -18058
rect -2794 -18098 -2306 -18092
rect -2584 -18160 -2524 -18098
rect -2794 -18166 -2306 -18160
rect -2794 -18200 -2747 -18166
rect -2713 -18200 -2675 -18166
rect -2641 -18200 -2603 -18166
rect -2569 -18200 -2531 -18166
rect -2497 -18200 -2459 -18166
rect -2425 -18200 -2387 -18166
rect -2353 -18200 -2306 -18166
rect -2794 -18206 -2306 -18200
rect -3086 -18274 -3076 -18269
rect -4060 -18303 -4054 -18274
rect -4100 -18341 -4054 -18303
rect -4100 -18375 -4094 -18341
rect -4060 -18375 -4054 -18341
rect -4100 -18413 -4054 -18375
rect -4100 -18447 -4094 -18413
rect -4060 -18447 -4054 -18413
rect -4100 -18485 -4054 -18447
rect -4100 -18519 -4094 -18485
rect -4060 -18519 -4054 -18485
rect -4100 -18557 -4054 -18519
rect -4100 -18591 -4094 -18557
rect -4060 -18591 -4054 -18557
rect -4100 -18629 -4054 -18591
rect -4100 -18663 -4094 -18629
rect -4060 -18663 -4054 -18629
rect -4100 -18701 -4054 -18663
rect -4100 -18735 -4094 -18701
rect -4060 -18735 -4054 -18701
rect -4100 -18773 -4054 -18735
rect -5078 -18807 -5066 -18778
rect -6866 -18876 -6378 -18870
rect -6866 -18910 -6819 -18876
rect -6785 -18910 -6747 -18876
rect -6713 -18910 -6675 -18876
rect -6641 -18910 -6603 -18876
rect -6569 -18910 -6531 -18876
rect -6497 -18910 -6459 -18876
rect -6425 -18910 -6378 -18876
rect -6866 -18916 -6378 -18910
rect -5848 -18876 -5360 -18870
rect -5848 -18910 -5801 -18876
rect -5767 -18910 -5729 -18876
rect -5695 -18910 -5657 -18876
rect -5623 -18910 -5585 -18876
rect -5551 -18910 -5513 -18876
rect -5479 -18910 -5441 -18876
rect -5407 -18910 -5360 -18876
rect -5848 -18916 -5360 -18910
rect -5126 -19000 -5066 -18807
rect -4100 -18807 -4094 -18773
rect -4060 -18807 -4054 -18773
rect -3082 -18303 -3076 -18274
rect -3042 -18274 -3026 -18269
rect -2066 -18269 -2006 -17989
rect -1050 -17989 -1040 -17980
rect -1006 -17980 -1000 -17955
rect -28 -17485 -22 -17451
rect 12 -17456 32 -17451
rect 12 -17485 18 -17456
rect -28 -17523 18 -17485
rect -28 -17557 -22 -17523
rect 12 -17557 18 -17523
rect -28 -17595 18 -17557
rect -28 -17629 -22 -17595
rect 12 -17629 18 -17595
rect -28 -17667 18 -17629
rect -28 -17701 -22 -17667
rect 12 -17701 18 -17667
rect -28 -17739 18 -17701
rect -28 -17773 -22 -17739
rect 12 -17773 18 -17739
rect -28 -17811 18 -17773
rect -28 -17845 -22 -17811
rect 12 -17845 18 -17811
rect -28 -17883 18 -17845
rect -28 -17917 -22 -17883
rect 12 -17917 18 -17883
rect -28 -17955 18 -17917
rect -1006 -17989 -990 -17980
rect -1776 -18058 -1288 -18052
rect -1776 -18092 -1729 -18058
rect -1695 -18092 -1657 -18058
rect -1623 -18092 -1585 -18058
rect -1551 -18092 -1513 -18058
rect -1479 -18092 -1441 -18058
rect -1407 -18092 -1369 -18058
rect -1335 -18092 -1288 -18058
rect -1776 -18098 -1288 -18092
rect -1572 -18160 -1512 -18098
rect -1776 -18166 -1288 -18160
rect -1776 -18200 -1729 -18166
rect -1695 -18200 -1657 -18166
rect -1623 -18200 -1585 -18166
rect -1551 -18200 -1513 -18166
rect -1479 -18200 -1441 -18166
rect -1407 -18200 -1369 -18166
rect -1335 -18200 -1288 -18166
rect -1776 -18206 -1288 -18200
rect -2066 -18274 -2058 -18269
rect -3042 -18303 -3036 -18274
rect -3082 -18341 -3036 -18303
rect -3082 -18375 -3076 -18341
rect -3042 -18375 -3036 -18341
rect -3082 -18413 -3036 -18375
rect -3082 -18447 -3076 -18413
rect -3042 -18447 -3036 -18413
rect -3082 -18485 -3036 -18447
rect -3082 -18519 -3076 -18485
rect -3042 -18519 -3036 -18485
rect -3082 -18557 -3036 -18519
rect -3082 -18591 -3076 -18557
rect -3042 -18591 -3036 -18557
rect -3082 -18629 -3036 -18591
rect -3082 -18663 -3076 -18629
rect -3042 -18663 -3036 -18629
rect -3082 -18701 -3036 -18663
rect -3082 -18735 -3076 -18701
rect -3042 -18735 -3036 -18701
rect -3082 -18773 -3036 -18735
rect -3082 -18782 -3076 -18773
rect -4100 -18838 -4054 -18807
rect -3090 -18807 -3076 -18782
rect -3042 -18782 -3036 -18773
rect -2064 -18303 -2058 -18274
rect -2024 -18274 -2006 -18269
rect -1050 -18269 -990 -17989
rect -28 -17989 -22 -17955
rect 12 -17984 18 -17955
rect 12 -17989 32 -17984
rect -758 -18058 -270 -18052
rect -758 -18092 -711 -18058
rect -677 -18092 -639 -18058
rect -605 -18092 -567 -18058
rect -533 -18092 -495 -18058
rect -461 -18092 -423 -18058
rect -389 -18092 -351 -18058
rect -317 -18092 -270 -18058
rect -758 -18098 -270 -18092
rect -552 -18160 -492 -18098
rect -758 -18166 -270 -18160
rect -758 -18200 -711 -18166
rect -677 -18200 -639 -18166
rect -605 -18200 -567 -18166
rect -533 -18200 -495 -18166
rect -461 -18200 -423 -18166
rect -389 -18200 -351 -18166
rect -317 -18200 -270 -18166
rect -758 -18206 -270 -18200
rect -1050 -18270 -1040 -18269
rect -2024 -18303 -2018 -18274
rect -2064 -18341 -2018 -18303
rect -2064 -18375 -2058 -18341
rect -2024 -18375 -2018 -18341
rect -2064 -18413 -2018 -18375
rect -2064 -18447 -2058 -18413
rect -2024 -18447 -2018 -18413
rect -2064 -18485 -2018 -18447
rect -2064 -18519 -2058 -18485
rect -2024 -18519 -2018 -18485
rect -2064 -18557 -2018 -18519
rect -2064 -18591 -2058 -18557
rect -2024 -18591 -2018 -18557
rect -2064 -18629 -2018 -18591
rect -2064 -18663 -2058 -18629
rect -2024 -18663 -2018 -18629
rect -2064 -18701 -2018 -18663
rect -2064 -18735 -2058 -18701
rect -2024 -18735 -2018 -18701
rect -2064 -18773 -2018 -18735
rect -3042 -18807 -3030 -18782
rect -4830 -18876 -4342 -18870
rect -4830 -18910 -4783 -18876
rect -4749 -18910 -4711 -18876
rect -4677 -18910 -4639 -18876
rect -4605 -18910 -4567 -18876
rect -4533 -18910 -4495 -18876
rect -4461 -18910 -4423 -18876
rect -4389 -18910 -4342 -18876
rect -4830 -18916 -4342 -18910
rect -3812 -18876 -3324 -18870
rect -3812 -18910 -3765 -18876
rect -3731 -18910 -3693 -18876
rect -3659 -18910 -3621 -18876
rect -3587 -18910 -3549 -18876
rect -3515 -18910 -3477 -18876
rect -3443 -18910 -3405 -18876
rect -3371 -18910 -3324 -18876
rect -3812 -18916 -3324 -18910
rect -3090 -19000 -3030 -18807
rect -2064 -18807 -2058 -18773
rect -2024 -18807 -2018 -18773
rect -1046 -18303 -1040 -18270
rect -1006 -18270 -990 -18269
rect -28 -18269 32 -17989
rect -1006 -18303 -1000 -18270
rect -1046 -18341 -1000 -18303
rect -1046 -18375 -1040 -18341
rect -1006 -18375 -1000 -18341
rect -1046 -18413 -1000 -18375
rect -1046 -18447 -1040 -18413
rect -1006 -18447 -1000 -18413
rect -1046 -18485 -1000 -18447
rect -1046 -18519 -1040 -18485
rect -1006 -18519 -1000 -18485
rect -1046 -18557 -1000 -18519
rect -1046 -18591 -1040 -18557
rect -1006 -18591 -1000 -18557
rect -1046 -18629 -1000 -18591
rect -1046 -18663 -1040 -18629
rect -1006 -18663 -1000 -18629
rect -1046 -18701 -1000 -18663
rect -1046 -18735 -1040 -18701
rect -1006 -18735 -1000 -18701
rect -1046 -18773 -1000 -18735
rect -28 -18303 -22 -18269
rect 12 -18274 32 -18269
rect 12 -18303 18 -18274
rect -28 -18341 18 -18303
rect -28 -18375 -22 -18341
rect 12 -18375 18 -18341
rect -28 -18413 18 -18375
rect -28 -18447 -22 -18413
rect 12 -18447 18 -18413
rect -28 -18485 18 -18447
rect -28 -18519 -22 -18485
rect 12 -18519 18 -18485
rect -28 -18557 18 -18519
rect -28 -18591 -22 -18557
rect 12 -18591 18 -18557
rect -28 -18629 18 -18591
rect -28 -18663 -22 -18629
rect 12 -18663 18 -18629
rect -28 -18701 18 -18663
rect -28 -18735 -22 -18701
rect 12 -18735 18 -18701
rect -28 -18772 18 -18735
rect -1046 -18784 -1040 -18773
rect -2064 -18838 -2018 -18807
rect -1054 -18807 -1040 -18784
rect -1006 -18784 -1000 -18773
rect -34 -18773 26 -18772
rect -1006 -18807 -994 -18784
rect -2794 -18876 -2306 -18870
rect -2794 -18910 -2747 -18876
rect -2713 -18910 -2675 -18876
rect -2641 -18910 -2603 -18876
rect -2569 -18910 -2531 -18876
rect -2497 -18910 -2459 -18876
rect -2425 -18910 -2387 -18876
rect -2353 -18910 -2306 -18876
rect -2794 -18916 -2306 -18910
rect -1776 -18876 -1288 -18870
rect -1776 -18910 -1729 -18876
rect -1695 -18910 -1657 -18876
rect -1623 -18910 -1585 -18876
rect -1551 -18910 -1513 -18876
rect -1479 -18910 -1441 -18876
rect -1407 -18910 -1369 -18876
rect -1335 -18910 -1288 -18876
rect -1776 -18916 -1288 -18910
rect -1054 -19000 -994 -18807
rect -34 -18807 -22 -18773
rect 12 -18807 26 -18773
rect -758 -18876 -270 -18870
rect -758 -18910 -711 -18876
rect -677 -18910 -639 -18876
rect -605 -18910 -567 -18876
rect -533 -18910 -495 -18876
rect -461 -18910 -423 -18876
rect -389 -18910 -351 -18876
rect -317 -18910 -270 -18876
rect -758 -18916 -270 -18910
rect -540 -19000 -480 -18916
rect -34 -19000 26 -18807
rect 1150 -18822 1210 -11682
rect 1144 -18826 1216 -18822
rect 1144 -18878 1154 -18826
rect 1206 -18878 1216 -18826
rect 1144 -18882 1216 -18878
rect -7164 -19060 1130 -19000
rect -12328 -19109 -12289 -19075
rect -12255 -19109 -12216 -19075
rect -12328 -19147 -12216 -19109
rect -12328 -19181 -12289 -19147
rect -12255 -19181 -12216 -19147
rect -12328 -19219 -12216 -19181
rect -12328 -19253 -12289 -19219
rect -12255 -19253 -12216 -19219
rect -12328 -19291 -12216 -19253
rect -12328 -19325 -12289 -19291
rect -12255 -19325 -12216 -19291
rect -12328 -19363 -12216 -19325
rect -12328 -19397 -12289 -19363
rect -12255 -19397 -12216 -19363
rect -12328 -19435 -12216 -19397
rect -12328 -19469 -12289 -19435
rect -12255 -19469 -12216 -19435
rect -12328 -19507 -12216 -19469
rect -12328 -19541 -12289 -19507
rect -12255 -19541 -12216 -19507
rect -12328 -19579 -12216 -19541
rect -12328 -19613 -12289 -19579
rect -12255 -19613 -12216 -19579
rect -12328 -19651 -12216 -19613
rect -12328 -19685 -12289 -19651
rect -12255 -19685 -12216 -19651
rect -12328 -19723 -12216 -19685
rect -12328 -19757 -12289 -19723
rect -12255 -19757 -12216 -19723
rect -12328 -19795 -12216 -19757
rect -12328 -19829 -12289 -19795
rect -12255 -19829 -12216 -19795
rect -3404 -19752 -3332 -19748
rect -3404 -19804 -3394 -19752
rect -3342 -19804 -3332 -19752
rect -3404 -19808 -3332 -19804
rect -12328 -19867 -12216 -19829
rect -12328 -19901 -12289 -19867
rect -12255 -19901 -12216 -19867
rect -12328 -19939 -12216 -19901
rect -12328 -19973 -12289 -19939
rect -12255 -19973 -12216 -19939
rect -12328 -20011 -12216 -19973
rect -12328 -20045 -12289 -20011
rect -12255 -20045 -12216 -20011
rect -9508 -19898 -9448 -19888
rect -9508 -19950 -9504 -19898
rect -9452 -19950 -9448 -19898
rect -12328 -20083 -12216 -20045
rect -10668 -20026 -10596 -20022
rect -10668 -20078 -10658 -20026
rect -10606 -20078 -10596 -20026
rect -10668 -20082 -10596 -20078
rect -12328 -20117 -12289 -20083
rect -12255 -20117 -12216 -20083
rect -12328 -20155 -12216 -20117
rect -12328 -20189 -12289 -20155
rect -12255 -20189 -12216 -20155
rect -12328 -20227 -12216 -20189
rect -12328 -20261 -12289 -20227
rect -12255 -20261 -12216 -20227
rect -12328 -20299 -12216 -20261
rect -12328 -20333 -12289 -20299
rect -12255 -20333 -12216 -20299
rect -12328 -20371 -12216 -20333
rect -12328 -20405 -12289 -20371
rect -12255 -20405 -12216 -20371
rect -12328 -20443 -12216 -20405
rect -12328 -20477 -12289 -20443
rect -12255 -20477 -12216 -20443
rect -12328 -20515 -12216 -20477
rect -12328 -20549 -12289 -20515
rect -12255 -20549 -12216 -20515
rect -12328 -20587 -12216 -20549
rect -12328 -20621 -12289 -20587
rect -12255 -20621 -12216 -20587
rect -12328 -20659 -12216 -20621
rect -12328 -20693 -12289 -20659
rect -12255 -20693 -12216 -20659
rect -12328 -20731 -12216 -20693
rect -12328 -20765 -12289 -20731
rect -12255 -20765 -12216 -20731
rect -12328 -20803 -12216 -20765
rect -12328 -20837 -12289 -20803
rect -12255 -20837 -12216 -20803
rect -12328 -20875 -12216 -20837
rect -12328 -20909 -12289 -20875
rect -12255 -20909 -12216 -20875
rect -12328 -20947 -12216 -20909
rect -12328 -20981 -12289 -20947
rect -12255 -20981 -12216 -20947
rect -12328 -21019 -12216 -20981
rect -12328 -21053 -12289 -21019
rect -12255 -21053 -12216 -21019
rect -12328 -21091 -12216 -21053
rect -12328 -21125 -12289 -21091
rect -12255 -21125 -12216 -21091
rect -12328 -21163 -12216 -21125
rect -12328 -21197 -12289 -21163
rect -12255 -21197 -12216 -21163
rect -12328 -21235 -12216 -21197
rect -12328 -21269 -12289 -21235
rect -12255 -21269 -12216 -21235
rect -12328 -21307 -12216 -21269
rect -12328 -21341 -12289 -21307
rect -12255 -21341 -12216 -21307
rect -12328 -21379 -12216 -21341
rect -12328 -21413 -12289 -21379
rect -12255 -21413 -12216 -21379
rect -12328 -21451 -12216 -21413
rect -12328 -21485 -12289 -21451
rect -12255 -21485 -12216 -21451
rect -12328 -21523 -12216 -21485
rect -12328 -21557 -12289 -21523
rect -12255 -21557 -12216 -21523
rect -12328 -21595 -12216 -21557
rect -12328 -21629 -12289 -21595
rect -12255 -21629 -12216 -21595
rect -12328 -21667 -12216 -21629
rect -12328 -21701 -12289 -21667
rect -12255 -21701 -12216 -21667
rect -12328 -21739 -12216 -21701
rect -12328 -21773 -12289 -21739
rect -12255 -21773 -12216 -21739
rect -12328 -21811 -12216 -21773
rect -12328 -21845 -12289 -21811
rect -12255 -21845 -12216 -21811
rect -12328 -21883 -12216 -21845
rect -12328 -21917 -12289 -21883
rect -12255 -21917 -12216 -21883
rect -12328 -21955 -12216 -21917
rect -12328 -21989 -12289 -21955
rect -12255 -21989 -12216 -21955
rect -12328 -22027 -12216 -21989
rect -12328 -22061 -12289 -22027
rect -12255 -22061 -12216 -22027
rect -12328 -22099 -12216 -22061
rect -12328 -22133 -12289 -22099
rect -12255 -22133 -12216 -22099
rect -12328 -22171 -12216 -22133
rect -12328 -22205 -12289 -22171
rect -12255 -22205 -12216 -22171
rect -12328 -22243 -12216 -22205
rect -12328 -22277 -12289 -22243
rect -12255 -22277 -12216 -22243
rect -10662 -22254 -10602 -20082
rect -9508 -20086 -9448 -19950
rect -5434 -19898 -5362 -19894
rect -5434 -19950 -5424 -19898
rect -5372 -19950 -5362 -19898
rect -5434 -19954 -5362 -19950
rect -7990 -20026 -7918 -20022
rect -7990 -20078 -7980 -20026
rect -7928 -20078 -7918 -20026
rect -7990 -20082 -7918 -20078
rect -6958 -20026 -6886 -20022
rect -6958 -20078 -6948 -20026
rect -6896 -20078 -6886 -20026
rect -6958 -20082 -6886 -20078
rect -10524 -20146 -9448 -20086
rect -10524 -20320 -10464 -20146
rect -10016 -20228 -9956 -20146
rect -9508 -20314 -9448 -20146
rect -7984 -20224 -7924 -20082
rect -6952 -20220 -6892 -20082
rect -5428 -20338 -5368 -19954
rect -3898 -20026 -3826 -20022
rect -3898 -20078 -3888 -20026
rect -3836 -20078 -3826 -20026
rect -3898 -20082 -3826 -20078
rect -3892 -20220 -3832 -20082
rect -9004 -20984 -8944 -20904
rect -9010 -20988 -8938 -20984
rect -9010 -21040 -9000 -20988
rect -8948 -21040 -8938 -20988
rect -9010 -21044 -8938 -21040
rect -9510 -21092 -9438 -21088
rect -9510 -21144 -9500 -21092
rect -9448 -21144 -9438 -21092
rect -9510 -21148 -9438 -21144
rect -9504 -21190 -9444 -21148
rect -10524 -21250 -9444 -21190
rect -10524 -21432 -10464 -21250
rect -10020 -21328 -9960 -21250
rect -12328 -22315 -12216 -22277
rect -10668 -22258 -10596 -22254
rect -10668 -22310 -10658 -22258
rect -10606 -22310 -10596 -22258
rect -10668 -22314 -10596 -22310
rect -12328 -22349 -12289 -22315
rect -12255 -22349 -12216 -22315
rect -12328 -22387 -12216 -22349
rect -12328 -22421 -12289 -22387
rect -12255 -22421 -12216 -22387
rect -12328 -22459 -12216 -22421
rect -12328 -22493 -12289 -22459
rect -12255 -22493 -12216 -22459
rect -12328 -22531 -12216 -22493
rect -12328 -22565 -12289 -22531
rect -12255 -22565 -12216 -22531
rect -12328 -22603 -12216 -22565
rect -12328 -22637 -12289 -22603
rect -12255 -22637 -12216 -22603
rect -12328 -22675 -12216 -22637
rect -12328 -22709 -12289 -22675
rect -12255 -22709 -12216 -22675
rect -12328 -22747 -12216 -22709
rect -12328 -22781 -12289 -22747
rect -12255 -22781 -12216 -22747
rect -12328 -22819 -12216 -22781
rect -12328 -22853 -12289 -22819
rect -12255 -22853 -12216 -22819
rect -12328 -22891 -12216 -22853
rect -12328 -22925 -12289 -22891
rect -12255 -22925 -12216 -22891
rect -12328 -22963 -12216 -22925
rect -12328 -22997 -12289 -22963
rect -12255 -22997 -12216 -22963
rect -12328 -23035 -12216 -22997
rect -12328 -23069 -12289 -23035
rect -12255 -23069 -12216 -23035
rect -12328 -23107 -12216 -23069
rect -12328 -23141 -12289 -23107
rect -12255 -23141 -12216 -23107
rect -12328 -23179 -12216 -23141
rect -12328 -23213 -12289 -23179
rect -12255 -23213 -12216 -23179
rect -12328 -23251 -12216 -23213
rect -12328 -23285 -12289 -23251
rect -12255 -23285 -12216 -23251
rect -12328 -23323 -12216 -23285
rect -12328 -23357 -12289 -23323
rect -12255 -23357 -12216 -23323
rect -12328 -23395 -12216 -23357
rect -12328 -23429 -12289 -23395
rect -12255 -23429 -12216 -23395
rect -12328 -23467 -12216 -23429
rect -12328 -23501 -12289 -23467
rect -12255 -23501 -12216 -23467
rect -12328 -23539 -12216 -23501
rect -12328 -23573 -12289 -23539
rect -12255 -23573 -12216 -23539
rect -12328 -23611 -12216 -23573
rect -12328 -23645 -12289 -23611
rect -12255 -23645 -12216 -23611
rect -12328 -23683 -12216 -23645
rect -12328 -23717 -12289 -23683
rect -12255 -23717 -12216 -23683
rect -12328 -23755 -12216 -23717
rect -12328 -23789 -12289 -23755
rect -12255 -23789 -12216 -23755
rect -12328 -23827 -12216 -23789
rect -12328 -23861 -12289 -23827
rect -12255 -23861 -12216 -23827
rect -12328 -23899 -12216 -23861
rect -12328 -23933 -12289 -23899
rect -12255 -23933 -12216 -23899
rect -12328 -23971 -12216 -23933
rect -12328 -24005 -12289 -23971
rect -12255 -24005 -12216 -23971
rect -12328 -24043 -12216 -24005
rect -12328 -24077 -12289 -24043
rect -12255 -24077 -12216 -24043
rect -12328 -24115 -12216 -24077
rect -12328 -24149 -12289 -24115
rect -12255 -24149 -12216 -24115
rect -12328 -24187 -12216 -24149
rect -12328 -24221 -12289 -24187
rect -12255 -24221 -12216 -24187
rect -12328 -24259 -12216 -24221
rect -12328 -24293 -12289 -24259
rect -12255 -24293 -12216 -24259
rect -12328 -24331 -12216 -24293
rect -12328 -24365 -12289 -24331
rect -12255 -24365 -12216 -24331
rect -12328 -24403 -12216 -24365
rect -10662 -24380 -10602 -22314
rect -9504 -22570 -9444 -21250
rect -8486 -21196 -8426 -20786
rect -7986 -20988 -7914 -20984
rect -7986 -21040 -7976 -20988
rect -7924 -21040 -7914 -20988
rect -7986 -21044 -7914 -21040
rect -8486 -21248 -8482 -21196
rect -8430 -21248 -8426 -21196
rect -9012 -22254 -8952 -22010
rect -9018 -22258 -8946 -22254
rect -9018 -22310 -9008 -22258
rect -8956 -22310 -8946 -22258
rect -9018 -22314 -8946 -22310
rect -9012 -22450 -8952 -22314
rect -10520 -23206 -10460 -23040
rect -10028 -23206 -9968 -23120
rect -9500 -23206 -9440 -23044
rect -10520 -23266 -9440 -23206
rect -9500 -23306 -9440 -23266
rect -8486 -23202 -8426 -21248
rect -7980 -21340 -7920 -21044
rect -7468 -21088 -7408 -20804
rect -6954 -20988 -6882 -20984
rect -6954 -21040 -6944 -20988
rect -6892 -21040 -6882 -20988
rect -6954 -21044 -6882 -21040
rect -7474 -21092 -7402 -21088
rect -7474 -21144 -7464 -21092
rect -7412 -21144 -7402 -21092
rect -7474 -21148 -7402 -21144
rect -6948 -21336 -6888 -21044
rect -6450 -21196 -6390 -20788
rect -5948 -20984 -5888 -20902
rect -4928 -20984 -4868 -20902
rect -5954 -20988 -5882 -20984
rect -5954 -21040 -5944 -20988
rect -5892 -21040 -5882 -20988
rect -5954 -21044 -5882 -21040
rect -4934 -20988 -4862 -20984
rect -4934 -21040 -4924 -20988
rect -4872 -21040 -4862 -20988
rect -4934 -21044 -4862 -21040
rect -5438 -21092 -5366 -21088
rect -5438 -21144 -5428 -21092
rect -5376 -21144 -5366 -21092
rect -5438 -21148 -5366 -21144
rect -6450 -21248 -6446 -21196
rect -6394 -21248 -6390 -21196
rect -7474 -22134 -7414 -21924
rect -7480 -22138 -7408 -22134
rect -7480 -22190 -7470 -22138
rect -7418 -22190 -7408 -22138
rect -7480 -22194 -7408 -22190
rect -7474 -22568 -7414 -22194
rect -8486 -23254 -8482 -23202
rect -8430 -23254 -8426 -23202
rect -9506 -23310 -9434 -23306
rect -9506 -23362 -9496 -23310
rect -9444 -23362 -9434 -23310
rect -9506 -23366 -9434 -23362
rect -9012 -23422 -8940 -23418
rect -9012 -23474 -9002 -23422
rect -8950 -23474 -8940 -23422
rect -9012 -23478 -8940 -23474
rect -9006 -23558 -8946 -23478
rect -8486 -23712 -8426 -23254
rect -7982 -23418 -7922 -23122
rect -7470 -23310 -7398 -23306
rect -7470 -23362 -7460 -23310
rect -7408 -23362 -7398 -23310
rect -7470 -23366 -7398 -23362
rect -7988 -23422 -7916 -23418
rect -7988 -23474 -7978 -23422
rect -7926 -23474 -7916 -23422
rect -7988 -23478 -7916 -23474
rect -7464 -23650 -7404 -23366
rect -6950 -23418 -6890 -23126
rect -6450 -23202 -6390 -21248
rect -5942 -22254 -5882 -22012
rect -5948 -22258 -5876 -22254
rect -5948 -22310 -5938 -22258
rect -5886 -22310 -5876 -22258
rect -5948 -22314 -5876 -22310
rect -5942 -22448 -5882 -22314
rect -5432 -22604 -5372 -21148
rect -4418 -21192 -4358 -20778
rect -3914 -20988 -3842 -20984
rect -3914 -21040 -3904 -20988
rect -3852 -21040 -3842 -20988
rect -3914 -21044 -3842 -21040
rect -4424 -21196 -4352 -21192
rect -4424 -21248 -4414 -21196
rect -4362 -21248 -4352 -21196
rect -4424 -21252 -4352 -21248
rect -4934 -22254 -4874 -22010
rect -4940 -22258 -4868 -22254
rect -4940 -22310 -4930 -22258
rect -4878 -22310 -4868 -22258
rect -4940 -22314 -4868 -22310
rect -4934 -22448 -4874 -22314
rect -6450 -23254 -6446 -23202
rect -6394 -23254 -6390 -23202
rect -6956 -23422 -6884 -23418
rect -6956 -23474 -6946 -23422
rect -6894 -23474 -6884 -23422
rect -6956 -23478 -6884 -23474
rect -6450 -23648 -6390 -23254
rect -5428 -23306 -5368 -23012
rect -4418 -23202 -4358 -21252
rect -3908 -21330 -3848 -21044
rect -3398 -21088 -3338 -19808
rect -1374 -19898 -1302 -19894
rect -1374 -19950 -1364 -19898
rect -1312 -19950 -1302 -19898
rect -1374 -19954 -1302 -19950
rect 810 -19898 882 -19894
rect 810 -19950 820 -19898
rect 872 -19950 882 -19898
rect 810 -19954 882 -19950
rect -2902 -20026 -2830 -20022
rect -2902 -20078 -2892 -20026
rect -2840 -20078 -2830 -20026
rect -2902 -20082 -2830 -20078
rect -2896 -20232 -2836 -20082
rect -1368 -20306 -1308 -19954
rect -2898 -20988 -2838 -20978
rect -2898 -21040 -2894 -20988
rect -2842 -21040 -2838 -20988
rect -3404 -21092 -3332 -21088
rect -3404 -21144 -3394 -21092
rect -3342 -21144 -3332 -21092
rect -3404 -21148 -3332 -21144
rect -2898 -21340 -2838 -21040
rect -2384 -21196 -2324 -20788
rect -1884 -20984 -1824 -20900
rect -1890 -20988 -1818 -20984
rect -1890 -21040 -1880 -20988
rect -1828 -21040 -1818 -20988
rect -1890 -21044 -1818 -21040
rect -866 -20988 -806 -20902
rect -866 -21040 -862 -20988
rect -810 -21040 -806 -20988
rect -866 -21050 -806 -21040
rect -340 -21078 -280 -20816
rect 164 -21078 224 -20896
rect 676 -21078 736 -20796
rect -1368 -21092 -1296 -21088
rect -1368 -21144 -1358 -21092
rect -1306 -21144 -1296 -21092
rect -1368 -21148 -1296 -21144
rect -340 -21138 736 -21078
rect -2384 -21248 -2380 -21196
rect -2328 -21248 -2324 -21196
rect -3398 -22134 -3338 -21906
rect -3404 -22138 -3332 -22134
rect -3404 -22190 -3394 -22138
rect -3342 -22190 -3332 -22138
rect -3404 -22194 -3332 -22190
rect -3398 -22540 -3338 -22194
rect -4418 -23254 -4414 -23202
rect -4362 -23254 -4358 -23202
rect -5434 -23310 -5362 -23306
rect -5434 -23362 -5424 -23310
rect -5372 -23362 -5362 -23310
rect -5434 -23366 -5362 -23362
rect -5956 -23422 -5884 -23418
rect -5956 -23474 -5946 -23422
rect -5894 -23474 -5884 -23422
rect -5956 -23478 -5884 -23474
rect -4936 -23422 -4864 -23418
rect -4936 -23474 -4926 -23422
rect -4874 -23474 -4864 -23422
rect -4936 -23478 -4864 -23474
rect -5950 -23560 -5890 -23478
rect -4930 -23560 -4870 -23478
rect -4418 -23670 -4358 -23254
rect -3910 -23418 -3850 -23132
rect -3400 -23310 -3328 -23306
rect -3400 -23362 -3390 -23310
rect -3338 -23362 -3328 -23310
rect -3400 -23366 -3328 -23362
rect -3916 -23422 -3844 -23418
rect -3916 -23474 -3906 -23422
rect -3854 -23474 -3844 -23422
rect -3916 -23478 -3844 -23474
rect -3394 -23656 -3334 -23366
rect -2900 -23422 -2840 -23122
rect -2900 -23474 -2896 -23422
rect -2844 -23474 -2840 -23422
rect -2900 -23484 -2840 -23474
rect -2384 -23202 -2324 -21248
rect -1872 -22254 -1812 -22018
rect -1878 -22258 -1806 -22254
rect -1878 -22310 -1868 -22258
rect -1816 -22310 -1806 -22258
rect -1878 -22314 -1806 -22310
rect -1872 -22444 -1812 -22314
rect -1362 -22554 -1302 -21148
rect -340 -21196 -280 -21138
rect -340 -21248 -336 -21196
rect -284 -21248 -280 -21196
rect -846 -22254 -786 -22010
rect -340 -22198 -280 -21248
rect 164 -21332 224 -21138
rect 160 -22198 220 -22012
rect 676 -22198 736 -21138
rect 816 -22134 876 -19954
rect 930 -20988 1002 -20984
rect 930 -21040 940 -20988
rect 992 -21040 1002 -20988
rect 930 -21044 1002 -21040
rect 810 -22138 882 -22134
rect 810 -22190 820 -22138
rect 872 -22190 882 -22138
rect 810 -22194 882 -22190
rect -852 -22258 -780 -22254
rect -852 -22310 -842 -22258
rect -790 -22310 -780 -22258
rect -852 -22314 -780 -22310
rect -340 -22258 736 -22198
rect -846 -22450 -786 -22314
rect -2384 -23254 -2380 -23202
rect -2328 -23254 -2324 -23202
rect -2384 -23652 -2324 -23254
rect -1358 -23306 -1298 -23028
rect -340 -23198 -280 -22258
rect 160 -22452 220 -22258
rect -346 -23202 -274 -23198
rect -346 -23254 -336 -23202
rect -284 -23254 -274 -23202
rect -346 -23258 -274 -23254
rect -1364 -23310 -1292 -23306
rect -1364 -23362 -1354 -23310
rect -1302 -23362 -1292 -23310
rect -1364 -23366 -1292 -23362
rect -340 -23310 -280 -23258
rect 168 -23310 228 -23120
rect 676 -23310 736 -22258
rect -340 -23370 736 -23310
rect -1892 -23422 -1820 -23418
rect -1892 -23474 -1882 -23422
rect -1830 -23474 -1820 -23422
rect -1892 -23478 -1820 -23474
rect -868 -23422 -808 -23412
rect -868 -23474 -864 -23422
rect -812 -23474 -808 -23422
rect -1886 -23562 -1826 -23478
rect -868 -23560 -808 -23474
rect -340 -23674 -280 -23370
rect 168 -23560 228 -23370
rect 676 -23652 736 -23370
rect -10524 -24330 -10464 -24144
rect -10020 -24330 -9960 -24244
rect -9506 -24330 -9446 -24150
rect -12328 -24437 -12289 -24403
rect -12255 -24437 -12216 -24403
rect -12328 -24475 -12216 -24437
rect -10668 -24384 -10596 -24380
rect -10668 -24436 -10658 -24384
rect -10606 -24436 -10596 -24384
rect -10524 -24390 -9446 -24330
rect -7992 -24380 -7932 -24238
rect -6960 -24380 -6900 -24242
rect -10668 -24440 -10596 -24436
rect -12328 -24509 -12289 -24475
rect -12255 -24509 -12216 -24475
rect -12328 -24547 -12216 -24509
rect -12328 -24581 -12289 -24547
rect -12255 -24581 -12216 -24547
rect -9506 -24514 -9446 -24390
rect -7998 -24384 -7926 -24380
rect -7998 -24436 -7988 -24384
rect -7936 -24436 -7926 -24384
rect -7998 -24440 -7926 -24436
rect -6966 -24384 -6894 -24380
rect -6966 -24436 -6956 -24384
rect -6904 -24436 -6894 -24384
rect -6966 -24440 -6894 -24436
rect -5426 -24510 -5366 -24126
rect -3900 -24380 -3840 -24242
rect -2904 -24380 -2844 -24230
rect -3906 -24384 -3834 -24380
rect -3906 -24436 -3896 -24384
rect -3844 -24436 -3834 -24384
rect -3906 -24440 -3834 -24436
rect -2910 -24384 -2838 -24380
rect -2910 -24436 -2900 -24384
rect -2848 -24436 -2838 -24384
rect -2910 -24440 -2838 -24436
rect -1366 -24510 -1306 -24158
rect 816 -24510 876 -22194
rect 936 -23418 996 -21044
rect 930 -23422 1002 -23418
rect 930 -23474 940 -23422
rect 992 -23474 1002 -23422
rect 930 -23478 1002 -23474
rect -9506 -24566 -9502 -24514
rect -9450 -24566 -9446 -24514
rect -9506 -24576 -9446 -24566
rect -5432 -24514 -5360 -24510
rect -5432 -24566 -5422 -24514
rect -5370 -24566 -5360 -24514
rect -5432 -24570 -5360 -24566
rect -1372 -24514 -1300 -24510
rect -1372 -24566 -1362 -24514
rect -1310 -24566 -1300 -24514
rect -1372 -24570 -1300 -24566
rect 810 -24514 882 -24510
rect 810 -24566 820 -24514
rect 872 -24566 882 -24514
rect 810 -24570 882 -24566
rect -12328 -24619 -12216 -24581
rect -12328 -24653 -12289 -24619
rect -12255 -24653 -12216 -24619
rect -12328 -24691 -12216 -24653
rect -12328 -24725 -12289 -24691
rect -12255 -24725 -12216 -24691
rect -12328 -24763 -12216 -24725
rect -12328 -24797 -12289 -24763
rect -12255 -24797 -12216 -24763
rect -12328 -24835 -12216 -24797
rect -12328 -24869 -12289 -24835
rect -12255 -24869 -12216 -24835
rect -12328 -24907 -12216 -24869
rect -12328 -24941 -12289 -24907
rect -12255 -24941 -12216 -24907
rect -12328 -24979 -12216 -24941
rect -12328 -25013 -12289 -24979
rect -12255 -25013 -12216 -24979
rect -12328 -25051 -12216 -25013
rect -12328 -25085 -12289 -25051
rect -12255 -25085 -12216 -25051
rect -12328 -25123 -12216 -25085
rect -12328 -25157 -12289 -25123
rect -12255 -25157 -12216 -25123
rect -12328 -25195 -12216 -25157
rect -10064 -24976 172 -24916
rect -10064 -25186 -10004 -24976
rect -9564 -25098 -9504 -24976
rect -12328 -25229 -12289 -25195
rect -12255 -25229 -12216 -25195
rect -9042 -25196 -8982 -24976
rect -8544 -25098 -8484 -24976
rect -7510 -25104 -7450 -24976
rect -6488 -25104 -6428 -24976
rect -5498 -25104 -5438 -24976
rect -4974 -25194 -4914 -24976
rect -4464 -25110 -4404 -24976
rect -3474 -25098 -3414 -24976
rect -2442 -25110 -2382 -24976
rect -1438 -25098 -1378 -24976
rect -898 -25220 -838 -24976
rect -418 -25104 -358 -24976
rect 112 -25192 172 -24976
rect -12328 -25267 -12216 -25229
rect -12328 -25301 -12289 -25267
rect -12255 -25301 -12216 -25267
rect -12328 -25339 -12216 -25301
rect -12328 -25373 -12289 -25339
rect -12255 -25373 -12216 -25339
rect -12328 -25411 -12216 -25373
rect -12328 -25445 -12289 -25411
rect -12255 -25445 -12216 -25411
rect -12328 -25483 -12216 -25445
rect -12328 -25517 -12289 -25483
rect -12255 -25517 -12216 -25483
rect -12328 -25555 -12216 -25517
rect -12328 -25589 -12289 -25555
rect -12255 -25589 -12216 -25555
rect -12328 -25627 -12216 -25589
rect -12328 -25661 -12289 -25627
rect -12255 -25661 -12216 -25627
rect -12328 -25699 -12216 -25661
rect -12328 -25733 -12289 -25699
rect -12255 -25733 -12216 -25699
rect -12328 -25771 -12216 -25733
rect -12328 -25805 -12289 -25771
rect -12255 -25805 -12216 -25771
rect -12328 -25843 -12216 -25805
rect -12328 -25877 -12289 -25843
rect -12255 -25877 -12216 -25843
rect -8028 -25876 -7968 -25670
rect -12328 -25915 -12216 -25877
rect -12328 -25949 -12289 -25915
rect -12255 -25949 -12216 -25915
rect -8034 -25880 -7962 -25876
rect -8034 -25932 -8024 -25880
rect -7972 -25932 -7962 -25880
rect -8034 -25936 -7962 -25932
rect -12328 -25987 -12216 -25949
rect -12328 -26021 -12289 -25987
rect -12255 -26021 -12216 -25987
rect -12328 -26059 -12216 -26021
rect -12328 -26093 -12289 -26059
rect -12255 -26093 -12216 -26059
rect -12328 -26131 -12216 -26093
rect -12328 -26165 -12289 -26131
rect -12255 -26165 -12216 -26131
rect -12328 -26203 -12216 -26165
rect -12328 -26237 -12289 -26203
rect -12255 -26237 -12216 -26203
rect -12328 -26275 -12216 -26237
rect -12328 -26309 -12289 -26275
rect -12255 -26309 -12216 -26275
rect -12328 -26816 -12216 -26309
rect -8028 -26430 -7968 -25936
rect -7010 -25988 -6950 -25694
rect -5990 -25876 -5930 -25682
rect -3954 -25876 -3894 -25682
rect -5996 -25880 -5924 -25876
rect -5996 -25932 -5986 -25880
rect -5934 -25932 -5924 -25880
rect -5996 -25936 -5924 -25932
rect -3960 -25880 -3888 -25876
rect -3960 -25932 -3950 -25880
rect -3898 -25932 -3888 -25880
rect -3960 -25936 -3888 -25932
rect -7016 -25992 -6944 -25988
rect -7016 -26044 -7006 -25992
rect -6954 -26044 -6944 -25992
rect -7016 -26048 -6944 -26044
rect -5990 -26430 -5930 -25936
rect -3954 -26430 -3894 -25936
rect -2936 -25988 -2876 -25690
rect -1918 -25876 -1858 -25696
rect -1924 -25880 -1852 -25876
rect -1924 -25932 -1914 -25880
rect -1862 -25932 -1852 -25880
rect -1924 -25936 -1852 -25932
rect -2942 -25992 -2870 -25988
rect -2942 -26044 -2932 -25992
rect -2880 -26044 -2870 -25992
rect -2942 -26048 -2870 -26044
rect -1918 -26430 -1858 -25936
rect 1070 -25988 1130 -19060
rect 1282 -19894 1342 -11554
rect 1276 -19898 1348 -19894
rect 1276 -19950 1286 -19898
rect 1338 -19950 1348 -19898
rect 1276 -19954 1348 -19950
rect 1402 -20022 1462 -11552
rect 1396 -20026 1468 -20022
rect 1396 -20078 1406 -20026
rect 1458 -20078 1468 -20026
rect 1396 -20082 1468 -20078
rect 1542 -20984 1602 -11534
rect 1654 -11616 1726 -11612
rect 1654 -11668 1664 -11616
rect 1716 -11668 1726 -11616
rect 1654 -11672 1726 -11668
rect 1660 -17740 1720 -11672
rect 1770 -12354 1830 -11518
rect 1764 -12358 1836 -12354
rect 1764 -12410 1774 -12358
rect 1826 -12410 1836 -12358
rect 1764 -12414 1836 -12410
rect 1888 -15274 1948 -11414
rect 2216 -12220 2276 -11408
rect 2336 -11412 2340 -11360
rect 2392 -11412 2396 -11360
rect 2210 -12224 2282 -12220
rect 2210 -12276 2220 -12224
rect 2272 -12276 2282 -12224
rect 2210 -12280 2282 -12276
rect 2006 -13582 2078 -13578
rect 2006 -13634 2016 -13582
rect 2068 -13634 2078 -13582
rect 2006 -13638 2078 -13634
rect 1886 -15284 1948 -15274
rect 1886 -15336 1890 -15284
rect 1942 -15336 1948 -15284
rect 1886 -15346 1948 -15336
rect 1654 -17744 1726 -17740
rect 1654 -17796 1664 -17744
rect 1716 -17796 1726 -17744
rect 1654 -17800 1726 -17796
rect 1536 -20988 1608 -20984
rect 1536 -21040 1546 -20988
rect 1598 -21040 1608 -20988
rect 1536 -21044 1608 -21040
rect 1888 -21342 1948 -15346
rect 2012 -16274 2072 -13638
rect 2218 -13918 2290 -13914
rect 2218 -13970 2228 -13918
rect 2280 -13970 2290 -13918
rect 2218 -13974 2290 -13970
rect 2114 -15178 2186 -15174
rect 2114 -15230 2124 -15178
rect 2176 -15230 2186 -15178
rect 2114 -15234 2186 -15230
rect 2006 -16278 2078 -16274
rect 2006 -16330 2016 -16278
rect 2068 -16330 2078 -16278
rect 2006 -16334 2078 -16330
rect 2120 -21192 2180 -15234
rect 2224 -16510 2284 -13974
rect 2336 -16396 2396 -11412
rect 2442 -11496 2502 -11486
rect 2442 -11548 2446 -11496
rect 2498 -11548 2502 -11496
rect 2442 -14036 2502 -11548
rect 13248 -11846 13320 -11842
rect 13248 -11848 13258 -11846
rect 2568 -11898 13258 -11848
rect 13310 -11848 13320 -11846
rect 18352 -11846 18424 -11842
rect 18352 -11848 18362 -11846
rect 13310 -11898 18362 -11848
rect 18414 -11848 18424 -11846
rect 22418 -11848 22478 -11842
rect 18414 -11852 22990 -11848
rect 18414 -11898 22422 -11852
rect 2568 -11904 22422 -11898
rect 22474 -11904 22990 -11852
rect 2568 -11908 22990 -11904
rect 2568 -13914 2628 -11908
rect 3090 -11996 3150 -11908
rect 4100 -12010 4160 -11908
rect 3080 -12828 3140 -12672
rect 3586 -13580 3646 -12590
rect 4086 -12822 4146 -12666
rect 4606 -12924 4666 -11908
rect 5130 -11992 5190 -11908
rect 6142 -12010 6202 -11908
rect 5098 -12816 5158 -12660
rect 5620 -13580 5680 -12578
rect 6120 -12828 6180 -12672
rect 6638 -12928 6698 -11908
rect 7154 -11992 7214 -11908
rect 8154 -11998 8214 -11908
rect 7132 -12828 7192 -12672
rect 7656 -13580 7716 -12584
rect 8162 -12828 8222 -12672
rect 8676 -12908 8736 -11908
rect 9188 -12004 9248 -11908
rect 10200 -12004 10260 -11908
rect 9168 -12822 9228 -12666
rect 9694 -13580 9754 -12584
rect 10190 -12822 10250 -12666
rect 10712 -12916 10772 -11908
rect 11224 -12004 11284 -11908
rect 12236 -11992 12296 -11908
rect 11214 -12828 11274 -12672
rect 11732 -13580 11792 -12578
rect 12220 -12822 12280 -12666
rect 12744 -12914 12804 -11908
rect 13258 -11998 13318 -11908
rect 14270 -12010 14330 -11908
rect 13244 -12816 13304 -12660
rect 13766 -13580 13826 -12578
rect 14266 -12822 14326 -12666
rect 14782 -12916 14842 -11908
rect 15294 -12010 15354 -11908
rect 16312 -11998 16372 -11908
rect 15278 -12822 15338 -12666
rect 15802 -13580 15862 -12578
rect 16290 -12828 16350 -12672
rect 16818 -12890 16878 -11908
rect 17334 -11992 17394 -11908
rect 18358 -11992 18418 -11908
rect 17314 -12816 17374 -12660
rect 17840 -13580 17900 -12554
rect 18336 -12834 18396 -12678
rect 18854 -12908 18914 -11908
rect 19376 -11998 19436 -11908
rect 20388 -11998 20448 -11908
rect 19354 -12822 19414 -12666
rect 19874 -13580 19934 -12514
rect 20384 -12810 20444 -12654
rect 20892 -12908 20952 -11908
rect 21398 -11992 21458 -11908
rect 22416 -11914 22478 -11908
rect 22416 -12004 22476 -11914
rect 21396 -12810 21456 -12654
rect 21910 -13580 21970 -12564
rect 22396 -12828 22456 -12672
rect 22930 -12716 22990 -11908
rect 24816 -12091 24928 -11284
rect 24816 -12125 24855 -12091
rect 24889 -12125 24928 -12091
rect 24816 -12163 24928 -12125
rect 24816 -12197 24855 -12163
rect 24889 -12197 24928 -12163
rect 24816 -12235 24928 -12197
rect 24816 -12269 24855 -12235
rect 24889 -12269 24928 -12235
rect 24816 -12307 24928 -12269
rect 24816 -12341 24855 -12307
rect 24889 -12341 24928 -12307
rect 24816 -12379 24928 -12341
rect 24816 -12413 24855 -12379
rect 24889 -12413 24928 -12379
rect 24816 -12451 24928 -12413
rect 24816 -12485 24855 -12451
rect 24889 -12485 24928 -12451
rect 24816 -12523 24928 -12485
rect 24816 -12557 24855 -12523
rect 24889 -12557 24928 -12523
rect 24816 -12595 24928 -12557
rect 24816 -12629 24855 -12595
rect 24889 -12629 24928 -12595
rect 24816 -12667 24928 -12629
rect 24816 -12701 24855 -12667
rect 24889 -12701 24928 -12667
rect 22930 -12776 23710 -12716
rect 22930 -12916 22990 -12776
rect 3586 -13582 23588 -13580
rect 3586 -13634 3590 -13582
rect 3642 -13634 23588 -13582
rect 3586 -13640 23588 -13634
rect 3586 -13644 3646 -13640
rect 4594 -13798 4666 -13794
rect 4594 -13850 4604 -13798
rect 4656 -13850 4666 -13798
rect 4594 -13854 4666 -13850
rect 6634 -13798 6706 -13794
rect 6634 -13850 6644 -13798
rect 6696 -13850 6706 -13798
rect 6634 -13854 6706 -13850
rect 8674 -13798 8746 -13794
rect 8674 -13850 8684 -13798
rect 8736 -13850 8746 -13798
rect 8674 -13854 8746 -13850
rect 10704 -13798 10776 -13794
rect 10704 -13850 10714 -13798
rect 10766 -13850 10776 -13798
rect 10704 -13854 10776 -13850
rect 12744 -13798 12816 -13794
rect 12744 -13850 12754 -13798
rect 12806 -13850 12816 -13798
rect 12744 -13854 12816 -13850
rect 14776 -13798 14848 -13794
rect 14776 -13850 14786 -13798
rect 14838 -13850 14848 -13798
rect 14776 -13854 14848 -13850
rect 16816 -13798 16888 -13794
rect 16816 -13850 16826 -13798
rect 16878 -13850 16888 -13798
rect 16816 -13854 16888 -13850
rect 18852 -13798 18924 -13794
rect 18852 -13850 18862 -13798
rect 18914 -13850 18924 -13798
rect 18852 -13854 18924 -13850
rect 20886 -13798 20958 -13794
rect 20886 -13850 20896 -13798
rect 20948 -13850 20958 -13798
rect 20886 -13854 20958 -13850
rect 2562 -13918 2634 -13914
rect 2562 -13970 2572 -13918
rect 2624 -13970 2634 -13918
rect 2562 -13974 2634 -13970
rect 4086 -13924 4158 -13920
rect 4086 -13976 4096 -13924
rect 4148 -13976 4158 -13924
rect 4086 -13980 4158 -13976
rect 2436 -14040 2508 -14036
rect 2436 -14092 2446 -14040
rect 2498 -14092 2508 -14040
rect 2436 -14096 2508 -14092
rect 2442 -16170 2502 -14096
rect 2864 -14160 3076 -14154
rect 3136 -14160 3352 -14154
rect 4092 -14160 4152 -13980
rect 2864 -14194 2911 -14160
rect 2945 -14194 2983 -14160
rect 3017 -14194 3055 -14160
rect 3089 -14194 3127 -14160
rect 3161 -14194 3199 -14160
rect 3233 -14194 3271 -14160
rect 3305 -14194 3352 -14160
rect 3894 -14194 3929 -14160
rect 3963 -14194 4001 -14160
rect 4035 -14194 4073 -14160
rect 4107 -14194 4145 -14160
rect 4179 -14194 4217 -14160
rect 4251 -14194 4289 -14160
rect 4323 -14194 4358 -14160
rect 2864 -14200 3352 -14194
rect 4600 -14244 4660 -13854
rect 5106 -13924 5166 -13914
rect 5106 -13976 5110 -13924
rect 5162 -13976 5166 -13924
rect 5106 -14160 5166 -13976
rect 6128 -13924 6188 -13914
rect 6128 -13976 6132 -13924
rect 6184 -13976 6188 -13924
rect 6128 -14160 6188 -13976
rect 4912 -14194 4947 -14160
rect 4981 -14194 5019 -14160
rect 5053 -14194 5091 -14160
rect 5125 -14194 5163 -14160
rect 5197 -14194 5235 -14160
rect 5269 -14194 5307 -14160
rect 5341 -14194 5376 -14160
rect 5930 -14194 5965 -14160
rect 5999 -14194 6037 -14160
rect 6071 -14194 6109 -14160
rect 6143 -14194 6181 -14160
rect 6215 -14194 6253 -14160
rect 6287 -14194 6325 -14160
rect 6359 -14194 6394 -14160
rect 2568 -14263 2628 -14244
rect 2568 -14278 2582 -14263
rect 2576 -14297 2582 -14278
rect 2616 -14278 2628 -14263
rect 3586 -14263 3646 -14244
rect 2616 -14297 2622 -14278
rect 3586 -14292 3600 -14263
rect 2576 -14335 2622 -14297
rect 2576 -14369 2582 -14335
rect 2616 -14369 2622 -14335
rect 2576 -14407 2622 -14369
rect 2576 -14441 2582 -14407
rect 2616 -14441 2622 -14407
rect 2576 -14479 2622 -14441
rect 2576 -14513 2582 -14479
rect 2616 -14513 2622 -14479
rect 2576 -14551 2622 -14513
rect 2576 -14585 2582 -14551
rect 2616 -14585 2622 -14551
rect 2576 -14623 2622 -14585
rect 2576 -14657 2582 -14623
rect 2616 -14657 2622 -14623
rect 2576 -14695 2622 -14657
rect 2576 -14729 2582 -14695
rect 2616 -14729 2622 -14695
rect 2576 -14767 2622 -14729
rect 2576 -14770 2582 -14767
rect 2568 -14801 2582 -14770
rect 2616 -14770 2622 -14767
rect 3594 -14297 3600 -14292
rect 3634 -14292 3646 -14263
rect 4600 -14263 4664 -14244
rect 3634 -14297 3640 -14292
rect 3594 -14335 3640 -14297
rect 4600 -14297 4618 -14263
rect 4652 -14276 4664 -14263
rect 5630 -14263 5676 -14232
rect 4652 -14297 4660 -14276
rect 4600 -14312 4660 -14297
rect 5630 -14297 5636 -14263
rect 5670 -14297 5676 -14263
rect 3594 -14369 3600 -14335
rect 3634 -14369 3640 -14335
rect 3594 -14407 3640 -14369
rect 3594 -14441 3600 -14407
rect 3634 -14441 3640 -14407
rect 3594 -14479 3640 -14441
rect 3594 -14513 3600 -14479
rect 3634 -14513 3640 -14479
rect 3594 -14551 3640 -14513
rect 3594 -14585 3600 -14551
rect 3634 -14585 3640 -14551
rect 3594 -14623 3640 -14585
rect 3594 -14657 3600 -14623
rect 3634 -14657 3640 -14623
rect 3594 -14695 3640 -14657
rect 3594 -14729 3600 -14695
rect 3634 -14729 3640 -14695
rect 3594 -14767 3640 -14729
rect 4612 -14335 4658 -14312
rect 4612 -14369 4618 -14335
rect 4652 -14369 4658 -14335
rect 4612 -14407 4658 -14369
rect 4612 -14441 4618 -14407
rect 4652 -14441 4658 -14407
rect 4612 -14479 4658 -14441
rect 4612 -14513 4618 -14479
rect 4652 -14513 4658 -14479
rect 4612 -14551 4658 -14513
rect 4612 -14585 4618 -14551
rect 4652 -14585 4658 -14551
rect 4612 -14623 4658 -14585
rect 4612 -14657 4618 -14623
rect 4652 -14657 4658 -14623
rect 4612 -14695 4658 -14657
rect 4612 -14729 4618 -14695
rect 4652 -14729 4658 -14695
rect 4612 -14756 4658 -14729
rect 5630 -14335 5676 -14297
rect 6640 -14263 6700 -13854
rect 7142 -13924 7202 -13914
rect 7142 -13974 7146 -13924
rect 7140 -13976 7146 -13974
rect 7198 -13976 7202 -13924
rect 8168 -13924 8228 -13914
rect 8168 -13974 8172 -13924
rect 7140 -13986 7202 -13976
rect 8166 -13976 8172 -13974
rect 8224 -13976 8228 -13924
rect 8166 -13986 8228 -13976
rect 7140 -14160 7200 -13986
rect 7650 -14040 7722 -14036
rect 7650 -14092 7660 -14040
rect 7712 -14092 7722 -14040
rect 7650 -14096 7722 -14092
rect 6948 -14194 6983 -14160
rect 7017 -14194 7055 -14160
rect 7089 -14194 7127 -14160
rect 7161 -14194 7199 -14160
rect 7233 -14194 7271 -14160
rect 7305 -14194 7343 -14160
rect 7377 -14194 7412 -14160
rect 6640 -14297 6654 -14263
rect 6688 -14297 6700 -14263
rect 7656 -14263 7716 -14096
rect 8166 -14160 8226 -13986
rect 7966 -14194 8001 -14160
rect 8035 -14194 8073 -14160
rect 8107 -14194 8145 -14160
rect 8179 -14194 8217 -14160
rect 8251 -14194 8289 -14160
rect 8323 -14194 8361 -14160
rect 8395 -14194 8430 -14160
rect 7656 -14286 7672 -14263
rect 6640 -14298 6700 -14297
rect 7666 -14297 7672 -14286
rect 7706 -14286 7716 -14263
rect 8680 -14263 8740 -13854
rect 9180 -13924 9240 -13914
rect 9180 -13976 9184 -13924
rect 9236 -13976 9240 -13924
rect 9180 -14160 9240 -13976
rect 10216 -13924 10276 -13914
rect 10216 -13976 10220 -13924
rect 10272 -13976 10276 -13924
rect 10216 -14160 10276 -13976
rect 8984 -14194 9019 -14160
rect 9053 -14194 9091 -14160
rect 9125 -14194 9163 -14160
rect 9197 -14194 9235 -14160
rect 9269 -14194 9307 -14160
rect 9341 -14194 9379 -14160
rect 9413 -14194 9448 -14160
rect 10002 -14194 10037 -14160
rect 10071 -14194 10109 -14160
rect 10143 -14194 10181 -14160
rect 10215 -14194 10253 -14160
rect 10287 -14194 10325 -14160
rect 10359 -14194 10397 -14160
rect 10431 -14194 10466 -14160
rect 7706 -14297 7712 -14286
rect 5630 -14369 5636 -14335
rect 5670 -14369 5676 -14335
rect 5630 -14407 5676 -14369
rect 5630 -14441 5636 -14407
rect 5670 -14441 5676 -14407
rect 5630 -14479 5676 -14441
rect 5630 -14513 5636 -14479
rect 5670 -14513 5676 -14479
rect 5630 -14551 5676 -14513
rect 5630 -14585 5636 -14551
rect 5670 -14585 5676 -14551
rect 5630 -14623 5676 -14585
rect 5630 -14657 5636 -14623
rect 5670 -14657 5676 -14623
rect 5630 -14695 5676 -14657
rect 5630 -14729 5636 -14695
rect 5670 -14729 5676 -14695
rect 2616 -14801 2628 -14770
rect 3594 -14784 3600 -14767
rect 2568 -14958 2628 -14801
rect 3586 -14801 3600 -14784
rect 3634 -14784 3640 -14767
rect 4604 -14767 4664 -14756
rect 3634 -14801 3646 -14784
rect 2864 -14870 3352 -14864
rect 2864 -14904 2911 -14870
rect 2945 -14904 2983 -14870
rect 3017 -14904 3055 -14870
rect 3089 -14904 3127 -14870
rect 3161 -14904 3199 -14870
rect 3233 -14904 3271 -14870
rect 3305 -14904 3352 -14870
rect 2864 -14910 3352 -14904
rect 3070 -14958 3130 -14910
rect 3586 -14958 3646 -14801
rect 4604 -14801 4618 -14767
rect 4652 -14801 4664 -14767
rect 5630 -14767 5676 -14729
rect 6648 -14335 6694 -14298
rect 6648 -14369 6654 -14335
rect 6688 -14369 6694 -14335
rect 6648 -14407 6694 -14369
rect 6648 -14441 6654 -14407
rect 6688 -14441 6694 -14407
rect 6648 -14479 6694 -14441
rect 6648 -14513 6654 -14479
rect 6688 -14513 6694 -14479
rect 6648 -14551 6694 -14513
rect 6648 -14585 6654 -14551
rect 6688 -14585 6694 -14551
rect 6648 -14623 6694 -14585
rect 6648 -14657 6654 -14623
rect 6688 -14657 6694 -14623
rect 6648 -14695 6694 -14657
rect 6648 -14729 6654 -14695
rect 6688 -14729 6694 -14695
rect 6648 -14748 6694 -14729
rect 7666 -14335 7712 -14297
rect 8680 -14297 8690 -14263
rect 8724 -14297 8740 -14263
rect 9696 -14263 9756 -14244
rect 9696 -14294 9708 -14263
rect 8680 -14318 8740 -14297
rect 9702 -14297 9708 -14294
rect 9742 -14294 9756 -14263
rect 10710 -14263 10770 -13854
rect 11222 -13924 11282 -13914
rect 11222 -13976 11226 -13924
rect 11278 -13976 11282 -13924
rect 11222 -14160 11282 -13976
rect 12230 -13924 12302 -13920
rect 12230 -13976 12240 -13924
rect 12292 -13976 12302 -13924
rect 12230 -13980 12302 -13976
rect 12236 -14160 12296 -13980
rect 11020 -14194 11055 -14160
rect 11089 -14194 11127 -14160
rect 11161 -14194 11199 -14160
rect 11233 -14194 11271 -14160
rect 11305 -14194 11343 -14160
rect 11377 -14194 11415 -14160
rect 11449 -14194 11484 -14160
rect 12038 -14194 12073 -14160
rect 12107 -14194 12145 -14160
rect 12179 -14194 12217 -14160
rect 12251 -14194 12289 -14160
rect 12323 -14194 12361 -14160
rect 12395 -14194 12433 -14160
rect 12467 -14194 12502 -14160
rect 9742 -14297 9748 -14294
rect 7666 -14369 7672 -14335
rect 7706 -14369 7712 -14335
rect 7666 -14407 7712 -14369
rect 7666 -14441 7672 -14407
rect 7706 -14441 7712 -14407
rect 7666 -14479 7712 -14441
rect 7666 -14513 7672 -14479
rect 7706 -14513 7712 -14479
rect 7666 -14551 7712 -14513
rect 7666 -14585 7672 -14551
rect 7706 -14585 7712 -14551
rect 7666 -14623 7712 -14585
rect 7666 -14657 7672 -14623
rect 7706 -14657 7712 -14623
rect 7666 -14695 7712 -14657
rect 7666 -14729 7672 -14695
rect 7706 -14729 7712 -14695
rect 7666 -14744 7712 -14729
rect 8684 -14335 8730 -14318
rect 8684 -14369 8690 -14335
rect 8724 -14369 8730 -14335
rect 8684 -14407 8730 -14369
rect 8684 -14441 8690 -14407
rect 8724 -14441 8730 -14407
rect 8684 -14479 8730 -14441
rect 8684 -14513 8690 -14479
rect 8724 -14513 8730 -14479
rect 8684 -14551 8730 -14513
rect 8684 -14585 8690 -14551
rect 8724 -14585 8730 -14551
rect 8684 -14623 8730 -14585
rect 8684 -14657 8690 -14623
rect 8724 -14657 8730 -14623
rect 8684 -14695 8730 -14657
rect 8684 -14729 8690 -14695
rect 8724 -14729 8730 -14695
rect 5630 -14774 5636 -14767
rect 5626 -14792 5636 -14774
rect 3882 -14870 4370 -14864
rect 3882 -14904 3929 -14870
rect 3963 -14904 4001 -14870
rect 4035 -14904 4073 -14870
rect 4107 -14904 4145 -14870
rect 4179 -14904 4217 -14870
rect 4251 -14904 4289 -14870
rect 4323 -14904 4370 -14870
rect 3882 -14910 4370 -14904
rect 2568 -15018 3646 -14958
rect 3586 -15174 3646 -15018
rect 4096 -15068 4156 -14910
rect 4604 -14958 4664 -14801
rect 5624 -14801 5636 -14792
rect 5670 -14774 5676 -14767
rect 6644 -14767 6704 -14748
rect 6644 -14772 6654 -14767
rect 5670 -14801 5686 -14774
rect 5624 -14820 5686 -14801
rect 6642 -14801 6654 -14772
rect 6688 -14801 6704 -14767
rect 6642 -14820 6704 -14801
rect 7656 -14760 7716 -14744
rect 7656 -14767 7720 -14760
rect 8684 -14764 8730 -14729
rect 9702 -14335 9748 -14297
rect 10710 -14297 10726 -14263
rect 10760 -14297 10770 -14263
rect 10710 -14312 10770 -14297
rect 11744 -14263 11778 -14244
rect 9702 -14369 9708 -14335
rect 9742 -14369 9748 -14335
rect 9702 -14407 9748 -14369
rect 9702 -14441 9708 -14407
rect 9742 -14441 9748 -14407
rect 9702 -14479 9748 -14441
rect 9702 -14513 9708 -14479
rect 9742 -14513 9748 -14479
rect 9702 -14551 9748 -14513
rect 9702 -14585 9708 -14551
rect 9742 -14585 9748 -14551
rect 9702 -14623 9748 -14585
rect 9702 -14657 9708 -14623
rect 9742 -14657 9748 -14623
rect 9702 -14695 9748 -14657
rect 9702 -14729 9708 -14695
rect 9742 -14729 9748 -14695
rect 9702 -14756 9748 -14729
rect 10720 -14335 10766 -14312
rect 11744 -14320 11778 -14297
rect 12750 -14263 12810 -13854
rect 13252 -13924 13312 -13914
rect 13252 -13976 13256 -13924
rect 13308 -13976 13312 -13924
rect 13252 -14160 13312 -13976
rect 14260 -13924 14320 -13914
rect 14260 -13976 14264 -13924
rect 14316 -13974 14320 -13924
rect 14316 -13976 14322 -13974
rect 14260 -13986 14322 -13976
rect 14262 -14160 14322 -13986
rect 13056 -14194 13091 -14160
rect 13125 -14194 13163 -14160
rect 13197 -14194 13235 -14160
rect 13269 -14194 13307 -14160
rect 13341 -14194 13379 -14160
rect 13413 -14194 13451 -14160
rect 13485 -14194 13520 -14160
rect 14074 -14194 14109 -14160
rect 14143 -14194 14181 -14160
rect 14215 -14194 14253 -14160
rect 14287 -14194 14325 -14160
rect 14359 -14194 14397 -14160
rect 14431 -14194 14469 -14160
rect 14503 -14194 14538 -14160
rect 12750 -14297 12762 -14263
rect 12796 -14297 12810 -14263
rect 13764 -14263 13824 -14244
rect 13764 -14278 13780 -14263
rect 12750 -14312 12810 -14297
rect 13774 -14297 13780 -14278
rect 13814 -14278 13824 -14263
rect 14782 -14263 14842 -13854
rect 15276 -13924 15336 -13914
rect 15276 -13976 15280 -13924
rect 15332 -13974 15336 -13924
rect 16300 -13924 16360 -13914
rect 15332 -13976 15338 -13974
rect 15276 -13986 15338 -13976
rect 15278 -14160 15338 -13986
rect 16300 -13976 16304 -13924
rect 16356 -13976 16360 -13924
rect 16300 -14160 16360 -13976
rect 15092 -14194 15127 -14160
rect 15161 -14194 15199 -14160
rect 15233 -14194 15271 -14160
rect 15305 -14194 15343 -14160
rect 15377 -14194 15415 -14160
rect 15449 -14194 15487 -14160
rect 15521 -14194 15556 -14160
rect 16110 -14194 16145 -14160
rect 16179 -14194 16217 -14160
rect 16251 -14194 16289 -14160
rect 16323 -14194 16361 -14160
rect 16395 -14194 16433 -14160
rect 16467 -14194 16505 -14160
rect 16539 -14194 16574 -14160
rect 13814 -14297 13820 -14278
rect 10720 -14369 10726 -14335
rect 10760 -14369 10766 -14335
rect 10720 -14407 10766 -14369
rect 10720 -14441 10726 -14407
rect 10760 -14441 10766 -14407
rect 10720 -14479 10766 -14441
rect 10720 -14513 10726 -14479
rect 10760 -14513 10766 -14479
rect 10720 -14551 10766 -14513
rect 10720 -14585 10726 -14551
rect 10760 -14585 10766 -14551
rect 10720 -14623 10766 -14585
rect 10720 -14657 10726 -14623
rect 10760 -14657 10766 -14623
rect 10720 -14695 10766 -14657
rect 10720 -14729 10726 -14695
rect 10760 -14729 10766 -14695
rect 10720 -14744 10766 -14729
rect 11738 -14335 11784 -14320
rect 11738 -14369 11744 -14335
rect 11778 -14369 11784 -14335
rect 11738 -14407 11784 -14369
rect 11738 -14441 11744 -14407
rect 11778 -14441 11784 -14407
rect 11738 -14479 11784 -14441
rect 11738 -14513 11744 -14479
rect 11778 -14513 11784 -14479
rect 11738 -14551 11784 -14513
rect 11738 -14585 11744 -14551
rect 11778 -14585 11784 -14551
rect 11738 -14623 11784 -14585
rect 11738 -14657 11744 -14623
rect 11778 -14657 11784 -14623
rect 11738 -14695 11784 -14657
rect 11738 -14729 11744 -14695
rect 11778 -14729 11784 -14695
rect 7656 -14801 7672 -14767
rect 7706 -14801 7720 -14767
rect 7656 -14820 7720 -14801
rect 8676 -14767 8736 -14764
rect 8676 -14801 8690 -14767
rect 8724 -14801 8736 -14767
rect 9696 -14767 9756 -14756
rect 9696 -14784 9708 -14767
rect 4900 -14870 5388 -14864
rect 4900 -14904 4947 -14870
rect 4981 -14904 5019 -14870
rect 5053 -14904 5091 -14870
rect 5125 -14904 5163 -14870
rect 5197 -14904 5235 -14870
rect 5269 -14904 5307 -14870
rect 5341 -14904 5388 -14870
rect 4900 -14910 5388 -14904
rect 4598 -14962 4670 -14958
rect 4598 -15014 4608 -14962
rect 4660 -15014 4670 -14962
rect 4598 -15018 4670 -15014
rect 4090 -15072 4162 -15068
rect 4090 -15124 4100 -15072
rect 4152 -15124 4162 -15072
rect 4090 -15128 4162 -15124
rect 3580 -15178 3652 -15174
rect 3580 -15230 3590 -15178
rect 3642 -15230 3652 -15178
rect 3580 -15234 3652 -15230
rect 2566 -15284 2638 -15280
rect 2566 -15336 2576 -15284
rect 2628 -15336 2638 -15284
rect 2566 -15340 2638 -15336
rect 3064 -15284 3136 -15280
rect 3064 -15336 3074 -15284
rect 3126 -15336 3136 -15284
rect 3064 -15340 3136 -15336
rect 3576 -15284 3648 -15280
rect 3576 -15336 3586 -15284
rect 3638 -15336 3648 -15284
rect 3576 -15340 3648 -15336
rect 2572 -15495 2632 -15340
rect 3070 -15386 3130 -15340
rect 2864 -15392 3352 -15386
rect 2864 -15426 2911 -15392
rect 2945 -15426 2983 -15392
rect 3017 -15426 3055 -15392
rect 3089 -15426 3127 -15392
rect 3161 -15426 3199 -15392
rect 3233 -15426 3271 -15392
rect 3305 -15426 3352 -15392
rect 2864 -15432 3352 -15426
rect 2572 -15516 2582 -15495
rect 2576 -15529 2582 -15516
rect 2616 -15516 2632 -15495
rect 3582 -15495 3642 -15340
rect 4096 -15386 4156 -15128
rect 3882 -15392 4370 -15386
rect 3882 -15426 3929 -15392
rect 3963 -15426 4001 -15392
rect 4035 -15426 4073 -15392
rect 4107 -15426 4145 -15392
rect 4179 -15426 4217 -15392
rect 4251 -15426 4289 -15392
rect 4323 -15426 4370 -15392
rect 3882 -15432 4370 -15426
rect 2616 -15529 2622 -15516
rect 3582 -15522 3600 -15495
rect 2576 -15567 2622 -15529
rect 2576 -15601 2582 -15567
rect 2616 -15601 2622 -15567
rect 2576 -15639 2622 -15601
rect 2576 -15673 2582 -15639
rect 2616 -15673 2622 -15639
rect 2576 -15711 2622 -15673
rect 2576 -15745 2582 -15711
rect 2616 -15745 2622 -15711
rect 2576 -15783 2622 -15745
rect 2576 -15817 2582 -15783
rect 2616 -15817 2622 -15783
rect 2576 -15855 2622 -15817
rect 2576 -15889 2582 -15855
rect 2616 -15889 2622 -15855
rect 2576 -15927 2622 -15889
rect 2576 -15961 2582 -15927
rect 2616 -15961 2622 -15927
rect 2576 -15999 2622 -15961
rect 2576 -16033 2582 -15999
rect 2616 -16033 2622 -15999
rect 2576 -16064 2622 -16033
rect 3594 -15529 3600 -15522
rect 3634 -15522 3642 -15495
rect 4604 -15495 4664 -15018
rect 5118 -15068 5178 -14910
rect 5112 -15072 5184 -15068
rect 5112 -15124 5122 -15072
rect 5174 -15124 5184 -15072
rect 5112 -15128 5184 -15124
rect 5118 -15386 5178 -15128
rect 5626 -15174 5686 -14820
rect 5918 -14870 6406 -14864
rect 5918 -14904 5965 -14870
rect 5999 -14904 6037 -14870
rect 6071 -14904 6109 -14870
rect 6143 -14904 6181 -14870
rect 6215 -14904 6253 -14870
rect 6287 -14904 6325 -14870
rect 6359 -14904 6406 -14870
rect 5918 -14910 6272 -14904
rect 6332 -14910 6406 -14904
rect 6132 -15068 6192 -14910
rect 6644 -14958 6704 -14820
rect 6936 -14870 7424 -14864
rect 6936 -14904 6983 -14870
rect 7017 -14904 7055 -14870
rect 7089 -14904 7127 -14870
rect 7161 -14904 7199 -14870
rect 7233 -14904 7271 -14870
rect 7305 -14904 7343 -14870
rect 7377 -14904 7424 -14870
rect 6936 -14910 7144 -14904
rect 7146 -14910 7424 -14904
rect 7954 -14870 8442 -14864
rect 7954 -14904 8001 -14870
rect 8035 -14904 8073 -14870
rect 8107 -14904 8145 -14870
rect 8179 -14904 8217 -14870
rect 8251 -14904 8289 -14870
rect 8323 -14904 8361 -14870
rect 8395 -14904 8442 -14870
rect 7954 -14910 8224 -14904
rect 8244 -14910 8442 -14904
rect 6638 -14962 6710 -14958
rect 6638 -15014 6648 -14962
rect 6700 -15014 6710 -14962
rect 6638 -15018 6710 -15014
rect 6126 -15072 6198 -15068
rect 6126 -15124 6136 -15072
rect 6188 -15124 6198 -15072
rect 6126 -15128 6198 -15124
rect 5620 -15178 5692 -15174
rect 5620 -15230 5630 -15178
rect 5682 -15230 5692 -15178
rect 5620 -15234 5692 -15230
rect 6132 -15386 6192 -15128
rect 4900 -15392 5388 -15386
rect 4900 -15426 4947 -15392
rect 4981 -15426 5019 -15392
rect 5053 -15426 5091 -15392
rect 5125 -15426 5163 -15392
rect 5197 -15426 5235 -15392
rect 5269 -15426 5307 -15392
rect 5341 -15426 5388 -15392
rect 4900 -15432 5388 -15426
rect 5918 -15392 6192 -15386
rect 6196 -15392 6406 -15386
rect 5918 -15426 5965 -15392
rect 5999 -15426 6037 -15392
rect 6071 -15426 6109 -15392
rect 6143 -15426 6181 -15392
rect 6215 -15426 6253 -15392
rect 6287 -15426 6325 -15392
rect 6359 -15426 6406 -15392
rect 5918 -15432 6406 -15426
rect 6644 -15476 6704 -15018
rect 7146 -15068 7206 -14910
rect 8164 -15068 8224 -14910
rect 8676 -14958 8736 -14801
rect 9694 -14801 9708 -14784
rect 9742 -14801 9756 -14767
rect 9694 -14820 9756 -14801
rect 8972 -14870 9460 -14864
rect 8972 -14904 9019 -14870
rect 9053 -14904 9091 -14870
rect 9125 -14904 9163 -14870
rect 9197 -14904 9235 -14870
rect 9269 -14904 9307 -14870
rect 9341 -14904 9379 -14870
rect 9413 -14904 9460 -14870
rect 8972 -14910 9460 -14904
rect 8670 -14962 8742 -14958
rect 8670 -15014 8680 -14962
rect 8732 -15014 8742 -14962
rect 8670 -15018 8742 -15014
rect 7140 -15072 7212 -15068
rect 7140 -15124 7150 -15072
rect 7202 -15124 7212 -15072
rect 7140 -15128 7212 -15124
rect 8158 -15072 8230 -15068
rect 8158 -15124 8168 -15072
rect 8220 -15124 8230 -15072
rect 8158 -15128 8230 -15124
rect 7146 -15386 7206 -15128
rect 7650 -15178 7722 -15174
rect 7650 -15230 7660 -15178
rect 7712 -15230 7722 -15178
rect 7650 -15234 7722 -15230
rect 6936 -15392 7138 -15386
rect 7146 -15392 7424 -15386
rect 6936 -15426 6983 -15392
rect 7017 -15426 7055 -15392
rect 7089 -15426 7127 -15392
rect 7161 -15426 7199 -15392
rect 7233 -15426 7271 -15392
rect 7305 -15426 7343 -15392
rect 7377 -15426 7424 -15392
rect 6936 -15432 7424 -15426
rect 4604 -15514 4618 -15495
rect 3634 -15529 3640 -15522
rect 3594 -15567 3640 -15529
rect 3594 -15601 3600 -15567
rect 3634 -15601 3640 -15567
rect 3594 -15639 3640 -15601
rect 3594 -15673 3600 -15639
rect 3634 -15673 3640 -15639
rect 3594 -15711 3640 -15673
rect 3594 -15745 3600 -15711
rect 3634 -15745 3640 -15711
rect 3594 -15783 3640 -15745
rect 3594 -15817 3600 -15783
rect 3634 -15817 3640 -15783
rect 3594 -15855 3640 -15817
rect 3594 -15889 3600 -15855
rect 3634 -15889 3640 -15855
rect 3594 -15927 3640 -15889
rect 3594 -15961 3600 -15927
rect 3634 -15961 3640 -15927
rect 3594 -15999 3640 -15961
rect 4612 -15529 4618 -15514
rect 4652 -15514 4664 -15495
rect 5624 -15495 5684 -15476
rect 4652 -15529 4658 -15514
rect 5624 -15528 5636 -15495
rect 4612 -15567 4658 -15529
rect 4612 -15601 4618 -15567
rect 4652 -15601 4658 -15567
rect 4612 -15639 4658 -15601
rect 4612 -15673 4618 -15639
rect 4652 -15673 4658 -15639
rect 4612 -15711 4658 -15673
rect 4612 -15745 4618 -15711
rect 4652 -15745 4658 -15711
rect 4612 -15783 4658 -15745
rect 4612 -15817 4618 -15783
rect 4652 -15817 4658 -15783
rect 4612 -15855 4658 -15817
rect 4612 -15889 4618 -15855
rect 4652 -15889 4658 -15855
rect 4612 -15927 4658 -15889
rect 4612 -15961 4618 -15927
rect 4652 -15961 4658 -15927
rect 4612 -15994 4658 -15961
rect 3594 -16033 3600 -15999
rect 3634 -16033 3640 -15999
rect 3594 -16064 3640 -16033
rect 4598 -15999 4658 -15994
rect 4598 -16033 4618 -15999
rect 4652 -16033 4658 -15999
rect 5630 -15529 5636 -15528
rect 5670 -15528 5684 -15495
rect 6642 -15495 6704 -15476
rect 5670 -15529 5676 -15528
rect 5630 -15567 5676 -15529
rect 6642 -15529 6654 -15495
rect 6688 -15510 6704 -15495
rect 7656 -15476 7716 -15234
rect 8164 -15386 8224 -15128
rect 7954 -15392 8158 -15386
rect 8164 -15392 8442 -15386
rect 7954 -15426 8001 -15392
rect 8035 -15426 8073 -15392
rect 8107 -15426 8145 -15392
rect 8179 -15426 8217 -15392
rect 8251 -15426 8289 -15392
rect 8323 -15426 8361 -15392
rect 8395 -15426 8442 -15392
rect 7954 -15432 8442 -15426
rect 7656 -15495 7718 -15476
rect 6688 -15529 6702 -15510
rect 7656 -15520 7672 -15495
rect 6642 -15540 6702 -15529
rect 7666 -15529 7672 -15520
rect 7706 -15510 7718 -15495
rect 8676 -15495 8736 -15018
rect 9190 -15068 9250 -14910
rect 9696 -15028 9756 -14820
rect 10708 -14767 10768 -14744
rect 11738 -14758 11784 -14729
rect 12756 -14335 12802 -14312
rect 12756 -14369 12762 -14335
rect 12796 -14369 12802 -14335
rect 12756 -14407 12802 -14369
rect 12756 -14441 12762 -14407
rect 12796 -14441 12802 -14407
rect 12756 -14479 12802 -14441
rect 12756 -14513 12762 -14479
rect 12796 -14513 12802 -14479
rect 12756 -14551 12802 -14513
rect 12756 -14585 12762 -14551
rect 12796 -14585 12802 -14551
rect 12756 -14623 12802 -14585
rect 12756 -14657 12762 -14623
rect 12796 -14657 12802 -14623
rect 12756 -14695 12802 -14657
rect 12756 -14729 12762 -14695
rect 12796 -14729 12802 -14695
rect 12756 -14754 12802 -14729
rect 13774 -14335 13820 -14297
rect 14782 -14297 14798 -14263
rect 14832 -14297 14842 -14263
rect 15802 -14263 15862 -14244
rect 15802 -14284 15816 -14263
rect 14782 -14298 14842 -14297
rect 15810 -14297 15816 -14284
rect 15850 -14284 15862 -14263
rect 16822 -14263 16882 -13854
rect 17322 -13924 17382 -13914
rect 17322 -13976 17326 -13924
rect 17378 -13976 17382 -13924
rect 18344 -13924 18404 -13914
rect 18344 -13974 18348 -13924
rect 17322 -14160 17382 -13976
rect 18342 -13976 18348 -13974
rect 18400 -13976 18404 -13924
rect 18342 -13986 18404 -13976
rect 17838 -14040 17910 -14036
rect 17838 -14092 17848 -14040
rect 17900 -14092 17910 -14040
rect 17838 -14096 17910 -14092
rect 17128 -14194 17163 -14160
rect 17197 -14194 17235 -14160
rect 17269 -14194 17307 -14160
rect 17341 -14194 17379 -14160
rect 17413 -14194 17451 -14160
rect 17485 -14194 17523 -14160
rect 17557 -14194 17592 -14160
rect 15850 -14297 15856 -14284
rect 13774 -14369 13780 -14335
rect 13814 -14369 13820 -14335
rect 13774 -14407 13820 -14369
rect 13774 -14441 13780 -14407
rect 13814 -14441 13820 -14407
rect 13774 -14479 13820 -14441
rect 13774 -14513 13780 -14479
rect 13814 -14513 13820 -14479
rect 13774 -14551 13820 -14513
rect 13774 -14585 13780 -14551
rect 13814 -14585 13820 -14551
rect 13774 -14623 13820 -14585
rect 13774 -14657 13780 -14623
rect 13814 -14657 13820 -14623
rect 13774 -14695 13820 -14657
rect 13774 -14729 13780 -14695
rect 13814 -14729 13820 -14695
rect 11732 -14760 11792 -14758
rect 10708 -14801 10726 -14767
rect 10760 -14801 10768 -14767
rect 9990 -14870 10478 -14864
rect 9990 -14904 10037 -14870
rect 10071 -14904 10109 -14870
rect 10143 -14904 10181 -14870
rect 10215 -14904 10253 -14870
rect 10287 -14904 10325 -14870
rect 10359 -14904 10397 -14870
rect 10431 -14904 10478 -14870
rect 9990 -14910 10478 -14904
rect 9184 -15072 9256 -15068
rect 9184 -15124 9194 -15072
rect 9246 -15124 9256 -15072
rect 9696 -15088 9922 -15028
rect 10210 -15068 10270 -14910
rect 10708 -14958 10768 -14801
rect 11730 -14767 11792 -14760
rect 11730 -14801 11744 -14767
rect 11778 -14801 11792 -14767
rect 11730 -14820 11792 -14801
rect 12744 -14767 12804 -14754
rect 12744 -14801 12762 -14767
rect 12796 -14801 12804 -14767
rect 13774 -14767 13820 -14729
rect 14792 -14335 14838 -14298
rect 14792 -14369 14798 -14335
rect 14832 -14369 14838 -14335
rect 14792 -14407 14838 -14369
rect 14792 -14441 14798 -14407
rect 14832 -14441 14838 -14407
rect 14792 -14479 14838 -14441
rect 14792 -14513 14798 -14479
rect 14832 -14513 14838 -14479
rect 14792 -14551 14838 -14513
rect 14792 -14585 14798 -14551
rect 14832 -14585 14838 -14551
rect 14792 -14623 14838 -14585
rect 14792 -14657 14798 -14623
rect 14832 -14657 14838 -14623
rect 14792 -14695 14838 -14657
rect 14792 -14729 14798 -14695
rect 14832 -14729 14838 -14695
rect 14792 -14760 14838 -14729
rect 15810 -14335 15856 -14297
rect 16822 -14297 16834 -14263
rect 16868 -14297 16882 -14263
rect 16822 -14298 16882 -14297
rect 17844 -14263 17904 -14096
rect 18342 -14160 18402 -13986
rect 18146 -14194 18181 -14160
rect 18215 -14194 18253 -14160
rect 18287 -14194 18325 -14160
rect 18359 -14194 18397 -14160
rect 18431 -14194 18469 -14160
rect 18503 -14194 18541 -14160
rect 18575 -14194 18610 -14160
rect 17844 -14297 17852 -14263
rect 17886 -14297 17904 -14263
rect 15810 -14369 15816 -14335
rect 15850 -14369 15856 -14335
rect 15810 -14407 15856 -14369
rect 15810 -14441 15816 -14407
rect 15850 -14441 15856 -14407
rect 15810 -14479 15856 -14441
rect 15810 -14513 15816 -14479
rect 15850 -14513 15856 -14479
rect 15810 -14551 15856 -14513
rect 15810 -14585 15816 -14551
rect 15850 -14585 15856 -14551
rect 15810 -14623 15856 -14585
rect 15810 -14657 15816 -14623
rect 15850 -14657 15856 -14623
rect 15810 -14695 15856 -14657
rect 15810 -14729 15816 -14695
rect 15850 -14729 15856 -14695
rect 15810 -14754 15856 -14729
rect 16828 -14335 16874 -14298
rect 17844 -14308 17904 -14297
rect 18858 -14263 18918 -13854
rect 19362 -13924 19422 -13914
rect 19362 -13976 19366 -13924
rect 19418 -13974 19422 -13924
rect 20376 -13924 20436 -13914
rect 19418 -13976 19424 -13974
rect 19362 -13986 19424 -13976
rect 20376 -13976 20380 -13924
rect 20432 -13974 20436 -13924
rect 20432 -13976 20438 -13974
rect 20376 -13986 20438 -13976
rect 19364 -14160 19424 -13986
rect 20378 -14160 20438 -13986
rect 19164 -14194 19199 -14160
rect 19233 -14194 19271 -14160
rect 19305 -14194 19343 -14160
rect 19377 -14194 19415 -14160
rect 19449 -14194 19487 -14160
rect 19521 -14194 19559 -14160
rect 19593 -14194 19628 -14160
rect 20182 -14194 20217 -14160
rect 20251 -14194 20289 -14160
rect 20323 -14194 20361 -14160
rect 20395 -14194 20433 -14160
rect 20467 -14194 20505 -14160
rect 20539 -14194 20577 -14160
rect 20611 -14194 20646 -14160
rect 20892 -14244 20952 -13854
rect 21400 -13924 21460 -13914
rect 21400 -13974 21404 -13924
rect 21398 -13976 21404 -13974
rect 21456 -13976 21460 -13924
rect 21398 -13986 21460 -13976
rect 21398 -14160 21458 -13986
rect 21910 -14040 21982 -14036
rect 21910 -14092 21920 -14040
rect 21972 -14092 21982 -14040
rect 21910 -14096 21982 -14092
rect 23042 -14040 23114 -14036
rect 23042 -14092 23052 -14040
rect 23104 -14092 23114 -14040
rect 23042 -14096 23114 -14092
rect 21200 -14194 21235 -14160
rect 21269 -14194 21307 -14160
rect 21341 -14194 21379 -14160
rect 21413 -14194 21451 -14160
rect 21485 -14194 21523 -14160
rect 21557 -14194 21595 -14160
rect 21629 -14194 21664 -14160
rect 21916 -14244 21976 -14096
rect 22206 -14160 22420 -14154
rect 22490 -14160 22694 -14154
rect 22206 -14194 22253 -14160
rect 22287 -14194 22325 -14160
rect 22359 -14194 22397 -14160
rect 22431 -14194 22469 -14160
rect 22503 -14194 22541 -14160
rect 22575 -14194 22613 -14160
rect 22647 -14194 22694 -14160
rect 22206 -14200 22694 -14194
rect 18858 -14297 18870 -14263
rect 18904 -14297 18918 -14263
rect 19874 -14263 19934 -14244
rect 19874 -14284 19888 -14263
rect 18858 -14304 18918 -14297
rect 19882 -14297 19888 -14284
rect 19922 -14284 19934 -14263
rect 20892 -14263 20954 -14244
rect 19922 -14297 19928 -14284
rect 16828 -14369 16834 -14335
rect 16868 -14369 16874 -14335
rect 16828 -14407 16874 -14369
rect 16828 -14441 16834 -14407
rect 16868 -14441 16874 -14407
rect 16828 -14479 16874 -14441
rect 16828 -14513 16834 -14479
rect 16868 -14513 16874 -14479
rect 16828 -14551 16874 -14513
rect 16828 -14585 16834 -14551
rect 16868 -14585 16874 -14551
rect 16828 -14623 16874 -14585
rect 16828 -14657 16834 -14623
rect 16868 -14657 16874 -14623
rect 16828 -14695 16874 -14657
rect 16828 -14729 16834 -14695
rect 16868 -14729 16874 -14695
rect 13774 -14772 13780 -14767
rect 11008 -14870 11496 -14864
rect 11008 -14904 11055 -14870
rect 11089 -14904 11127 -14870
rect 11161 -14904 11199 -14870
rect 11233 -14904 11271 -14870
rect 11305 -14904 11343 -14870
rect 11377 -14904 11415 -14870
rect 11449 -14904 11496 -14870
rect 11008 -14910 11496 -14904
rect 10702 -14962 10774 -14958
rect 10702 -15014 10712 -14962
rect 10764 -15014 10774 -14962
rect 10702 -15018 10774 -15014
rect 9184 -15128 9256 -15124
rect 9190 -15386 9250 -15128
rect 9690 -15178 9762 -15174
rect 9690 -15230 9700 -15178
rect 9752 -15230 9762 -15178
rect 9690 -15234 9762 -15230
rect 8972 -15392 9460 -15386
rect 8972 -15426 9019 -15392
rect 9053 -15426 9091 -15392
rect 9125 -15426 9163 -15392
rect 9197 -15426 9235 -15392
rect 9269 -15426 9307 -15392
rect 9341 -15426 9379 -15392
rect 9413 -15426 9460 -15392
rect 8972 -15432 9460 -15426
rect 9696 -15476 9756 -15234
rect 9862 -15280 9922 -15088
rect 10204 -15072 10276 -15068
rect 10204 -15124 10214 -15072
rect 10266 -15124 10276 -15072
rect 10204 -15128 10276 -15124
rect 9856 -15284 9928 -15280
rect 9856 -15336 9866 -15284
rect 9918 -15336 9928 -15284
rect 9856 -15340 9928 -15336
rect 10210 -15386 10270 -15128
rect 9990 -15392 10478 -15386
rect 9990 -15426 10037 -15392
rect 10071 -15426 10109 -15392
rect 10143 -15426 10181 -15392
rect 10215 -15426 10253 -15392
rect 10287 -15426 10325 -15392
rect 10359 -15426 10397 -15392
rect 10431 -15426 10478 -15392
rect 9990 -15432 10478 -15426
rect 7706 -15520 7716 -15510
rect 8676 -15518 8690 -15495
rect 7706 -15529 7712 -15520
rect 5630 -15601 5636 -15567
rect 5670 -15601 5676 -15567
rect 5630 -15639 5676 -15601
rect 5630 -15673 5636 -15639
rect 5670 -15673 5676 -15639
rect 5630 -15711 5676 -15673
rect 5630 -15745 5636 -15711
rect 5670 -15745 5676 -15711
rect 5630 -15783 5676 -15745
rect 5630 -15817 5636 -15783
rect 5670 -15817 5676 -15783
rect 5630 -15855 5676 -15817
rect 5630 -15889 5636 -15855
rect 5670 -15889 5676 -15855
rect 5630 -15927 5676 -15889
rect 5630 -15961 5636 -15927
rect 5670 -15961 5676 -15927
rect 5630 -15999 5676 -15961
rect 6648 -15567 6694 -15540
rect 6648 -15601 6654 -15567
rect 6688 -15601 6694 -15567
rect 6648 -15639 6694 -15601
rect 6648 -15673 6654 -15639
rect 6688 -15673 6694 -15639
rect 6648 -15711 6694 -15673
rect 6648 -15745 6654 -15711
rect 6688 -15745 6694 -15711
rect 6648 -15783 6694 -15745
rect 6648 -15817 6654 -15783
rect 6688 -15817 6694 -15783
rect 6648 -15855 6694 -15817
rect 6648 -15889 6654 -15855
rect 6688 -15889 6694 -15855
rect 6648 -15927 6694 -15889
rect 6648 -15961 6654 -15927
rect 6688 -15961 6694 -15927
rect 6648 -15988 6694 -15961
rect 5630 -16032 5636 -15999
rect 2864 -16102 3352 -16096
rect 2864 -16136 2911 -16102
rect 2945 -16136 2983 -16102
rect 3017 -16136 3055 -16102
rect 3089 -16136 3127 -16102
rect 3161 -16136 3199 -16102
rect 3233 -16136 3271 -16102
rect 3305 -16136 3352 -16102
rect 2864 -16142 3352 -16136
rect 3882 -16102 4370 -16096
rect 3882 -16136 3929 -16102
rect 3963 -16136 4001 -16102
rect 4035 -16136 4073 -16102
rect 4107 -16136 4145 -16102
rect 4179 -16136 4217 -16102
rect 4251 -16136 4289 -16102
rect 4323 -16136 4370 -16102
rect 3882 -16142 4370 -16136
rect 2436 -16174 2508 -16170
rect 2436 -16226 2446 -16174
rect 2498 -16226 2508 -16174
rect 2436 -16230 2508 -16226
rect 4598 -16274 4658 -16033
rect 5620 -16033 5636 -16032
rect 5670 -16032 5676 -15999
rect 6634 -15999 6694 -15988
rect 5670 -16033 5680 -16032
rect 4900 -16102 5388 -16096
rect 4900 -16136 4947 -16102
rect 4981 -16136 5019 -16102
rect 5053 -16136 5091 -16102
rect 5125 -16136 5163 -16102
rect 5197 -16136 5235 -16102
rect 5269 -16136 5307 -16102
rect 5341 -16136 5388 -16102
rect 4900 -16142 5388 -16136
rect 2560 -16278 2632 -16274
rect 2560 -16330 2570 -16278
rect 2622 -16330 2632 -16278
rect 2560 -16334 2632 -16330
rect 4080 -16278 4152 -16274
rect 4080 -16330 4090 -16278
rect 4142 -16330 4152 -16278
rect 4080 -16334 4152 -16330
rect 4592 -16278 4664 -16274
rect 4592 -16330 4602 -16278
rect 4654 -16330 4664 -16278
rect 4592 -16334 4664 -16330
rect 2330 -16400 2402 -16396
rect 2330 -16452 2340 -16400
rect 2392 -16452 2402 -16400
rect 2330 -16456 2402 -16452
rect 2218 -16514 2290 -16510
rect 2218 -16566 2228 -16514
rect 2280 -16566 2290 -16514
rect 2218 -16570 2290 -16566
rect 2336 -17638 2396 -16456
rect 2566 -16729 2626 -16334
rect 3066 -16514 3138 -16510
rect 3066 -16566 3076 -16514
rect 3128 -16566 3138 -16514
rect 3066 -16570 3138 -16566
rect 3072 -16620 3132 -16570
rect 4086 -16620 4146 -16334
rect 4598 -16512 4670 -16508
rect 4598 -16564 4608 -16512
rect 4660 -16564 4670 -16512
rect 4598 -16568 4670 -16564
rect 2862 -16626 3132 -16620
rect 3136 -16626 3350 -16620
rect 2862 -16660 2909 -16626
rect 2943 -16660 2981 -16626
rect 3015 -16660 3053 -16626
rect 3087 -16660 3125 -16626
rect 3159 -16660 3197 -16626
rect 3231 -16660 3269 -16626
rect 3303 -16660 3350 -16626
rect 2862 -16666 3350 -16660
rect 3880 -16626 4368 -16620
rect 3880 -16660 3927 -16626
rect 3961 -16660 3999 -16626
rect 4033 -16660 4071 -16626
rect 4105 -16660 4143 -16626
rect 4177 -16660 4215 -16626
rect 4249 -16660 4287 -16626
rect 4321 -16660 4368 -16626
rect 3880 -16666 4368 -16660
rect 2566 -16763 2580 -16729
rect 2614 -16763 2626 -16729
rect 3586 -16729 3646 -16710
rect 3586 -16742 3598 -16729
rect 2566 -16766 2626 -16763
rect 3592 -16763 3598 -16742
rect 3632 -16742 3646 -16729
rect 4604 -16729 4664 -16568
rect 5102 -16620 5162 -16142
rect 5620 -16170 5680 -16033
rect 6634 -16033 6654 -15999
rect 6688 -16033 6694 -15999
rect 5918 -16102 6120 -16096
rect 6122 -16102 6406 -16096
rect 5918 -16136 5965 -16102
rect 5999 -16136 6037 -16102
rect 6071 -16136 6109 -16102
rect 6143 -16136 6181 -16102
rect 6215 -16136 6253 -16102
rect 6287 -16136 6325 -16102
rect 6359 -16136 6406 -16102
rect 5918 -16142 6120 -16136
rect 6122 -16142 6406 -16136
rect 5614 -16174 5686 -16170
rect 5614 -16226 5624 -16174
rect 5676 -16226 5686 -16174
rect 5614 -16230 5686 -16226
rect 5616 -16278 5688 -16274
rect 5616 -16330 5626 -16278
rect 5678 -16330 5688 -16278
rect 5616 -16334 5688 -16330
rect 4898 -16626 5386 -16620
rect 4898 -16660 4945 -16626
rect 4979 -16660 5017 -16626
rect 5051 -16660 5089 -16626
rect 5123 -16660 5161 -16626
rect 5195 -16660 5233 -16626
rect 5267 -16660 5305 -16626
rect 5339 -16660 5386 -16626
rect 4898 -16666 5386 -16660
rect 4604 -16736 4616 -16729
rect 3632 -16763 3638 -16742
rect 2580 -16798 2614 -16766
rect 2574 -16801 2620 -16798
rect 2574 -16835 2580 -16801
rect 2614 -16835 2620 -16801
rect 2574 -16873 2620 -16835
rect 2574 -16907 2580 -16873
rect 2614 -16907 2620 -16873
rect 2574 -16945 2620 -16907
rect 2574 -16979 2580 -16945
rect 2614 -16979 2620 -16945
rect 2574 -17017 2620 -16979
rect 2574 -17051 2580 -17017
rect 2614 -17051 2620 -17017
rect 2574 -17089 2620 -17051
rect 2574 -17123 2580 -17089
rect 2614 -17123 2620 -17089
rect 2574 -17161 2620 -17123
rect 2574 -17195 2580 -17161
rect 2614 -17195 2620 -17161
rect 2574 -17233 2620 -17195
rect 2574 -17267 2580 -17233
rect 2614 -17267 2620 -17233
rect 3592 -16801 3638 -16763
rect 3592 -16835 3598 -16801
rect 3632 -16835 3638 -16801
rect 3592 -16873 3638 -16835
rect 3592 -16907 3598 -16873
rect 3632 -16907 3638 -16873
rect 3592 -16945 3638 -16907
rect 3592 -16979 3598 -16945
rect 3632 -16979 3638 -16945
rect 3592 -17017 3638 -16979
rect 3592 -17051 3598 -17017
rect 3632 -17051 3638 -17017
rect 3592 -17089 3638 -17051
rect 3592 -17123 3598 -17089
rect 3632 -17123 3638 -17089
rect 3592 -17161 3638 -17123
rect 3592 -17195 3598 -17161
rect 3632 -17195 3638 -17161
rect 3592 -17233 3638 -17195
rect 3592 -17242 3598 -17233
rect 2574 -17298 2620 -17267
rect 3586 -17267 3598 -17242
rect 3632 -17242 3638 -17233
rect 4610 -16763 4616 -16736
rect 4650 -16736 4664 -16729
rect 5622 -16729 5682 -16334
rect 6122 -16620 6182 -16142
rect 6634 -16274 6694 -16033
rect 7666 -15567 7712 -15529
rect 7666 -15601 7672 -15567
rect 7706 -15601 7712 -15567
rect 7666 -15639 7712 -15601
rect 7666 -15673 7672 -15639
rect 7706 -15673 7712 -15639
rect 7666 -15711 7712 -15673
rect 7666 -15745 7672 -15711
rect 7706 -15745 7712 -15711
rect 7666 -15783 7712 -15745
rect 7666 -15817 7672 -15783
rect 7706 -15817 7712 -15783
rect 7666 -15855 7712 -15817
rect 7666 -15889 7672 -15855
rect 7706 -15889 7712 -15855
rect 7666 -15927 7712 -15889
rect 7666 -15961 7672 -15927
rect 7706 -15961 7712 -15927
rect 7666 -15999 7712 -15961
rect 7666 -16033 7672 -15999
rect 7706 -16033 7712 -15999
rect 8684 -15529 8690 -15518
rect 8724 -15518 8736 -15495
rect 9692 -15495 9756 -15476
rect 8724 -15529 8730 -15518
rect 8684 -15567 8730 -15529
rect 9692 -15529 9708 -15495
rect 9742 -15516 9756 -15495
rect 10708 -15495 10768 -15018
rect 11230 -15068 11290 -14910
rect 11224 -15072 11296 -15068
rect 11224 -15124 11234 -15072
rect 11286 -15124 11296 -15072
rect 11224 -15128 11296 -15124
rect 11230 -15386 11290 -15128
rect 11730 -15174 11790 -14820
rect 12026 -14870 12514 -14864
rect 12026 -14904 12073 -14870
rect 12107 -14904 12145 -14870
rect 12179 -14904 12217 -14870
rect 12251 -14904 12289 -14870
rect 12323 -14904 12361 -14870
rect 12395 -14904 12433 -14870
rect 12467 -14904 12514 -14870
rect 12026 -14910 12372 -14904
rect 12432 -14910 12514 -14904
rect 12232 -15068 12292 -14910
rect 12744 -14958 12804 -14801
rect 13766 -14801 13780 -14772
rect 13814 -14772 13820 -14767
rect 14780 -14767 14840 -14760
rect 13814 -14801 13826 -14772
rect 13044 -14870 13532 -14864
rect 13044 -14904 13091 -14870
rect 13125 -14904 13163 -14870
rect 13197 -14904 13235 -14870
rect 13269 -14904 13307 -14870
rect 13341 -14904 13379 -14870
rect 13413 -14904 13451 -14870
rect 13485 -14904 13532 -14870
rect 13044 -14910 13380 -14904
rect 13440 -14910 13532 -14904
rect 12738 -14962 12810 -14958
rect 12738 -15014 12748 -14962
rect 12800 -15014 12810 -14962
rect 12738 -15018 12810 -15014
rect 12226 -15072 12298 -15068
rect 12226 -15124 12236 -15072
rect 12288 -15124 12298 -15072
rect 12226 -15128 12298 -15124
rect 11724 -15178 11796 -15174
rect 11724 -15230 11734 -15178
rect 11786 -15230 11796 -15178
rect 11724 -15234 11796 -15230
rect 11724 -15284 11796 -15280
rect 11724 -15336 11734 -15284
rect 11786 -15336 11796 -15284
rect 11724 -15340 11796 -15336
rect 11008 -15392 11496 -15386
rect 11008 -15426 11055 -15392
rect 11089 -15426 11127 -15392
rect 11161 -15426 11199 -15392
rect 11233 -15426 11271 -15392
rect 11305 -15426 11343 -15392
rect 11377 -15426 11415 -15392
rect 11449 -15426 11496 -15392
rect 11008 -15432 11496 -15426
rect 11730 -15476 11790 -15340
rect 12232 -15386 12292 -15128
rect 12026 -15392 12514 -15386
rect 12026 -15426 12073 -15392
rect 12107 -15426 12145 -15392
rect 12179 -15426 12217 -15392
rect 12251 -15426 12289 -15392
rect 12323 -15426 12361 -15392
rect 12395 -15426 12433 -15392
rect 12467 -15426 12514 -15392
rect 12026 -15432 12514 -15426
rect 9742 -15529 9752 -15516
rect 9692 -15538 9752 -15529
rect 10708 -15529 10726 -15495
rect 10760 -15529 10768 -15495
rect 11728 -15495 11792 -15476
rect 11728 -15528 11744 -15495
rect 10708 -15532 10768 -15529
rect 11738 -15529 11744 -15528
rect 11778 -15520 11792 -15495
rect 12744 -15495 12804 -15018
rect 13258 -15068 13318 -14910
rect 13252 -15072 13324 -15068
rect 13252 -15124 13262 -15072
rect 13314 -15124 13324 -15072
rect 13252 -15128 13324 -15124
rect 13258 -15386 13318 -15128
rect 13766 -15174 13826 -14801
rect 14780 -14801 14798 -14767
rect 14832 -14801 14840 -14767
rect 15806 -14767 15866 -14754
rect 15806 -14780 15816 -14767
rect 14062 -14870 14422 -14864
rect 14482 -14870 14550 -14864
rect 14062 -14904 14109 -14870
rect 14143 -14904 14181 -14870
rect 14215 -14904 14253 -14870
rect 14287 -14904 14325 -14870
rect 14359 -14904 14397 -14870
rect 14431 -14904 14469 -14870
rect 14503 -14904 14550 -14870
rect 14062 -14910 14422 -14904
rect 14482 -14910 14550 -14904
rect 14276 -15068 14336 -14910
rect 14780 -14958 14840 -14801
rect 15804 -14801 15816 -14780
rect 15850 -14801 15866 -14767
rect 16828 -14767 16874 -14729
rect 17846 -14335 17892 -14308
rect 17846 -14369 17852 -14335
rect 17886 -14369 17892 -14335
rect 17846 -14407 17892 -14369
rect 17846 -14441 17852 -14407
rect 17886 -14441 17892 -14407
rect 17846 -14479 17892 -14441
rect 17846 -14513 17852 -14479
rect 17886 -14513 17892 -14479
rect 17846 -14551 17892 -14513
rect 17846 -14585 17852 -14551
rect 17886 -14585 17892 -14551
rect 17846 -14623 17892 -14585
rect 17846 -14657 17852 -14623
rect 17886 -14657 17892 -14623
rect 17846 -14695 17892 -14657
rect 17846 -14729 17852 -14695
rect 17886 -14729 17892 -14695
rect 17846 -14764 17892 -14729
rect 18864 -14335 18910 -14304
rect 18864 -14369 18870 -14335
rect 18904 -14369 18910 -14335
rect 18864 -14407 18910 -14369
rect 18864 -14441 18870 -14407
rect 18904 -14441 18910 -14407
rect 18864 -14479 18910 -14441
rect 18864 -14513 18870 -14479
rect 18904 -14513 18910 -14479
rect 18864 -14551 18910 -14513
rect 18864 -14585 18870 -14551
rect 18904 -14585 18910 -14551
rect 18864 -14623 18910 -14585
rect 18864 -14657 18870 -14623
rect 18904 -14657 18910 -14623
rect 18864 -14695 18910 -14657
rect 18864 -14729 18870 -14695
rect 18904 -14729 18910 -14695
rect 16828 -14770 16834 -14767
rect 15804 -14820 15866 -14801
rect 16818 -14801 16834 -14770
rect 16868 -14770 16874 -14767
rect 17838 -14766 17898 -14764
rect 17838 -14767 17900 -14766
rect 16868 -14801 16878 -14770
rect 15080 -14870 15568 -14864
rect 15080 -14904 15127 -14870
rect 15161 -14904 15199 -14870
rect 15233 -14904 15271 -14870
rect 15305 -14904 15343 -14870
rect 15377 -14904 15415 -14870
rect 15449 -14904 15487 -14870
rect 15521 -14904 15568 -14870
rect 15080 -14910 15568 -14904
rect 14774 -14962 14846 -14958
rect 14774 -15014 14784 -14962
rect 14836 -15014 14846 -14962
rect 14774 -15018 14846 -15014
rect 14270 -15072 14342 -15068
rect 14270 -15124 14280 -15072
rect 14332 -15124 14342 -15072
rect 14270 -15128 14342 -15124
rect 13760 -15178 13832 -15174
rect 13760 -15230 13770 -15178
rect 13822 -15230 13832 -15178
rect 13760 -15234 13832 -15230
rect 13762 -15284 13834 -15280
rect 13762 -15336 13772 -15284
rect 13824 -15336 13834 -15284
rect 13762 -15340 13834 -15336
rect 13044 -15392 13532 -15386
rect 13044 -15426 13091 -15392
rect 13125 -15426 13163 -15392
rect 13197 -15426 13235 -15392
rect 13269 -15426 13307 -15392
rect 13341 -15426 13379 -15392
rect 13413 -15426 13451 -15392
rect 13485 -15426 13532 -15392
rect 13044 -15432 13532 -15426
rect 13768 -15476 13828 -15340
rect 14276 -15386 14336 -15128
rect 14062 -15392 14550 -15386
rect 14062 -15426 14109 -15392
rect 14143 -15426 14181 -15392
rect 14215 -15426 14253 -15392
rect 14287 -15426 14325 -15392
rect 14359 -15426 14397 -15392
rect 14431 -15426 14469 -15392
rect 14503 -15426 14550 -15392
rect 14062 -15432 14550 -15426
rect 11778 -15528 11788 -15520
rect 12744 -15524 12762 -15495
rect 11778 -15529 11784 -15528
rect 8684 -15601 8690 -15567
rect 8724 -15601 8730 -15567
rect 8684 -15639 8730 -15601
rect 8684 -15673 8690 -15639
rect 8724 -15673 8730 -15639
rect 8684 -15711 8730 -15673
rect 8684 -15745 8690 -15711
rect 8724 -15745 8730 -15711
rect 8684 -15783 8730 -15745
rect 8684 -15817 8690 -15783
rect 8724 -15817 8730 -15783
rect 8684 -15855 8730 -15817
rect 8684 -15889 8690 -15855
rect 8724 -15889 8730 -15855
rect 8684 -15927 8730 -15889
rect 8684 -15961 8690 -15927
rect 8724 -15961 8730 -15927
rect 8684 -15999 8730 -15961
rect 8684 -16010 8690 -15999
rect 7666 -16064 7712 -16033
rect 8676 -16033 8690 -16010
rect 8724 -16010 8730 -15999
rect 9702 -15567 9748 -15538
rect 9702 -15601 9708 -15567
rect 9742 -15601 9748 -15567
rect 9702 -15639 9748 -15601
rect 9702 -15673 9708 -15639
rect 9742 -15673 9748 -15639
rect 9702 -15711 9748 -15673
rect 9702 -15745 9708 -15711
rect 9742 -15745 9748 -15711
rect 9702 -15783 9748 -15745
rect 9702 -15817 9708 -15783
rect 9742 -15817 9748 -15783
rect 9702 -15855 9748 -15817
rect 9702 -15889 9708 -15855
rect 9742 -15889 9748 -15855
rect 9702 -15927 9748 -15889
rect 9702 -15961 9708 -15927
rect 9742 -15961 9748 -15927
rect 9702 -15999 9748 -15961
rect 8724 -16033 8736 -16010
rect 8676 -16052 8736 -16033
rect 9702 -16033 9708 -15999
rect 9742 -16033 9748 -15999
rect 10720 -15567 10766 -15532
rect 10720 -15601 10726 -15567
rect 10760 -15601 10766 -15567
rect 10720 -15639 10766 -15601
rect 10720 -15673 10726 -15639
rect 10760 -15673 10766 -15639
rect 10720 -15711 10766 -15673
rect 10720 -15745 10726 -15711
rect 10760 -15745 10766 -15711
rect 10720 -15783 10766 -15745
rect 10720 -15817 10726 -15783
rect 10760 -15817 10766 -15783
rect 10720 -15855 10766 -15817
rect 10720 -15889 10726 -15855
rect 10760 -15889 10766 -15855
rect 10720 -15927 10766 -15889
rect 10720 -15961 10726 -15927
rect 10760 -15961 10766 -15927
rect 11738 -15567 11784 -15529
rect 11738 -15601 11744 -15567
rect 11778 -15601 11784 -15567
rect 11738 -15639 11784 -15601
rect 11738 -15673 11744 -15639
rect 11778 -15673 11784 -15639
rect 11738 -15711 11784 -15673
rect 11738 -15745 11744 -15711
rect 11778 -15745 11784 -15711
rect 11738 -15783 11784 -15745
rect 11738 -15817 11744 -15783
rect 11778 -15817 11784 -15783
rect 11738 -15855 11784 -15817
rect 11738 -15889 11744 -15855
rect 11778 -15889 11784 -15855
rect 11738 -15927 11784 -15889
rect 11738 -15928 11744 -15927
rect 10720 -15999 10766 -15961
rect 10720 -16010 10726 -15999
rect 9702 -16064 9748 -16033
rect 10712 -16033 10726 -16010
rect 10760 -16010 10766 -15999
rect 11778 -15928 11784 -15927
rect 12756 -15529 12762 -15524
rect 12796 -15524 12804 -15495
rect 13764 -15495 13830 -15476
rect 13764 -15516 13780 -15495
rect 12796 -15529 12802 -15524
rect 12756 -15567 12802 -15529
rect 12756 -15601 12762 -15567
rect 12796 -15601 12802 -15567
rect 12756 -15639 12802 -15601
rect 12756 -15673 12762 -15639
rect 12796 -15673 12802 -15639
rect 12756 -15711 12802 -15673
rect 12756 -15745 12762 -15711
rect 12796 -15745 12802 -15711
rect 12756 -15783 12802 -15745
rect 12756 -15817 12762 -15783
rect 12796 -15817 12802 -15783
rect 12756 -15855 12802 -15817
rect 12756 -15889 12762 -15855
rect 12796 -15889 12802 -15855
rect 12756 -15927 12802 -15889
rect 11744 -15999 11778 -15961
rect 10760 -16033 10772 -16010
rect 6936 -16102 7424 -16096
rect 6936 -16136 6983 -16102
rect 7017 -16136 7055 -16102
rect 7089 -16136 7127 -16102
rect 7161 -16136 7199 -16102
rect 7233 -16136 7271 -16102
rect 7305 -16136 7343 -16102
rect 7377 -16136 7424 -16102
rect 6936 -16142 7132 -16136
rect 7134 -16142 7424 -16136
rect 7954 -16102 8442 -16096
rect 7954 -16136 8001 -16102
rect 8035 -16136 8073 -16102
rect 8107 -16136 8145 -16102
rect 8179 -16136 8217 -16102
rect 8251 -16136 8289 -16102
rect 8323 -16136 8361 -16102
rect 8395 -16136 8442 -16102
rect 7954 -16142 8442 -16136
rect 8972 -16102 9460 -16096
rect 8972 -16136 9019 -16102
rect 9053 -16136 9091 -16102
rect 9125 -16136 9163 -16102
rect 9197 -16136 9235 -16102
rect 9269 -16136 9307 -16102
rect 9341 -16136 9379 -16102
rect 9413 -16136 9460 -16102
rect 8972 -16142 9460 -16136
rect 9990 -16102 10478 -16096
rect 9990 -16136 10037 -16102
rect 10071 -16136 10109 -16102
rect 10143 -16136 10181 -16102
rect 10215 -16136 10253 -16102
rect 10287 -16136 10325 -16102
rect 10359 -16136 10397 -16102
rect 10431 -16136 10478 -16102
rect 9990 -16142 10478 -16136
rect 6628 -16278 6700 -16274
rect 6628 -16330 6638 -16278
rect 6690 -16330 6700 -16278
rect 6628 -16334 6700 -16330
rect 6634 -16512 6706 -16508
rect 6634 -16564 6644 -16512
rect 6696 -16564 6706 -16512
rect 6634 -16568 6706 -16564
rect 5916 -16626 6120 -16620
rect 6122 -16626 6404 -16620
rect 5916 -16660 5963 -16626
rect 5997 -16660 6035 -16626
rect 6069 -16660 6107 -16626
rect 6141 -16660 6179 -16626
rect 6213 -16660 6251 -16626
rect 6285 -16660 6323 -16626
rect 6357 -16660 6404 -16626
rect 5916 -16666 6404 -16660
rect 4650 -16763 4656 -16736
rect 5622 -16742 5634 -16729
rect 4610 -16801 4656 -16763
rect 4610 -16835 4616 -16801
rect 4650 -16835 4656 -16801
rect 4610 -16873 4656 -16835
rect 4610 -16907 4616 -16873
rect 4650 -16907 4656 -16873
rect 4610 -16945 4656 -16907
rect 4610 -16979 4616 -16945
rect 4650 -16979 4656 -16945
rect 4610 -17017 4656 -16979
rect 4610 -17051 4616 -17017
rect 4650 -17051 4656 -17017
rect 4610 -17089 4656 -17051
rect 4610 -17123 4616 -17089
rect 4650 -17123 4656 -17089
rect 4610 -17161 4656 -17123
rect 4610 -17195 4616 -17161
rect 4650 -17195 4656 -17161
rect 4610 -17233 4656 -17195
rect 3632 -17267 3646 -17242
rect 2862 -17336 3350 -17330
rect 2862 -17370 2909 -17336
rect 2943 -17370 2981 -17336
rect 3015 -17370 3053 -17336
rect 3087 -17370 3125 -17336
rect 3159 -17370 3197 -17336
rect 3231 -17370 3269 -17336
rect 3303 -17370 3350 -17336
rect 2862 -17376 3350 -17370
rect 3586 -17438 3646 -17267
rect 4610 -17267 4616 -17233
rect 4650 -17267 4656 -17233
rect 5628 -16763 5634 -16742
rect 5668 -16742 5682 -16729
rect 6640 -16729 6700 -16568
rect 7134 -16620 7194 -16142
rect 7648 -16278 7720 -16274
rect 7648 -16330 7658 -16278
rect 7710 -16330 7720 -16278
rect 7648 -16334 7720 -16330
rect 6934 -16626 7132 -16620
rect 7134 -16626 7422 -16620
rect 6934 -16660 6981 -16626
rect 7015 -16660 7053 -16626
rect 7087 -16660 7125 -16626
rect 7159 -16660 7197 -16626
rect 7231 -16660 7269 -16626
rect 7303 -16660 7341 -16626
rect 7375 -16660 7422 -16626
rect 6934 -16666 7422 -16660
rect 6640 -16740 6652 -16729
rect 5668 -16763 5674 -16742
rect 5628 -16801 5674 -16763
rect 5628 -16835 5634 -16801
rect 5668 -16835 5674 -16801
rect 5628 -16873 5674 -16835
rect 5628 -16907 5634 -16873
rect 5668 -16907 5674 -16873
rect 5628 -16945 5674 -16907
rect 5628 -16979 5634 -16945
rect 5668 -16979 5674 -16945
rect 5628 -17017 5674 -16979
rect 5628 -17051 5634 -17017
rect 5668 -17051 5674 -17017
rect 5628 -17089 5674 -17051
rect 5628 -17123 5634 -17089
rect 5668 -17123 5674 -17089
rect 5628 -17161 5674 -17123
rect 5628 -17195 5634 -17161
rect 5668 -17195 5674 -17161
rect 5628 -17233 5674 -17195
rect 5628 -17246 5634 -17233
rect 4610 -17298 4656 -17267
rect 5620 -17267 5634 -17246
rect 5668 -17246 5674 -17233
rect 6646 -16763 6652 -16740
rect 6686 -16740 6700 -16729
rect 7654 -16729 7714 -16334
rect 8160 -16620 8220 -16142
rect 8670 -16174 8742 -16170
rect 8670 -16226 8680 -16174
rect 8732 -16226 8742 -16174
rect 8670 -16230 8742 -16226
rect 7952 -16626 8440 -16620
rect 7952 -16660 7999 -16626
rect 8033 -16660 8071 -16626
rect 8105 -16660 8143 -16626
rect 8177 -16660 8215 -16626
rect 8249 -16660 8287 -16626
rect 8321 -16660 8359 -16626
rect 8393 -16660 8440 -16626
rect 7952 -16666 8440 -16660
rect 6686 -16763 6692 -16740
rect 7654 -16754 7670 -16729
rect 6646 -16801 6692 -16763
rect 6646 -16835 6652 -16801
rect 6686 -16835 6692 -16801
rect 6646 -16873 6692 -16835
rect 6646 -16907 6652 -16873
rect 6686 -16907 6692 -16873
rect 6646 -16945 6692 -16907
rect 6646 -16979 6652 -16945
rect 6686 -16979 6692 -16945
rect 6646 -17017 6692 -16979
rect 6646 -17051 6652 -17017
rect 6686 -17051 6692 -17017
rect 6646 -17089 6692 -17051
rect 6646 -17123 6652 -17089
rect 6686 -17123 6692 -17089
rect 6646 -17161 6692 -17123
rect 6646 -17195 6652 -17161
rect 6686 -17195 6692 -17161
rect 6646 -17233 6692 -17195
rect 5668 -17267 5680 -17246
rect 3880 -17336 4368 -17330
rect 3880 -17370 3927 -17336
rect 3961 -17370 3999 -17336
rect 4033 -17370 4071 -17336
rect 4105 -17370 4143 -17336
rect 4177 -17370 4215 -17336
rect 4249 -17370 4287 -17336
rect 4321 -17370 4368 -17336
rect 3880 -17376 4368 -17370
rect 4898 -17336 5386 -17330
rect 4898 -17370 4945 -17336
rect 4979 -17370 5017 -17336
rect 5051 -17370 5089 -17336
rect 5123 -17370 5161 -17336
rect 5195 -17370 5233 -17336
rect 5267 -17370 5305 -17336
rect 5339 -17370 5386 -17336
rect 4898 -17376 5386 -17370
rect 2442 -17442 2514 -17438
rect 2442 -17494 2452 -17442
rect 2504 -17494 2514 -17442
rect 2442 -17498 2514 -17494
rect 3580 -17442 3652 -17438
rect 3580 -17494 3590 -17442
rect 3642 -17494 3652 -17442
rect 3580 -17498 3652 -17494
rect 2330 -17642 2402 -17638
rect 2330 -17694 2340 -17642
rect 2392 -17694 2402 -17642
rect 2330 -17698 2402 -17694
rect 2224 -17744 2296 -17740
rect 2224 -17796 2234 -17744
rect 2286 -17796 2296 -17744
rect 2224 -17800 2296 -17796
rect 2114 -21196 2186 -21192
rect 2114 -21248 2124 -21196
rect 2176 -21248 2186 -21196
rect 2230 -21230 2290 -17800
rect 2336 -18874 2396 -17698
rect 2330 -18878 2402 -18874
rect 2330 -18930 2340 -18878
rect 2392 -18930 2402 -18878
rect 2330 -18934 2402 -18930
rect 2114 -21252 2186 -21248
rect 2224 -21234 2296 -21230
rect 1882 -21346 1954 -21342
rect 1882 -21398 1892 -21346
rect 1944 -21398 1954 -21346
rect 1882 -21402 1954 -21398
rect 2120 -24928 2180 -21252
rect 2224 -21286 2234 -21234
rect 2286 -21286 2296 -21234
rect 2224 -21290 2296 -21286
rect 2230 -23720 2290 -21290
rect 2336 -23594 2396 -18934
rect 2448 -20212 2508 -17498
rect 3578 -17642 3650 -17638
rect 3578 -17694 3588 -17642
rect 3640 -17694 3650 -17642
rect 3578 -17698 3650 -17694
rect 3584 -17742 3644 -17698
rect 2568 -17802 3644 -17742
rect 2568 -17804 3132 -17802
rect 2568 -17963 2628 -17804
rect 3072 -17854 3132 -17804
rect 2862 -17860 3350 -17854
rect 2862 -17894 2909 -17860
rect 2943 -17894 2981 -17860
rect 3015 -17894 3053 -17860
rect 3087 -17894 3125 -17860
rect 3159 -17894 3197 -17860
rect 3231 -17894 3269 -17860
rect 3303 -17894 3350 -17860
rect 2862 -17900 3350 -17894
rect 2568 -17976 2580 -17963
rect 2574 -17997 2580 -17976
rect 2614 -17976 2628 -17963
rect 3584 -17963 3644 -17802
rect 4088 -17854 4148 -17376
rect 4596 -17522 4668 -17518
rect 4596 -17574 4606 -17522
rect 4658 -17574 4668 -17522
rect 4596 -17578 4668 -17574
rect 3880 -17860 4368 -17854
rect 3880 -17894 3927 -17860
rect 3961 -17894 3999 -17860
rect 4033 -17894 4071 -17860
rect 4105 -17894 4143 -17860
rect 4177 -17894 4215 -17860
rect 4249 -17894 4287 -17860
rect 4321 -17894 4368 -17860
rect 3880 -17900 4368 -17894
rect 2614 -17997 2620 -17976
rect 3584 -17980 3598 -17963
rect 2574 -18035 2620 -17997
rect 2574 -18069 2580 -18035
rect 2614 -18069 2620 -18035
rect 2574 -18107 2620 -18069
rect 2574 -18141 2580 -18107
rect 2614 -18141 2620 -18107
rect 2574 -18179 2620 -18141
rect 2574 -18213 2580 -18179
rect 2614 -18213 2620 -18179
rect 2574 -18251 2620 -18213
rect 2574 -18285 2580 -18251
rect 2614 -18285 2620 -18251
rect 2574 -18323 2620 -18285
rect 2574 -18357 2580 -18323
rect 2614 -18357 2620 -18323
rect 2574 -18395 2620 -18357
rect 2574 -18429 2580 -18395
rect 2614 -18429 2620 -18395
rect 2574 -18467 2620 -18429
rect 2574 -18501 2580 -18467
rect 2614 -18501 2620 -18467
rect 2574 -18532 2620 -18501
rect 3592 -17997 3598 -17980
rect 3632 -17980 3644 -17963
rect 4602 -17963 4662 -17578
rect 5116 -17632 5176 -17376
rect 5620 -17414 5680 -17267
rect 6646 -17267 6652 -17233
rect 6686 -17267 6692 -17233
rect 7664 -16763 7670 -16754
rect 7704 -16754 7714 -16729
rect 8676 -16729 8736 -16230
rect 10712 -16274 10772 -16033
rect 12756 -15961 12762 -15927
rect 12796 -15961 12802 -15927
rect 13774 -15529 13780 -15516
rect 13814 -15514 13830 -15495
rect 14780 -15495 14840 -15018
rect 15284 -15068 15344 -14910
rect 15804 -15036 15864 -14820
rect 16296 -14864 16356 -14862
rect 16098 -14870 16586 -14864
rect 16098 -14904 16145 -14870
rect 16179 -14904 16217 -14870
rect 16251 -14904 16289 -14870
rect 16323 -14904 16361 -14870
rect 16395 -14904 16433 -14870
rect 16467 -14904 16505 -14870
rect 16539 -14904 16586 -14870
rect 16098 -14910 16586 -14904
rect 15278 -15072 15350 -15068
rect 15278 -15124 15288 -15072
rect 15340 -15124 15350 -15072
rect 15278 -15128 15350 -15124
rect 15648 -15096 15864 -15036
rect 16296 -15068 16356 -14910
rect 16818 -14958 16878 -14801
rect 17838 -14801 17852 -14767
rect 17886 -14801 17900 -14767
rect 18864 -14767 18910 -14729
rect 19882 -14335 19928 -14297
rect 19882 -14369 19888 -14335
rect 19922 -14369 19928 -14335
rect 19882 -14407 19928 -14369
rect 19882 -14441 19888 -14407
rect 19922 -14441 19928 -14407
rect 19882 -14479 19928 -14441
rect 19882 -14513 19888 -14479
rect 19922 -14513 19928 -14479
rect 19882 -14551 19928 -14513
rect 19882 -14585 19888 -14551
rect 19922 -14585 19928 -14551
rect 19882 -14623 19928 -14585
rect 19882 -14657 19888 -14623
rect 19922 -14657 19928 -14623
rect 19882 -14695 19928 -14657
rect 19882 -14729 19888 -14695
rect 19922 -14729 19928 -14695
rect 19882 -14764 19928 -14729
rect 20892 -14297 20906 -14263
rect 20940 -14276 20954 -14263
rect 21912 -14263 21976 -14244
rect 21912 -14272 21924 -14263
rect 20940 -14297 20952 -14276
rect 20892 -14335 20952 -14297
rect 21916 -14297 21924 -14272
rect 21958 -14297 21976 -14263
rect 22942 -14263 22976 -14244
rect 21916 -14308 21976 -14297
rect 22936 -14297 22942 -14284
rect 22976 -14297 22982 -14284
rect 20892 -14369 20906 -14335
rect 20940 -14369 20952 -14335
rect 20892 -14407 20952 -14369
rect 20892 -14441 20906 -14407
rect 20940 -14441 20952 -14407
rect 20892 -14479 20952 -14441
rect 20892 -14513 20906 -14479
rect 20940 -14513 20952 -14479
rect 20892 -14551 20952 -14513
rect 20892 -14585 20906 -14551
rect 20940 -14585 20952 -14551
rect 20892 -14623 20952 -14585
rect 20892 -14657 20906 -14623
rect 20940 -14657 20952 -14623
rect 20892 -14695 20952 -14657
rect 20892 -14729 20906 -14695
rect 20940 -14729 20952 -14695
rect 18864 -14784 18870 -14767
rect 17838 -14820 17900 -14801
rect 18856 -14801 18870 -14784
rect 18904 -14784 18910 -14767
rect 19872 -14767 19932 -14764
rect 18904 -14801 18916 -14784
rect 17328 -14864 17388 -14862
rect 17116 -14870 17604 -14864
rect 17116 -14904 17163 -14870
rect 17197 -14904 17235 -14870
rect 17269 -14904 17307 -14870
rect 17341 -14904 17379 -14870
rect 17413 -14904 17451 -14870
rect 17485 -14904 17523 -14870
rect 17557 -14904 17604 -14870
rect 17116 -14910 17604 -14904
rect 18134 -14870 18622 -14864
rect 18134 -14904 18181 -14870
rect 18215 -14904 18253 -14870
rect 18287 -14904 18325 -14870
rect 18359 -14904 18397 -14870
rect 18431 -14904 18469 -14870
rect 18503 -14904 18541 -14870
rect 18575 -14904 18622 -14870
rect 18134 -14910 18622 -14904
rect 16812 -14962 16884 -14958
rect 16812 -15014 16822 -14962
rect 16874 -15014 16884 -14962
rect 16812 -15018 16884 -15014
rect 16290 -15072 16362 -15068
rect 15284 -15386 15344 -15128
rect 15648 -15280 15708 -15096
rect 16290 -15124 16300 -15072
rect 16352 -15124 16362 -15072
rect 16290 -15128 16362 -15124
rect 15796 -15178 15868 -15174
rect 15796 -15230 15806 -15178
rect 15858 -15230 15868 -15178
rect 15796 -15234 15868 -15230
rect 15642 -15284 15714 -15280
rect 15642 -15336 15652 -15284
rect 15704 -15336 15714 -15284
rect 15642 -15340 15714 -15336
rect 15080 -15392 15568 -15386
rect 15080 -15426 15127 -15392
rect 15161 -15426 15199 -15392
rect 15233 -15426 15271 -15392
rect 15305 -15426 15343 -15392
rect 15377 -15426 15415 -15392
rect 15449 -15426 15487 -15392
rect 15521 -15426 15568 -15392
rect 15080 -15432 15568 -15426
rect 13814 -15516 13828 -15514
rect 13814 -15529 13820 -15516
rect 14780 -15522 14798 -15495
rect 13774 -15567 13820 -15529
rect 13774 -15601 13780 -15567
rect 13814 -15601 13820 -15567
rect 13774 -15639 13820 -15601
rect 13774 -15673 13780 -15639
rect 13814 -15673 13820 -15639
rect 13774 -15711 13820 -15673
rect 13774 -15745 13780 -15711
rect 13814 -15745 13820 -15711
rect 13774 -15783 13820 -15745
rect 13774 -15817 13780 -15783
rect 13814 -15817 13820 -15783
rect 13774 -15855 13820 -15817
rect 13774 -15889 13780 -15855
rect 13814 -15889 13820 -15855
rect 13774 -15927 13820 -15889
rect 13774 -15938 13780 -15927
rect 12756 -15999 12802 -15961
rect 12756 -16004 12762 -15999
rect 11744 -16052 11778 -16033
rect 12750 -16033 12762 -16004
rect 12796 -16004 12802 -15999
rect 13814 -15938 13820 -15927
rect 14792 -15529 14798 -15522
rect 14832 -15522 14840 -15495
rect 15802 -15476 15862 -15234
rect 16296 -15386 16356 -15128
rect 16098 -15392 16586 -15386
rect 16098 -15426 16145 -15392
rect 16179 -15426 16217 -15392
rect 16251 -15426 16289 -15392
rect 16323 -15426 16361 -15392
rect 16395 -15426 16433 -15392
rect 16467 -15426 16505 -15392
rect 16539 -15426 16586 -15392
rect 16098 -15432 16586 -15426
rect 15802 -15495 15866 -15476
rect 14832 -15529 14838 -15522
rect 15802 -15528 15816 -15495
rect 14792 -15567 14838 -15529
rect 14792 -15601 14798 -15567
rect 14832 -15601 14838 -15567
rect 14792 -15639 14838 -15601
rect 14792 -15673 14798 -15639
rect 14832 -15673 14838 -15639
rect 14792 -15711 14838 -15673
rect 14792 -15745 14798 -15711
rect 14832 -15745 14838 -15711
rect 14792 -15783 14838 -15745
rect 14792 -15817 14798 -15783
rect 14832 -15817 14838 -15783
rect 14792 -15855 14838 -15817
rect 14792 -15889 14798 -15855
rect 14832 -15889 14838 -15855
rect 14792 -15927 14838 -15889
rect 13780 -15999 13814 -15961
rect 14792 -15961 14798 -15927
rect 14832 -15961 14838 -15927
rect 14792 -15998 14838 -15961
rect 15810 -15529 15816 -15528
rect 15850 -15518 15866 -15495
rect 16818 -15495 16878 -15018
rect 17328 -15068 17388 -14910
rect 18342 -15068 18402 -14910
rect 18856 -14958 18916 -14801
rect 19872 -14801 19888 -14767
rect 19922 -14801 19932 -14767
rect 19152 -14870 19640 -14864
rect 19152 -14904 19199 -14870
rect 19233 -14904 19271 -14870
rect 19305 -14904 19343 -14870
rect 19377 -14904 19415 -14870
rect 19449 -14904 19487 -14870
rect 19521 -14904 19559 -14870
rect 19593 -14904 19640 -14870
rect 19152 -14910 19420 -14904
rect 19424 -14910 19640 -14904
rect 18850 -14962 18922 -14958
rect 18850 -15014 18860 -14962
rect 18912 -15014 18922 -14962
rect 18850 -15018 18922 -15014
rect 17322 -15072 17394 -15068
rect 17322 -15124 17332 -15072
rect 17384 -15124 17394 -15072
rect 17322 -15128 17394 -15124
rect 18336 -15072 18408 -15068
rect 18336 -15124 18346 -15072
rect 18398 -15124 18408 -15072
rect 18336 -15128 18408 -15124
rect 17328 -15386 17388 -15128
rect 17836 -15178 17908 -15174
rect 17836 -15230 17846 -15178
rect 17898 -15230 17908 -15178
rect 17836 -15234 17908 -15230
rect 17116 -15392 17314 -15386
rect 17328 -15392 17604 -15386
rect 17116 -15426 17163 -15392
rect 17197 -15426 17235 -15392
rect 17269 -15426 17307 -15392
rect 17341 -15426 17379 -15392
rect 17413 -15426 17451 -15392
rect 17485 -15426 17523 -15392
rect 17557 -15426 17604 -15392
rect 17116 -15432 17604 -15426
rect 17842 -15476 17902 -15234
rect 18342 -15386 18402 -15128
rect 18134 -15392 18402 -15386
rect 18412 -15392 18622 -15386
rect 18134 -15426 18181 -15392
rect 18215 -15426 18253 -15392
rect 18287 -15426 18325 -15392
rect 18359 -15426 18397 -15392
rect 18431 -15426 18469 -15392
rect 18503 -15426 18541 -15392
rect 18575 -15426 18622 -15392
rect 18134 -15432 18622 -15426
rect 15850 -15528 15862 -15518
rect 15850 -15529 15856 -15528
rect 15810 -15567 15856 -15529
rect 15810 -15601 15816 -15567
rect 15850 -15601 15856 -15567
rect 15810 -15639 15856 -15601
rect 15810 -15673 15816 -15639
rect 15850 -15673 15856 -15639
rect 15810 -15711 15856 -15673
rect 15810 -15745 15816 -15711
rect 15850 -15745 15856 -15711
rect 15810 -15783 15856 -15745
rect 15810 -15817 15816 -15783
rect 15850 -15817 15856 -15783
rect 15810 -15855 15856 -15817
rect 15810 -15889 15816 -15855
rect 15850 -15889 15856 -15855
rect 15810 -15927 15856 -15889
rect 15810 -15961 15816 -15927
rect 15850 -15961 15856 -15927
rect 12796 -16033 12810 -16004
rect 11008 -16102 11176 -16096
rect 12424 -16102 12514 -16096
rect 11008 -16136 11055 -16102
rect 11089 -16136 11127 -16102
rect 11161 -16136 11199 -16102
rect 11233 -16136 11271 -16102
rect 11305 -16136 11343 -16102
rect 11377 -16136 11415 -16102
rect 11449 -16136 11484 -16102
rect 12038 -16136 12073 -16102
rect 12107 -16136 12145 -16102
rect 12179 -16136 12217 -16102
rect 12251 -16136 12289 -16102
rect 12323 -16136 12361 -16102
rect 12395 -16136 12433 -16102
rect 12467 -16136 12514 -16102
rect 11008 -16142 11176 -16136
rect 12424 -16142 12514 -16136
rect 12750 -16274 12810 -16033
rect 13780 -16052 13814 -16033
rect 14780 -15999 14840 -15998
rect 14780 -16033 14798 -15999
rect 14832 -16033 14840 -15999
rect 14780 -16052 14840 -16033
rect 15810 -15999 15856 -15961
rect 15810 -16033 15816 -15999
rect 15850 -16033 15856 -15999
rect 15810 -16064 15856 -16033
rect 16818 -15529 16834 -15495
rect 16868 -15529 16878 -15495
rect 17838 -15495 17902 -15476
rect 17838 -15518 17852 -15495
rect 16818 -15567 16878 -15529
rect 17842 -15529 17852 -15518
rect 17886 -15529 17902 -15495
rect 17842 -15538 17902 -15529
rect 18856 -15495 18916 -15018
rect 19360 -15068 19420 -14910
rect 19354 -15072 19426 -15068
rect 19354 -15124 19364 -15072
rect 19416 -15124 19426 -15072
rect 19354 -15128 19426 -15124
rect 19360 -15386 19420 -15128
rect 19872 -15174 19932 -14801
rect 20892 -14767 20952 -14729
rect 21918 -14335 21964 -14308
rect 21918 -14369 21924 -14335
rect 21958 -14369 21964 -14335
rect 21918 -14407 21964 -14369
rect 21918 -14441 21924 -14407
rect 21958 -14441 21964 -14407
rect 21918 -14479 21964 -14441
rect 21918 -14513 21924 -14479
rect 21958 -14513 21964 -14479
rect 21918 -14551 21964 -14513
rect 21918 -14585 21924 -14551
rect 21958 -14585 21964 -14551
rect 21918 -14623 21964 -14585
rect 21918 -14657 21924 -14623
rect 21958 -14657 21964 -14623
rect 21918 -14695 21964 -14657
rect 21918 -14729 21924 -14695
rect 21958 -14729 21964 -14695
rect 21918 -14760 21964 -14729
rect 22936 -14335 22982 -14297
rect 22936 -14369 22942 -14335
rect 22976 -14369 22982 -14335
rect 22936 -14407 22982 -14369
rect 22936 -14441 22942 -14407
rect 22976 -14441 22982 -14407
rect 22936 -14479 22982 -14441
rect 22936 -14513 22942 -14479
rect 22976 -14513 22982 -14479
rect 22936 -14551 22982 -14513
rect 22936 -14585 22942 -14551
rect 22976 -14585 22982 -14551
rect 22936 -14623 22982 -14585
rect 22936 -14657 22942 -14623
rect 22976 -14657 22982 -14623
rect 22936 -14695 22982 -14657
rect 22936 -14729 22942 -14695
rect 22976 -14729 22982 -14695
rect 20892 -14801 20906 -14767
rect 20940 -14801 20952 -14767
rect 20170 -14870 20658 -14864
rect 20170 -14904 20217 -14870
rect 20251 -14904 20289 -14870
rect 20323 -14904 20361 -14870
rect 20395 -14904 20433 -14870
rect 20467 -14904 20505 -14870
rect 20539 -14904 20577 -14870
rect 20611 -14904 20658 -14870
rect 20170 -14910 20658 -14904
rect 20384 -15068 20444 -14910
rect 20892 -14958 20952 -14801
rect 21912 -14767 21972 -14760
rect 21912 -14801 21924 -14767
rect 21958 -14801 21972 -14767
rect 22936 -14767 22982 -14729
rect 22936 -14772 22942 -14767
rect 21188 -14870 21676 -14864
rect 21188 -14904 21235 -14870
rect 21269 -14904 21307 -14870
rect 21341 -14904 21379 -14870
rect 21413 -14904 21451 -14870
rect 21485 -14904 21523 -14870
rect 21557 -14904 21595 -14870
rect 21629 -14904 21676 -14870
rect 21188 -14910 21676 -14904
rect 20886 -14962 20958 -14958
rect 20886 -15014 20896 -14962
rect 20948 -15014 20958 -14962
rect 20886 -15018 20958 -15014
rect 20378 -15072 20450 -15068
rect 20378 -15124 20388 -15072
rect 20440 -15124 20450 -15072
rect 20378 -15128 20450 -15124
rect 19866 -15178 19938 -15174
rect 19866 -15230 19876 -15178
rect 19928 -15230 19938 -15178
rect 19866 -15234 19938 -15230
rect 19866 -15282 19938 -15278
rect 19866 -15334 19876 -15282
rect 19928 -15334 19938 -15282
rect 19866 -15338 19938 -15334
rect 19152 -15392 19352 -15386
rect 19360 -15392 19640 -15386
rect 19152 -15426 19199 -15392
rect 19233 -15426 19271 -15392
rect 19305 -15426 19343 -15392
rect 19377 -15426 19415 -15392
rect 19449 -15426 19487 -15392
rect 19521 -15426 19559 -15392
rect 19593 -15426 19640 -15392
rect 19152 -15432 19640 -15426
rect 19352 -15444 19412 -15432
rect 19872 -15476 19932 -15338
rect 20384 -15386 20444 -15128
rect 20170 -15392 20658 -15386
rect 20170 -15426 20217 -15392
rect 20251 -15426 20289 -15392
rect 20323 -15426 20361 -15392
rect 20395 -15426 20433 -15392
rect 20467 -15426 20505 -15392
rect 20539 -15426 20577 -15392
rect 20611 -15426 20658 -15392
rect 20170 -15432 20658 -15426
rect 18856 -15529 18870 -15495
rect 18904 -15529 18916 -15495
rect 19870 -15495 19932 -15476
rect 19870 -15522 19888 -15495
rect 18856 -15534 18916 -15529
rect 19872 -15529 19888 -15522
rect 19922 -15529 19932 -15495
rect 20892 -15495 20952 -15018
rect 21404 -15068 21464 -14910
rect 21912 -14968 21972 -14801
rect 22928 -14801 22942 -14772
rect 22976 -14772 22982 -14767
rect 22976 -14801 22988 -14772
rect 22206 -14870 22694 -14864
rect 22206 -14904 22253 -14870
rect 22287 -14904 22325 -14870
rect 22359 -14904 22397 -14870
rect 22431 -14904 22469 -14870
rect 22503 -14904 22541 -14870
rect 22575 -14904 22613 -14870
rect 22647 -14904 22694 -14870
rect 22206 -14910 22694 -14904
rect 22422 -14968 22482 -14910
rect 22928 -14968 22988 -14801
rect 23048 -14968 23108 -14096
rect 21912 -15028 23108 -14968
rect 21398 -15072 21470 -15068
rect 21398 -15124 21408 -15072
rect 21460 -15124 21470 -15072
rect 21398 -15128 21470 -15124
rect 21404 -15386 21464 -15128
rect 21906 -15178 21978 -15174
rect 21906 -15230 21916 -15178
rect 21968 -15230 21978 -15178
rect 21906 -15234 21978 -15230
rect 21912 -15276 21972 -15234
rect 21912 -15336 22990 -15276
rect 23048 -15278 23108 -15028
rect 21188 -15392 21676 -15386
rect 21188 -15426 21235 -15392
rect 21269 -15426 21307 -15392
rect 21341 -15426 21379 -15392
rect 21413 -15426 21451 -15392
rect 21485 -15426 21523 -15392
rect 21557 -15426 21595 -15392
rect 21629 -15426 21676 -15392
rect 21188 -15432 21676 -15426
rect 20892 -15502 20906 -15495
rect 16818 -15601 16834 -15567
rect 16868 -15601 16878 -15567
rect 16818 -15639 16878 -15601
rect 16818 -15673 16834 -15639
rect 16868 -15673 16878 -15639
rect 16818 -15711 16878 -15673
rect 16818 -15745 16834 -15711
rect 16868 -15745 16878 -15711
rect 16818 -15783 16878 -15745
rect 16818 -15817 16834 -15783
rect 16868 -15817 16878 -15783
rect 16818 -15855 16878 -15817
rect 16818 -15889 16834 -15855
rect 16868 -15889 16878 -15855
rect 16818 -15927 16878 -15889
rect 16818 -15961 16834 -15927
rect 16868 -15961 16878 -15927
rect 16818 -15999 16878 -15961
rect 16818 -16033 16834 -15999
rect 16868 -16033 16878 -15999
rect 13044 -16102 13236 -16096
rect 14480 -16102 14550 -16096
rect 13044 -16136 13091 -16102
rect 13125 -16136 13163 -16102
rect 13197 -16136 13235 -16102
rect 13269 -16136 13307 -16102
rect 13341 -16136 13379 -16102
rect 13413 -16136 13451 -16102
rect 13485 -16136 13520 -16102
rect 14074 -16136 14109 -16102
rect 14143 -16136 14181 -16102
rect 14215 -16136 14253 -16102
rect 14287 -16136 14325 -16102
rect 14359 -16136 14397 -16102
rect 14431 -16136 14469 -16102
rect 14503 -16136 14550 -16102
rect 13044 -16142 13236 -16136
rect 14480 -16142 14550 -16136
rect 15080 -16102 15568 -16096
rect 15080 -16136 15127 -16102
rect 15161 -16136 15199 -16102
rect 15233 -16136 15271 -16102
rect 15305 -16136 15343 -16102
rect 15377 -16136 15415 -16102
rect 15449 -16136 15487 -16102
rect 15521 -16136 15568 -16102
rect 15080 -16142 15568 -16136
rect 16098 -16102 16586 -16096
rect 16098 -16136 16145 -16102
rect 16179 -16136 16217 -16102
rect 16251 -16136 16289 -16102
rect 16323 -16136 16361 -16102
rect 16395 -16136 16433 -16102
rect 16467 -16136 16505 -16102
rect 16539 -16136 16586 -16102
rect 16098 -16142 16586 -16136
rect 14776 -16174 14848 -16170
rect 14776 -16226 14786 -16174
rect 14838 -16226 14848 -16174
rect 14776 -16230 14848 -16226
rect 10706 -16278 10778 -16274
rect 10706 -16330 10716 -16278
rect 10768 -16330 10778 -16278
rect 10706 -16334 10778 -16330
rect 12744 -16278 12816 -16274
rect 12744 -16330 12754 -16278
rect 12806 -16330 12816 -16278
rect 12744 -16334 12816 -16330
rect 9690 -16400 9762 -16396
rect 9690 -16452 9700 -16400
rect 9752 -16452 9762 -16400
rect 9690 -16456 9762 -16452
rect 11724 -16400 11796 -16396
rect 11724 -16452 11734 -16400
rect 11786 -16452 11796 -16400
rect 11724 -16456 11796 -16452
rect 13754 -16400 13826 -16396
rect 13754 -16452 13764 -16400
rect 13816 -16452 13826 -16400
rect 13754 -16456 13826 -16452
rect 8970 -16626 9458 -16620
rect 8970 -16660 9017 -16626
rect 9051 -16660 9089 -16626
rect 9123 -16660 9161 -16626
rect 9195 -16660 9233 -16626
rect 9267 -16660 9305 -16626
rect 9339 -16660 9377 -16626
rect 9411 -16660 9458 -16626
rect 8970 -16666 9458 -16660
rect 7704 -16763 7710 -16754
rect 7664 -16801 7710 -16763
rect 8676 -16763 8688 -16729
rect 8722 -16763 8736 -16729
rect 8676 -16772 8736 -16763
rect 9696 -16729 9756 -16456
rect 9988 -16626 10476 -16620
rect 9988 -16660 10035 -16626
rect 10069 -16660 10107 -16626
rect 10141 -16660 10179 -16626
rect 10213 -16660 10251 -16626
rect 10285 -16660 10323 -16626
rect 10357 -16660 10395 -16626
rect 10429 -16660 10476 -16626
rect 9988 -16666 10476 -16660
rect 11006 -16626 11494 -16620
rect 11006 -16660 11053 -16626
rect 11087 -16660 11125 -16626
rect 11159 -16660 11197 -16626
rect 11231 -16660 11269 -16626
rect 11303 -16660 11341 -16626
rect 11375 -16660 11413 -16626
rect 11447 -16660 11494 -16626
rect 11006 -16666 11494 -16660
rect 9696 -16763 9706 -16729
rect 9740 -16763 9756 -16729
rect 9696 -16766 9756 -16763
rect 10718 -16729 10764 -16698
rect 10718 -16763 10724 -16729
rect 10758 -16763 10764 -16729
rect 11730 -16729 11790 -16456
rect 12024 -16626 12512 -16620
rect 12024 -16660 12071 -16626
rect 12105 -16660 12143 -16626
rect 12177 -16660 12215 -16626
rect 12249 -16660 12287 -16626
rect 12321 -16660 12359 -16626
rect 12393 -16660 12431 -16626
rect 12465 -16660 12512 -16626
rect 12024 -16666 12512 -16660
rect 13042 -16626 13530 -16620
rect 13042 -16660 13089 -16626
rect 13123 -16660 13161 -16626
rect 13195 -16660 13233 -16626
rect 13267 -16660 13305 -16626
rect 13339 -16660 13377 -16626
rect 13411 -16660 13449 -16626
rect 13483 -16660 13530 -16626
rect 13042 -16666 13530 -16660
rect 11730 -16760 11742 -16729
rect 7664 -16835 7670 -16801
rect 7704 -16835 7710 -16801
rect 7664 -16873 7710 -16835
rect 7664 -16907 7670 -16873
rect 7704 -16907 7710 -16873
rect 7664 -16945 7710 -16907
rect 7664 -16979 7670 -16945
rect 7704 -16979 7710 -16945
rect 7664 -17017 7710 -16979
rect 7664 -17051 7670 -17017
rect 7704 -17051 7710 -17017
rect 7664 -17089 7710 -17051
rect 7664 -17123 7670 -17089
rect 7704 -17123 7710 -17089
rect 7664 -17161 7710 -17123
rect 7664 -17195 7670 -17161
rect 7704 -17195 7710 -17161
rect 7664 -17233 7710 -17195
rect 7664 -17236 7670 -17233
rect 6646 -17298 6692 -17267
rect 7656 -17267 7670 -17236
rect 7704 -17236 7710 -17233
rect 8682 -16801 8728 -16772
rect 8682 -16835 8688 -16801
rect 8722 -16835 8728 -16801
rect 8682 -16873 8728 -16835
rect 8682 -16907 8688 -16873
rect 8722 -16907 8728 -16873
rect 8682 -16945 8728 -16907
rect 8682 -16979 8688 -16945
rect 8722 -16979 8728 -16945
rect 8682 -17017 8728 -16979
rect 8682 -17051 8688 -17017
rect 8722 -17051 8728 -17017
rect 8682 -17089 8728 -17051
rect 8682 -17123 8688 -17089
rect 8722 -17123 8728 -17089
rect 8682 -17161 8728 -17123
rect 8682 -17195 8688 -17161
rect 8722 -17195 8728 -17161
rect 8682 -17233 8728 -17195
rect 7704 -17267 7716 -17236
rect 8682 -17250 8688 -17233
rect 5916 -17336 6404 -17330
rect 5916 -17370 5963 -17336
rect 5997 -17370 6035 -17336
rect 6069 -17370 6107 -17336
rect 6141 -17370 6179 -17336
rect 6213 -17370 6251 -17336
rect 6285 -17370 6323 -17336
rect 6357 -17370 6404 -17336
rect 5916 -17376 6404 -17370
rect 6934 -17336 7422 -17330
rect 6934 -17370 6981 -17336
rect 7015 -17370 7053 -17336
rect 7087 -17370 7125 -17336
rect 7159 -17370 7197 -17336
rect 7231 -17370 7269 -17336
rect 7303 -17370 7341 -17336
rect 7375 -17370 7422 -17336
rect 6934 -17376 7422 -17370
rect 5614 -17418 5686 -17414
rect 5614 -17470 5624 -17418
rect 5676 -17470 5686 -17418
rect 5614 -17474 5686 -17470
rect 5110 -17636 5182 -17632
rect 5110 -17688 5120 -17636
rect 5172 -17688 5182 -17636
rect 5110 -17692 5182 -17688
rect 5116 -17854 5176 -17692
rect 4898 -17860 5386 -17854
rect 4898 -17894 4945 -17860
rect 4979 -17894 5017 -17860
rect 5051 -17894 5089 -17860
rect 5123 -17894 5161 -17860
rect 5195 -17894 5233 -17860
rect 5267 -17894 5305 -17860
rect 5339 -17894 5386 -17860
rect 4898 -17900 5386 -17894
rect 3632 -17997 3638 -17980
rect 4602 -17986 4616 -17963
rect 3592 -18035 3638 -17997
rect 3592 -18069 3598 -18035
rect 3632 -18069 3638 -18035
rect 3592 -18107 3638 -18069
rect 3592 -18141 3598 -18107
rect 3632 -18141 3638 -18107
rect 3592 -18179 3638 -18141
rect 3592 -18213 3598 -18179
rect 3632 -18213 3638 -18179
rect 3592 -18251 3638 -18213
rect 3592 -18285 3598 -18251
rect 3632 -18285 3638 -18251
rect 3592 -18323 3638 -18285
rect 3592 -18357 3598 -18323
rect 3632 -18357 3638 -18323
rect 3592 -18395 3638 -18357
rect 3592 -18429 3598 -18395
rect 3632 -18429 3638 -18395
rect 3592 -18467 3638 -18429
rect 4610 -17997 4616 -17986
rect 4650 -17986 4662 -17963
rect 5620 -17963 5680 -17474
rect 6118 -17626 6178 -17376
rect 6636 -17522 6708 -17518
rect 6636 -17574 6646 -17522
rect 6698 -17574 6708 -17522
rect 6636 -17578 6708 -17574
rect 6118 -17636 6180 -17626
rect 6118 -17688 6124 -17636
rect 6176 -17688 6180 -17636
rect 6118 -17698 6180 -17688
rect 6118 -17854 6178 -17698
rect 5916 -17860 6404 -17854
rect 5916 -17894 5963 -17860
rect 5997 -17894 6035 -17860
rect 6069 -17894 6107 -17860
rect 6141 -17894 6179 -17860
rect 6213 -17894 6251 -17860
rect 6285 -17894 6323 -17860
rect 6357 -17894 6404 -17860
rect 5916 -17900 6404 -17894
rect 4650 -17997 4656 -17986
rect 5620 -17988 5634 -17963
rect 4610 -18035 4656 -17997
rect 4610 -18069 4616 -18035
rect 4650 -18069 4656 -18035
rect 4610 -18107 4656 -18069
rect 4610 -18141 4616 -18107
rect 4650 -18141 4656 -18107
rect 4610 -18179 4656 -18141
rect 4610 -18213 4616 -18179
rect 4650 -18213 4656 -18179
rect 4610 -18251 4656 -18213
rect 4610 -18285 4616 -18251
rect 4650 -18285 4656 -18251
rect 4610 -18323 4656 -18285
rect 4610 -18357 4616 -18323
rect 4650 -18357 4656 -18323
rect 4610 -18395 4656 -18357
rect 4610 -18429 4616 -18395
rect 4650 -18429 4656 -18395
rect 4610 -18462 4656 -18429
rect 5628 -17997 5634 -17988
rect 5668 -17988 5680 -17963
rect 6642 -17963 6702 -17578
rect 7134 -17626 7194 -17376
rect 7656 -17414 7716 -17267
rect 8674 -17267 8688 -17250
rect 8722 -17250 8728 -17233
rect 9700 -16801 9746 -16766
rect 9700 -16835 9706 -16801
rect 9740 -16835 9746 -16801
rect 9700 -16873 9746 -16835
rect 9700 -16907 9706 -16873
rect 9740 -16907 9746 -16873
rect 9700 -16945 9746 -16907
rect 9700 -16979 9706 -16945
rect 9740 -16979 9746 -16945
rect 9700 -17017 9746 -16979
rect 9700 -17051 9706 -17017
rect 9740 -17051 9746 -17017
rect 9700 -17089 9746 -17051
rect 9700 -17123 9706 -17089
rect 9740 -17123 9746 -17089
rect 9700 -17161 9746 -17123
rect 9700 -17195 9706 -17161
rect 9740 -17195 9746 -17161
rect 9700 -17233 9746 -17195
rect 8722 -17267 8734 -17250
rect 7952 -17336 8440 -17330
rect 7952 -17370 7999 -17336
rect 8033 -17370 8071 -17336
rect 8105 -17370 8143 -17336
rect 8177 -17370 8215 -17336
rect 8249 -17370 8287 -17336
rect 8321 -17370 8359 -17336
rect 8393 -17370 8440 -17336
rect 7952 -17376 8440 -17370
rect 7650 -17418 7722 -17414
rect 7650 -17470 7660 -17418
rect 7712 -17470 7722 -17418
rect 7650 -17474 7722 -17470
rect 7132 -17636 7194 -17626
rect 7132 -17688 7136 -17636
rect 7188 -17688 7194 -17636
rect 7132 -17698 7194 -17688
rect 7134 -17854 7194 -17698
rect 6934 -17860 7422 -17854
rect 6934 -17894 6981 -17860
rect 7015 -17894 7053 -17860
rect 7087 -17894 7125 -17860
rect 7159 -17894 7197 -17860
rect 7231 -17894 7269 -17860
rect 7303 -17894 7341 -17860
rect 7375 -17894 7422 -17860
rect 6934 -17900 7422 -17894
rect 6642 -17986 6652 -17963
rect 5668 -17997 5674 -17988
rect 5628 -18035 5674 -17997
rect 5628 -18069 5634 -18035
rect 5668 -18069 5674 -18035
rect 5628 -18107 5674 -18069
rect 5628 -18141 5634 -18107
rect 5668 -18141 5674 -18107
rect 5628 -18179 5674 -18141
rect 5628 -18213 5634 -18179
rect 5668 -18213 5674 -18179
rect 5628 -18251 5674 -18213
rect 5628 -18285 5634 -18251
rect 5668 -18285 5674 -18251
rect 5628 -18323 5674 -18285
rect 5628 -18357 5634 -18323
rect 5668 -18357 5674 -18323
rect 5628 -18395 5674 -18357
rect 5628 -18429 5634 -18395
rect 5668 -18429 5674 -18395
rect 3592 -18501 3598 -18467
rect 3632 -18501 3638 -18467
rect 3592 -18532 3638 -18501
rect 4604 -18467 4664 -18462
rect 4604 -18501 4616 -18467
rect 4650 -18501 4664 -18467
rect 5628 -18467 5674 -18429
rect 5628 -18472 5634 -18467
rect 2862 -18570 3350 -18564
rect 2862 -18604 2909 -18570
rect 2943 -18604 2981 -18570
rect 3015 -18604 3053 -18570
rect 3087 -18604 3125 -18570
rect 3159 -18604 3197 -18570
rect 3231 -18604 3269 -18570
rect 3303 -18604 3350 -18570
rect 2862 -18610 3350 -18604
rect 3880 -18570 4368 -18564
rect 3880 -18604 3927 -18570
rect 3961 -18604 3999 -18570
rect 4033 -18604 4071 -18570
rect 4105 -18604 4143 -18570
rect 4177 -18604 4215 -18570
rect 4249 -18604 4287 -18570
rect 4321 -18604 4368 -18570
rect 3880 -18610 4368 -18604
rect 3578 -18674 3650 -18670
rect 3578 -18726 3588 -18674
rect 3640 -18726 3650 -18674
rect 3578 -18730 3650 -18726
rect 2862 -19092 3350 -19086
rect 2862 -19126 2909 -19092
rect 2943 -19126 2981 -19092
rect 3015 -19126 3053 -19092
rect 3087 -19126 3125 -19092
rect 3159 -19126 3197 -19092
rect 3231 -19126 3269 -19092
rect 3303 -19126 3350 -19092
rect 2862 -19132 3350 -19126
rect 2574 -19195 2620 -19164
rect 2574 -19229 2580 -19195
rect 2614 -19229 2620 -19195
rect 3584 -19195 3644 -18730
rect 4090 -18772 4150 -18610
rect 4084 -18776 4156 -18772
rect 4084 -18828 4094 -18776
rect 4146 -18828 4156 -18776
rect 4084 -18832 4156 -18828
rect 4604 -18974 4664 -18501
rect 5622 -18501 5634 -18472
rect 5668 -18472 5674 -18467
rect 6646 -17997 6652 -17986
rect 6686 -17986 6702 -17963
rect 7656 -17963 7716 -17474
rect 8152 -17636 8212 -17376
rect 8674 -17518 8734 -17267
rect 9700 -17267 9706 -17233
rect 9740 -17267 9746 -17233
rect 10718 -16801 10764 -16763
rect 10718 -16835 10724 -16801
rect 10758 -16835 10764 -16801
rect 10718 -16873 10764 -16835
rect 10718 -16907 10724 -16873
rect 10758 -16907 10764 -16873
rect 10718 -16945 10764 -16907
rect 10718 -16979 10724 -16945
rect 10758 -16979 10764 -16945
rect 10718 -17017 10764 -16979
rect 10718 -17051 10724 -17017
rect 10758 -17051 10764 -17017
rect 10718 -17089 10764 -17051
rect 10718 -17123 10724 -17089
rect 10758 -17123 10764 -17089
rect 10718 -17161 10764 -17123
rect 10718 -17195 10724 -17161
rect 10758 -17195 10764 -17161
rect 10718 -17233 10764 -17195
rect 10718 -17256 10724 -17233
rect 9700 -17298 9746 -17267
rect 10708 -17267 10724 -17256
rect 10758 -17256 10764 -17233
rect 11736 -16763 11742 -16760
rect 11776 -16760 11790 -16729
rect 12754 -16729 12800 -16698
rect 11776 -16763 11782 -16760
rect 11736 -16801 11782 -16763
rect 11736 -16835 11742 -16801
rect 11776 -16835 11782 -16801
rect 11736 -16873 11782 -16835
rect 11736 -16907 11742 -16873
rect 11776 -16907 11782 -16873
rect 11736 -16945 11782 -16907
rect 11736 -16979 11742 -16945
rect 11776 -16979 11782 -16945
rect 11736 -17017 11782 -16979
rect 11736 -17051 11742 -17017
rect 11776 -17051 11782 -17017
rect 11736 -17089 11782 -17051
rect 11736 -17123 11742 -17089
rect 11776 -17123 11782 -17089
rect 11736 -17161 11782 -17123
rect 11736 -17195 11742 -17161
rect 11776 -17195 11782 -17161
rect 11736 -17233 11782 -17195
rect 10758 -17267 10768 -17256
rect 8970 -17336 9458 -17330
rect 8970 -17370 9017 -17336
rect 9051 -17370 9089 -17336
rect 9123 -17370 9161 -17336
rect 9195 -17370 9233 -17336
rect 9267 -17370 9305 -17336
rect 9339 -17370 9377 -17336
rect 9411 -17370 9458 -17336
rect 8970 -17376 9458 -17370
rect 9988 -17336 10476 -17330
rect 9988 -17370 10035 -17336
rect 10069 -17370 10107 -17336
rect 10141 -17370 10179 -17336
rect 10213 -17370 10251 -17336
rect 10285 -17370 10323 -17336
rect 10357 -17370 10395 -17336
rect 10429 -17370 10476 -17336
rect 9988 -17376 10476 -17370
rect 8668 -17522 8740 -17518
rect 8668 -17574 8678 -17522
rect 8730 -17574 8740 -17522
rect 8668 -17578 8740 -17574
rect 9164 -17574 9224 -17376
rect 10206 -17574 10266 -17376
rect 10708 -17518 10768 -17267
rect 11736 -17267 11742 -17233
rect 11776 -17267 11782 -17233
rect 12754 -16763 12760 -16729
rect 12794 -16763 12800 -16729
rect 13760 -16729 13820 -16456
rect 14060 -16626 14548 -16620
rect 14060 -16660 14107 -16626
rect 14141 -16660 14179 -16626
rect 14213 -16660 14251 -16626
rect 14285 -16660 14323 -16626
rect 14357 -16660 14395 -16626
rect 14429 -16660 14467 -16626
rect 14501 -16660 14548 -16626
rect 14060 -16666 14548 -16660
rect 13760 -16754 13778 -16729
rect 12754 -16801 12800 -16763
rect 12754 -16835 12760 -16801
rect 12794 -16835 12800 -16801
rect 12754 -16873 12800 -16835
rect 12754 -16907 12760 -16873
rect 12794 -16907 12800 -16873
rect 12754 -16945 12800 -16907
rect 12754 -16979 12760 -16945
rect 12794 -16979 12800 -16945
rect 12754 -17017 12800 -16979
rect 12754 -17051 12760 -17017
rect 12794 -17051 12800 -17017
rect 12754 -17089 12800 -17051
rect 12754 -17123 12760 -17089
rect 12794 -17123 12800 -17089
rect 12754 -17161 12800 -17123
rect 12754 -17195 12760 -17161
rect 12794 -17195 12800 -17161
rect 12754 -17233 12800 -17195
rect 12754 -17244 12760 -17233
rect 11736 -17298 11782 -17267
rect 12748 -17267 12760 -17244
rect 12794 -17244 12800 -17233
rect 13772 -16763 13778 -16754
rect 13812 -16754 13820 -16729
rect 14782 -16729 14842 -16230
rect 15304 -16620 15364 -16142
rect 15794 -16278 15866 -16274
rect 15794 -16330 15804 -16278
rect 15856 -16330 15866 -16278
rect 15794 -16334 15866 -16330
rect 15078 -16626 15566 -16620
rect 15078 -16660 15125 -16626
rect 15159 -16660 15197 -16626
rect 15231 -16660 15269 -16626
rect 15303 -16660 15341 -16626
rect 15375 -16660 15413 -16626
rect 15447 -16660 15485 -16626
rect 15519 -16660 15566 -16626
rect 15078 -16666 15566 -16660
rect 13812 -16763 13818 -16754
rect 14782 -16762 14796 -16729
rect 13772 -16801 13818 -16763
rect 13772 -16835 13778 -16801
rect 13812 -16835 13818 -16801
rect 13772 -16873 13818 -16835
rect 13772 -16907 13778 -16873
rect 13812 -16907 13818 -16873
rect 13772 -16945 13818 -16907
rect 13772 -16979 13778 -16945
rect 13812 -16979 13818 -16945
rect 13772 -17017 13818 -16979
rect 13772 -17051 13778 -17017
rect 13812 -17051 13818 -17017
rect 13772 -17089 13818 -17051
rect 13772 -17123 13778 -17089
rect 13812 -17123 13818 -17089
rect 13772 -17161 13818 -17123
rect 13772 -17195 13778 -17161
rect 13812 -17195 13818 -17161
rect 13772 -17233 13818 -17195
rect 12794 -17267 12808 -17244
rect 11006 -17336 11494 -17330
rect 11006 -17370 11053 -17336
rect 11087 -17370 11125 -17336
rect 11159 -17370 11197 -17336
rect 11231 -17370 11269 -17336
rect 11303 -17370 11341 -17336
rect 11375 -17370 11413 -17336
rect 11447 -17370 11494 -17336
rect 11006 -17376 11494 -17370
rect 12024 -17336 12512 -17330
rect 12024 -17370 12071 -17336
rect 12105 -17370 12143 -17336
rect 12177 -17370 12215 -17336
rect 12249 -17370 12287 -17336
rect 12321 -17370 12359 -17336
rect 12393 -17370 12431 -17336
rect 12465 -17370 12512 -17336
rect 12024 -17376 12512 -17370
rect 8152 -17688 8156 -17636
rect 8208 -17688 8212 -17636
rect 8152 -17854 8212 -17688
rect 8668 -17634 8740 -17630
rect 8668 -17686 8678 -17634
rect 8730 -17686 8740 -17634
rect 8668 -17690 8740 -17686
rect 9164 -17634 10266 -17574
rect 10702 -17522 10774 -17518
rect 10702 -17574 10712 -17522
rect 10764 -17574 10774 -17522
rect 10702 -17578 10774 -17574
rect 7952 -17860 8440 -17854
rect 7952 -17894 7999 -17860
rect 8033 -17894 8071 -17860
rect 8105 -17894 8143 -17860
rect 8177 -17894 8215 -17860
rect 8249 -17894 8287 -17860
rect 8321 -17894 8359 -17860
rect 8393 -17894 8440 -17860
rect 7952 -17900 8440 -17894
rect 6686 -17997 6692 -17986
rect 7656 -17992 7670 -17963
rect 6646 -18035 6692 -17997
rect 6646 -18069 6652 -18035
rect 6686 -18069 6692 -18035
rect 6646 -18107 6692 -18069
rect 6646 -18141 6652 -18107
rect 6686 -18141 6692 -18107
rect 6646 -18179 6692 -18141
rect 6646 -18213 6652 -18179
rect 6686 -18213 6692 -18179
rect 6646 -18251 6692 -18213
rect 6646 -18285 6652 -18251
rect 6686 -18285 6692 -18251
rect 6646 -18323 6692 -18285
rect 6646 -18357 6652 -18323
rect 6686 -18357 6692 -18323
rect 6646 -18395 6692 -18357
rect 6646 -18429 6652 -18395
rect 6686 -18429 6692 -18395
rect 6646 -18467 6692 -18429
rect 5668 -18501 5682 -18472
rect 4898 -18570 5386 -18564
rect 4898 -18604 4945 -18570
rect 4979 -18604 5017 -18570
rect 5051 -18604 5089 -18570
rect 5123 -18604 5161 -18570
rect 5195 -18604 5233 -18570
rect 5267 -18604 5305 -18570
rect 5339 -18604 5386 -18570
rect 4898 -18610 5386 -18604
rect 5622 -18670 5682 -18501
rect 6646 -18501 6652 -18467
rect 6686 -18501 6692 -18467
rect 7664 -17997 7670 -17992
rect 7704 -17992 7716 -17963
rect 8674 -17963 8734 -17690
rect 9164 -17854 9224 -17634
rect 9686 -17744 9758 -17740
rect 9686 -17796 9696 -17744
rect 9748 -17796 9758 -17744
rect 9686 -17800 9758 -17796
rect 8970 -17860 9458 -17854
rect 8970 -17894 9017 -17860
rect 9051 -17894 9089 -17860
rect 9123 -17894 9161 -17860
rect 9195 -17894 9233 -17860
rect 9267 -17894 9305 -17860
rect 9339 -17894 9377 -17860
rect 9411 -17894 9458 -17860
rect 8970 -17900 9458 -17894
rect 7704 -17997 7710 -17992
rect 7664 -18035 7710 -17997
rect 8674 -17997 8688 -17963
rect 8722 -17997 8734 -17963
rect 9692 -17963 9752 -17800
rect 10206 -17854 10266 -17634
rect 10704 -17634 10776 -17630
rect 10704 -17686 10714 -17634
rect 10766 -17686 10776 -17634
rect 10704 -17690 10776 -17686
rect 9988 -17860 10476 -17854
rect 9988 -17894 10035 -17860
rect 10069 -17894 10107 -17860
rect 10141 -17894 10179 -17860
rect 10213 -17894 10251 -17860
rect 10285 -17894 10323 -17860
rect 10357 -17894 10395 -17860
rect 10429 -17894 10476 -17860
rect 9988 -17900 10476 -17894
rect 9692 -17990 9706 -17963
rect 8674 -18002 8734 -17997
rect 9700 -17997 9706 -17990
rect 9740 -17990 9752 -17963
rect 10710 -17963 10770 -17690
rect 11206 -17854 11266 -17376
rect 11720 -17744 11792 -17740
rect 11720 -17796 11730 -17744
rect 11782 -17796 11792 -17744
rect 11720 -17800 11792 -17796
rect 11006 -17860 11494 -17854
rect 11006 -17894 11053 -17860
rect 11087 -17894 11125 -17860
rect 11159 -17894 11197 -17860
rect 11231 -17894 11269 -17860
rect 11303 -17894 11341 -17860
rect 11375 -17894 11413 -17860
rect 11447 -17894 11494 -17860
rect 11006 -17900 11494 -17894
rect 9740 -17997 9746 -17990
rect 7664 -18069 7670 -18035
rect 7704 -18069 7710 -18035
rect 7664 -18107 7710 -18069
rect 7664 -18141 7670 -18107
rect 7704 -18141 7710 -18107
rect 7664 -18179 7710 -18141
rect 7664 -18213 7670 -18179
rect 7704 -18213 7710 -18179
rect 7664 -18251 7710 -18213
rect 7664 -18285 7670 -18251
rect 7704 -18285 7710 -18251
rect 7664 -18323 7710 -18285
rect 7664 -18357 7670 -18323
rect 7704 -18357 7710 -18323
rect 7664 -18395 7710 -18357
rect 7664 -18429 7670 -18395
rect 7704 -18429 7710 -18395
rect 7664 -18467 7710 -18429
rect 7664 -18470 7670 -18467
rect 6646 -18532 6692 -18501
rect 7658 -18501 7670 -18470
rect 7704 -18470 7710 -18467
rect 8682 -18035 8728 -18002
rect 8682 -18069 8688 -18035
rect 8722 -18069 8728 -18035
rect 8682 -18107 8728 -18069
rect 8682 -18141 8688 -18107
rect 8722 -18141 8728 -18107
rect 8682 -18179 8728 -18141
rect 8682 -18213 8688 -18179
rect 8722 -18213 8728 -18179
rect 8682 -18251 8728 -18213
rect 8682 -18285 8688 -18251
rect 8722 -18285 8728 -18251
rect 8682 -18323 8728 -18285
rect 8682 -18357 8688 -18323
rect 8722 -18357 8728 -18323
rect 8682 -18395 8728 -18357
rect 8682 -18429 8688 -18395
rect 8722 -18429 8728 -18395
rect 8682 -18467 8728 -18429
rect 7704 -18501 7718 -18470
rect 5916 -18570 6404 -18564
rect 5916 -18604 5963 -18570
rect 5997 -18604 6035 -18570
rect 6069 -18604 6107 -18570
rect 6141 -18604 6179 -18570
rect 6213 -18604 6251 -18570
rect 6285 -18604 6323 -18570
rect 6357 -18604 6404 -18570
rect 5916 -18610 6404 -18604
rect 6934 -18570 7422 -18564
rect 6934 -18604 6981 -18570
rect 7015 -18604 7053 -18570
rect 7087 -18604 7125 -18570
rect 7159 -18604 7197 -18570
rect 7231 -18604 7269 -18570
rect 7303 -18604 7341 -18570
rect 7375 -18604 7422 -18570
rect 6934 -18610 7422 -18604
rect 5616 -18674 5688 -18670
rect 5616 -18726 5626 -18674
rect 5678 -18726 5688 -18674
rect 5616 -18730 5688 -18726
rect 5614 -18878 5686 -18874
rect 5614 -18930 5624 -18878
rect 5676 -18930 5686 -18878
rect 6128 -18880 6188 -18610
rect 7150 -18880 7210 -18610
rect 7658 -18670 7718 -18501
rect 8682 -18501 8688 -18467
rect 8722 -18501 8728 -18467
rect 8682 -18532 8728 -18501
rect 9700 -18035 9746 -17997
rect 10710 -17997 10724 -17963
rect 10758 -17997 10770 -17963
rect 11726 -17963 11786 -17800
rect 12240 -17854 12300 -17376
rect 12748 -17518 12808 -17267
rect 13772 -17267 13778 -17233
rect 13812 -17267 13818 -17233
rect 14790 -16763 14796 -16762
rect 14830 -16762 14842 -16729
rect 15800 -16729 15860 -16334
rect 16306 -16620 16366 -16142
rect 16818 -16274 16878 -16033
rect 17846 -15567 17892 -15538
rect 17846 -15601 17852 -15567
rect 17886 -15601 17892 -15567
rect 17846 -15639 17892 -15601
rect 17846 -15673 17852 -15639
rect 17886 -15673 17892 -15639
rect 17846 -15711 17892 -15673
rect 17846 -15745 17852 -15711
rect 17886 -15745 17892 -15711
rect 17846 -15783 17892 -15745
rect 17846 -15817 17852 -15783
rect 17886 -15817 17892 -15783
rect 17846 -15855 17892 -15817
rect 17846 -15889 17852 -15855
rect 17886 -15889 17892 -15855
rect 17846 -15927 17892 -15889
rect 17846 -15961 17852 -15927
rect 17886 -15961 17892 -15927
rect 17846 -15999 17892 -15961
rect 17846 -16033 17852 -15999
rect 17886 -16033 17892 -15999
rect 18864 -15567 18910 -15534
rect 19872 -15550 19932 -15529
rect 20900 -15529 20906 -15502
rect 20940 -15502 20952 -15495
rect 21912 -15495 21972 -15336
rect 22398 -15386 22458 -15336
rect 22206 -15392 22458 -15386
rect 22476 -15392 22694 -15386
rect 22206 -15426 22253 -15392
rect 22287 -15426 22325 -15392
rect 22359 -15426 22397 -15392
rect 22431 -15426 22469 -15392
rect 22503 -15426 22541 -15392
rect 22575 -15426 22613 -15392
rect 22647 -15426 22694 -15392
rect 22206 -15432 22694 -15426
rect 22930 -15476 22990 -15336
rect 23042 -15282 23114 -15278
rect 23042 -15334 23052 -15282
rect 23104 -15334 23114 -15282
rect 23042 -15338 23114 -15334
rect 20940 -15529 20946 -15502
rect 18864 -15601 18870 -15567
rect 18904 -15601 18910 -15567
rect 18864 -15639 18910 -15601
rect 18864 -15673 18870 -15639
rect 18904 -15673 18910 -15639
rect 18864 -15711 18910 -15673
rect 18864 -15745 18870 -15711
rect 18904 -15745 18910 -15711
rect 18864 -15783 18910 -15745
rect 18864 -15817 18870 -15783
rect 18904 -15817 18910 -15783
rect 18864 -15855 18910 -15817
rect 18864 -15889 18870 -15855
rect 18904 -15889 18910 -15855
rect 18864 -15927 18910 -15889
rect 18864 -15961 18870 -15927
rect 18904 -15961 18910 -15927
rect 18864 -15999 18910 -15961
rect 19882 -15567 19928 -15550
rect 19882 -15601 19888 -15567
rect 19922 -15601 19928 -15567
rect 19882 -15639 19928 -15601
rect 19882 -15673 19888 -15639
rect 19922 -15673 19928 -15639
rect 19882 -15711 19928 -15673
rect 19882 -15745 19888 -15711
rect 19922 -15745 19928 -15711
rect 19882 -15783 19928 -15745
rect 19882 -15817 19888 -15783
rect 19922 -15817 19928 -15783
rect 19882 -15855 19928 -15817
rect 19882 -15889 19888 -15855
rect 19922 -15889 19928 -15855
rect 19882 -15927 19928 -15889
rect 19882 -15961 19888 -15927
rect 19922 -15961 19928 -15927
rect 19882 -15998 19928 -15961
rect 20900 -15567 20946 -15529
rect 21912 -15529 21924 -15495
rect 21958 -15529 21972 -15495
rect 22926 -15495 22990 -15476
rect 22926 -15512 22942 -15495
rect 22930 -15518 22942 -15512
rect 21912 -15532 21972 -15529
rect 22936 -15529 22942 -15518
rect 22976 -15518 22990 -15495
rect 22976 -15529 22982 -15518
rect 20900 -15601 20906 -15567
rect 20940 -15601 20946 -15567
rect 20900 -15639 20946 -15601
rect 20900 -15673 20906 -15639
rect 20940 -15673 20946 -15639
rect 20900 -15711 20946 -15673
rect 20900 -15745 20906 -15711
rect 20940 -15745 20946 -15711
rect 20900 -15783 20946 -15745
rect 20900 -15817 20906 -15783
rect 20940 -15817 20946 -15783
rect 20900 -15855 20946 -15817
rect 20900 -15889 20906 -15855
rect 20940 -15889 20946 -15855
rect 20900 -15927 20946 -15889
rect 20900 -15961 20906 -15927
rect 20940 -15961 20946 -15927
rect 20900 -15994 20946 -15961
rect 21918 -15567 21964 -15532
rect 21918 -15601 21924 -15567
rect 21958 -15601 21964 -15567
rect 21918 -15639 21964 -15601
rect 21918 -15673 21924 -15639
rect 21958 -15673 21964 -15639
rect 21918 -15711 21964 -15673
rect 21918 -15745 21924 -15711
rect 21958 -15745 21964 -15711
rect 21918 -15783 21964 -15745
rect 21918 -15817 21924 -15783
rect 21958 -15817 21964 -15783
rect 21918 -15855 21964 -15817
rect 21918 -15889 21924 -15855
rect 21958 -15889 21964 -15855
rect 21918 -15927 21964 -15889
rect 21918 -15961 21924 -15927
rect 21958 -15961 21964 -15927
rect 18864 -16004 18870 -15999
rect 17846 -16064 17892 -16033
rect 18854 -16033 18870 -16004
rect 18904 -16004 18910 -15999
rect 19876 -15999 19936 -15998
rect 18904 -16033 18914 -16004
rect 17116 -16102 17604 -16096
rect 17116 -16136 17163 -16102
rect 17197 -16136 17235 -16102
rect 17269 -16136 17379 -16102
rect 17413 -16136 17451 -16102
rect 17485 -16136 17523 -16102
rect 17557 -16136 17604 -16102
rect 17116 -16142 17604 -16136
rect 18134 -16102 18622 -16096
rect 18134 -16136 18181 -16102
rect 18215 -16136 18253 -16102
rect 18287 -16136 18469 -16102
rect 18503 -16136 18541 -16102
rect 18575 -16136 18622 -16102
rect 18134 -16142 18622 -16136
rect 16812 -16278 16884 -16274
rect 16812 -16330 16822 -16278
rect 16874 -16330 16884 -16278
rect 16812 -16334 16884 -16330
rect 17318 -16620 17378 -16142
rect 17832 -16278 17904 -16274
rect 17832 -16330 17842 -16278
rect 17894 -16330 17904 -16278
rect 17832 -16334 17904 -16330
rect 16096 -16626 16584 -16620
rect 16096 -16660 16143 -16626
rect 16177 -16660 16215 -16626
rect 16249 -16660 16287 -16626
rect 16321 -16660 16359 -16626
rect 16393 -16660 16431 -16626
rect 16465 -16660 16503 -16626
rect 16537 -16660 16584 -16626
rect 16096 -16666 16584 -16660
rect 17114 -16626 17602 -16620
rect 17114 -16660 17161 -16626
rect 17195 -16660 17233 -16626
rect 17267 -16660 17305 -16626
rect 17339 -16660 17377 -16626
rect 17411 -16660 17449 -16626
rect 17483 -16660 17521 -16626
rect 17555 -16660 17602 -16626
rect 17114 -16666 17602 -16660
rect 15800 -16758 15814 -16729
rect 14830 -16763 14836 -16762
rect 14790 -16801 14836 -16763
rect 14790 -16835 14796 -16801
rect 14830 -16835 14836 -16801
rect 14790 -16873 14836 -16835
rect 14790 -16907 14796 -16873
rect 14830 -16907 14836 -16873
rect 14790 -16945 14836 -16907
rect 14790 -16979 14796 -16945
rect 14830 -16979 14836 -16945
rect 14790 -17017 14836 -16979
rect 14790 -17051 14796 -17017
rect 14830 -17051 14836 -17017
rect 14790 -17089 14836 -17051
rect 14790 -17123 14796 -17089
rect 14830 -17123 14836 -17089
rect 14790 -17161 14836 -17123
rect 14790 -17195 14796 -17161
rect 14830 -17195 14836 -17161
rect 14790 -17233 14836 -17195
rect 14790 -17234 14796 -17233
rect 13772 -17298 13818 -17267
rect 14782 -17267 14796 -17234
rect 14830 -17234 14836 -17233
rect 15808 -16763 15814 -16758
rect 15848 -16758 15860 -16729
rect 16826 -16729 16872 -16698
rect 15848 -16763 15854 -16758
rect 15808 -16801 15854 -16763
rect 15808 -16835 15814 -16801
rect 15848 -16835 15854 -16801
rect 15808 -16873 15854 -16835
rect 15808 -16907 15814 -16873
rect 15848 -16907 15854 -16873
rect 15808 -16945 15854 -16907
rect 15808 -16979 15814 -16945
rect 15848 -16979 15854 -16945
rect 15808 -17017 15854 -16979
rect 15808 -17051 15814 -17017
rect 15848 -17051 15854 -17017
rect 15808 -17089 15854 -17051
rect 15808 -17123 15814 -17089
rect 15848 -17123 15854 -17089
rect 15808 -17161 15854 -17123
rect 15808 -17195 15814 -17161
rect 15848 -17195 15854 -17161
rect 15808 -17233 15854 -17195
rect 14830 -17267 14842 -17234
rect 15808 -17254 15814 -17233
rect 13042 -17336 13530 -17330
rect 13042 -17370 13089 -17336
rect 13123 -17370 13161 -17336
rect 13195 -17370 13233 -17336
rect 13267 -17370 13305 -17336
rect 13339 -17370 13377 -17336
rect 13411 -17370 13449 -17336
rect 13483 -17370 13530 -17336
rect 13042 -17376 13530 -17370
rect 14060 -17336 14548 -17330
rect 14060 -17370 14107 -17336
rect 14141 -17370 14179 -17336
rect 14213 -17370 14251 -17336
rect 14285 -17370 14323 -17336
rect 14357 -17370 14395 -17336
rect 14429 -17370 14467 -17336
rect 14501 -17370 14548 -17336
rect 14060 -17376 14548 -17370
rect 12742 -17522 12814 -17518
rect 12742 -17574 12752 -17522
rect 12804 -17574 12814 -17522
rect 12742 -17578 12814 -17574
rect 13262 -17574 13322 -17376
rect 14270 -17574 14330 -17376
rect 14782 -17518 14842 -17267
rect 15800 -17267 15814 -17254
rect 15848 -17254 15854 -17233
rect 16826 -16763 16832 -16729
rect 16866 -16763 16872 -16729
rect 16826 -16801 16872 -16763
rect 17838 -16729 17898 -16334
rect 18352 -16620 18412 -16142
rect 18854 -16274 18914 -16033
rect 19876 -16033 19888 -15999
rect 19922 -16033 19936 -15999
rect 19152 -16102 19640 -16096
rect 19152 -16136 19199 -16102
rect 19233 -16136 19271 -16102
rect 19305 -16136 19343 -16102
rect 19377 -16136 19415 -16102
rect 19449 -16136 19487 -16102
rect 19521 -16136 19559 -16102
rect 19593 -16136 19640 -16102
rect 19152 -16142 19368 -16136
rect 19428 -16142 19640 -16136
rect 19876 -16170 19936 -16033
rect 20890 -15999 20950 -15994
rect 20890 -16033 20906 -15999
rect 20940 -16033 20950 -15999
rect 20170 -16102 20658 -16096
rect 20170 -16136 20217 -16102
rect 20251 -16136 20289 -16102
rect 20323 -16136 20361 -16102
rect 20395 -16136 20433 -16102
rect 20467 -16136 20505 -16102
rect 20539 -16136 20577 -16102
rect 20611 -16136 20658 -16102
rect 20170 -16142 20658 -16136
rect 19870 -16174 19942 -16170
rect 19870 -16226 19880 -16174
rect 19932 -16226 19942 -16174
rect 19870 -16230 19942 -16226
rect 20890 -16274 20950 -16033
rect 21918 -15999 21964 -15961
rect 22936 -15567 22982 -15529
rect 22936 -15601 22942 -15567
rect 22976 -15601 22982 -15567
rect 22936 -15639 22982 -15601
rect 22936 -15673 22942 -15639
rect 22976 -15673 22982 -15639
rect 22936 -15711 22982 -15673
rect 22936 -15745 22942 -15711
rect 22976 -15745 22982 -15711
rect 22936 -15783 22982 -15745
rect 22936 -15817 22942 -15783
rect 22976 -15817 22982 -15783
rect 22936 -15855 22982 -15817
rect 22936 -15889 22942 -15855
rect 22976 -15889 22982 -15855
rect 22936 -15927 22982 -15889
rect 22936 -15961 22942 -15927
rect 22976 -15961 22982 -15927
rect 22936 -15970 22982 -15961
rect 21918 -16033 21924 -15999
rect 21958 -16033 21964 -15999
rect 22942 -15999 22976 -15970
rect 21918 -16064 21964 -16033
rect 22932 -16033 22942 -16008
rect 22976 -16033 22992 -16008
rect 21188 -16102 21676 -16096
rect 21188 -16136 21235 -16102
rect 21269 -16136 21307 -16102
rect 21341 -16136 21379 -16102
rect 21413 -16136 21451 -16102
rect 21485 -16136 21523 -16102
rect 21557 -16136 21595 -16102
rect 21629 -16136 21676 -16102
rect 21188 -16142 21676 -16136
rect 22206 -16102 22694 -16096
rect 22206 -16136 22253 -16102
rect 22287 -16136 22325 -16102
rect 22359 -16136 22397 -16102
rect 22431 -16136 22469 -16102
rect 22503 -16136 22541 -16102
rect 22575 -16136 22613 -16102
rect 22647 -16136 22694 -16102
rect 22206 -16142 22694 -16136
rect 18848 -16278 18920 -16274
rect 18848 -16330 18858 -16278
rect 18910 -16330 18920 -16278
rect 18848 -16334 18920 -16330
rect 20884 -16278 20956 -16274
rect 20884 -16330 20894 -16278
rect 20946 -16330 20956 -16278
rect 20884 -16334 20956 -16330
rect 21380 -16620 21440 -16142
rect 22932 -16178 22992 -16033
rect 22932 -16238 23222 -16178
rect 22418 -16544 22986 -16484
rect 22418 -16620 22478 -16544
rect 18132 -16626 18620 -16620
rect 18132 -16660 18179 -16626
rect 18213 -16660 18251 -16626
rect 18285 -16660 18323 -16626
rect 18357 -16660 18395 -16626
rect 18429 -16660 18467 -16626
rect 18501 -16660 18539 -16626
rect 18573 -16660 18620 -16626
rect 18132 -16666 18620 -16660
rect 19150 -16626 19638 -16620
rect 19150 -16660 19197 -16626
rect 19231 -16660 19269 -16626
rect 19303 -16660 19341 -16626
rect 19375 -16660 19413 -16626
rect 19447 -16660 19485 -16626
rect 19519 -16660 19557 -16626
rect 19591 -16660 19638 -16626
rect 19150 -16666 19638 -16660
rect 20168 -16626 20656 -16620
rect 20168 -16660 20215 -16626
rect 20249 -16660 20287 -16626
rect 20321 -16660 20359 -16626
rect 20393 -16660 20431 -16626
rect 20465 -16660 20503 -16626
rect 20537 -16660 20575 -16626
rect 20609 -16660 20656 -16626
rect 20168 -16666 20656 -16660
rect 21186 -16626 21674 -16620
rect 21186 -16660 21233 -16626
rect 21267 -16660 21305 -16626
rect 21339 -16660 21377 -16626
rect 21411 -16660 21449 -16626
rect 21483 -16660 21521 -16626
rect 21555 -16660 21593 -16626
rect 21627 -16660 21674 -16626
rect 21186 -16666 21674 -16660
rect 22204 -16626 22692 -16620
rect 22204 -16660 22251 -16626
rect 22285 -16660 22323 -16626
rect 22357 -16660 22395 -16626
rect 22429 -16660 22467 -16626
rect 22501 -16660 22539 -16626
rect 22573 -16660 22611 -16626
rect 22645 -16660 22692 -16626
rect 22204 -16666 22692 -16660
rect 17838 -16763 17850 -16729
rect 17884 -16763 17898 -16729
rect 17838 -16768 17898 -16763
rect 18862 -16729 18908 -16698
rect 18862 -16763 18868 -16729
rect 18902 -16763 18908 -16729
rect 16826 -16835 16832 -16801
rect 16866 -16835 16872 -16801
rect 16826 -16873 16872 -16835
rect 16826 -16907 16832 -16873
rect 16866 -16907 16872 -16873
rect 16826 -16945 16872 -16907
rect 16826 -16979 16832 -16945
rect 16866 -16979 16872 -16945
rect 16826 -17017 16872 -16979
rect 16826 -17051 16832 -17017
rect 16866 -17051 16872 -17017
rect 16826 -17089 16872 -17051
rect 16826 -17123 16832 -17089
rect 16866 -17123 16872 -17089
rect 16826 -17161 16872 -17123
rect 16826 -17195 16832 -17161
rect 16866 -17195 16872 -17161
rect 16826 -17233 16872 -17195
rect 16826 -17250 16832 -17233
rect 15848 -17267 15860 -17254
rect 15078 -17336 15566 -17330
rect 15078 -17370 15125 -17336
rect 15159 -17370 15197 -17336
rect 15231 -17370 15269 -17336
rect 15303 -17370 15341 -17336
rect 15375 -17370 15413 -17336
rect 15447 -17370 15485 -17336
rect 15519 -17370 15566 -17336
rect 15078 -17376 15566 -17370
rect 12740 -17634 12812 -17630
rect 12740 -17686 12750 -17634
rect 12802 -17686 12812 -17634
rect 12740 -17690 12812 -17686
rect 13262 -17634 14330 -17574
rect 14776 -17522 14848 -17518
rect 14776 -17574 14786 -17522
rect 14838 -17574 14848 -17522
rect 14776 -17578 14848 -17574
rect 14972 -17526 15044 -17522
rect 14972 -17578 14982 -17526
rect 15034 -17578 15044 -17526
rect 14972 -17582 15044 -17578
rect 12024 -17860 12512 -17854
rect 12024 -17894 12071 -17860
rect 12105 -17894 12143 -17860
rect 12177 -17894 12215 -17860
rect 12249 -17894 12287 -17860
rect 12321 -17894 12359 -17860
rect 12393 -17894 12431 -17860
rect 12465 -17894 12512 -17860
rect 12024 -17900 12512 -17894
rect 11726 -17992 11742 -17963
rect 10710 -18012 10770 -17997
rect 11736 -17997 11742 -17992
rect 11776 -17992 11786 -17963
rect 12746 -17963 12806 -17690
rect 13262 -17854 13322 -17634
rect 13760 -17744 13832 -17740
rect 13760 -17796 13770 -17744
rect 13822 -17796 13832 -17744
rect 13760 -17800 13832 -17796
rect 13042 -17860 13530 -17854
rect 13042 -17894 13089 -17860
rect 13123 -17894 13161 -17860
rect 13195 -17894 13233 -17860
rect 13267 -17894 13305 -17860
rect 13339 -17894 13377 -17860
rect 13411 -17894 13449 -17860
rect 13483 -17894 13530 -17860
rect 13042 -17900 13530 -17894
rect 11776 -17997 11782 -17992
rect 12746 -17994 12760 -17963
rect 9700 -18069 9706 -18035
rect 9740 -18069 9746 -18035
rect 9700 -18107 9746 -18069
rect 9700 -18141 9706 -18107
rect 9740 -18141 9746 -18107
rect 9700 -18179 9746 -18141
rect 9700 -18213 9706 -18179
rect 9740 -18213 9746 -18179
rect 9700 -18251 9746 -18213
rect 9700 -18285 9706 -18251
rect 9740 -18285 9746 -18251
rect 9700 -18323 9746 -18285
rect 9700 -18357 9706 -18323
rect 9740 -18357 9746 -18323
rect 9700 -18395 9746 -18357
rect 9700 -18429 9706 -18395
rect 9740 -18429 9746 -18395
rect 9700 -18467 9746 -18429
rect 9700 -18501 9706 -18467
rect 9740 -18501 9746 -18467
rect 9700 -18532 9746 -18501
rect 10718 -18035 10764 -18012
rect 10718 -18069 10724 -18035
rect 10758 -18069 10764 -18035
rect 10718 -18107 10764 -18069
rect 10718 -18141 10724 -18107
rect 10758 -18141 10764 -18107
rect 10718 -18179 10764 -18141
rect 10718 -18213 10724 -18179
rect 10758 -18213 10764 -18179
rect 10718 -18251 10764 -18213
rect 10718 -18285 10724 -18251
rect 10758 -18285 10764 -18251
rect 10718 -18323 10764 -18285
rect 10718 -18357 10724 -18323
rect 10758 -18357 10764 -18323
rect 10718 -18395 10764 -18357
rect 10718 -18429 10724 -18395
rect 10758 -18429 10764 -18395
rect 10718 -18467 10764 -18429
rect 10718 -18501 10724 -18467
rect 10758 -18501 10764 -18467
rect 10718 -18532 10764 -18501
rect 11736 -18035 11782 -17997
rect 11736 -18069 11742 -18035
rect 11776 -18069 11782 -18035
rect 11736 -18107 11782 -18069
rect 11736 -18141 11742 -18107
rect 11776 -18141 11782 -18107
rect 11736 -18179 11782 -18141
rect 11736 -18213 11742 -18179
rect 11776 -18213 11782 -18179
rect 11736 -18251 11782 -18213
rect 11736 -18285 11742 -18251
rect 11776 -18285 11782 -18251
rect 11736 -18323 11782 -18285
rect 11736 -18357 11742 -18323
rect 11776 -18357 11782 -18323
rect 11736 -18395 11782 -18357
rect 11736 -18429 11742 -18395
rect 11776 -18429 11782 -18395
rect 11736 -18467 11782 -18429
rect 11736 -18501 11742 -18467
rect 11776 -18501 11782 -18467
rect 11736 -18532 11782 -18501
rect 12754 -17997 12760 -17994
rect 12794 -17994 12806 -17963
rect 13766 -17963 13826 -17800
rect 14270 -17854 14330 -17634
rect 14776 -17634 14848 -17630
rect 14776 -17686 14786 -17634
rect 14838 -17686 14848 -17634
rect 14776 -17690 14848 -17686
rect 14060 -17860 14548 -17854
rect 14060 -17894 14107 -17860
rect 14141 -17894 14179 -17860
rect 14213 -17894 14251 -17860
rect 14285 -17894 14323 -17860
rect 14357 -17894 14395 -17860
rect 14429 -17894 14467 -17860
rect 14501 -17894 14548 -17860
rect 14060 -17900 14548 -17894
rect 13766 -17982 13778 -17963
rect 12794 -17997 12800 -17994
rect 12754 -18035 12800 -17997
rect 12754 -18069 12760 -18035
rect 12794 -18069 12800 -18035
rect 12754 -18107 12800 -18069
rect 12754 -18141 12760 -18107
rect 12794 -18141 12800 -18107
rect 12754 -18179 12800 -18141
rect 12754 -18213 12760 -18179
rect 12794 -18213 12800 -18179
rect 12754 -18251 12800 -18213
rect 12754 -18285 12760 -18251
rect 12794 -18285 12800 -18251
rect 12754 -18323 12800 -18285
rect 12754 -18357 12760 -18323
rect 12794 -18357 12800 -18323
rect 12754 -18395 12800 -18357
rect 12754 -18429 12760 -18395
rect 12794 -18429 12800 -18395
rect 12754 -18467 12800 -18429
rect 12754 -18501 12760 -18467
rect 12794 -18501 12800 -18467
rect 13772 -17997 13778 -17982
rect 13812 -17982 13826 -17963
rect 14782 -17963 14842 -17690
rect 14978 -17740 15038 -17582
rect 15272 -17738 15332 -17376
rect 15800 -17414 15860 -17267
rect 16816 -17267 16832 -17250
rect 16866 -17250 16872 -17233
rect 17844 -16801 17890 -16768
rect 17844 -16835 17850 -16801
rect 17884 -16835 17890 -16801
rect 17844 -16873 17890 -16835
rect 17844 -16907 17850 -16873
rect 17884 -16907 17890 -16873
rect 17844 -16945 17890 -16907
rect 17844 -16979 17850 -16945
rect 17884 -16979 17890 -16945
rect 17844 -17017 17890 -16979
rect 17844 -17051 17850 -17017
rect 17884 -17051 17890 -17017
rect 17844 -17089 17890 -17051
rect 17844 -17123 17850 -17089
rect 17884 -17123 17890 -17089
rect 17844 -17161 17890 -17123
rect 17844 -17195 17850 -17161
rect 17884 -17195 17890 -17161
rect 17844 -17233 17890 -17195
rect 18862 -16801 18908 -16763
rect 18862 -16835 18868 -16801
rect 18902 -16835 18908 -16801
rect 18862 -16873 18908 -16835
rect 18862 -16907 18868 -16873
rect 18902 -16907 18908 -16873
rect 18862 -16945 18908 -16907
rect 18862 -16979 18868 -16945
rect 18902 -16979 18908 -16945
rect 18862 -17017 18908 -16979
rect 18862 -17051 18868 -17017
rect 18902 -17051 18908 -17017
rect 18862 -17089 18908 -17051
rect 18862 -17123 18868 -17089
rect 18902 -17123 18908 -17089
rect 18862 -17161 18908 -17123
rect 18862 -17195 18868 -17161
rect 18902 -17195 18908 -17161
rect 18862 -17230 18908 -17195
rect 19880 -16729 19926 -16698
rect 19880 -16763 19886 -16729
rect 19920 -16763 19926 -16729
rect 19880 -16801 19926 -16763
rect 19880 -16835 19886 -16801
rect 19920 -16835 19926 -16801
rect 19880 -16873 19926 -16835
rect 19880 -16907 19886 -16873
rect 19920 -16907 19926 -16873
rect 19880 -16945 19926 -16907
rect 19880 -16979 19886 -16945
rect 19920 -16979 19926 -16945
rect 19880 -17017 19926 -16979
rect 19880 -17051 19886 -17017
rect 19920 -17051 19926 -17017
rect 19880 -17089 19926 -17051
rect 19880 -17123 19886 -17089
rect 19920 -17123 19926 -17089
rect 19880 -17161 19926 -17123
rect 19880 -17195 19886 -17161
rect 19920 -17195 19926 -17161
rect 17844 -17240 17850 -17233
rect 16866 -17267 16876 -17250
rect 16096 -17336 16584 -17330
rect 16096 -17370 16143 -17336
rect 16177 -17370 16215 -17336
rect 16249 -17370 16287 -17336
rect 16321 -17370 16359 -17336
rect 16393 -17370 16431 -17336
rect 16465 -17370 16503 -17336
rect 16537 -17370 16584 -17336
rect 16096 -17376 16584 -17370
rect 15794 -17418 15866 -17414
rect 15794 -17470 15804 -17418
rect 15856 -17470 15866 -17418
rect 15794 -17474 15866 -17470
rect 14972 -17744 15044 -17740
rect 14972 -17796 14982 -17744
rect 15034 -17796 15044 -17744
rect 14972 -17800 15044 -17796
rect 15266 -17742 15338 -17738
rect 15266 -17794 15276 -17742
rect 15328 -17794 15338 -17742
rect 15266 -17798 15338 -17794
rect 15272 -17854 15332 -17798
rect 15078 -17860 15566 -17854
rect 15078 -17894 15125 -17860
rect 15159 -17894 15197 -17860
rect 15231 -17894 15269 -17860
rect 15303 -17894 15341 -17860
rect 15375 -17894 15413 -17860
rect 15447 -17894 15485 -17860
rect 15519 -17894 15566 -17860
rect 15078 -17900 15566 -17894
rect 13812 -17997 13818 -17982
rect 14782 -17988 14796 -17963
rect 13772 -18035 13818 -17997
rect 13772 -18069 13778 -18035
rect 13812 -18069 13818 -18035
rect 13772 -18107 13818 -18069
rect 13772 -18141 13778 -18107
rect 13812 -18141 13818 -18107
rect 13772 -18179 13818 -18141
rect 13772 -18213 13778 -18179
rect 13812 -18213 13818 -18179
rect 13772 -18251 13818 -18213
rect 13772 -18285 13778 -18251
rect 13812 -18285 13818 -18251
rect 13772 -18323 13818 -18285
rect 13772 -18357 13778 -18323
rect 13812 -18357 13818 -18323
rect 13772 -18395 13818 -18357
rect 13772 -18429 13778 -18395
rect 13812 -18429 13818 -18395
rect 13772 -18467 13818 -18429
rect 13772 -18474 13778 -18467
rect 12754 -18532 12800 -18501
rect 13766 -18501 13778 -18474
rect 13812 -18474 13818 -18467
rect 14790 -17997 14796 -17988
rect 14830 -17988 14842 -17963
rect 15800 -17963 15860 -17474
rect 16302 -17732 16362 -17376
rect 16816 -17630 16876 -17267
rect 17836 -17267 17850 -17240
rect 17884 -17240 17890 -17233
rect 18854 -17233 18914 -17230
rect 17884 -17267 17896 -17240
rect 17114 -17336 17602 -17330
rect 17114 -17370 17161 -17336
rect 17195 -17370 17233 -17336
rect 17267 -17370 17305 -17336
rect 17339 -17370 17377 -17336
rect 17411 -17370 17449 -17336
rect 17483 -17370 17521 -17336
rect 17555 -17370 17602 -17336
rect 17114 -17376 17602 -17370
rect 16810 -17634 16882 -17630
rect 16810 -17686 16820 -17634
rect 16872 -17686 16882 -17634
rect 16810 -17690 16882 -17686
rect 16300 -17742 16362 -17732
rect 16300 -17794 16304 -17742
rect 16356 -17794 16362 -17742
rect 16300 -17804 16362 -17794
rect 16812 -17748 16884 -17744
rect 16812 -17800 16822 -17748
rect 16874 -17800 16884 -17748
rect 16812 -17804 16884 -17800
rect 16302 -17854 16362 -17804
rect 16096 -17860 16584 -17854
rect 16096 -17894 16143 -17860
rect 16177 -17894 16215 -17860
rect 16249 -17894 16287 -17860
rect 16321 -17894 16359 -17860
rect 16393 -17894 16431 -17860
rect 16465 -17894 16503 -17860
rect 16537 -17894 16584 -17860
rect 16096 -17900 16584 -17894
rect 15800 -17988 15814 -17963
rect 14830 -17997 14836 -17988
rect 14790 -18035 14836 -17997
rect 14790 -18069 14796 -18035
rect 14830 -18069 14836 -18035
rect 14790 -18107 14836 -18069
rect 14790 -18141 14796 -18107
rect 14830 -18141 14836 -18107
rect 14790 -18179 14836 -18141
rect 14790 -18213 14796 -18179
rect 14830 -18213 14836 -18179
rect 14790 -18251 14836 -18213
rect 14790 -18285 14796 -18251
rect 14830 -18285 14836 -18251
rect 14790 -18323 14836 -18285
rect 14790 -18357 14796 -18323
rect 14830 -18357 14836 -18323
rect 14790 -18395 14836 -18357
rect 14790 -18429 14796 -18395
rect 14830 -18429 14836 -18395
rect 14790 -18467 14836 -18429
rect 13812 -18501 13826 -18474
rect 7952 -18570 8440 -18564
rect 7952 -18604 7999 -18570
rect 8033 -18604 8071 -18570
rect 8105 -18604 8143 -18570
rect 8177 -18604 8215 -18570
rect 8249 -18604 8287 -18570
rect 8321 -18604 8359 -18570
rect 8393 -18604 8440 -18570
rect 7952 -18610 8440 -18604
rect 8970 -18570 9458 -18564
rect 8970 -18604 9017 -18570
rect 9051 -18604 9089 -18570
rect 9123 -18604 9161 -18570
rect 9195 -18604 9233 -18570
rect 9267 -18604 9305 -18570
rect 9339 -18604 9377 -18570
rect 9411 -18604 9458 -18570
rect 8970 -18610 9458 -18604
rect 9988 -18570 10476 -18564
rect 9988 -18604 10035 -18570
rect 10069 -18604 10107 -18570
rect 10141 -18604 10179 -18570
rect 10213 -18604 10251 -18570
rect 10285 -18604 10323 -18570
rect 10357 -18604 10395 -18570
rect 10429 -18604 10476 -18570
rect 9988 -18610 10476 -18604
rect 11006 -18570 11494 -18564
rect 11006 -18604 11053 -18570
rect 11087 -18604 11125 -18570
rect 11159 -18604 11197 -18570
rect 11231 -18604 11269 -18570
rect 11303 -18604 11341 -18570
rect 11375 -18604 11413 -18570
rect 11447 -18604 11494 -18570
rect 11006 -18610 11494 -18604
rect 12024 -18570 12512 -18564
rect 12024 -18604 12071 -18570
rect 12105 -18604 12143 -18570
rect 12177 -18604 12215 -18570
rect 12249 -18604 12287 -18570
rect 12321 -18604 12359 -18570
rect 12393 -18604 12431 -18570
rect 12465 -18604 12512 -18570
rect 12024 -18610 12238 -18604
rect 12240 -18610 12512 -18604
rect 13042 -18570 13530 -18564
rect 13042 -18604 13089 -18570
rect 13123 -18604 13161 -18570
rect 13195 -18604 13233 -18570
rect 13267 -18604 13305 -18570
rect 13339 -18604 13377 -18570
rect 13411 -18604 13449 -18570
rect 13483 -18604 13530 -18570
rect 13042 -18610 13264 -18604
rect 13268 -18610 13530 -18604
rect 7652 -18674 7724 -18670
rect 7652 -18726 7662 -18674
rect 7714 -18726 7724 -18674
rect 7652 -18730 7724 -18726
rect 5614 -18934 5686 -18930
rect 6122 -18884 6194 -18880
rect 4598 -18978 4670 -18974
rect 4598 -19030 4608 -18978
rect 4660 -19030 4670 -18978
rect 4598 -19034 4670 -19030
rect 3880 -19092 4368 -19086
rect 3880 -19126 3927 -19092
rect 3961 -19126 3999 -19092
rect 4033 -19126 4071 -19092
rect 4105 -19126 4143 -19092
rect 4177 -19126 4215 -19092
rect 4249 -19126 4287 -19092
rect 4321 -19126 4368 -19092
rect 3880 -19132 4368 -19126
rect 3584 -19214 3598 -19195
rect 2574 -19267 2620 -19229
rect 2574 -19301 2580 -19267
rect 2614 -19301 2620 -19267
rect 2574 -19339 2620 -19301
rect 2574 -19373 2580 -19339
rect 2614 -19373 2620 -19339
rect 2574 -19411 2620 -19373
rect 2574 -19445 2580 -19411
rect 2614 -19445 2620 -19411
rect 2574 -19483 2620 -19445
rect 2574 -19517 2580 -19483
rect 2614 -19517 2620 -19483
rect 2574 -19555 2620 -19517
rect 2574 -19589 2580 -19555
rect 2614 -19589 2620 -19555
rect 2574 -19627 2620 -19589
rect 2574 -19661 2580 -19627
rect 2614 -19661 2620 -19627
rect 2574 -19699 2620 -19661
rect 2574 -19706 2580 -19699
rect 2564 -19733 2580 -19706
rect 2614 -19706 2620 -19699
rect 3592 -19229 3598 -19214
rect 3632 -19214 3644 -19195
rect 4604 -19195 4664 -19034
rect 4898 -19092 5386 -19086
rect 4898 -19126 4945 -19092
rect 4979 -19126 5017 -19092
rect 5051 -19126 5089 -19092
rect 5123 -19126 5161 -19092
rect 5195 -19126 5233 -19092
rect 5267 -19126 5305 -19092
rect 5339 -19126 5386 -19092
rect 4898 -19132 5386 -19126
rect 3632 -19229 3638 -19214
rect 4604 -19216 4616 -19195
rect 3592 -19267 3638 -19229
rect 3592 -19301 3598 -19267
rect 3632 -19301 3638 -19267
rect 3592 -19339 3638 -19301
rect 3592 -19373 3598 -19339
rect 3632 -19373 3638 -19339
rect 3592 -19411 3638 -19373
rect 3592 -19445 3598 -19411
rect 3632 -19445 3638 -19411
rect 3592 -19483 3638 -19445
rect 3592 -19517 3598 -19483
rect 3632 -19517 3638 -19483
rect 3592 -19555 3638 -19517
rect 3592 -19589 3598 -19555
rect 3632 -19589 3638 -19555
rect 3592 -19627 3638 -19589
rect 3592 -19661 3598 -19627
rect 3632 -19661 3638 -19627
rect 3592 -19699 3638 -19661
rect 2614 -19733 2624 -19706
rect 3592 -19710 3598 -19699
rect 2564 -19914 2624 -19733
rect 3582 -19733 3598 -19710
rect 3632 -19710 3638 -19699
rect 4610 -19229 4616 -19216
rect 4650 -19216 4664 -19195
rect 5620 -19195 5680 -18934
rect 6122 -18936 6132 -18884
rect 6184 -18936 6194 -18884
rect 6122 -18940 6194 -18936
rect 7144 -18884 7216 -18880
rect 7144 -18936 7154 -18884
rect 7206 -18936 7216 -18884
rect 7144 -18940 7216 -18936
rect 6632 -18978 6704 -18974
rect 6632 -19030 6642 -18978
rect 6694 -19030 6704 -18978
rect 6632 -19034 6704 -19030
rect 5916 -19092 6404 -19086
rect 5916 -19126 5963 -19092
rect 5997 -19126 6035 -19092
rect 6069 -19126 6107 -19092
rect 6141 -19126 6179 -19092
rect 6213 -19126 6251 -19092
rect 6285 -19126 6323 -19092
rect 6357 -19126 6404 -19092
rect 5916 -19132 6404 -19126
rect 4650 -19229 4656 -19216
rect 5620 -19228 5634 -19195
rect 4610 -19267 4656 -19229
rect 4610 -19301 4616 -19267
rect 4650 -19301 4656 -19267
rect 4610 -19339 4656 -19301
rect 4610 -19373 4616 -19339
rect 4650 -19373 4656 -19339
rect 4610 -19411 4656 -19373
rect 4610 -19445 4616 -19411
rect 4650 -19445 4656 -19411
rect 4610 -19483 4656 -19445
rect 4610 -19517 4616 -19483
rect 4650 -19517 4656 -19483
rect 4610 -19555 4656 -19517
rect 4610 -19589 4616 -19555
rect 4650 -19589 4656 -19555
rect 4610 -19627 4656 -19589
rect 4610 -19661 4616 -19627
rect 4650 -19661 4656 -19627
rect 4610 -19699 4656 -19661
rect 3632 -19733 3642 -19710
rect 2862 -19802 3350 -19796
rect 2862 -19836 2909 -19802
rect 2943 -19836 2981 -19802
rect 3015 -19836 3053 -19802
rect 3087 -19836 3125 -19802
rect 3159 -19836 3197 -19802
rect 3231 -19836 3269 -19802
rect 3303 -19836 3350 -19802
rect 2862 -19842 3350 -19836
rect 3076 -19914 3136 -19842
rect 3582 -19914 3642 -19733
rect 4610 -19733 4616 -19699
rect 4650 -19733 4656 -19699
rect 4610 -19764 4656 -19733
rect 5628 -19229 5634 -19228
rect 5668 -19228 5680 -19195
rect 6638 -19195 6698 -19034
rect 7150 -19086 7210 -18940
rect 6934 -19092 7422 -19086
rect 6934 -19126 6981 -19092
rect 7015 -19126 7053 -19092
rect 7087 -19126 7125 -19092
rect 7159 -19126 7197 -19092
rect 7231 -19126 7269 -19092
rect 7303 -19126 7341 -19092
rect 7375 -19126 7422 -19092
rect 6934 -19132 7422 -19126
rect 6638 -19220 6652 -19195
rect 5668 -19229 5674 -19228
rect 5628 -19267 5674 -19229
rect 5628 -19301 5634 -19267
rect 5668 -19301 5674 -19267
rect 5628 -19339 5674 -19301
rect 5628 -19373 5634 -19339
rect 5668 -19373 5674 -19339
rect 5628 -19411 5674 -19373
rect 5628 -19445 5634 -19411
rect 5668 -19445 5674 -19411
rect 5628 -19483 5674 -19445
rect 5628 -19517 5634 -19483
rect 5668 -19517 5674 -19483
rect 5628 -19555 5674 -19517
rect 5628 -19589 5634 -19555
rect 5668 -19589 5674 -19555
rect 5628 -19627 5674 -19589
rect 5628 -19661 5634 -19627
rect 5668 -19661 5674 -19627
rect 5628 -19699 5674 -19661
rect 5628 -19733 5634 -19699
rect 5668 -19733 5674 -19699
rect 6646 -19229 6652 -19220
rect 6686 -19220 6698 -19195
rect 7658 -19195 7718 -18730
rect 8164 -18880 8224 -18610
rect 9182 -18772 9242 -18610
rect 10202 -18660 10262 -18610
rect 11202 -18660 11262 -18610
rect 12240 -18660 12300 -18610
rect 13268 -18660 13328 -18610
rect 9684 -18674 9756 -18670
rect 9684 -18726 9694 -18674
rect 9746 -18726 9756 -18674
rect 10202 -18720 13328 -18660
rect 9684 -18730 9756 -18726
rect 9176 -18776 9248 -18772
rect 9176 -18828 9186 -18776
rect 9238 -18828 9248 -18776
rect 9176 -18832 9248 -18828
rect 8158 -18884 8230 -18880
rect 8158 -18936 8168 -18884
rect 8220 -18936 8230 -18884
rect 8158 -18940 8230 -18936
rect 9176 -18884 9248 -18880
rect 9176 -18936 9186 -18884
rect 9238 -18936 9248 -18884
rect 9176 -18940 9248 -18936
rect 8164 -19086 8224 -18940
rect 8668 -18978 8740 -18974
rect 8668 -19030 8678 -18978
rect 8730 -19030 8740 -18978
rect 8668 -19034 8740 -19030
rect 7952 -19092 8440 -19086
rect 7952 -19126 7999 -19092
rect 8033 -19126 8071 -19092
rect 8105 -19126 8143 -19092
rect 8177 -19126 8215 -19092
rect 8249 -19126 8287 -19092
rect 8321 -19126 8359 -19092
rect 8393 -19126 8440 -19092
rect 7952 -19132 8440 -19126
rect 6686 -19229 6692 -19220
rect 6646 -19267 6692 -19229
rect 6646 -19301 6652 -19267
rect 6686 -19301 6692 -19267
rect 6646 -19339 6692 -19301
rect 6646 -19373 6652 -19339
rect 6686 -19373 6692 -19339
rect 6646 -19411 6692 -19373
rect 6646 -19445 6652 -19411
rect 6686 -19445 6692 -19411
rect 6646 -19483 6692 -19445
rect 6646 -19517 6652 -19483
rect 6686 -19517 6692 -19483
rect 6646 -19555 6692 -19517
rect 6646 -19589 6652 -19555
rect 6686 -19589 6692 -19555
rect 6646 -19627 6692 -19589
rect 6646 -19661 6652 -19627
rect 6686 -19661 6692 -19627
rect 6646 -19699 6692 -19661
rect 6646 -19716 6652 -19699
rect 5628 -19764 5674 -19733
rect 6638 -19733 6652 -19716
rect 6686 -19716 6692 -19699
rect 7658 -19229 7670 -19195
rect 7704 -19229 7718 -19195
rect 8674 -19195 8734 -19034
rect 9182 -19086 9242 -18940
rect 8970 -19092 9458 -19086
rect 8970 -19126 9017 -19092
rect 9051 -19126 9089 -19092
rect 9123 -19126 9161 -19092
rect 9195 -19126 9233 -19092
rect 9267 -19126 9305 -19092
rect 9339 -19126 9377 -19092
rect 9411 -19126 9458 -19092
rect 8970 -19132 9458 -19126
rect 8674 -19212 8688 -19195
rect 7658 -19267 7718 -19229
rect 7658 -19301 7670 -19267
rect 7704 -19301 7718 -19267
rect 7658 -19339 7718 -19301
rect 7658 -19373 7670 -19339
rect 7704 -19373 7718 -19339
rect 7658 -19411 7718 -19373
rect 7658 -19445 7670 -19411
rect 7704 -19445 7718 -19411
rect 7658 -19483 7718 -19445
rect 7658 -19517 7670 -19483
rect 7704 -19517 7718 -19483
rect 7658 -19555 7718 -19517
rect 7658 -19589 7670 -19555
rect 7704 -19589 7718 -19555
rect 7658 -19627 7718 -19589
rect 7658 -19661 7670 -19627
rect 7704 -19661 7718 -19627
rect 7658 -19699 7718 -19661
rect 6686 -19733 6698 -19716
rect 3880 -19802 4368 -19796
rect 3880 -19836 3927 -19802
rect 3961 -19836 3999 -19802
rect 4033 -19836 4071 -19802
rect 4105 -19836 4143 -19802
rect 4177 -19836 4215 -19802
rect 4249 -19836 4287 -19802
rect 4321 -19836 4368 -19802
rect 3880 -19842 4368 -19836
rect 4898 -19802 5386 -19796
rect 4898 -19836 4945 -19802
rect 4979 -19836 5017 -19802
rect 5051 -19836 5089 -19802
rect 5123 -19836 5161 -19802
rect 5195 -19836 5233 -19802
rect 5267 -19836 5305 -19802
rect 5339 -19836 5386 -19802
rect 4898 -19842 5386 -19836
rect 5916 -19802 6404 -19796
rect 5916 -19836 5963 -19802
rect 5997 -19836 6035 -19802
rect 6069 -19836 6107 -19802
rect 6141 -19836 6179 -19802
rect 6213 -19836 6251 -19802
rect 6285 -19836 6323 -19802
rect 6357 -19836 6404 -19802
rect 5916 -19842 6404 -19836
rect 4086 -19898 4146 -19842
rect 2564 -19974 3642 -19914
rect 4080 -19902 4152 -19898
rect 4080 -19954 4090 -19902
rect 4142 -19954 4152 -19902
rect 4080 -19958 4152 -19954
rect 4990 -19902 5062 -19898
rect 4990 -19954 5000 -19902
rect 5052 -19954 5062 -19902
rect 4990 -19958 5062 -19954
rect 4080 -20118 4152 -20114
rect 4080 -20170 4090 -20118
rect 4142 -20170 4152 -20118
rect 4080 -20174 4152 -20170
rect 4086 -20180 4148 -20174
rect 2448 -20222 2510 -20212
rect 2448 -20274 2454 -20222
rect 2506 -20274 2510 -20222
rect 2448 -20284 2510 -20274
rect 2448 -22462 2508 -20284
rect 4088 -20320 4148 -20180
rect 4996 -20320 5056 -19958
rect 5124 -20118 5184 -19842
rect 5992 -19902 6064 -19898
rect 5992 -19954 6002 -19902
rect 6054 -19954 6064 -19902
rect 5992 -19958 6064 -19954
rect 5124 -20170 5128 -20118
rect 5180 -20170 5184 -20118
rect 5124 -20180 5184 -20170
rect 5998 -20320 6058 -19958
rect 6138 -20114 6198 -19842
rect 6638 -20000 6698 -19733
rect 7658 -19733 7670 -19699
rect 7704 -19733 7718 -19699
rect 6934 -19802 7422 -19796
rect 6934 -19836 6981 -19802
rect 7015 -19836 7053 -19802
rect 7087 -19836 7125 -19802
rect 7159 -19836 7197 -19802
rect 7231 -19836 7269 -19802
rect 7303 -19836 7341 -19802
rect 7375 -19836 7422 -19802
rect 6934 -19842 7126 -19836
rect 7150 -19842 7422 -19836
rect 7150 -19898 7210 -19842
rect 7144 -19902 7216 -19898
rect 7144 -19954 7154 -19902
rect 7206 -19954 7216 -19902
rect 7144 -19958 7216 -19954
rect 6632 -20004 6704 -20000
rect 6632 -20056 6642 -20004
rect 6694 -20056 6704 -20004
rect 6632 -20060 6704 -20056
rect 6132 -20118 6204 -20114
rect 6132 -20170 6142 -20118
rect 6194 -20170 6204 -20118
rect 6132 -20174 6204 -20170
rect 7150 -20320 7210 -19958
rect 2862 -20326 3350 -20320
rect 2862 -20360 2909 -20326
rect 2943 -20360 2981 -20326
rect 3015 -20360 3053 -20326
rect 3087 -20360 3125 -20326
rect 3159 -20360 3197 -20326
rect 3231 -20360 3269 -20326
rect 3303 -20360 3350 -20326
rect 2862 -20366 3350 -20360
rect 3880 -20326 4368 -20320
rect 3880 -20360 3927 -20326
rect 3961 -20360 3999 -20326
rect 4033 -20360 4071 -20326
rect 4105 -20360 4143 -20326
rect 4177 -20360 4215 -20326
rect 4249 -20360 4287 -20326
rect 4321 -20360 4368 -20326
rect 3880 -20366 4368 -20360
rect 4898 -20326 5386 -20320
rect 4898 -20360 4945 -20326
rect 4979 -20360 5017 -20326
rect 5051 -20360 5089 -20326
rect 5123 -20360 5161 -20326
rect 5195 -20360 5233 -20326
rect 5267 -20360 5305 -20326
rect 5339 -20360 5386 -20326
rect 4898 -20366 5386 -20360
rect 5916 -20326 6404 -20320
rect 5916 -20360 5963 -20326
rect 5997 -20360 6035 -20326
rect 6069 -20360 6107 -20326
rect 6141 -20360 6179 -20326
rect 6213 -20360 6251 -20326
rect 6285 -20360 6323 -20326
rect 6357 -20360 6404 -20326
rect 5916 -20366 6404 -20360
rect 6934 -20326 7422 -20320
rect 6934 -20360 6981 -20326
rect 7015 -20360 7053 -20326
rect 7087 -20360 7125 -20326
rect 7159 -20360 7197 -20326
rect 7231 -20360 7269 -20326
rect 7303 -20360 7341 -20326
rect 7375 -20360 7422 -20326
rect 6934 -20366 7422 -20360
rect 2574 -20429 2620 -20398
rect 2574 -20463 2580 -20429
rect 2614 -20463 2620 -20429
rect 2574 -20501 2620 -20463
rect 2574 -20535 2580 -20501
rect 2614 -20535 2620 -20501
rect 2574 -20573 2620 -20535
rect 2574 -20607 2580 -20573
rect 2614 -20607 2620 -20573
rect 2574 -20645 2620 -20607
rect 2574 -20679 2580 -20645
rect 2614 -20679 2620 -20645
rect 2574 -20717 2620 -20679
rect 2574 -20751 2580 -20717
rect 2614 -20751 2620 -20717
rect 2574 -20789 2620 -20751
rect 2574 -20823 2580 -20789
rect 2614 -20823 2620 -20789
rect 2574 -20861 2620 -20823
rect 2574 -20895 2580 -20861
rect 2614 -20895 2620 -20861
rect 2574 -20933 2620 -20895
rect 2574 -20948 2580 -20933
rect 2568 -20967 2580 -20948
rect 2614 -20948 2620 -20933
rect 3592 -20429 3638 -20398
rect 3592 -20463 3598 -20429
rect 3632 -20463 3638 -20429
rect 3592 -20501 3638 -20463
rect 3592 -20535 3598 -20501
rect 3632 -20535 3638 -20501
rect 3592 -20573 3638 -20535
rect 3592 -20607 3598 -20573
rect 3632 -20607 3638 -20573
rect 3592 -20645 3638 -20607
rect 3592 -20679 3598 -20645
rect 3632 -20679 3638 -20645
rect 3592 -20717 3638 -20679
rect 3592 -20751 3598 -20717
rect 3632 -20751 3638 -20717
rect 3592 -20789 3638 -20751
rect 3592 -20823 3598 -20789
rect 3632 -20823 3638 -20789
rect 3592 -20861 3638 -20823
rect 3592 -20895 3598 -20861
rect 3632 -20895 3638 -20861
rect 3592 -20933 3638 -20895
rect 3592 -20948 3598 -20933
rect 2614 -20967 2628 -20948
rect 2568 -21116 2628 -20967
rect 3586 -20967 3598 -20948
rect 3632 -20948 3638 -20933
rect 4610 -20429 4656 -20398
rect 4610 -20463 4616 -20429
rect 4650 -20463 4656 -20429
rect 4610 -20501 4656 -20463
rect 4610 -20535 4616 -20501
rect 4650 -20535 4656 -20501
rect 4610 -20573 4656 -20535
rect 4610 -20607 4616 -20573
rect 4650 -20607 4656 -20573
rect 4610 -20645 4656 -20607
rect 4610 -20679 4616 -20645
rect 4650 -20679 4656 -20645
rect 4610 -20717 4656 -20679
rect 4610 -20751 4616 -20717
rect 4650 -20751 4656 -20717
rect 4610 -20789 4656 -20751
rect 4610 -20823 4616 -20789
rect 4650 -20823 4656 -20789
rect 4610 -20861 4656 -20823
rect 4610 -20895 4616 -20861
rect 4650 -20895 4656 -20861
rect 4610 -20933 4656 -20895
rect 5628 -20429 5674 -20398
rect 5628 -20463 5634 -20429
rect 5668 -20463 5674 -20429
rect 5628 -20501 5674 -20463
rect 5628 -20535 5634 -20501
rect 5668 -20535 5674 -20501
rect 5628 -20573 5674 -20535
rect 5628 -20607 5634 -20573
rect 5668 -20607 5674 -20573
rect 5628 -20645 5674 -20607
rect 5628 -20679 5634 -20645
rect 5668 -20679 5674 -20645
rect 5628 -20717 5674 -20679
rect 5628 -20751 5634 -20717
rect 5668 -20751 5674 -20717
rect 5628 -20789 5674 -20751
rect 5628 -20823 5634 -20789
rect 5668 -20823 5674 -20789
rect 5628 -20861 5674 -20823
rect 5628 -20895 5634 -20861
rect 5668 -20895 5674 -20861
rect 5628 -20928 5674 -20895
rect 6646 -20429 6692 -20398
rect 6646 -20463 6652 -20429
rect 6686 -20463 6692 -20429
rect 6646 -20501 6692 -20463
rect 7658 -20429 7718 -19733
rect 8682 -19229 8688 -19212
rect 8722 -19212 8734 -19195
rect 9690 -19195 9750 -18730
rect 10196 -18884 10268 -18880
rect 10196 -18936 10206 -18884
rect 10258 -18936 10268 -18884
rect 10196 -18940 10268 -18936
rect 13268 -18896 13328 -18720
rect 13766 -18786 13826 -18501
rect 14790 -18501 14796 -18467
rect 14830 -18501 14836 -18467
rect 14790 -18532 14836 -18501
rect 15808 -17997 15814 -17988
rect 15848 -17988 15860 -17963
rect 16818 -17963 16878 -17804
rect 17326 -17854 17386 -17376
rect 17836 -17414 17896 -17267
rect 18854 -17267 18868 -17233
rect 18902 -17267 18914 -17233
rect 19880 -17233 19926 -17195
rect 19880 -17242 19886 -17233
rect 18132 -17336 18620 -17330
rect 18132 -17370 18179 -17336
rect 18213 -17370 18251 -17336
rect 18285 -17370 18323 -17336
rect 18357 -17370 18395 -17336
rect 18429 -17370 18467 -17336
rect 18501 -17370 18539 -17336
rect 18573 -17370 18620 -17336
rect 18132 -17376 18620 -17370
rect 17830 -17418 17902 -17414
rect 17830 -17470 17840 -17418
rect 17892 -17470 17902 -17418
rect 17830 -17474 17902 -17470
rect 17114 -17860 17602 -17854
rect 17114 -17894 17161 -17860
rect 17195 -17894 17233 -17860
rect 17267 -17894 17305 -17860
rect 17339 -17894 17377 -17860
rect 17411 -17894 17449 -17860
rect 17483 -17894 17521 -17860
rect 17555 -17894 17602 -17860
rect 17114 -17900 17602 -17894
rect 16818 -17974 16832 -17963
rect 15848 -17997 15854 -17988
rect 15808 -18035 15854 -17997
rect 15808 -18069 15814 -18035
rect 15848 -18069 15854 -18035
rect 15808 -18107 15854 -18069
rect 15808 -18141 15814 -18107
rect 15848 -18141 15854 -18107
rect 15808 -18179 15854 -18141
rect 15808 -18213 15814 -18179
rect 15848 -18213 15854 -18179
rect 15808 -18251 15854 -18213
rect 15808 -18285 15814 -18251
rect 15848 -18285 15854 -18251
rect 15808 -18323 15854 -18285
rect 15808 -18357 15814 -18323
rect 15848 -18357 15854 -18323
rect 15808 -18395 15854 -18357
rect 15808 -18429 15814 -18395
rect 15848 -18429 15854 -18395
rect 15808 -18467 15854 -18429
rect 15808 -18501 15814 -18467
rect 15848 -18501 15854 -18467
rect 16826 -17997 16832 -17974
rect 16866 -17974 16878 -17963
rect 17836 -17963 17896 -17474
rect 18352 -17854 18412 -17376
rect 18854 -17630 18914 -17267
rect 19870 -17267 19886 -17242
rect 19920 -17242 19926 -17233
rect 20898 -16729 20944 -16698
rect 20898 -16763 20904 -16729
rect 20938 -16763 20944 -16729
rect 20898 -16801 20944 -16763
rect 20898 -16835 20904 -16801
rect 20938 -16835 20944 -16801
rect 20898 -16873 20944 -16835
rect 20898 -16907 20904 -16873
rect 20938 -16907 20944 -16873
rect 20898 -16945 20944 -16907
rect 20898 -16979 20904 -16945
rect 20938 -16979 20944 -16945
rect 20898 -17017 20944 -16979
rect 20898 -17051 20904 -17017
rect 20938 -17051 20944 -17017
rect 20898 -17089 20944 -17051
rect 20898 -17123 20904 -17089
rect 20938 -17123 20944 -17089
rect 20898 -17161 20944 -17123
rect 20898 -17195 20904 -17161
rect 20938 -17195 20944 -17161
rect 20898 -17233 20944 -17195
rect 20898 -17242 20904 -17233
rect 19920 -17267 19930 -17242
rect 19150 -17336 19638 -17330
rect 19150 -17370 19197 -17336
rect 19231 -17370 19269 -17336
rect 19303 -17370 19341 -17336
rect 19375 -17370 19413 -17336
rect 19447 -17370 19485 -17336
rect 19519 -17370 19557 -17336
rect 19591 -17370 19638 -17336
rect 19150 -17376 19638 -17370
rect 18848 -17634 18920 -17630
rect 18848 -17686 18858 -17634
rect 18910 -17686 18920 -17634
rect 18848 -17690 18920 -17686
rect 19360 -17680 19420 -17376
rect 19870 -17522 19930 -17267
rect 20894 -17267 20904 -17242
rect 20938 -17242 20944 -17233
rect 21916 -16729 21962 -16698
rect 21916 -16763 21922 -16729
rect 21956 -16763 21962 -16729
rect 22926 -16729 22986 -16544
rect 23028 -16512 23100 -16508
rect 23028 -16564 23038 -16512
rect 23090 -16564 23100 -16512
rect 23162 -16526 23222 -16238
rect 23028 -16568 23100 -16564
rect 23156 -16530 23228 -16526
rect 22926 -16738 22940 -16729
rect 21916 -16801 21962 -16763
rect 21916 -16835 21922 -16801
rect 21956 -16835 21962 -16801
rect 21916 -16873 21962 -16835
rect 21916 -16907 21922 -16873
rect 21956 -16907 21962 -16873
rect 21916 -16945 21962 -16907
rect 21916 -16979 21922 -16945
rect 21956 -16979 21962 -16945
rect 21916 -17017 21962 -16979
rect 21916 -17051 21922 -17017
rect 21956 -17051 21962 -17017
rect 21916 -17089 21962 -17051
rect 21916 -17123 21922 -17089
rect 21956 -17123 21962 -17089
rect 21916 -17161 21962 -17123
rect 21916 -17195 21922 -17161
rect 21956 -17195 21962 -17161
rect 21916 -17233 21962 -17195
rect 22934 -16763 22940 -16738
rect 22974 -16738 22986 -16729
rect 22974 -16763 22980 -16738
rect 22934 -16801 22980 -16763
rect 22934 -16835 22940 -16801
rect 22974 -16835 22980 -16801
rect 22934 -16873 22980 -16835
rect 22934 -16907 22940 -16873
rect 22974 -16907 22980 -16873
rect 22934 -16945 22980 -16907
rect 22934 -16979 22940 -16945
rect 22974 -16979 22980 -16945
rect 22934 -17017 22980 -16979
rect 22934 -17051 22940 -17017
rect 22974 -17051 22980 -17017
rect 22934 -17089 22980 -17051
rect 22934 -17123 22940 -17089
rect 22974 -17123 22980 -17089
rect 22934 -17161 22980 -17123
rect 22934 -17195 22940 -17161
rect 22974 -17195 22980 -17161
rect 22934 -17228 22980 -17195
rect 21916 -17236 21922 -17233
rect 20938 -17267 20954 -17242
rect 20168 -17336 20656 -17330
rect 20168 -17370 20215 -17336
rect 20249 -17370 20287 -17336
rect 20321 -17370 20359 -17336
rect 20393 -17370 20431 -17336
rect 20465 -17370 20503 -17336
rect 20537 -17370 20575 -17336
rect 20609 -17370 20656 -17336
rect 20168 -17376 20656 -17370
rect 20376 -17520 20436 -17376
rect 19864 -17526 19936 -17522
rect 19864 -17578 19874 -17526
rect 19926 -17578 19936 -17526
rect 19864 -17582 19936 -17578
rect 20374 -17530 20436 -17520
rect 20374 -17582 20378 -17530
rect 20430 -17582 20436 -17530
rect 20374 -17592 20436 -17582
rect 20376 -17680 20436 -17592
rect 20894 -17630 20954 -17267
rect 21910 -17267 21922 -17236
rect 21956 -17236 21962 -17233
rect 22928 -17233 22988 -17228
rect 21956 -17267 21970 -17236
rect 21186 -17336 21674 -17330
rect 21186 -17370 21233 -17336
rect 21267 -17370 21305 -17336
rect 21339 -17370 21377 -17336
rect 21411 -17370 21449 -17336
rect 21483 -17370 21521 -17336
rect 21555 -17370 21593 -17336
rect 21627 -17370 21674 -17336
rect 21186 -17376 21674 -17370
rect 19360 -17740 20436 -17680
rect 20888 -17634 20960 -17630
rect 20888 -17686 20898 -17634
rect 20950 -17686 20960 -17634
rect 20888 -17690 20960 -17686
rect 18848 -17748 18920 -17744
rect 18848 -17800 18858 -17748
rect 18910 -17800 18920 -17748
rect 18848 -17804 18920 -17800
rect 18132 -17860 18620 -17854
rect 18132 -17894 18179 -17860
rect 18213 -17894 18251 -17860
rect 18285 -17894 18323 -17860
rect 18357 -17894 18395 -17860
rect 18429 -17894 18467 -17860
rect 18501 -17894 18539 -17860
rect 18573 -17894 18620 -17860
rect 18132 -17900 18620 -17894
rect 16866 -17997 16872 -17974
rect 17836 -17984 17850 -17963
rect 16826 -18035 16872 -17997
rect 16826 -18069 16832 -18035
rect 16866 -18069 16872 -18035
rect 16826 -18107 16872 -18069
rect 16826 -18141 16832 -18107
rect 16866 -18141 16872 -18107
rect 16826 -18179 16872 -18141
rect 16826 -18213 16832 -18179
rect 16866 -18213 16872 -18179
rect 16826 -18251 16872 -18213
rect 16826 -18285 16832 -18251
rect 16866 -18285 16872 -18251
rect 16826 -18323 16872 -18285
rect 16826 -18357 16832 -18323
rect 16866 -18357 16872 -18323
rect 16826 -18395 16872 -18357
rect 16826 -18429 16832 -18395
rect 16866 -18429 16872 -18395
rect 16826 -18467 16872 -18429
rect 16826 -18480 16832 -18467
rect 15808 -18532 15854 -18501
rect 16818 -18501 16832 -18480
rect 16866 -18480 16872 -18467
rect 17844 -17997 17850 -17984
rect 17884 -17984 17896 -17963
rect 18854 -17963 18914 -17804
rect 19360 -17854 19420 -17740
rect 20376 -17854 20436 -17740
rect 20886 -17748 20958 -17744
rect 20886 -17800 20896 -17748
rect 20948 -17800 20958 -17748
rect 20886 -17804 20958 -17800
rect 19150 -17860 19638 -17854
rect 19150 -17894 19197 -17860
rect 19231 -17894 19269 -17860
rect 19303 -17894 19341 -17860
rect 19375 -17894 19413 -17860
rect 19447 -17894 19485 -17860
rect 19519 -17894 19557 -17860
rect 19591 -17894 19638 -17860
rect 19150 -17900 19638 -17894
rect 20168 -17860 20656 -17854
rect 20168 -17894 20215 -17860
rect 20249 -17894 20287 -17860
rect 20321 -17894 20359 -17860
rect 20393 -17894 20431 -17860
rect 20465 -17894 20503 -17860
rect 20537 -17894 20575 -17860
rect 20609 -17894 20656 -17860
rect 20168 -17900 20656 -17894
rect 17884 -17997 17890 -17984
rect 18854 -17986 18868 -17963
rect 17844 -18035 17890 -17997
rect 17844 -18069 17850 -18035
rect 17884 -18069 17890 -18035
rect 17844 -18107 17890 -18069
rect 17844 -18141 17850 -18107
rect 17884 -18141 17890 -18107
rect 17844 -18179 17890 -18141
rect 17844 -18213 17850 -18179
rect 17884 -18213 17890 -18179
rect 17844 -18251 17890 -18213
rect 17844 -18285 17850 -18251
rect 17884 -18285 17890 -18251
rect 17844 -18323 17890 -18285
rect 17844 -18357 17850 -18323
rect 17884 -18357 17890 -18323
rect 17844 -18395 17890 -18357
rect 17844 -18429 17850 -18395
rect 17884 -18429 17890 -18395
rect 17844 -18467 17890 -18429
rect 16866 -18501 16878 -18480
rect 17844 -18486 17850 -18467
rect 14060 -18570 14548 -18564
rect 14060 -18604 14107 -18570
rect 14141 -18604 14179 -18570
rect 14213 -18604 14251 -18570
rect 14285 -18604 14323 -18570
rect 14357 -18604 14395 -18570
rect 14429 -18604 14467 -18570
rect 14501 -18604 14548 -18570
rect 14060 -18610 14548 -18604
rect 15078 -18570 15566 -18564
rect 15078 -18604 15125 -18570
rect 15159 -18604 15197 -18570
rect 15231 -18604 15269 -18570
rect 15303 -18604 15341 -18570
rect 15375 -18604 15413 -18570
rect 15447 -18604 15485 -18570
rect 15519 -18604 15566 -18570
rect 15078 -18610 15566 -18604
rect 16096 -18570 16584 -18564
rect 16096 -18604 16143 -18570
rect 16177 -18604 16215 -18570
rect 16249 -18604 16287 -18570
rect 16321 -18604 16359 -18570
rect 16393 -18604 16431 -18570
rect 16465 -18604 16503 -18570
rect 16537 -18604 16584 -18570
rect 16096 -18610 16584 -18604
rect 14272 -18662 14332 -18610
rect 14272 -18714 14276 -18662
rect 14328 -18714 14332 -18662
rect 13760 -18790 13832 -18786
rect 13760 -18842 13770 -18790
rect 13822 -18842 13832 -18790
rect 13760 -18846 13832 -18842
rect 14272 -18896 14332 -18714
rect 10202 -19086 10262 -18940
rect 13268 -18956 14332 -18896
rect 15796 -18988 15868 -18984
rect 15796 -19040 15806 -18988
rect 15858 -19040 15868 -18988
rect 15796 -19044 15868 -19040
rect 9988 -19092 10476 -19086
rect 9988 -19126 10035 -19092
rect 10069 -19126 10107 -19092
rect 10141 -19126 10179 -19092
rect 10213 -19126 10251 -19092
rect 10285 -19126 10323 -19092
rect 10357 -19126 10395 -19092
rect 10429 -19126 10476 -19092
rect 9988 -19132 10476 -19126
rect 11006 -19092 11494 -19086
rect 11006 -19126 11053 -19092
rect 11087 -19126 11125 -19092
rect 11159 -19126 11197 -19092
rect 11231 -19126 11269 -19092
rect 11303 -19126 11341 -19092
rect 11375 -19126 11413 -19092
rect 11447 -19126 11494 -19092
rect 11006 -19132 11494 -19126
rect 12024 -19092 12512 -19086
rect 12024 -19126 12071 -19092
rect 12105 -19126 12143 -19092
rect 12177 -19126 12215 -19092
rect 12249 -19126 12287 -19092
rect 12321 -19126 12359 -19092
rect 12393 -19126 12431 -19092
rect 12465 -19126 12512 -19092
rect 12024 -19132 12512 -19126
rect 13042 -19092 13530 -19086
rect 13042 -19126 13089 -19092
rect 13123 -19126 13161 -19092
rect 13195 -19126 13233 -19092
rect 13267 -19126 13305 -19092
rect 13339 -19126 13377 -19092
rect 13411 -19126 13449 -19092
rect 13483 -19126 13530 -19092
rect 13042 -19132 13530 -19126
rect 14060 -19092 14548 -19086
rect 14060 -19126 14107 -19092
rect 14141 -19126 14179 -19092
rect 14213 -19126 14251 -19092
rect 14285 -19126 14323 -19092
rect 14357 -19126 14395 -19092
rect 14429 -19126 14467 -19092
rect 14501 -19126 14548 -19092
rect 14060 -19132 14548 -19126
rect 15078 -19092 15566 -19086
rect 15078 -19126 15125 -19092
rect 15159 -19126 15197 -19092
rect 15231 -19126 15269 -19092
rect 15303 -19126 15341 -19092
rect 15375 -19126 15413 -19092
rect 15447 -19126 15485 -19092
rect 15519 -19126 15566 -19092
rect 15078 -19132 15566 -19126
rect 8722 -19229 8728 -19212
rect 9690 -19214 9706 -19195
rect 8682 -19267 8728 -19229
rect 8682 -19301 8688 -19267
rect 8722 -19301 8728 -19267
rect 8682 -19339 8728 -19301
rect 8682 -19373 8688 -19339
rect 8722 -19373 8728 -19339
rect 8682 -19411 8728 -19373
rect 8682 -19445 8688 -19411
rect 8722 -19445 8728 -19411
rect 8682 -19483 8728 -19445
rect 8682 -19517 8688 -19483
rect 8722 -19517 8728 -19483
rect 8682 -19555 8728 -19517
rect 8682 -19589 8688 -19555
rect 8722 -19589 8728 -19555
rect 8682 -19627 8728 -19589
rect 8682 -19661 8688 -19627
rect 8722 -19661 8728 -19627
rect 8682 -19699 8728 -19661
rect 8682 -19733 8688 -19699
rect 8722 -19733 8728 -19699
rect 8682 -19764 8728 -19733
rect 9700 -19229 9706 -19214
rect 9740 -19214 9750 -19195
rect 10718 -19195 10764 -19164
rect 9740 -19229 9746 -19214
rect 9700 -19267 9746 -19229
rect 9700 -19301 9706 -19267
rect 9740 -19301 9746 -19267
rect 9700 -19339 9746 -19301
rect 9700 -19373 9706 -19339
rect 9740 -19373 9746 -19339
rect 9700 -19411 9746 -19373
rect 9700 -19445 9706 -19411
rect 9740 -19445 9746 -19411
rect 9700 -19483 9746 -19445
rect 9700 -19517 9706 -19483
rect 9740 -19517 9746 -19483
rect 9700 -19555 9746 -19517
rect 9700 -19589 9706 -19555
rect 9740 -19589 9746 -19555
rect 9700 -19627 9746 -19589
rect 9700 -19661 9706 -19627
rect 9740 -19661 9746 -19627
rect 9700 -19699 9746 -19661
rect 9700 -19733 9706 -19699
rect 9740 -19733 9746 -19699
rect 10718 -19229 10724 -19195
rect 10758 -19229 10764 -19195
rect 10718 -19267 10764 -19229
rect 10718 -19301 10724 -19267
rect 10758 -19301 10764 -19267
rect 10718 -19339 10764 -19301
rect 10718 -19373 10724 -19339
rect 10758 -19373 10764 -19339
rect 10718 -19411 10764 -19373
rect 10718 -19445 10724 -19411
rect 10758 -19445 10764 -19411
rect 10718 -19483 10764 -19445
rect 10718 -19517 10724 -19483
rect 10758 -19517 10764 -19483
rect 10718 -19555 10764 -19517
rect 10718 -19589 10724 -19555
rect 10758 -19589 10764 -19555
rect 10718 -19627 10764 -19589
rect 10718 -19661 10724 -19627
rect 10758 -19661 10764 -19627
rect 10718 -19699 10764 -19661
rect 10718 -19710 10724 -19699
rect 9700 -19764 9746 -19733
rect 10710 -19733 10724 -19710
rect 10758 -19710 10764 -19699
rect 11736 -19195 11782 -19164
rect 11736 -19229 11742 -19195
rect 11776 -19229 11782 -19195
rect 11736 -19267 11782 -19229
rect 11736 -19301 11742 -19267
rect 11776 -19301 11782 -19267
rect 11736 -19339 11782 -19301
rect 11736 -19373 11742 -19339
rect 11776 -19373 11782 -19339
rect 11736 -19411 11782 -19373
rect 11736 -19445 11742 -19411
rect 11776 -19445 11782 -19411
rect 11736 -19483 11782 -19445
rect 11736 -19517 11742 -19483
rect 11776 -19517 11782 -19483
rect 11736 -19555 11782 -19517
rect 11736 -19589 11742 -19555
rect 11776 -19589 11782 -19555
rect 11736 -19627 11782 -19589
rect 11736 -19661 11742 -19627
rect 11776 -19661 11782 -19627
rect 11736 -19699 11782 -19661
rect 10758 -19733 10770 -19710
rect 11736 -19714 11742 -19699
rect 7952 -19802 8440 -19796
rect 7952 -19836 7999 -19802
rect 8033 -19836 8071 -19802
rect 8105 -19836 8143 -19802
rect 8177 -19836 8215 -19802
rect 8249 -19836 8287 -19802
rect 8321 -19836 8359 -19802
rect 8393 -19836 8440 -19802
rect 7952 -19842 8220 -19836
rect 8224 -19842 8440 -19836
rect 8970 -19802 9458 -19796
rect 8970 -19836 9017 -19802
rect 9051 -19836 9089 -19802
rect 9123 -19836 9161 -19802
rect 9195 -19836 9233 -19802
rect 9267 -19836 9305 -19802
rect 9339 -19836 9377 -19802
rect 9411 -19836 9458 -19802
rect 8970 -19842 9458 -19836
rect 9988 -19802 10476 -19796
rect 9988 -19836 10035 -19802
rect 10069 -19836 10107 -19802
rect 10141 -19836 10179 -19802
rect 10213 -19836 10251 -19802
rect 10285 -19836 10323 -19802
rect 10357 -19836 10395 -19802
rect 10429 -19836 10476 -19802
rect 9988 -19842 10476 -19836
rect 8160 -19898 8220 -19842
rect 9166 -19898 9226 -19842
rect 10210 -19898 10270 -19842
rect 10710 -19892 10770 -19733
rect 11730 -19733 11742 -19714
rect 11776 -19714 11782 -19699
rect 12754 -19195 12800 -19164
rect 12754 -19229 12760 -19195
rect 12794 -19229 12800 -19195
rect 12754 -19267 12800 -19229
rect 12754 -19301 12760 -19267
rect 12794 -19301 12800 -19267
rect 12754 -19339 12800 -19301
rect 12754 -19373 12760 -19339
rect 12794 -19373 12800 -19339
rect 12754 -19411 12800 -19373
rect 12754 -19445 12760 -19411
rect 12794 -19445 12800 -19411
rect 12754 -19483 12800 -19445
rect 12754 -19517 12760 -19483
rect 12794 -19517 12800 -19483
rect 12754 -19555 12800 -19517
rect 12754 -19589 12760 -19555
rect 12794 -19589 12800 -19555
rect 12754 -19627 12800 -19589
rect 12754 -19661 12760 -19627
rect 12794 -19661 12800 -19627
rect 12754 -19699 12800 -19661
rect 11776 -19733 11790 -19714
rect 12754 -19720 12760 -19699
rect 11006 -19802 11494 -19796
rect 11006 -19836 11053 -19802
rect 11087 -19836 11125 -19802
rect 11159 -19836 11197 -19802
rect 11231 -19836 11269 -19802
rect 11303 -19836 11341 -19802
rect 11375 -19836 11413 -19802
rect 11447 -19836 11494 -19802
rect 11006 -19842 11494 -19836
rect 10704 -19896 10776 -19892
rect 8154 -19902 8226 -19898
rect 8154 -19954 8164 -19902
rect 8216 -19954 8226 -19902
rect 8154 -19958 8226 -19954
rect 9160 -19902 9232 -19898
rect 9160 -19954 9170 -19902
rect 9222 -19954 9232 -19902
rect 9160 -19958 9232 -19954
rect 10204 -19902 10276 -19898
rect 10204 -19954 10214 -19902
rect 10266 -19954 10276 -19902
rect 10704 -19948 10714 -19896
rect 10766 -19948 10776 -19896
rect 10704 -19952 10776 -19948
rect 10204 -19958 10276 -19954
rect 8160 -20320 8220 -19958
rect 9158 -20118 9230 -20114
rect 9158 -20170 9168 -20118
rect 9220 -20170 9230 -20118
rect 9158 -20174 9230 -20170
rect 10198 -20118 10270 -20114
rect 10198 -20170 10208 -20118
rect 10260 -20170 10270 -20118
rect 10198 -20174 10270 -20170
rect 9164 -20320 9224 -20174
rect 9682 -20222 9754 -20218
rect 9682 -20274 9692 -20222
rect 9744 -20274 9754 -20222
rect 9682 -20278 9754 -20274
rect 7952 -20326 8440 -20320
rect 7952 -20360 7999 -20326
rect 8033 -20360 8071 -20326
rect 8105 -20360 8143 -20326
rect 8177 -20360 8215 -20326
rect 8249 -20360 8287 -20326
rect 8321 -20360 8359 -20326
rect 8393 -20360 8440 -20326
rect 7952 -20366 8440 -20360
rect 8970 -20326 9458 -20320
rect 8970 -20360 9017 -20326
rect 9051 -20360 9089 -20326
rect 9123 -20360 9161 -20326
rect 9195 -20360 9233 -20326
rect 9267 -20360 9305 -20326
rect 9339 -20360 9377 -20326
rect 9411 -20360 9458 -20326
rect 8970 -20366 9458 -20360
rect 7658 -20463 7670 -20429
rect 7704 -20463 7718 -20429
rect 7658 -20492 7718 -20463
rect 8682 -20429 8728 -20398
rect 8682 -20463 8688 -20429
rect 8722 -20463 8728 -20429
rect 6646 -20535 6652 -20501
rect 6686 -20535 6692 -20501
rect 6646 -20573 6692 -20535
rect 6646 -20607 6652 -20573
rect 6686 -20607 6692 -20573
rect 6646 -20645 6692 -20607
rect 6646 -20679 6652 -20645
rect 6686 -20679 6692 -20645
rect 6646 -20717 6692 -20679
rect 6646 -20751 6652 -20717
rect 6686 -20751 6692 -20717
rect 6646 -20789 6692 -20751
rect 6646 -20823 6652 -20789
rect 6686 -20823 6692 -20789
rect 6646 -20861 6692 -20823
rect 6646 -20895 6652 -20861
rect 6686 -20895 6692 -20861
rect 4610 -20936 4616 -20933
rect 3632 -20967 3646 -20948
rect 2862 -21036 3350 -21030
rect 2862 -21070 2909 -21036
rect 2943 -21070 2981 -21036
rect 3015 -21070 3053 -21036
rect 3087 -21070 3125 -21036
rect 3159 -21070 3197 -21036
rect 3231 -21070 3269 -21036
rect 3303 -21070 3350 -21036
rect 2862 -21076 3350 -21070
rect 3066 -21116 3126 -21076
rect 3586 -21116 3646 -20967
rect 4602 -20967 4616 -20936
rect 4650 -20936 4656 -20933
rect 5620 -20933 5680 -20928
rect 4650 -20967 4662 -20936
rect 3880 -21036 4368 -21030
rect 3880 -21070 3927 -21036
rect 3961 -21070 3999 -21036
rect 4033 -21070 4071 -21036
rect 4105 -21070 4143 -21036
rect 4177 -21070 4215 -21036
rect 4249 -21070 4287 -21036
rect 4321 -21070 4368 -21036
rect 3880 -21076 4368 -21070
rect 2568 -21176 3646 -21116
rect 3586 -21230 3646 -21176
rect 4078 -21130 4150 -21126
rect 4078 -21182 4088 -21130
rect 4140 -21182 4150 -21130
rect 4078 -21186 4150 -21182
rect 3580 -21234 3652 -21230
rect 3580 -21286 3590 -21234
rect 3642 -21286 3652 -21234
rect 3580 -21290 3652 -21286
rect 3576 -21444 3648 -21440
rect 3576 -21496 3586 -21444
rect 3638 -21496 3648 -21444
rect 3576 -21500 3648 -21496
rect 2862 -21560 3350 -21554
rect 2862 -21594 2909 -21560
rect 2943 -21594 2981 -21560
rect 3015 -21594 3053 -21560
rect 3087 -21594 3125 -21560
rect 3159 -21594 3197 -21560
rect 3231 -21594 3269 -21560
rect 3303 -21594 3350 -21560
rect 2862 -21600 3350 -21594
rect 2574 -21663 2620 -21632
rect 2574 -21697 2580 -21663
rect 2614 -21697 2620 -21663
rect 2574 -21735 2620 -21697
rect 3582 -21663 3642 -21500
rect 4084 -21554 4144 -21186
rect 4602 -21342 4662 -20967
rect 5620 -20967 5634 -20933
rect 5668 -20967 5680 -20933
rect 6646 -20933 6692 -20895
rect 6646 -20940 6652 -20933
rect 4898 -21036 5386 -21030
rect 4898 -21070 4945 -21036
rect 4979 -21070 5017 -21036
rect 5051 -21070 5089 -21036
rect 5123 -21070 5161 -21036
rect 5195 -21070 5233 -21036
rect 5267 -21070 5305 -21036
rect 5339 -21070 5386 -21036
rect 4898 -21076 5386 -21070
rect 5092 -21126 5152 -21076
rect 5086 -21130 5158 -21126
rect 5086 -21182 5096 -21130
rect 5148 -21182 5158 -21130
rect 5086 -21186 5158 -21182
rect 4596 -21346 4668 -21342
rect 4596 -21398 4606 -21346
rect 4658 -21398 4668 -21346
rect 4596 -21402 4668 -21398
rect 5620 -21440 5680 -20967
rect 6640 -20967 6652 -20940
rect 6686 -20940 6692 -20933
rect 7664 -20501 7710 -20492
rect 7664 -20535 7670 -20501
rect 7704 -20535 7710 -20501
rect 7664 -20573 7710 -20535
rect 7664 -20607 7670 -20573
rect 7704 -20607 7710 -20573
rect 7664 -20645 7710 -20607
rect 7664 -20679 7670 -20645
rect 7704 -20679 7710 -20645
rect 7664 -20717 7710 -20679
rect 7664 -20751 7670 -20717
rect 7704 -20751 7710 -20717
rect 7664 -20789 7710 -20751
rect 7664 -20823 7670 -20789
rect 7704 -20823 7710 -20789
rect 7664 -20861 7710 -20823
rect 7664 -20895 7670 -20861
rect 7704 -20895 7710 -20861
rect 7664 -20933 7710 -20895
rect 7664 -20940 7670 -20933
rect 6686 -20967 6700 -20940
rect 5916 -21036 6404 -21030
rect 5916 -21070 5963 -21036
rect 5997 -21070 6035 -21036
rect 6069 -21070 6107 -21036
rect 6141 -21070 6179 -21036
rect 6213 -21070 6251 -21036
rect 6285 -21070 6323 -21036
rect 6357 -21070 6404 -21036
rect 5916 -21076 6404 -21070
rect 6106 -21126 6166 -21076
rect 6100 -21130 6172 -21126
rect 6100 -21182 6110 -21130
rect 6162 -21182 6172 -21130
rect 6100 -21186 6172 -21182
rect 6640 -21342 6700 -20967
rect 7660 -20967 7670 -20940
rect 7704 -20940 7710 -20933
rect 8682 -20501 8728 -20463
rect 9688 -20429 9748 -20278
rect 10204 -20320 10264 -20174
rect 9988 -20326 10476 -20320
rect 9988 -20360 10035 -20326
rect 10069 -20360 10107 -20326
rect 10141 -20360 10179 -20326
rect 10213 -20360 10251 -20326
rect 10285 -20360 10323 -20326
rect 10357 -20360 10395 -20326
rect 10429 -20360 10476 -20326
rect 9988 -20366 10476 -20360
rect 9688 -20463 9706 -20429
rect 9740 -20463 9748 -20429
rect 10710 -20429 10770 -19952
rect 11218 -20114 11278 -19842
rect 11212 -20118 11284 -20114
rect 11212 -20170 11222 -20118
rect 11274 -20170 11284 -20118
rect 11212 -20174 11284 -20170
rect 11218 -20320 11278 -20174
rect 11730 -20218 11790 -19733
rect 12746 -19733 12760 -19720
rect 12794 -19720 12800 -19699
rect 13772 -19195 13818 -19164
rect 13772 -19229 13778 -19195
rect 13812 -19229 13818 -19195
rect 13772 -19267 13818 -19229
rect 13772 -19301 13778 -19267
rect 13812 -19301 13818 -19267
rect 13772 -19339 13818 -19301
rect 13772 -19373 13778 -19339
rect 13812 -19373 13818 -19339
rect 13772 -19411 13818 -19373
rect 13772 -19445 13778 -19411
rect 13812 -19445 13818 -19411
rect 13772 -19483 13818 -19445
rect 13772 -19517 13778 -19483
rect 13812 -19517 13818 -19483
rect 13772 -19555 13818 -19517
rect 13772 -19589 13778 -19555
rect 13812 -19589 13818 -19555
rect 13772 -19627 13818 -19589
rect 13772 -19661 13778 -19627
rect 13812 -19661 13818 -19627
rect 13772 -19699 13818 -19661
rect 13772 -19718 13778 -19699
rect 12794 -19733 12806 -19720
rect 12024 -19802 12512 -19796
rect 12024 -19836 12071 -19802
rect 12105 -19836 12143 -19802
rect 12177 -19836 12215 -19802
rect 12249 -19836 12287 -19802
rect 12321 -19836 12359 -19802
rect 12393 -19836 12431 -19802
rect 12465 -19836 12512 -19802
rect 12024 -19842 12512 -19836
rect 12226 -20114 12286 -19842
rect 12746 -19892 12806 -19733
rect 13768 -19733 13778 -19718
rect 13812 -19718 13818 -19699
rect 14790 -19195 14836 -19164
rect 14790 -19229 14796 -19195
rect 14830 -19229 14836 -19195
rect 14790 -19267 14836 -19229
rect 14790 -19301 14796 -19267
rect 14830 -19301 14836 -19267
rect 14790 -19339 14836 -19301
rect 14790 -19373 14796 -19339
rect 14830 -19373 14836 -19339
rect 14790 -19411 14836 -19373
rect 14790 -19445 14796 -19411
rect 14830 -19445 14836 -19411
rect 14790 -19483 14836 -19445
rect 14790 -19517 14796 -19483
rect 14830 -19517 14836 -19483
rect 14790 -19555 14836 -19517
rect 14790 -19589 14796 -19555
rect 14830 -19589 14836 -19555
rect 14790 -19627 14836 -19589
rect 14790 -19661 14796 -19627
rect 14830 -19661 14836 -19627
rect 14790 -19699 14836 -19661
rect 13812 -19733 13828 -19718
rect 14790 -19720 14796 -19699
rect 13042 -19802 13530 -19796
rect 13042 -19836 13089 -19802
rect 13123 -19836 13161 -19802
rect 13195 -19836 13233 -19802
rect 13267 -19836 13305 -19802
rect 13339 -19836 13377 -19802
rect 13411 -19836 13449 -19802
rect 13483 -19836 13530 -19802
rect 13042 -19842 13530 -19836
rect 12740 -19896 12812 -19892
rect 12740 -19948 12750 -19896
rect 12802 -19948 12812 -19896
rect 12740 -19952 12812 -19948
rect 13270 -20114 13330 -19842
rect 12220 -20118 12292 -20114
rect 12220 -20170 12230 -20118
rect 12282 -20170 12292 -20118
rect 12220 -20174 12292 -20170
rect 13264 -20118 13336 -20114
rect 13264 -20170 13274 -20118
rect 13326 -20170 13336 -20118
rect 13264 -20174 13336 -20170
rect 11724 -20222 11796 -20218
rect 11724 -20274 11734 -20222
rect 11786 -20274 11796 -20222
rect 11724 -20278 11796 -20274
rect 11006 -20326 11494 -20320
rect 11006 -20360 11053 -20326
rect 11087 -20360 11125 -20326
rect 11159 -20360 11197 -20326
rect 11231 -20360 11269 -20326
rect 11303 -20360 11341 -20326
rect 11375 -20360 11413 -20326
rect 11447 -20360 11494 -20326
rect 11006 -20366 11494 -20360
rect 10710 -20446 10724 -20429
rect 9688 -20474 9748 -20463
rect 10718 -20463 10724 -20446
rect 10758 -20446 10770 -20429
rect 11730 -20429 11790 -20278
rect 12226 -20320 12286 -20174
rect 13270 -20320 13330 -20174
rect 13768 -20218 13828 -19733
rect 14782 -19733 14796 -19720
rect 14830 -19720 14836 -19699
rect 15802 -19195 15862 -19044
rect 16096 -19092 16584 -19086
rect 16096 -19126 16143 -19092
rect 16177 -19126 16215 -19092
rect 16249 -19126 16287 -19092
rect 16321 -19126 16359 -19092
rect 16393 -19126 16431 -19092
rect 16465 -19126 16503 -19092
rect 16537 -19126 16584 -19092
rect 16096 -19132 16584 -19126
rect 15802 -19229 15814 -19195
rect 15848 -19229 15862 -19195
rect 16818 -19195 16878 -18501
rect 17838 -18501 17850 -18486
rect 17884 -18486 17890 -18467
rect 18862 -17997 18868 -17986
rect 18902 -17986 18914 -17963
rect 19880 -17963 19926 -17932
rect 18902 -17997 18908 -17986
rect 18862 -18035 18908 -17997
rect 18862 -18069 18868 -18035
rect 18902 -18069 18908 -18035
rect 18862 -18107 18908 -18069
rect 18862 -18141 18868 -18107
rect 18902 -18141 18908 -18107
rect 18862 -18179 18908 -18141
rect 18862 -18213 18868 -18179
rect 18902 -18213 18908 -18179
rect 18862 -18251 18908 -18213
rect 18862 -18285 18868 -18251
rect 18902 -18285 18908 -18251
rect 18862 -18323 18908 -18285
rect 18862 -18357 18868 -18323
rect 18902 -18357 18908 -18323
rect 18862 -18395 18908 -18357
rect 18862 -18429 18868 -18395
rect 18902 -18429 18908 -18395
rect 18862 -18467 18908 -18429
rect 19880 -17997 19886 -17963
rect 19920 -17997 19926 -17963
rect 20892 -17963 20952 -17804
rect 21394 -17854 21454 -17376
rect 21910 -17414 21970 -17267
rect 22928 -17267 22940 -17233
rect 22974 -17267 22988 -17233
rect 22204 -17336 22692 -17330
rect 22204 -17370 22251 -17336
rect 22285 -17370 22323 -17336
rect 22357 -17370 22395 -17336
rect 22429 -17370 22467 -17336
rect 22501 -17370 22539 -17336
rect 22573 -17370 22611 -17336
rect 22645 -17370 22692 -17336
rect 22204 -17376 22692 -17370
rect 22928 -17396 22988 -17267
rect 22922 -17400 22994 -17396
rect 21904 -17418 21976 -17414
rect 21904 -17470 21914 -17418
rect 21966 -17470 21976 -17418
rect 22922 -17452 22932 -17400
rect 22984 -17452 22994 -17400
rect 22922 -17456 22994 -17452
rect 21904 -17474 21976 -17470
rect 21910 -17692 21970 -17474
rect 21910 -17752 22984 -17692
rect 23034 -17744 23094 -16568
rect 23156 -16582 23166 -16530
rect 23218 -16582 23228 -16530
rect 23156 -16586 23228 -16582
rect 23528 -17526 23588 -13640
rect 23522 -17530 23594 -17526
rect 23522 -17582 23532 -17530
rect 23584 -17582 23594 -17530
rect 23522 -17586 23594 -17582
rect 23272 -17634 23344 -17630
rect 23272 -17686 23282 -17634
rect 23334 -17686 23344 -17634
rect 23272 -17690 23344 -17686
rect 21186 -17860 21674 -17854
rect 21186 -17894 21233 -17860
rect 21267 -17894 21305 -17860
rect 21339 -17894 21377 -17860
rect 21411 -17894 21449 -17860
rect 21483 -17894 21521 -17860
rect 21555 -17894 21593 -17860
rect 21627 -17894 21674 -17860
rect 21186 -17900 21674 -17894
rect 20892 -17986 20904 -17963
rect 19880 -18035 19926 -17997
rect 19880 -18069 19886 -18035
rect 19920 -18069 19926 -18035
rect 19880 -18107 19926 -18069
rect 19880 -18141 19886 -18107
rect 19920 -18141 19926 -18107
rect 19880 -18179 19926 -18141
rect 19880 -18213 19886 -18179
rect 19920 -18213 19926 -18179
rect 19880 -18251 19926 -18213
rect 19880 -18285 19886 -18251
rect 19920 -18285 19926 -18251
rect 19880 -18323 19926 -18285
rect 19880 -18357 19886 -18323
rect 19920 -18357 19926 -18323
rect 19880 -18395 19926 -18357
rect 19880 -18429 19886 -18395
rect 19920 -18429 19926 -18395
rect 19880 -18462 19926 -18429
rect 20898 -17997 20904 -17986
rect 20938 -17986 20952 -17963
rect 21910 -17963 21970 -17752
rect 22414 -17854 22474 -17752
rect 22204 -17860 22692 -17854
rect 22204 -17894 22251 -17860
rect 22285 -17894 22323 -17860
rect 22357 -17894 22395 -17860
rect 22429 -17894 22467 -17860
rect 22501 -17894 22539 -17860
rect 22573 -17894 22611 -17860
rect 22645 -17894 22692 -17860
rect 22204 -17900 22692 -17894
rect 21910 -17978 21922 -17963
rect 20938 -17997 20944 -17986
rect 20898 -18035 20944 -17997
rect 20898 -18069 20904 -18035
rect 20938 -18069 20944 -18035
rect 20898 -18107 20944 -18069
rect 20898 -18141 20904 -18107
rect 20938 -18141 20944 -18107
rect 20898 -18179 20944 -18141
rect 20898 -18213 20904 -18179
rect 20938 -18213 20944 -18179
rect 20898 -18251 20944 -18213
rect 20898 -18285 20904 -18251
rect 20938 -18285 20944 -18251
rect 20898 -18323 20944 -18285
rect 20898 -18357 20904 -18323
rect 20938 -18357 20944 -18323
rect 20898 -18395 20944 -18357
rect 20898 -18429 20904 -18395
rect 20938 -18429 20944 -18395
rect 17884 -18501 17898 -18486
rect 17114 -18570 17602 -18564
rect 17114 -18604 17161 -18570
rect 17195 -18604 17233 -18570
rect 17267 -18604 17305 -18570
rect 17339 -18604 17377 -18570
rect 17411 -18604 17449 -18570
rect 17483 -18604 17521 -18570
rect 17555 -18604 17602 -18570
rect 17114 -18610 17602 -18604
rect 17314 -18880 17374 -18610
rect 17308 -18884 17380 -18880
rect 17308 -18936 17318 -18884
rect 17370 -18936 17380 -18884
rect 17308 -18940 17380 -18936
rect 17314 -19086 17374 -18940
rect 17114 -19092 17602 -19086
rect 17114 -19126 17161 -19092
rect 17195 -19126 17233 -19092
rect 17267 -19126 17305 -19092
rect 17339 -19126 17377 -19092
rect 17411 -19126 17449 -19092
rect 17483 -19126 17521 -19092
rect 17555 -19126 17602 -19092
rect 17114 -19132 17602 -19126
rect 16818 -19216 16832 -19195
rect 15802 -19267 15862 -19229
rect 15802 -19301 15814 -19267
rect 15848 -19301 15862 -19267
rect 15802 -19339 15862 -19301
rect 15802 -19373 15814 -19339
rect 15848 -19373 15862 -19339
rect 15802 -19411 15862 -19373
rect 15802 -19445 15814 -19411
rect 15848 -19445 15862 -19411
rect 15802 -19483 15862 -19445
rect 15802 -19517 15814 -19483
rect 15848 -19517 15862 -19483
rect 15802 -19555 15862 -19517
rect 15802 -19589 15814 -19555
rect 15848 -19589 15862 -19555
rect 15802 -19627 15862 -19589
rect 15802 -19661 15814 -19627
rect 15848 -19661 15862 -19627
rect 15802 -19699 15862 -19661
rect 14830 -19733 14842 -19720
rect 14060 -19802 14548 -19796
rect 14060 -19836 14107 -19802
rect 14141 -19836 14179 -19802
rect 14213 -19836 14251 -19802
rect 14285 -19836 14323 -19802
rect 14357 -19836 14395 -19802
rect 14429 -19836 14467 -19802
rect 14501 -19836 14548 -19802
rect 14060 -19842 14548 -19836
rect 14260 -20114 14320 -19842
rect 14782 -19892 14842 -19733
rect 15802 -19733 15814 -19699
rect 15848 -19733 15862 -19699
rect 16826 -19229 16832 -19216
rect 16866 -19216 16878 -19195
rect 17838 -19195 17898 -18501
rect 18862 -18501 18868 -18467
rect 18902 -18501 18908 -18467
rect 18862 -18532 18908 -18501
rect 19872 -18467 19932 -18462
rect 19872 -18501 19886 -18467
rect 19920 -18501 19932 -18467
rect 18344 -18564 18404 -18562
rect 18132 -18570 18620 -18564
rect 18132 -18604 18179 -18570
rect 18213 -18604 18251 -18570
rect 18285 -18604 18323 -18570
rect 18357 -18604 18395 -18570
rect 18429 -18604 18467 -18570
rect 18501 -18604 18539 -18570
rect 18573 -18604 18620 -18570
rect 18132 -18610 18620 -18604
rect 19150 -18570 19638 -18564
rect 19150 -18604 19197 -18570
rect 19231 -18604 19269 -18570
rect 19303 -18604 19341 -18570
rect 19375 -18604 19413 -18570
rect 19447 -18604 19485 -18570
rect 19519 -18604 19557 -18570
rect 19591 -18604 19638 -18570
rect 19150 -18610 19638 -18604
rect 18344 -18880 18404 -18610
rect 19366 -18658 19426 -18610
rect 19498 -18658 19570 -18654
rect 19360 -18662 19432 -18658
rect 19360 -18714 19370 -18662
rect 19422 -18714 19432 -18662
rect 19498 -18710 19508 -18658
rect 19560 -18710 19570 -18658
rect 19498 -18714 19570 -18710
rect 19360 -18718 19432 -18714
rect 19504 -18880 19564 -18714
rect 19872 -18880 19932 -18501
rect 20898 -18467 20944 -18429
rect 20898 -18501 20904 -18467
rect 20938 -18501 20944 -18467
rect 21916 -17997 21922 -17978
rect 21956 -17978 21970 -17963
rect 22924 -17963 22984 -17752
rect 23028 -17748 23100 -17744
rect 23028 -17800 23038 -17748
rect 23090 -17800 23100 -17748
rect 23028 -17804 23100 -17800
rect 22924 -17968 22940 -17963
rect 21956 -17997 21962 -17978
rect 21916 -18035 21962 -17997
rect 21916 -18069 21922 -18035
rect 21956 -18069 21962 -18035
rect 21916 -18107 21962 -18069
rect 21916 -18141 21922 -18107
rect 21956 -18141 21962 -18107
rect 21916 -18179 21962 -18141
rect 21916 -18213 21922 -18179
rect 21956 -18213 21962 -18179
rect 21916 -18251 21962 -18213
rect 21916 -18285 21922 -18251
rect 21956 -18285 21962 -18251
rect 21916 -18323 21962 -18285
rect 21916 -18357 21922 -18323
rect 21956 -18357 21962 -18323
rect 21916 -18395 21962 -18357
rect 21916 -18429 21922 -18395
rect 21956 -18429 21962 -18395
rect 21916 -18467 21962 -18429
rect 21916 -18480 21922 -18467
rect 20898 -18532 20944 -18501
rect 21910 -18501 21922 -18480
rect 21956 -18480 21962 -18467
rect 22934 -17997 22940 -17968
rect 22974 -17968 22984 -17963
rect 22974 -17997 22980 -17968
rect 22934 -18035 22980 -17997
rect 22934 -18069 22940 -18035
rect 22974 -18069 22980 -18035
rect 22934 -18107 22980 -18069
rect 22934 -18141 22940 -18107
rect 22974 -18141 22980 -18107
rect 22934 -18179 22980 -18141
rect 22934 -18213 22940 -18179
rect 22974 -18213 22980 -18179
rect 22934 -18251 22980 -18213
rect 22934 -18285 22940 -18251
rect 22974 -18285 22980 -18251
rect 22934 -18323 22980 -18285
rect 22934 -18357 22940 -18323
rect 22974 -18357 22980 -18323
rect 22934 -18395 22980 -18357
rect 22934 -18429 22940 -18395
rect 22974 -18429 22980 -18395
rect 22934 -18467 22980 -18429
rect 21956 -18501 21970 -18480
rect 20168 -18570 20656 -18564
rect 20168 -18604 20215 -18570
rect 20249 -18604 20287 -18570
rect 20321 -18604 20359 -18570
rect 20393 -18604 20431 -18570
rect 20465 -18604 20503 -18570
rect 20537 -18604 20575 -18570
rect 20609 -18604 20656 -18570
rect 20168 -18610 20656 -18604
rect 21186 -18570 21674 -18564
rect 21186 -18604 21233 -18570
rect 21267 -18604 21305 -18570
rect 21339 -18604 21377 -18570
rect 21411 -18604 21449 -18570
rect 21483 -18604 21521 -18570
rect 21555 -18604 21593 -18570
rect 21627 -18604 21674 -18570
rect 21186 -18610 21674 -18604
rect 21392 -18654 21452 -18610
rect 20380 -18658 20452 -18654
rect 20380 -18710 20390 -18658
rect 20442 -18710 20452 -18658
rect 20380 -18714 20452 -18710
rect 21386 -18658 21458 -18654
rect 21910 -18658 21970 -18501
rect 22934 -18501 22940 -18467
rect 22974 -18501 22980 -18467
rect 22934 -18532 22980 -18501
rect 22204 -18570 22692 -18564
rect 22204 -18604 22251 -18570
rect 22285 -18604 22323 -18570
rect 22357 -18604 22395 -18570
rect 22429 -18604 22467 -18570
rect 22501 -18604 22539 -18570
rect 22573 -18604 22611 -18570
rect 22645 -18604 22692 -18570
rect 22204 -18610 22692 -18604
rect 21386 -18710 21396 -18658
rect 21448 -18710 21458 -18658
rect 21386 -18714 21458 -18710
rect 21904 -18662 21976 -18658
rect 21904 -18714 21914 -18662
rect 21966 -18714 21976 -18662
rect 18338 -18884 18410 -18880
rect 18338 -18936 18348 -18884
rect 18400 -18936 18410 -18884
rect 18338 -18940 18410 -18936
rect 19498 -18884 19570 -18880
rect 19498 -18936 19508 -18884
rect 19560 -18936 19570 -18884
rect 19498 -18940 19570 -18936
rect 19866 -18884 19938 -18880
rect 19866 -18936 19876 -18884
rect 19928 -18936 19938 -18884
rect 19866 -18940 19938 -18936
rect 18344 -19086 18404 -18940
rect 19504 -19086 19564 -18940
rect 19872 -18984 19932 -18940
rect 19866 -18988 19938 -18984
rect 19866 -19040 19876 -18988
rect 19928 -19040 19938 -18988
rect 19866 -19044 19938 -19040
rect 20386 -19086 20446 -18714
rect 21904 -18718 21976 -18714
rect 21904 -18790 21976 -18786
rect 21904 -18842 21914 -18790
rect 21966 -18842 21976 -18790
rect 21904 -18846 21976 -18842
rect 20882 -18986 20954 -18982
rect 20882 -19038 20892 -18986
rect 20944 -19038 20954 -18986
rect 20882 -19042 20954 -19038
rect 18132 -19092 18620 -19086
rect 18132 -19126 18179 -19092
rect 18213 -19126 18251 -19092
rect 18285 -19126 18323 -19092
rect 18357 -19126 18395 -19092
rect 18429 -19126 18467 -19092
rect 18501 -19126 18539 -19092
rect 18573 -19126 18620 -19092
rect 18132 -19132 18620 -19126
rect 19150 -19092 19638 -19086
rect 19150 -19126 19197 -19092
rect 19231 -19126 19269 -19092
rect 19303 -19126 19341 -19092
rect 19375 -19126 19413 -19092
rect 19447 -19126 19485 -19092
rect 19519 -19126 19557 -19092
rect 19591 -19126 19638 -19092
rect 19150 -19132 19638 -19126
rect 20168 -19092 20656 -19086
rect 20168 -19126 20215 -19092
rect 20249 -19126 20287 -19092
rect 20321 -19126 20359 -19092
rect 20393 -19126 20431 -19092
rect 20465 -19126 20503 -19092
rect 20537 -19126 20575 -19092
rect 20609 -19126 20656 -19092
rect 20168 -19132 20656 -19126
rect 20386 -19134 20446 -19132
rect 16866 -19229 16872 -19216
rect 17838 -19222 17850 -19195
rect 16826 -19267 16872 -19229
rect 16826 -19301 16832 -19267
rect 16866 -19301 16872 -19267
rect 16826 -19339 16872 -19301
rect 16826 -19373 16832 -19339
rect 16866 -19373 16872 -19339
rect 16826 -19411 16872 -19373
rect 16826 -19445 16832 -19411
rect 16866 -19445 16872 -19411
rect 16826 -19483 16872 -19445
rect 16826 -19517 16832 -19483
rect 16866 -19517 16872 -19483
rect 16826 -19555 16872 -19517
rect 16826 -19589 16832 -19555
rect 16866 -19589 16872 -19555
rect 16826 -19627 16872 -19589
rect 16826 -19661 16832 -19627
rect 16866 -19661 16872 -19627
rect 16826 -19699 16872 -19661
rect 16826 -19720 16832 -19699
rect 15078 -19802 15566 -19796
rect 15078 -19836 15125 -19802
rect 15159 -19836 15197 -19802
rect 15231 -19836 15269 -19802
rect 15303 -19836 15341 -19802
rect 15375 -19836 15413 -19802
rect 15447 -19836 15485 -19802
rect 15519 -19836 15566 -19802
rect 15078 -19842 15566 -19836
rect 14776 -19896 14848 -19892
rect 14776 -19948 14786 -19896
rect 14838 -19948 14848 -19896
rect 14776 -19952 14848 -19948
rect 15278 -20114 15338 -19842
rect 14254 -20118 14326 -20114
rect 14254 -20170 14264 -20118
rect 14316 -20170 14326 -20118
rect 14254 -20174 14326 -20170
rect 15272 -20118 15344 -20114
rect 15272 -20170 15282 -20118
rect 15334 -20170 15344 -20118
rect 15272 -20174 15344 -20170
rect 13762 -20222 13834 -20218
rect 13762 -20274 13772 -20222
rect 13824 -20274 13834 -20222
rect 13762 -20278 13834 -20274
rect 12024 -20326 12512 -20320
rect 12024 -20360 12071 -20326
rect 12105 -20360 12143 -20326
rect 12177 -20360 12215 -20326
rect 12249 -20360 12287 -20326
rect 12321 -20360 12359 -20326
rect 12393 -20360 12431 -20326
rect 12465 -20360 12512 -20326
rect 12024 -20366 12512 -20360
rect 13042 -20326 13530 -20320
rect 13042 -20360 13089 -20326
rect 13123 -20360 13161 -20326
rect 13195 -20360 13233 -20326
rect 13267 -20360 13305 -20326
rect 13339 -20360 13377 -20326
rect 13411 -20360 13449 -20326
rect 13483 -20360 13530 -20326
rect 13042 -20366 13530 -20360
rect 10758 -20463 10764 -20446
rect 11730 -20448 11742 -20429
rect 8682 -20535 8688 -20501
rect 8722 -20535 8728 -20501
rect 8682 -20573 8728 -20535
rect 8682 -20607 8688 -20573
rect 8722 -20607 8728 -20573
rect 8682 -20645 8728 -20607
rect 8682 -20679 8688 -20645
rect 8722 -20679 8728 -20645
rect 8682 -20717 8728 -20679
rect 8682 -20751 8688 -20717
rect 8722 -20751 8728 -20717
rect 8682 -20789 8728 -20751
rect 8682 -20823 8688 -20789
rect 8722 -20823 8728 -20789
rect 8682 -20861 8728 -20823
rect 8682 -20895 8688 -20861
rect 8722 -20895 8728 -20861
rect 8682 -20933 8728 -20895
rect 7704 -20967 7720 -20940
rect 8682 -20942 8688 -20933
rect 6934 -21036 7422 -21030
rect 6934 -21070 6981 -21036
rect 7015 -21070 7053 -21036
rect 7087 -21070 7125 -21036
rect 7159 -21070 7197 -21036
rect 7231 -21070 7269 -21036
rect 7303 -21070 7341 -21036
rect 7375 -21070 7422 -21036
rect 6934 -21076 7422 -21070
rect 7144 -21126 7204 -21076
rect 7138 -21130 7210 -21126
rect 7138 -21182 7148 -21130
rect 7200 -21182 7210 -21130
rect 7138 -21186 7210 -21182
rect 6634 -21346 6706 -21342
rect 6634 -21398 6644 -21346
rect 6696 -21398 6706 -21346
rect 6634 -21402 6706 -21398
rect 5614 -21444 5686 -21440
rect 5614 -21496 5624 -21444
rect 5676 -21496 5686 -21444
rect 5614 -21500 5686 -21496
rect 7144 -21554 7204 -21186
rect 7660 -21440 7720 -20967
rect 8678 -20967 8688 -20942
rect 8722 -20942 8728 -20933
rect 9700 -20501 9746 -20474
rect 9700 -20535 9706 -20501
rect 9740 -20535 9746 -20501
rect 9700 -20573 9746 -20535
rect 9700 -20607 9706 -20573
rect 9740 -20607 9746 -20573
rect 9700 -20645 9746 -20607
rect 9700 -20679 9706 -20645
rect 9740 -20679 9746 -20645
rect 9700 -20717 9746 -20679
rect 9700 -20751 9706 -20717
rect 9740 -20751 9746 -20717
rect 9700 -20789 9746 -20751
rect 9700 -20823 9706 -20789
rect 9740 -20823 9746 -20789
rect 9700 -20861 9746 -20823
rect 9700 -20895 9706 -20861
rect 9740 -20895 9746 -20861
rect 9700 -20933 9746 -20895
rect 10718 -20501 10764 -20463
rect 10718 -20535 10724 -20501
rect 10758 -20535 10764 -20501
rect 10718 -20573 10764 -20535
rect 10718 -20607 10724 -20573
rect 10758 -20607 10764 -20573
rect 10718 -20645 10764 -20607
rect 10718 -20679 10724 -20645
rect 10758 -20679 10764 -20645
rect 10718 -20717 10764 -20679
rect 10718 -20751 10724 -20717
rect 10758 -20751 10764 -20717
rect 10718 -20789 10764 -20751
rect 10718 -20823 10724 -20789
rect 10758 -20823 10764 -20789
rect 10718 -20861 10764 -20823
rect 10718 -20895 10724 -20861
rect 10758 -20895 10764 -20861
rect 10718 -20928 10764 -20895
rect 11736 -20463 11742 -20448
rect 11776 -20448 11790 -20429
rect 12754 -20429 12800 -20398
rect 11776 -20463 11782 -20448
rect 11736 -20501 11782 -20463
rect 11736 -20535 11742 -20501
rect 11776 -20535 11782 -20501
rect 11736 -20573 11782 -20535
rect 11736 -20607 11742 -20573
rect 11776 -20607 11782 -20573
rect 11736 -20645 11782 -20607
rect 11736 -20679 11742 -20645
rect 11776 -20679 11782 -20645
rect 11736 -20717 11782 -20679
rect 11736 -20751 11742 -20717
rect 11776 -20751 11782 -20717
rect 11736 -20789 11782 -20751
rect 11736 -20823 11742 -20789
rect 11776 -20823 11782 -20789
rect 11736 -20861 11782 -20823
rect 11736 -20895 11742 -20861
rect 11776 -20895 11782 -20861
rect 8722 -20967 8738 -20942
rect 7952 -21036 8440 -21030
rect 7952 -21070 7999 -21036
rect 8033 -21070 8071 -21036
rect 8105 -21070 8143 -21036
rect 8177 -21070 8215 -21036
rect 8249 -21070 8287 -21036
rect 8321 -21070 8359 -21036
rect 8393 -21070 8440 -21036
rect 7952 -21076 8222 -21070
rect 8230 -21076 8440 -21070
rect 8162 -21126 8222 -21076
rect 8678 -21120 8738 -20967
rect 9700 -20967 9706 -20933
rect 9740 -20967 9746 -20933
rect 9700 -20998 9746 -20967
rect 10714 -20933 10774 -20928
rect 10714 -20967 10724 -20933
rect 10758 -20967 10774 -20933
rect 8970 -21036 9458 -21030
rect 8970 -21070 9017 -21036
rect 9051 -21070 9089 -21036
rect 9123 -21070 9161 -21036
rect 9195 -21070 9233 -21036
rect 9267 -21070 9305 -21036
rect 9339 -21070 9377 -21036
rect 9411 -21070 9458 -21036
rect 8970 -21076 9458 -21070
rect 9988 -21036 10476 -21030
rect 9988 -21070 10035 -21036
rect 10069 -21070 10107 -21036
rect 10141 -21070 10179 -21036
rect 10213 -21070 10251 -21036
rect 10285 -21070 10323 -21036
rect 10357 -21070 10395 -21036
rect 10429 -21070 10476 -21036
rect 9988 -21076 10476 -21070
rect 8672 -21124 8744 -21120
rect 8156 -21130 8228 -21126
rect 8156 -21182 8166 -21130
rect 8218 -21182 8228 -21130
rect 8672 -21176 8682 -21124
rect 8734 -21176 8744 -21124
rect 8672 -21180 8744 -21176
rect 10714 -21124 10774 -20967
rect 11736 -20933 11782 -20895
rect 11736 -20967 11742 -20933
rect 11776 -20967 11782 -20933
rect 12754 -20463 12760 -20429
rect 12794 -20463 12800 -20429
rect 13768 -20429 13828 -20278
rect 14260 -20320 14320 -20174
rect 15802 -20218 15862 -19733
rect 16820 -19733 16832 -19720
rect 16866 -19720 16872 -19699
rect 17844 -19229 17850 -19222
rect 17884 -19222 17898 -19195
rect 18862 -19195 18908 -19164
rect 17884 -19229 17890 -19222
rect 17844 -19267 17890 -19229
rect 17844 -19301 17850 -19267
rect 17884 -19301 17890 -19267
rect 17844 -19339 17890 -19301
rect 17844 -19373 17850 -19339
rect 17884 -19373 17890 -19339
rect 17844 -19411 17890 -19373
rect 17844 -19445 17850 -19411
rect 17884 -19445 17890 -19411
rect 17844 -19483 17890 -19445
rect 17844 -19517 17850 -19483
rect 17884 -19517 17890 -19483
rect 17844 -19555 17890 -19517
rect 17844 -19589 17850 -19555
rect 17884 -19589 17890 -19555
rect 17844 -19627 17890 -19589
rect 17844 -19661 17850 -19627
rect 17884 -19661 17890 -19627
rect 17844 -19699 17890 -19661
rect 17844 -19708 17850 -19699
rect 16866 -19733 16880 -19720
rect 16096 -19802 16584 -19796
rect 16096 -19836 16143 -19802
rect 16177 -19836 16215 -19802
rect 16249 -19836 16287 -19802
rect 16321 -19836 16359 -19802
rect 16393 -19836 16431 -19802
rect 16465 -19836 16503 -19802
rect 16537 -19836 16584 -19802
rect 16096 -19842 16584 -19836
rect 16312 -20114 16372 -19842
rect 16820 -19892 16880 -19733
rect 17836 -19733 17850 -19708
rect 17884 -19708 17890 -19699
rect 18862 -19229 18868 -19195
rect 18902 -19229 18908 -19195
rect 18862 -19267 18908 -19229
rect 18862 -19301 18868 -19267
rect 18902 -19301 18908 -19267
rect 18862 -19339 18908 -19301
rect 18862 -19373 18868 -19339
rect 18902 -19373 18908 -19339
rect 18862 -19411 18908 -19373
rect 18862 -19445 18868 -19411
rect 18902 -19445 18908 -19411
rect 18862 -19483 18908 -19445
rect 18862 -19517 18868 -19483
rect 18902 -19517 18908 -19483
rect 18862 -19555 18908 -19517
rect 18862 -19589 18868 -19555
rect 18902 -19589 18908 -19555
rect 18862 -19627 18908 -19589
rect 18862 -19661 18868 -19627
rect 18902 -19661 18908 -19627
rect 18862 -19699 18908 -19661
rect 17884 -19733 17896 -19708
rect 18862 -19712 18868 -19699
rect 17114 -19802 17602 -19796
rect 17114 -19836 17161 -19802
rect 17195 -19836 17233 -19802
rect 17267 -19836 17305 -19802
rect 17339 -19836 17377 -19802
rect 17411 -19836 17449 -19802
rect 17483 -19836 17521 -19802
rect 17555 -19836 17602 -19802
rect 17114 -19842 17602 -19836
rect 16814 -19896 16886 -19892
rect 16814 -19948 16824 -19896
rect 16876 -19948 16886 -19896
rect 16814 -19952 16886 -19948
rect 16806 -20004 16878 -20000
rect 16806 -20056 16816 -20004
rect 16868 -20056 16878 -20004
rect 16806 -20060 16878 -20056
rect 16306 -20118 16378 -20114
rect 16306 -20170 16316 -20118
rect 16368 -20170 16378 -20118
rect 16306 -20174 16378 -20170
rect 15796 -20222 15868 -20218
rect 15796 -20274 15806 -20222
rect 15858 -20274 15868 -20222
rect 15796 -20278 15868 -20274
rect 16308 -20226 16380 -20222
rect 16308 -20278 16318 -20226
rect 16370 -20278 16380 -20226
rect 16308 -20282 16380 -20278
rect 16314 -20320 16374 -20282
rect 14060 -20326 14548 -20320
rect 14060 -20360 14107 -20326
rect 14141 -20360 14179 -20326
rect 14213 -20360 14251 -20326
rect 14285 -20360 14323 -20326
rect 14357 -20360 14395 -20326
rect 14429 -20360 14467 -20326
rect 14501 -20360 14548 -20326
rect 14060 -20366 14548 -20360
rect 15078 -20326 15566 -20320
rect 15078 -20360 15125 -20326
rect 15159 -20360 15197 -20326
rect 15231 -20360 15269 -20326
rect 15303 -20360 15341 -20326
rect 15375 -20360 15413 -20326
rect 15447 -20360 15485 -20326
rect 15519 -20360 15566 -20326
rect 15078 -20366 15566 -20360
rect 16096 -20326 16584 -20320
rect 16096 -20360 16143 -20326
rect 16177 -20360 16215 -20326
rect 16249 -20360 16287 -20326
rect 16321 -20360 16359 -20326
rect 16393 -20360 16431 -20326
rect 16465 -20360 16503 -20326
rect 16537 -20360 16584 -20326
rect 16096 -20366 16584 -20360
rect 13768 -20446 13778 -20429
rect 12754 -20501 12800 -20463
rect 12754 -20535 12760 -20501
rect 12794 -20535 12800 -20501
rect 12754 -20573 12800 -20535
rect 12754 -20607 12760 -20573
rect 12794 -20607 12800 -20573
rect 12754 -20645 12800 -20607
rect 12754 -20679 12760 -20645
rect 12794 -20679 12800 -20645
rect 12754 -20717 12800 -20679
rect 12754 -20751 12760 -20717
rect 12794 -20751 12800 -20717
rect 12754 -20789 12800 -20751
rect 12754 -20823 12760 -20789
rect 12794 -20823 12800 -20789
rect 12754 -20861 12800 -20823
rect 12754 -20895 12760 -20861
rect 12794 -20895 12800 -20861
rect 12754 -20933 12800 -20895
rect 12754 -20936 12760 -20933
rect 11736 -20998 11782 -20967
rect 12746 -20967 12760 -20936
rect 12794 -20936 12800 -20933
rect 13772 -20463 13778 -20446
rect 13812 -20446 13828 -20429
rect 14790 -20429 14836 -20398
rect 13812 -20463 13818 -20446
rect 13772 -20501 13818 -20463
rect 13772 -20535 13778 -20501
rect 13812 -20535 13818 -20501
rect 13772 -20573 13818 -20535
rect 13772 -20607 13778 -20573
rect 13812 -20607 13818 -20573
rect 13772 -20645 13818 -20607
rect 13772 -20679 13778 -20645
rect 13812 -20679 13818 -20645
rect 13772 -20717 13818 -20679
rect 13772 -20751 13778 -20717
rect 13812 -20751 13818 -20717
rect 13772 -20789 13818 -20751
rect 13772 -20823 13778 -20789
rect 13812 -20823 13818 -20789
rect 13772 -20861 13818 -20823
rect 13772 -20895 13778 -20861
rect 13812 -20895 13818 -20861
rect 13772 -20933 13818 -20895
rect 14790 -20463 14796 -20429
rect 14830 -20463 14836 -20429
rect 14790 -20501 14836 -20463
rect 14790 -20535 14796 -20501
rect 14830 -20535 14836 -20501
rect 14790 -20573 14836 -20535
rect 14790 -20607 14796 -20573
rect 14830 -20607 14836 -20573
rect 14790 -20645 14836 -20607
rect 14790 -20679 14796 -20645
rect 14830 -20679 14836 -20645
rect 14790 -20717 14836 -20679
rect 14790 -20751 14796 -20717
rect 14830 -20751 14836 -20717
rect 14790 -20789 14836 -20751
rect 14790 -20823 14796 -20789
rect 14830 -20823 14836 -20789
rect 14790 -20861 14836 -20823
rect 14790 -20895 14796 -20861
rect 14830 -20895 14836 -20861
rect 14790 -20924 14836 -20895
rect 15808 -20429 15854 -20398
rect 15808 -20463 15814 -20429
rect 15848 -20463 15854 -20429
rect 16812 -20429 16872 -20060
rect 17336 -20222 17396 -19842
rect 17836 -20216 17896 -19733
rect 18856 -19733 18868 -19712
rect 18902 -19712 18908 -19699
rect 19880 -19195 19926 -19164
rect 19880 -19229 19886 -19195
rect 19920 -19229 19926 -19195
rect 20888 -19195 20948 -19042
rect 21186 -19092 21674 -19086
rect 21186 -19126 21233 -19092
rect 21267 -19126 21305 -19092
rect 21339 -19126 21377 -19092
rect 21411 -19126 21449 -19092
rect 21483 -19126 21521 -19092
rect 21555 -19126 21593 -19092
rect 21627 -19126 21674 -19092
rect 21186 -19132 21674 -19126
rect 20888 -19226 20904 -19195
rect 19880 -19267 19926 -19229
rect 19880 -19301 19886 -19267
rect 19920 -19301 19926 -19267
rect 19880 -19339 19926 -19301
rect 19880 -19373 19886 -19339
rect 19920 -19373 19926 -19339
rect 19880 -19411 19926 -19373
rect 19880 -19445 19886 -19411
rect 19920 -19445 19926 -19411
rect 19880 -19483 19926 -19445
rect 19880 -19517 19886 -19483
rect 19920 -19517 19926 -19483
rect 19880 -19555 19926 -19517
rect 19880 -19589 19886 -19555
rect 19920 -19589 19926 -19555
rect 19880 -19627 19926 -19589
rect 19880 -19661 19886 -19627
rect 19920 -19661 19926 -19627
rect 19880 -19699 19926 -19661
rect 19880 -19708 19886 -19699
rect 18902 -19733 18916 -19712
rect 18132 -19802 18620 -19796
rect 18132 -19836 18179 -19802
rect 18213 -19836 18251 -19802
rect 18285 -19836 18323 -19802
rect 18357 -19836 18395 -19802
rect 18429 -19836 18467 -19802
rect 18501 -19836 18539 -19802
rect 18573 -19836 18620 -19802
rect 18132 -19842 18620 -19836
rect 17830 -20220 17902 -20216
rect 17330 -20226 17402 -20222
rect 17330 -20278 17340 -20226
rect 17392 -20278 17402 -20226
rect 17830 -20272 17840 -20220
rect 17892 -20272 17902 -20220
rect 17830 -20276 17902 -20272
rect 17330 -20282 17402 -20278
rect 17336 -20320 17396 -20282
rect 17114 -20326 17602 -20320
rect 17114 -20360 17161 -20326
rect 17195 -20360 17233 -20326
rect 17267 -20360 17305 -20326
rect 17339 -20360 17377 -20326
rect 17411 -20360 17449 -20326
rect 17483 -20360 17521 -20326
rect 17555 -20360 17602 -20326
rect 17114 -20366 17602 -20360
rect 16812 -20446 16832 -20429
rect 15808 -20501 15854 -20463
rect 15808 -20535 15814 -20501
rect 15848 -20535 15854 -20501
rect 15808 -20573 15854 -20535
rect 15808 -20607 15814 -20573
rect 15848 -20607 15854 -20573
rect 15808 -20645 15854 -20607
rect 15808 -20679 15814 -20645
rect 15848 -20679 15854 -20645
rect 15808 -20717 15854 -20679
rect 15808 -20751 15814 -20717
rect 15848 -20751 15854 -20717
rect 15808 -20789 15854 -20751
rect 15808 -20823 15814 -20789
rect 15848 -20823 15854 -20789
rect 15808 -20861 15854 -20823
rect 15808 -20895 15814 -20861
rect 15848 -20895 15854 -20861
rect 12794 -20967 12806 -20936
rect 11006 -21036 11494 -21030
rect 11006 -21070 11053 -21036
rect 11087 -21070 11125 -21036
rect 11159 -21070 11197 -21036
rect 11231 -21070 11269 -21036
rect 11303 -21070 11341 -21036
rect 11375 -21070 11413 -21036
rect 11447 -21070 11494 -21036
rect 11006 -21076 11494 -21070
rect 12024 -21036 12512 -21030
rect 12024 -21070 12071 -21036
rect 12105 -21070 12143 -21036
rect 12177 -21070 12215 -21036
rect 12249 -21070 12287 -21036
rect 12321 -21070 12359 -21036
rect 12393 -21070 12431 -21036
rect 12465 -21070 12512 -21036
rect 12024 -21076 12512 -21070
rect 12746 -21120 12806 -20967
rect 13772 -20967 13778 -20933
rect 13812 -20967 13818 -20933
rect 13772 -20998 13818 -20967
rect 14780 -20933 14840 -20924
rect 14780 -20967 14796 -20933
rect 14830 -20967 14840 -20933
rect 15808 -20933 15854 -20895
rect 15808 -20944 15814 -20933
rect 13042 -21036 13530 -21030
rect 13042 -21070 13089 -21036
rect 13123 -21070 13161 -21036
rect 13195 -21070 13233 -21036
rect 13267 -21070 13305 -21036
rect 13339 -21070 13377 -21036
rect 13411 -21070 13449 -21036
rect 13483 -21070 13530 -21036
rect 13042 -21076 13530 -21070
rect 14060 -21036 14548 -21030
rect 14060 -21070 14107 -21036
rect 14141 -21070 14179 -21036
rect 14213 -21070 14251 -21036
rect 14285 -21070 14323 -21036
rect 14357 -21070 14395 -21036
rect 14429 -21070 14467 -21036
rect 14501 -21070 14548 -21036
rect 14060 -21076 14548 -21070
rect 14780 -21120 14840 -20967
rect 15802 -20967 15814 -20944
rect 15848 -20944 15854 -20933
rect 16826 -20463 16832 -20446
rect 16866 -20463 16872 -20429
rect 16826 -20501 16872 -20463
rect 16826 -20535 16832 -20501
rect 16866 -20535 16872 -20501
rect 17836 -20429 17896 -20276
rect 18314 -20320 18374 -19842
rect 18856 -19892 18916 -19733
rect 19870 -19733 19886 -19708
rect 19920 -19708 19926 -19699
rect 20898 -19229 20904 -19226
rect 20938 -19226 20948 -19195
rect 21910 -19195 21970 -18846
rect 22204 -19092 22692 -19086
rect 22204 -19126 22251 -19092
rect 22285 -19126 22323 -19092
rect 22357 -19126 22395 -19092
rect 22429 -19126 22467 -19092
rect 22501 -19126 22539 -19092
rect 22573 -19126 22611 -19092
rect 22645 -19126 22692 -19092
rect 22204 -19132 22692 -19126
rect 20938 -19229 20944 -19226
rect 21910 -19228 21922 -19195
rect 20898 -19267 20944 -19229
rect 20898 -19301 20904 -19267
rect 20938 -19301 20944 -19267
rect 20898 -19339 20944 -19301
rect 20898 -19373 20904 -19339
rect 20938 -19373 20944 -19339
rect 20898 -19411 20944 -19373
rect 20898 -19445 20904 -19411
rect 20938 -19445 20944 -19411
rect 20898 -19483 20944 -19445
rect 20898 -19517 20904 -19483
rect 20938 -19517 20944 -19483
rect 20898 -19555 20944 -19517
rect 20898 -19589 20904 -19555
rect 20938 -19589 20944 -19555
rect 20898 -19627 20944 -19589
rect 20898 -19661 20904 -19627
rect 20938 -19661 20944 -19627
rect 20898 -19699 20944 -19661
rect 19920 -19733 19930 -19708
rect 20898 -19724 20904 -19699
rect 19150 -19802 19638 -19796
rect 19150 -19836 19197 -19802
rect 19231 -19836 19269 -19802
rect 19303 -19836 19341 -19802
rect 19375 -19836 19413 -19802
rect 19447 -19836 19485 -19802
rect 19519 -19836 19557 -19802
rect 19591 -19836 19638 -19802
rect 19150 -19842 19638 -19836
rect 18850 -19896 18922 -19892
rect 18850 -19948 18860 -19896
rect 18912 -19948 18922 -19896
rect 18850 -19952 18922 -19948
rect 18846 -20004 18918 -20000
rect 18846 -20056 18856 -20004
rect 18908 -20056 18918 -20004
rect 18846 -20060 18918 -20056
rect 18132 -20326 18620 -20320
rect 18132 -20360 18179 -20326
rect 18213 -20360 18251 -20326
rect 18285 -20360 18323 -20326
rect 18357 -20360 18395 -20326
rect 18429 -20360 18467 -20326
rect 18501 -20360 18539 -20326
rect 18573 -20360 18620 -20326
rect 18132 -20366 18620 -20360
rect 17836 -20463 17850 -20429
rect 17884 -20463 17896 -20429
rect 17836 -20501 17896 -20463
rect 18852 -20429 18912 -20060
rect 19338 -20118 19410 -20114
rect 19338 -20170 19348 -20118
rect 19400 -20170 19410 -20118
rect 19338 -20174 19410 -20170
rect 19344 -20320 19404 -20174
rect 19870 -20216 19930 -19733
rect 20894 -19733 20904 -19724
rect 20938 -19724 20944 -19699
rect 21916 -19229 21922 -19228
rect 21956 -19228 21970 -19195
rect 22934 -19195 22980 -19164
rect 21956 -19229 21962 -19228
rect 21916 -19267 21962 -19229
rect 21916 -19301 21922 -19267
rect 21956 -19301 21962 -19267
rect 21916 -19339 21962 -19301
rect 21916 -19373 21922 -19339
rect 21956 -19373 21962 -19339
rect 21916 -19411 21962 -19373
rect 21916 -19445 21922 -19411
rect 21956 -19445 21962 -19411
rect 21916 -19483 21962 -19445
rect 21916 -19517 21922 -19483
rect 21956 -19517 21962 -19483
rect 21916 -19555 21962 -19517
rect 21916 -19589 21922 -19555
rect 21956 -19589 21962 -19555
rect 21916 -19627 21962 -19589
rect 21916 -19661 21922 -19627
rect 21956 -19661 21962 -19627
rect 21916 -19699 21962 -19661
rect 21916 -19724 21922 -19699
rect 20938 -19733 20954 -19724
rect 20168 -19802 20656 -19796
rect 20168 -19836 20215 -19802
rect 20249 -19836 20287 -19802
rect 20321 -19836 20359 -19802
rect 20393 -19836 20431 -19802
rect 20465 -19836 20503 -19802
rect 20537 -19836 20575 -19802
rect 20609 -19836 20656 -19802
rect 20168 -19842 20656 -19836
rect 20894 -19892 20954 -19733
rect 21910 -19733 21922 -19724
rect 21956 -19724 21962 -19699
rect 22934 -19229 22940 -19195
rect 22974 -19229 22980 -19195
rect 22934 -19267 22980 -19229
rect 22934 -19301 22940 -19267
rect 22974 -19301 22980 -19267
rect 22934 -19339 22980 -19301
rect 22934 -19373 22940 -19339
rect 22974 -19373 22980 -19339
rect 22934 -19411 22980 -19373
rect 22934 -19445 22940 -19411
rect 22974 -19445 22980 -19411
rect 22934 -19483 22980 -19445
rect 22934 -19517 22940 -19483
rect 22974 -19517 22980 -19483
rect 22934 -19555 22980 -19517
rect 22934 -19589 22940 -19555
rect 22974 -19589 22980 -19555
rect 22934 -19627 22980 -19589
rect 22934 -19661 22940 -19627
rect 22974 -19661 22980 -19627
rect 22934 -19699 22980 -19661
rect 22934 -19718 22940 -19699
rect 21956 -19733 21970 -19724
rect 21186 -19802 21674 -19796
rect 21186 -19836 21233 -19802
rect 21267 -19836 21305 -19802
rect 21339 -19836 21377 -19802
rect 21411 -19836 21449 -19802
rect 21483 -19836 21521 -19802
rect 21555 -19836 21593 -19802
rect 21627 -19836 21674 -19802
rect 21186 -19842 21674 -19836
rect 20888 -19896 20960 -19892
rect 20888 -19948 20898 -19896
rect 20950 -19948 20960 -19896
rect 20888 -19952 20960 -19948
rect 20884 -20004 20956 -20000
rect 20884 -20056 20894 -20004
rect 20946 -20056 20956 -20004
rect 20884 -20060 20956 -20056
rect 20376 -20118 20448 -20114
rect 20376 -20170 20386 -20118
rect 20438 -20170 20448 -20118
rect 20376 -20174 20448 -20170
rect 19864 -20220 19936 -20216
rect 19864 -20272 19874 -20220
rect 19926 -20272 19936 -20220
rect 19864 -20276 19936 -20272
rect 20382 -20320 20442 -20174
rect 19150 -20326 19638 -20320
rect 19150 -20360 19197 -20326
rect 19231 -20360 19269 -20326
rect 19303 -20360 19341 -20326
rect 19375 -20360 19413 -20326
rect 19447 -20360 19485 -20326
rect 19519 -20360 19557 -20326
rect 19591 -20360 19638 -20326
rect 19150 -20366 19638 -20360
rect 20168 -20326 20656 -20320
rect 20168 -20360 20215 -20326
rect 20249 -20360 20287 -20326
rect 20321 -20360 20359 -20326
rect 20393 -20360 20431 -20326
rect 20465 -20360 20503 -20326
rect 20537 -20360 20575 -20326
rect 20609 -20360 20656 -20326
rect 20168 -20366 20656 -20360
rect 18852 -20463 18868 -20429
rect 18902 -20463 18912 -20429
rect 18852 -20476 18912 -20463
rect 19880 -20429 19926 -20398
rect 19880 -20463 19886 -20429
rect 19920 -20463 19926 -20429
rect 20890 -20429 20950 -20060
rect 21408 -20114 21468 -19842
rect 21910 -19934 21970 -19733
rect 22924 -19733 22940 -19718
rect 22974 -19718 22980 -19699
rect 22974 -19733 22984 -19718
rect 22204 -19802 22692 -19796
rect 22204 -19836 22251 -19802
rect 22285 -19836 22323 -19802
rect 22357 -19836 22395 -19802
rect 22429 -19836 22467 -19802
rect 22501 -19836 22539 -19802
rect 22573 -19836 22611 -19802
rect 22645 -19836 22692 -19802
rect 22204 -19842 22692 -19836
rect 22418 -19934 22478 -19842
rect 22924 -19934 22984 -19733
rect 21910 -19994 22984 -19934
rect 21402 -20118 21474 -20114
rect 21402 -20170 21412 -20118
rect 21464 -20170 21474 -20118
rect 21402 -20174 21474 -20170
rect 21906 -20220 21978 -20216
rect 21906 -20272 21916 -20220
rect 21968 -20272 21978 -20220
rect 21906 -20276 21978 -20272
rect 21186 -20326 21674 -20320
rect 21186 -20360 21233 -20326
rect 21267 -20360 21305 -20326
rect 21339 -20360 21377 -20326
rect 21411 -20360 21449 -20326
rect 21483 -20360 21521 -20326
rect 21555 -20360 21593 -20326
rect 21627 -20360 21674 -20326
rect 21186 -20366 21674 -20360
rect 20890 -20462 20904 -20429
rect 17836 -20504 17850 -20501
rect 16826 -20573 16872 -20535
rect 16826 -20607 16832 -20573
rect 16866 -20607 16872 -20573
rect 16826 -20645 16872 -20607
rect 16826 -20679 16832 -20645
rect 16866 -20679 16872 -20645
rect 16826 -20717 16872 -20679
rect 16826 -20751 16832 -20717
rect 16866 -20751 16872 -20717
rect 16826 -20789 16872 -20751
rect 16826 -20823 16832 -20789
rect 16866 -20823 16872 -20789
rect 16826 -20861 16872 -20823
rect 16826 -20895 16832 -20861
rect 16866 -20895 16872 -20861
rect 16826 -20933 16872 -20895
rect 15848 -20967 15862 -20944
rect 15078 -21036 15566 -21030
rect 15078 -21070 15125 -21036
rect 15159 -21070 15197 -21036
rect 15231 -21070 15269 -21036
rect 15303 -21070 15341 -21036
rect 15375 -21070 15413 -21036
rect 15447 -21070 15485 -21036
rect 15519 -21070 15566 -21036
rect 15078 -21076 15566 -21070
rect 10714 -21176 10718 -21124
rect 10770 -21176 10774 -21124
rect 8156 -21186 8228 -21182
rect 7654 -21444 7726 -21440
rect 7654 -21496 7664 -21444
rect 7716 -21496 7726 -21444
rect 7654 -21500 7726 -21496
rect 3880 -21560 4368 -21554
rect 3880 -21594 3927 -21560
rect 3961 -21594 3999 -21560
rect 4033 -21594 4071 -21560
rect 4105 -21594 4143 -21560
rect 4177 -21594 4215 -21560
rect 4249 -21594 4287 -21560
rect 4321 -21594 4368 -21560
rect 3880 -21600 4368 -21594
rect 4898 -21560 5386 -21554
rect 4898 -21594 4945 -21560
rect 4979 -21594 5017 -21560
rect 5051 -21594 5089 -21560
rect 5123 -21594 5161 -21560
rect 5195 -21594 5233 -21560
rect 5267 -21594 5305 -21560
rect 5339 -21594 5386 -21560
rect 4898 -21600 5386 -21594
rect 5916 -21560 6404 -21554
rect 5916 -21594 5963 -21560
rect 5997 -21594 6035 -21560
rect 6069 -21594 6107 -21560
rect 6141 -21594 6179 -21560
rect 6213 -21594 6251 -21560
rect 6285 -21594 6323 -21560
rect 6357 -21594 6404 -21560
rect 5916 -21600 6404 -21594
rect 6934 -21560 7422 -21554
rect 6934 -21594 6981 -21560
rect 7015 -21594 7053 -21560
rect 7087 -21594 7125 -21560
rect 7159 -21594 7197 -21560
rect 7231 -21594 7269 -21560
rect 7303 -21594 7341 -21560
rect 7375 -21594 7422 -21560
rect 6934 -21600 7422 -21594
rect 3582 -21697 3598 -21663
rect 3632 -21697 3642 -21663
rect 3582 -21698 3642 -21697
rect 4610 -21663 4656 -21632
rect 4610 -21697 4616 -21663
rect 4650 -21697 4656 -21663
rect 2574 -21769 2580 -21735
rect 2614 -21769 2620 -21735
rect 2574 -21807 2620 -21769
rect 2574 -21841 2580 -21807
rect 2614 -21841 2620 -21807
rect 2574 -21879 2620 -21841
rect 2574 -21913 2580 -21879
rect 2614 -21913 2620 -21879
rect 2574 -21951 2620 -21913
rect 2574 -21985 2580 -21951
rect 2614 -21985 2620 -21951
rect 2574 -22023 2620 -21985
rect 2574 -22057 2580 -22023
rect 2614 -22057 2620 -22023
rect 2574 -22095 2620 -22057
rect 2574 -22129 2580 -22095
rect 2614 -22129 2620 -22095
rect 2574 -22167 2620 -22129
rect 2574 -22186 2580 -22167
rect 2564 -22201 2580 -22186
rect 2614 -22186 2620 -22167
rect 3592 -21735 3638 -21698
rect 3592 -21769 3598 -21735
rect 3632 -21769 3638 -21735
rect 3592 -21807 3638 -21769
rect 3592 -21841 3598 -21807
rect 3632 -21841 3638 -21807
rect 3592 -21879 3638 -21841
rect 3592 -21913 3598 -21879
rect 3632 -21913 3638 -21879
rect 3592 -21951 3638 -21913
rect 3592 -21985 3598 -21951
rect 3632 -21985 3638 -21951
rect 3592 -22023 3638 -21985
rect 3592 -22057 3598 -22023
rect 3632 -22057 3638 -22023
rect 3592 -22095 3638 -22057
rect 3592 -22129 3598 -22095
rect 3632 -22129 3638 -22095
rect 3592 -22167 3638 -22129
rect 2614 -22201 2624 -22186
rect 3592 -22190 3598 -22167
rect 2564 -22352 2624 -22201
rect 3588 -22201 3598 -22190
rect 3632 -22190 3638 -22167
rect 4610 -21735 4656 -21697
rect 4610 -21769 4616 -21735
rect 4650 -21769 4656 -21735
rect 4610 -21807 4656 -21769
rect 4610 -21841 4616 -21807
rect 4650 -21841 4656 -21807
rect 4610 -21879 4656 -21841
rect 4610 -21913 4616 -21879
rect 4650 -21913 4656 -21879
rect 4610 -21951 4656 -21913
rect 4610 -21985 4616 -21951
rect 4650 -21985 4656 -21951
rect 4610 -22023 4656 -21985
rect 4610 -22057 4616 -22023
rect 4650 -22057 4656 -22023
rect 4610 -22095 4656 -22057
rect 4610 -22129 4616 -22095
rect 4650 -22129 4656 -22095
rect 4610 -22167 4656 -22129
rect 4610 -22174 4616 -22167
rect 3632 -22201 3648 -22190
rect 2862 -22270 3350 -22264
rect 2862 -22304 2909 -22270
rect 2943 -22304 2981 -22270
rect 3015 -22304 3053 -22270
rect 3087 -22304 3125 -22270
rect 3159 -22304 3197 -22270
rect 3231 -22304 3269 -22270
rect 3303 -22304 3350 -22270
rect 2862 -22310 3350 -22304
rect 3084 -22352 3144 -22310
rect 3588 -22352 3648 -22201
rect 4602 -22201 4616 -22174
rect 4650 -22174 4656 -22167
rect 5628 -21663 5674 -21632
rect 5628 -21697 5634 -21663
rect 5668 -21697 5674 -21663
rect 5628 -21735 5674 -21697
rect 5628 -21769 5634 -21735
rect 5668 -21769 5674 -21735
rect 5628 -21807 5674 -21769
rect 5628 -21841 5634 -21807
rect 5668 -21841 5674 -21807
rect 5628 -21879 5674 -21841
rect 5628 -21913 5634 -21879
rect 5668 -21913 5674 -21879
rect 5628 -21951 5674 -21913
rect 5628 -21985 5634 -21951
rect 5668 -21985 5674 -21951
rect 5628 -22023 5674 -21985
rect 5628 -22057 5634 -22023
rect 5668 -22057 5674 -22023
rect 5628 -22095 5674 -22057
rect 5628 -22129 5634 -22095
rect 5668 -22129 5674 -22095
rect 5628 -22167 5674 -22129
rect 4650 -22201 4662 -22174
rect 5628 -22190 5634 -22167
rect 3880 -22270 4368 -22264
rect 3880 -22304 3927 -22270
rect 3961 -22304 3999 -22270
rect 4033 -22304 4071 -22270
rect 4105 -22304 4143 -22270
rect 4177 -22304 4215 -22270
rect 4249 -22304 4287 -22270
rect 4321 -22304 4368 -22270
rect 3880 -22310 4368 -22304
rect 2564 -22412 3648 -22352
rect 2442 -22466 2514 -22462
rect 2442 -22518 2452 -22466
rect 2504 -22518 2514 -22466
rect 2442 -22522 2514 -22518
rect 3588 -22558 3648 -22412
rect 2564 -22618 3648 -22558
rect 2564 -22895 2624 -22618
rect 3076 -22786 3136 -22618
rect 3588 -22678 3648 -22618
rect 3582 -22682 3654 -22678
rect 3582 -22734 3592 -22682
rect 3644 -22734 3654 -22682
rect 3582 -22738 3654 -22734
rect 2862 -22792 3350 -22786
rect 2862 -22826 2909 -22792
rect 2943 -22826 2981 -22792
rect 3015 -22826 3053 -22792
rect 3087 -22826 3125 -22792
rect 3159 -22826 3197 -22792
rect 3231 -22826 3269 -22792
rect 3303 -22826 3350 -22792
rect 2862 -22832 3350 -22826
rect 2564 -22912 2580 -22895
rect 2574 -22929 2580 -22912
rect 2614 -22912 2624 -22895
rect 3588 -22895 3648 -22738
rect 4080 -22786 4140 -22310
rect 4602 -22364 4662 -22201
rect 5620 -22201 5634 -22190
rect 5668 -22190 5674 -22167
rect 6646 -21663 6692 -21632
rect 6646 -21697 6652 -21663
rect 6686 -21697 6692 -21663
rect 7660 -21663 7720 -21500
rect 8162 -21554 8222 -21186
rect 7952 -21560 8440 -21554
rect 7952 -21594 7999 -21560
rect 8033 -21594 8071 -21560
rect 8105 -21594 8143 -21560
rect 8177 -21594 8215 -21560
rect 8249 -21594 8287 -21560
rect 8321 -21594 8359 -21560
rect 8393 -21594 8440 -21560
rect 7952 -21600 8440 -21594
rect 7660 -21674 7670 -21663
rect 6646 -21735 6692 -21697
rect 6646 -21769 6652 -21735
rect 6686 -21769 6692 -21735
rect 6646 -21807 6692 -21769
rect 6646 -21841 6652 -21807
rect 6686 -21841 6692 -21807
rect 6646 -21879 6692 -21841
rect 6646 -21913 6652 -21879
rect 6686 -21913 6692 -21879
rect 6646 -21951 6692 -21913
rect 6646 -21985 6652 -21951
rect 6686 -21985 6692 -21951
rect 6646 -22023 6692 -21985
rect 6646 -22057 6652 -22023
rect 6686 -22057 6692 -22023
rect 6646 -22095 6692 -22057
rect 6646 -22129 6652 -22095
rect 6686 -22129 6692 -22095
rect 6646 -22167 6692 -22129
rect 7664 -21697 7670 -21674
rect 7704 -21674 7720 -21663
rect 8678 -21663 8738 -21180
rect 10714 -21186 10774 -21176
rect 12740 -21124 12812 -21120
rect 12740 -21176 12750 -21124
rect 12802 -21176 12812 -21124
rect 12740 -21180 12812 -21176
rect 14774 -21124 14846 -21120
rect 14774 -21176 14784 -21124
rect 14836 -21176 14846 -21124
rect 14774 -21180 14846 -21176
rect 11724 -21234 11796 -21230
rect 11724 -21286 11734 -21234
rect 11786 -21286 11796 -21234
rect 11724 -21290 11796 -21286
rect 13760 -21234 13832 -21230
rect 13760 -21286 13770 -21234
rect 13822 -21286 13832 -21234
rect 13760 -21290 13832 -21286
rect 10706 -21346 10778 -21342
rect 10706 -21398 10716 -21346
rect 10768 -21398 10778 -21346
rect 10706 -21402 10778 -21398
rect 9690 -21444 9762 -21440
rect 9690 -21496 9700 -21444
rect 9752 -21496 9762 -21444
rect 9690 -21500 9762 -21496
rect 8970 -21560 9458 -21554
rect 8970 -21594 9017 -21560
rect 9051 -21594 9089 -21560
rect 9123 -21594 9161 -21560
rect 9195 -21594 9233 -21560
rect 9267 -21594 9305 -21560
rect 9339 -21594 9377 -21560
rect 9411 -21594 9458 -21560
rect 8970 -21600 9458 -21594
rect 7704 -21697 7710 -21674
rect 8678 -21686 8688 -21663
rect 7664 -21735 7710 -21697
rect 7664 -21769 7670 -21735
rect 7704 -21769 7710 -21735
rect 7664 -21807 7710 -21769
rect 7664 -21841 7670 -21807
rect 7704 -21841 7710 -21807
rect 7664 -21879 7710 -21841
rect 7664 -21913 7670 -21879
rect 7704 -21913 7710 -21879
rect 7664 -21951 7710 -21913
rect 7664 -21985 7670 -21951
rect 7704 -21985 7710 -21951
rect 7664 -22023 7710 -21985
rect 7664 -22057 7670 -22023
rect 7704 -22057 7710 -22023
rect 7664 -22095 7710 -22057
rect 7664 -22129 7670 -22095
rect 7704 -22129 7710 -22095
rect 7664 -22156 7710 -22129
rect 8682 -21697 8688 -21686
rect 8722 -21686 8738 -21663
rect 9696 -21663 9756 -21500
rect 9988 -21560 10476 -21554
rect 9988 -21594 10035 -21560
rect 10069 -21594 10107 -21560
rect 10141 -21594 10179 -21560
rect 10213 -21594 10251 -21560
rect 10285 -21594 10323 -21560
rect 10357 -21594 10395 -21560
rect 10429 -21594 10476 -21560
rect 9988 -21600 10476 -21594
rect 9696 -21680 9706 -21663
rect 8722 -21697 8728 -21686
rect 8682 -21735 8728 -21697
rect 8682 -21769 8688 -21735
rect 8722 -21769 8728 -21735
rect 8682 -21807 8728 -21769
rect 8682 -21841 8688 -21807
rect 8722 -21841 8728 -21807
rect 8682 -21879 8728 -21841
rect 8682 -21913 8688 -21879
rect 8722 -21913 8728 -21879
rect 8682 -21951 8728 -21913
rect 8682 -21985 8688 -21951
rect 8722 -21985 8728 -21951
rect 8682 -22023 8728 -21985
rect 8682 -22057 8688 -22023
rect 8722 -22057 8728 -22023
rect 8682 -22095 8728 -22057
rect 8682 -22129 8688 -22095
rect 8722 -22129 8728 -22095
rect 6646 -22178 6652 -22167
rect 5668 -22201 5680 -22190
rect 4898 -22270 5386 -22264
rect 4898 -22304 4945 -22270
rect 4979 -22304 5017 -22270
rect 5051 -22304 5089 -22270
rect 5123 -22304 5161 -22270
rect 5195 -22304 5233 -22270
rect 5267 -22304 5305 -22270
rect 5339 -22304 5386 -22270
rect 4898 -22310 5386 -22304
rect 4596 -22368 4668 -22364
rect 4596 -22420 4606 -22368
rect 4658 -22420 4668 -22368
rect 4596 -22424 4668 -22420
rect 4600 -22562 4672 -22558
rect 4600 -22614 4610 -22562
rect 4662 -22614 4672 -22562
rect 4600 -22618 4672 -22614
rect 3880 -22792 4368 -22786
rect 3880 -22826 3927 -22792
rect 3961 -22826 3999 -22792
rect 4033 -22826 4071 -22792
rect 4105 -22826 4143 -22792
rect 4177 -22826 4215 -22792
rect 4249 -22826 4287 -22792
rect 4321 -22826 4368 -22792
rect 3880 -22832 4368 -22826
rect 2614 -22929 2620 -22912
rect 3588 -22916 3598 -22895
rect 2574 -22967 2620 -22929
rect 2574 -23001 2580 -22967
rect 2614 -23001 2620 -22967
rect 2574 -23039 2620 -23001
rect 2574 -23073 2580 -23039
rect 2614 -23073 2620 -23039
rect 2574 -23111 2620 -23073
rect 2574 -23145 2580 -23111
rect 2614 -23145 2620 -23111
rect 2574 -23183 2620 -23145
rect 2574 -23217 2580 -23183
rect 2614 -23217 2620 -23183
rect 2574 -23255 2620 -23217
rect 2574 -23289 2580 -23255
rect 2614 -23289 2620 -23255
rect 2574 -23327 2620 -23289
rect 2574 -23361 2580 -23327
rect 2614 -23361 2620 -23327
rect 2574 -23399 2620 -23361
rect 2574 -23433 2580 -23399
rect 2614 -23433 2620 -23399
rect 2574 -23464 2620 -23433
rect 3592 -22929 3598 -22916
rect 3632 -22916 3648 -22895
rect 4606 -22895 4666 -22618
rect 5100 -22622 5160 -22310
rect 5620 -22462 5680 -22201
rect 6638 -22201 6652 -22178
rect 6686 -22178 6692 -22167
rect 7656 -22167 7716 -22156
rect 6686 -22201 6698 -22178
rect 5916 -22270 6404 -22264
rect 5916 -22304 5963 -22270
rect 5997 -22304 6035 -22270
rect 6069 -22304 6107 -22270
rect 6141 -22304 6179 -22270
rect 6213 -22304 6251 -22270
rect 6285 -22304 6323 -22270
rect 6357 -22304 6404 -22270
rect 5916 -22310 6404 -22304
rect 5614 -22466 5686 -22462
rect 5614 -22518 5624 -22466
rect 5676 -22518 5686 -22466
rect 5614 -22522 5686 -22518
rect 6134 -22622 6194 -22310
rect 6638 -22364 6698 -22201
rect 7656 -22201 7670 -22167
rect 7704 -22201 7716 -22167
rect 8682 -22167 8728 -22129
rect 8682 -22180 8688 -22167
rect 6934 -22270 7422 -22264
rect 6934 -22304 6981 -22270
rect 7015 -22304 7053 -22270
rect 7087 -22304 7125 -22270
rect 7159 -22304 7197 -22270
rect 7231 -22304 7269 -22270
rect 7303 -22304 7341 -22270
rect 7375 -22304 7422 -22270
rect 6934 -22310 7422 -22304
rect 6632 -22368 6704 -22364
rect 6632 -22420 6642 -22368
rect 6694 -22420 6704 -22368
rect 6632 -22424 6704 -22420
rect 7144 -22462 7204 -22310
rect 7138 -22466 7210 -22462
rect 7138 -22518 7148 -22466
rect 7200 -22518 7210 -22466
rect 7138 -22522 7210 -22518
rect 6636 -22562 6708 -22558
rect 6636 -22614 6646 -22562
rect 6698 -22614 6708 -22562
rect 6636 -22618 6708 -22614
rect 5100 -22682 6194 -22622
rect 5100 -22786 5160 -22682
rect 6134 -22786 6194 -22682
rect 4898 -22792 5386 -22786
rect 4898 -22826 4945 -22792
rect 4979 -22826 5017 -22792
rect 5051 -22826 5089 -22792
rect 5123 -22826 5161 -22792
rect 5195 -22826 5233 -22792
rect 5267 -22826 5305 -22792
rect 5339 -22826 5386 -22792
rect 4898 -22832 5386 -22826
rect 5916 -22792 6404 -22786
rect 5916 -22826 5963 -22792
rect 5997 -22826 6035 -22792
rect 6069 -22826 6107 -22792
rect 6141 -22826 6179 -22792
rect 6213 -22826 6251 -22792
rect 6285 -22826 6323 -22792
rect 6357 -22826 6404 -22792
rect 5916 -22832 6404 -22826
rect 3632 -22929 3638 -22916
rect 4606 -22920 4616 -22895
rect 3592 -22967 3638 -22929
rect 3592 -23001 3598 -22967
rect 3632 -23001 3638 -22967
rect 3592 -23039 3638 -23001
rect 3592 -23073 3598 -23039
rect 3632 -23073 3638 -23039
rect 3592 -23111 3638 -23073
rect 3592 -23145 3598 -23111
rect 3632 -23145 3638 -23111
rect 3592 -23183 3638 -23145
rect 3592 -23217 3598 -23183
rect 3632 -23217 3638 -23183
rect 3592 -23255 3638 -23217
rect 3592 -23289 3598 -23255
rect 3632 -23289 3638 -23255
rect 3592 -23327 3638 -23289
rect 3592 -23361 3598 -23327
rect 3632 -23361 3638 -23327
rect 3592 -23399 3638 -23361
rect 3592 -23433 3598 -23399
rect 3632 -23433 3638 -23399
rect 3592 -23464 3638 -23433
rect 4610 -22929 4616 -22920
rect 4650 -22920 4666 -22895
rect 5628 -22895 5674 -22864
rect 4650 -22929 4656 -22920
rect 4610 -22967 4656 -22929
rect 4610 -23001 4616 -22967
rect 4650 -23001 4656 -22967
rect 4610 -23039 4656 -23001
rect 4610 -23073 4616 -23039
rect 4650 -23073 4656 -23039
rect 4610 -23111 4656 -23073
rect 4610 -23145 4616 -23111
rect 4650 -23145 4656 -23111
rect 4610 -23183 4656 -23145
rect 4610 -23217 4616 -23183
rect 4650 -23217 4656 -23183
rect 4610 -23255 4656 -23217
rect 4610 -23289 4616 -23255
rect 4650 -23289 4656 -23255
rect 4610 -23327 4656 -23289
rect 4610 -23361 4616 -23327
rect 4650 -23361 4656 -23327
rect 4610 -23399 4656 -23361
rect 4610 -23433 4616 -23399
rect 4650 -23433 4656 -23399
rect 5628 -22929 5634 -22895
rect 5668 -22929 5674 -22895
rect 6642 -22895 6702 -22618
rect 7144 -22786 7204 -22522
rect 7656 -22678 7716 -22201
rect 8676 -22201 8688 -22180
rect 8722 -22180 8728 -22167
rect 9700 -21697 9706 -21680
rect 9740 -21680 9756 -21663
rect 10712 -21663 10772 -21402
rect 11006 -21560 11494 -21554
rect 11006 -21594 11053 -21560
rect 11087 -21594 11125 -21560
rect 11159 -21594 11197 -21560
rect 11231 -21594 11269 -21560
rect 11303 -21594 11341 -21560
rect 11375 -21594 11413 -21560
rect 11447 -21594 11494 -21560
rect 11006 -21600 11494 -21594
rect 10712 -21670 10724 -21663
rect 9740 -21697 9746 -21680
rect 9700 -21735 9746 -21697
rect 9700 -21769 9706 -21735
rect 9740 -21769 9746 -21735
rect 9700 -21807 9746 -21769
rect 9700 -21841 9706 -21807
rect 9740 -21841 9746 -21807
rect 9700 -21879 9746 -21841
rect 9700 -21913 9706 -21879
rect 9740 -21913 9746 -21879
rect 9700 -21951 9746 -21913
rect 9700 -21985 9706 -21951
rect 9740 -21985 9746 -21951
rect 9700 -22023 9746 -21985
rect 9700 -22057 9706 -22023
rect 9740 -22057 9746 -22023
rect 9700 -22095 9746 -22057
rect 9700 -22129 9706 -22095
rect 9740 -22129 9746 -22095
rect 9700 -22167 9746 -22129
rect 10718 -21697 10724 -21670
rect 10758 -21670 10772 -21663
rect 11730 -21663 11790 -21290
rect 12024 -21560 12512 -21554
rect 12024 -21594 12071 -21560
rect 12105 -21594 12143 -21560
rect 12177 -21594 12215 -21560
rect 12249 -21594 12287 -21560
rect 12321 -21594 12359 -21560
rect 12393 -21594 12431 -21560
rect 12465 -21594 12512 -21560
rect 12024 -21600 12512 -21594
rect 13042 -21560 13530 -21554
rect 13042 -21594 13089 -21560
rect 13123 -21594 13161 -21560
rect 13195 -21594 13233 -21560
rect 13267 -21594 13305 -21560
rect 13339 -21594 13377 -21560
rect 13411 -21594 13449 -21560
rect 13483 -21594 13530 -21560
rect 13042 -21600 13530 -21594
rect 10758 -21697 10764 -21670
rect 11730 -21676 11742 -21663
rect 10718 -21735 10764 -21697
rect 10718 -21769 10724 -21735
rect 10758 -21769 10764 -21735
rect 10718 -21807 10764 -21769
rect 10718 -21841 10724 -21807
rect 10758 -21841 10764 -21807
rect 10718 -21879 10764 -21841
rect 10718 -21913 10724 -21879
rect 10758 -21913 10764 -21879
rect 10718 -21951 10764 -21913
rect 10718 -21985 10724 -21951
rect 10758 -21985 10764 -21951
rect 10718 -22023 10764 -21985
rect 10718 -22057 10724 -22023
rect 10758 -22057 10764 -22023
rect 10718 -22095 10764 -22057
rect 10718 -22129 10724 -22095
rect 10758 -22129 10764 -22095
rect 10718 -22164 10764 -22129
rect 11736 -21697 11742 -21676
rect 11776 -21676 11790 -21663
rect 12754 -21663 12800 -21632
rect 11776 -21697 11782 -21676
rect 11736 -21735 11782 -21697
rect 11736 -21769 11742 -21735
rect 11776 -21769 11782 -21735
rect 11736 -21807 11782 -21769
rect 11736 -21841 11742 -21807
rect 11776 -21841 11782 -21807
rect 11736 -21879 11782 -21841
rect 11736 -21913 11742 -21879
rect 11776 -21913 11782 -21879
rect 11736 -21951 11782 -21913
rect 11736 -21985 11742 -21951
rect 11776 -21985 11782 -21951
rect 11736 -22023 11782 -21985
rect 11736 -22057 11742 -22023
rect 11776 -22057 11782 -22023
rect 11736 -22095 11782 -22057
rect 11736 -22129 11742 -22095
rect 11776 -22129 11782 -22095
rect 8722 -22201 8736 -22180
rect 9700 -22186 9706 -22167
rect 7952 -22270 8440 -22264
rect 7952 -22304 7999 -22270
rect 8033 -22304 8071 -22270
rect 8105 -22304 8143 -22270
rect 8177 -22304 8215 -22270
rect 8249 -22304 8287 -22270
rect 8321 -22304 8359 -22270
rect 8393 -22304 8440 -22270
rect 7952 -22310 8440 -22304
rect 8166 -22466 8226 -22310
rect 8676 -22364 8736 -22201
rect 9690 -22201 9706 -22186
rect 9740 -22186 9746 -22167
rect 10708 -22167 10768 -22164
rect 9740 -22201 9750 -22186
rect 8970 -22270 9458 -22264
rect 8970 -22304 9017 -22270
rect 9051 -22304 9089 -22270
rect 9123 -22304 9161 -22270
rect 9195 -22304 9233 -22270
rect 9267 -22304 9305 -22270
rect 9339 -22304 9377 -22270
rect 9411 -22304 9458 -22270
rect 8970 -22310 9458 -22304
rect 8670 -22368 8742 -22364
rect 8670 -22420 8680 -22368
rect 8732 -22420 8742 -22368
rect 8670 -22424 8742 -22420
rect 9190 -22456 9250 -22310
rect 8166 -22518 8170 -22466
rect 8222 -22518 8226 -22466
rect 7650 -22682 7722 -22678
rect 7650 -22734 7660 -22682
rect 7712 -22734 7722 -22682
rect 7650 -22738 7722 -22734
rect 6934 -22792 7422 -22786
rect 6934 -22826 6981 -22792
rect 7015 -22826 7053 -22792
rect 7087 -22826 7125 -22792
rect 7159 -22826 7197 -22792
rect 7231 -22826 7269 -22792
rect 7303 -22826 7341 -22792
rect 7375 -22826 7422 -22792
rect 6934 -22832 7422 -22826
rect 6642 -22928 6652 -22895
rect 5628 -22967 5674 -22929
rect 5628 -23001 5634 -22967
rect 5668 -23001 5674 -22967
rect 5628 -23039 5674 -23001
rect 5628 -23073 5634 -23039
rect 5668 -23073 5674 -23039
rect 5628 -23111 5674 -23073
rect 5628 -23145 5634 -23111
rect 5668 -23145 5674 -23111
rect 5628 -23183 5674 -23145
rect 5628 -23217 5634 -23183
rect 5668 -23217 5674 -23183
rect 5628 -23255 5674 -23217
rect 5628 -23289 5634 -23255
rect 5668 -23289 5674 -23255
rect 5628 -23327 5674 -23289
rect 5628 -23361 5634 -23327
rect 5668 -23361 5674 -23327
rect 5628 -23399 5674 -23361
rect 5628 -23410 5634 -23399
rect 4610 -23464 4656 -23433
rect 5620 -23433 5634 -23410
rect 5668 -23410 5674 -23399
rect 6646 -22929 6652 -22928
rect 6686 -22928 6702 -22895
rect 7656 -22895 7716 -22738
rect 8166 -22786 8226 -22518
rect 9188 -22466 9250 -22456
rect 9188 -22518 9192 -22466
rect 9244 -22518 9250 -22466
rect 9188 -22528 9250 -22518
rect 8664 -22562 8736 -22558
rect 8664 -22614 8674 -22562
rect 8726 -22614 8736 -22562
rect 8664 -22618 8736 -22614
rect 7952 -22792 8440 -22786
rect 7952 -22826 7999 -22792
rect 8033 -22826 8071 -22792
rect 8105 -22826 8143 -22792
rect 8177 -22826 8215 -22792
rect 8249 -22826 8287 -22792
rect 8321 -22826 8359 -22792
rect 8393 -22826 8440 -22792
rect 7952 -22832 8440 -22826
rect 7656 -22916 7670 -22895
rect 6686 -22929 6692 -22928
rect 6646 -22967 6692 -22929
rect 6646 -23001 6652 -22967
rect 6686 -23001 6692 -22967
rect 6646 -23039 6692 -23001
rect 6646 -23073 6652 -23039
rect 6686 -23073 6692 -23039
rect 6646 -23111 6692 -23073
rect 6646 -23145 6652 -23111
rect 6686 -23145 6692 -23111
rect 6646 -23183 6692 -23145
rect 6646 -23217 6652 -23183
rect 6686 -23217 6692 -23183
rect 6646 -23255 6692 -23217
rect 6646 -23289 6652 -23255
rect 6686 -23289 6692 -23255
rect 6646 -23327 6692 -23289
rect 6646 -23361 6652 -23327
rect 6686 -23361 6692 -23327
rect 6646 -23399 6692 -23361
rect 7664 -22929 7670 -22916
rect 7704 -22916 7716 -22895
rect 8670 -22895 8730 -22618
rect 9190 -22786 9250 -22528
rect 9690 -22678 9750 -22201
rect 10708 -22201 10724 -22167
rect 10758 -22201 10768 -22167
rect 9988 -22270 10476 -22264
rect 9988 -22304 10035 -22270
rect 10069 -22304 10107 -22270
rect 10141 -22304 10179 -22270
rect 10213 -22304 10251 -22270
rect 10285 -22304 10323 -22270
rect 10357 -22304 10395 -22270
rect 10429 -22304 10476 -22270
rect 9988 -22310 10252 -22304
rect 10264 -22310 10476 -22304
rect 10192 -22462 10252 -22310
rect 10538 -22348 10598 -22338
rect 10708 -22344 10768 -22201
rect 11736 -22167 11782 -22129
rect 12754 -21697 12760 -21663
rect 12794 -21697 12800 -21663
rect 13766 -21663 13826 -21290
rect 15308 -21328 15368 -21076
rect 15802 -21118 15862 -20967
rect 16826 -20967 16832 -20933
rect 16866 -20967 16872 -20933
rect 17844 -20535 17850 -20504
rect 17884 -20504 17896 -20501
rect 18862 -20501 18908 -20476
rect 17884 -20535 17890 -20504
rect 17844 -20573 17890 -20535
rect 17844 -20607 17850 -20573
rect 17884 -20607 17890 -20573
rect 17844 -20645 17890 -20607
rect 17844 -20679 17850 -20645
rect 17884 -20679 17890 -20645
rect 17844 -20717 17890 -20679
rect 17844 -20751 17850 -20717
rect 17884 -20751 17890 -20717
rect 17844 -20789 17890 -20751
rect 17844 -20823 17850 -20789
rect 17884 -20823 17890 -20789
rect 17844 -20861 17890 -20823
rect 17844 -20895 17850 -20861
rect 17884 -20895 17890 -20861
rect 17844 -20933 17890 -20895
rect 17844 -20944 17850 -20933
rect 16826 -20998 16872 -20967
rect 17836 -20967 17850 -20944
rect 17884 -20944 17890 -20933
rect 18862 -20535 18868 -20501
rect 18902 -20535 18908 -20501
rect 18862 -20573 18908 -20535
rect 18862 -20607 18868 -20573
rect 18902 -20607 18908 -20573
rect 18862 -20645 18908 -20607
rect 18862 -20679 18868 -20645
rect 18902 -20679 18908 -20645
rect 18862 -20717 18908 -20679
rect 18862 -20751 18868 -20717
rect 18902 -20751 18908 -20717
rect 18862 -20789 18908 -20751
rect 18862 -20823 18868 -20789
rect 18902 -20823 18908 -20789
rect 18862 -20861 18908 -20823
rect 18862 -20895 18868 -20861
rect 18902 -20895 18908 -20861
rect 18862 -20933 18908 -20895
rect 17884 -20967 17896 -20944
rect 16096 -21036 16584 -21030
rect 16096 -21070 16143 -21036
rect 16177 -21070 16215 -21036
rect 16249 -21070 16287 -21036
rect 16321 -21070 16359 -21036
rect 16393 -21070 16431 -21036
rect 16465 -21070 16503 -21036
rect 16537 -21070 16584 -21036
rect 16096 -21076 16584 -21070
rect 17114 -21036 17602 -21030
rect 17114 -21070 17161 -21036
rect 17195 -21070 17233 -21036
rect 17267 -21070 17305 -21036
rect 17339 -21070 17377 -21036
rect 17411 -21070 17449 -21036
rect 17483 -21070 17521 -21036
rect 17555 -21070 17602 -21036
rect 17114 -21076 17602 -21070
rect 15796 -21122 15868 -21118
rect 15796 -21174 15806 -21122
rect 15858 -21174 15868 -21122
rect 15796 -21178 15868 -21174
rect 16150 -21122 16222 -21118
rect 16150 -21174 16160 -21122
rect 16212 -21174 16222 -21122
rect 16150 -21178 16222 -21174
rect 15792 -21234 15864 -21230
rect 15792 -21286 15802 -21234
rect 15854 -21286 15864 -21234
rect 15792 -21290 15864 -21286
rect 15302 -21332 15374 -21328
rect 15302 -21384 15312 -21332
rect 15364 -21384 15374 -21332
rect 15302 -21388 15374 -21384
rect 14060 -21560 14548 -21554
rect 14060 -21594 14107 -21560
rect 14141 -21594 14179 -21560
rect 14213 -21594 14251 -21560
rect 14285 -21594 14323 -21560
rect 14357 -21594 14395 -21560
rect 14429 -21594 14467 -21560
rect 14501 -21594 14548 -21560
rect 14060 -21600 14548 -21594
rect 15078 -21560 15566 -21554
rect 15078 -21594 15125 -21560
rect 15159 -21594 15197 -21560
rect 15231 -21594 15269 -21560
rect 15303 -21594 15341 -21560
rect 15375 -21594 15413 -21560
rect 15447 -21594 15485 -21560
rect 15519 -21594 15566 -21560
rect 15078 -21600 15566 -21594
rect 13766 -21682 13778 -21663
rect 12754 -21735 12800 -21697
rect 12754 -21769 12760 -21735
rect 12794 -21769 12800 -21735
rect 12754 -21807 12800 -21769
rect 12754 -21841 12760 -21807
rect 12794 -21841 12800 -21807
rect 12754 -21879 12800 -21841
rect 12754 -21913 12760 -21879
rect 12794 -21913 12800 -21879
rect 12754 -21951 12800 -21913
rect 12754 -21985 12760 -21951
rect 12794 -21985 12800 -21951
rect 12754 -22023 12800 -21985
rect 12754 -22057 12760 -22023
rect 12794 -22057 12800 -22023
rect 12754 -22095 12800 -22057
rect 12754 -22129 12760 -22095
rect 12794 -22129 12800 -22095
rect 12754 -22150 12800 -22129
rect 13772 -21697 13778 -21682
rect 13812 -21682 13826 -21663
rect 14790 -21663 14836 -21632
rect 13812 -21697 13818 -21682
rect 13772 -21735 13818 -21697
rect 13772 -21769 13778 -21735
rect 13812 -21769 13818 -21735
rect 13772 -21807 13818 -21769
rect 13772 -21841 13778 -21807
rect 13812 -21841 13818 -21807
rect 13772 -21879 13818 -21841
rect 13772 -21913 13778 -21879
rect 13812 -21913 13818 -21879
rect 13772 -21951 13818 -21913
rect 13772 -21985 13778 -21951
rect 13812 -21985 13818 -21951
rect 13772 -22023 13818 -21985
rect 13772 -22057 13778 -22023
rect 13812 -22057 13818 -22023
rect 13772 -22095 13818 -22057
rect 13772 -22129 13778 -22095
rect 13812 -22129 13818 -22095
rect 11736 -22201 11742 -22167
rect 11776 -22201 11782 -22167
rect 11736 -22232 11782 -22201
rect 12750 -22167 12810 -22150
rect 12750 -22201 12760 -22167
rect 12794 -22201 12810 -22167
rect 11006 -22270 11494 -22264
rect 11006 -22304 11053 -22270
rect 11087 -22304 11125 -22270
rect 11159 -22304 11197 -22270
rect 11231 -22304 11269 -22270
rect 11303 -22304 11341 -22270
rect 11375 -22304 11413 -22270
rect 11447 -22304 11494 -22270
rect 11006 -22310 11494 -22304
rect 12024 -22270 12512 -22264
rect 12024 -22304 12071 -22270
rect 12105 -22304 12143 -22270
rect 12177 -22304 12215 -22270
rect 12249 -22304 12287 -22270
rect 12321 -22304 12359 -22270
rect 12393 -22304 12431 -22270
rect 12465 -22304 12512 -22270
rect 12024 -22310 12512 -22304
rect 10538 -22400 10542 -22348
rect 10594 -22400 10598 -22348
rect 10186 -22466 10258 -22462
rect 10186 -22518 10196 -22466
rect 10248 -22518 10258 -22466
rect 10186 -22522 10258 -22518
rect 9684 -22682 9756 -22678
rect 9684 -22734 9694 -22682
rect 9746 -22734 9756 -22682
rect 9684 -22738 9756 -22734
rect 8970 -22792 9458 -22786
rect 8970 -22826 9017 -22792
rect 9051 -22826 9089 -22792
rect 9123 -22826 9161 -22792
rect 9195 -22826 9233 -22792
rect 9267 -22826 9305 -22792
rect 9339 -22826 9377 -22792
rect 9411 -22826 9458 -22792
rect 8970 -22832 9458 -22826
rect 7704 -22929 7710 -22916
rect 7664 -22967 7710 -22929
rect 8670 -22929 8688 -22895
rect 8722 -22929 8730 -22895
rect 9690 -22895 9750 -22738
rect 10192 -22786 10252 -22522
rect 10538 -22558 10598 -22400
rect 10702 -22348 10774 -22344
rect 10702 -22400 10712 -22348
rect 10764 -22400 10774 -22348
rect 10702 -22404 10774 -22400
rect 10708 -22556 10780 -22552
rect 10532 -22562 10604 -22558
rect 10532 -22614 10542 -22562
rect 10594 -22614 10604 -22562
rect 10708 -22608 10718 -22556
rect 10770 -22608 10780 -22556
rect 10708 -22612 10780 -22608
rect 10532 -22618 10604 -22614
rect 9988 -22792 10252 -22786
rect 10264 -22792 10476 -22786
rect 9988 -22826 10035 -22792
rect 10069 -22826 10107 -22792
rect 10141 -22826 10179 -22792
rect 10213 -22826 10251 -22792
rect 10285 -22826 10323 -22792
rect 10357 -22826 10395 -22792
rect 10429 -22826 10476 -22792
rect 9988 -22832 10476 -22826
rect 9690 -22916 9706 -22895
rect 8670 -22936 8730 -22929
rect 9700 -22929 9706 -22916
rect 9740 -22916 9750 -22895
rect 10714 -22895 10774 -22612
rect 11230 -22614 11290 -22310
rect 12244 -22450 12304 -22310
rect 12750 -22344 12810 -22201
rect 13772 -22167 13818 -22129
rect 14790 -21697 14796 -21663
rect 14830 -21697 14836 -21663
rect 15798 -21663 15858 -21290
rect 16156 -21440 16216 -21178
rect 16346 -21328 16406 -21076
rect 17322 -21328 17382 -21076
rect 16340 -21332 16412 -21328
rect 16340 -21384 16350 -21332
rect 16402 -21384 16412 -21332
rect 16340 -21388 16412 -21384
rect 17316 -21332 17388 -21328
rect 17316 -21384 17326 -21332
rect 17378 -21384 17388 -21332
rect 17316 -21388 17388 -21384
rect 17836 -21440 17896 -20967
rect 18862 -20967 18868 -20933
rect 18902 -20967 18908 -20933
rect 19880 -20501 19926 -20463
rect 19880 -20535 19886 -20501
rect 19920 -20535 19926 -20501
rect 19880 -20573 19926 -20535
rect 19880 -20607 19886 -20573
rect 19920 -20607 19926 -20573
rect 19880 -20645 19926 -20607
rect 19880 -20679 19886 -20645
rect 19920 -20679 19926 -20645
rect 19880 -20717 19926 -20679
rect 19880 -20751 19886 -20717
rect 19920 -20751 19926 -20717
rect 19880 -20789 19926 -20751
rect 19880 -20823 19886 -20789
rect 19920 -20823 19926 -20789
rect 19880 -20861 19926 -20823
rect 19880 -20895 19886 -20861
rect 19920 -20895 19926 -20861
rect 19880 -20933 19926 -20895
rect 19880 -20942 19886 -20933
rect 18862 -20998 18908 -20967
rect 19874 -20967 19886 -20942
rect 19920 -20942 19926 -20933
rect 20898 -20463 20904 -20462
rect 20938 -20462 20950 -20429
rect 21912 -20429 21972 -20276
rect 22204 -20326 22692 -20320
rect 22204 -20360 22251 -20326
rect 22285 -20360 22323 -20326
rect 22357 -20360 22395 -20326
rect 22429 -20360 22467 -20326
rect 22501 -20360 22539 -20326
rect 22573 -20360 22611 -20326
rect 22645 -20360 22692 -20326
rect 22204 -20366 22692 -20360
rect 21912 -20444 21922 -20429
rect 20938 -20463 20944 -20462
rect 20898 -20501 20944 -20463
rect 20898 -20535 20904 -20501
rect 20938 -20535 20944 -20501
rect 20898 -20573 20944 -20535
rect 20898 -20607 20904 -20573
rect 20938 -20607 20944 -20573
rect 20898 -20645 20944 -20607
rect 20898 -20679 20904 -20645
rect 20938 -20679 20944 -20645
rect 20898 -20717 20944 -20679
rect 20898 -20751 20904 -20717
rect 20938 -20751 20944 -20717
rect 20898 -20789 20944 -20751
rect 20898 -20823 20904 -20789
rect 20938 -20823 20944 -20789
rect 20898 -20861 20944 -20823
rect 20898 -20895 20904 -20861
rect 20938 -20895 20944 -20861
rect 20898 -20933 20944 -20895
rect 20898 -20936 20904 -20933
rect 19920 -20967 19934 -20942
rect 18132 -21036 18620 -21030
rect 18132 -21070 18179 -21036
rect 18213 -21070 18251 -21036
rect 18285 -21070 18323 -21036
rect 18357 -21070 18395 -21036
rect 18429 -21070 18467 -21036
rect 18501 -21070 18539 -21036
rect 18573 -21070 18620 -21036
rect 18132 -21076 18620 -21070
rect 19150 -21036 19638 -21030
rect 19150 -21070 19197 -21036
rect 19231 -21070 19269 -21036
rect 19303 -21070 19341 -21036
rect 19375 -21070 19413 -21036
rect 19447 -21070 19485 -21036
rect 19519 -21070 19557 -21036
rect 19591 -21070 19638 -21036
rect 19150 -21076 19638 -21070
rect 18338 -21328 18398 -21076
rect 19874 -21118 19934 -20967
rect 20892 -20967 20904 -20936
rect 20938 -20936 20944 -20933
rect 21916 -20463 21922 -20444
rect 21956 -20444 21972 -20429
rect 22934 -20429 22980 -20398
rect 21956 -20463 21962 -20444
rect 21916 -20501 21962 -20463
rect 21916 -20535 21922 -20501
rect 21956 -20535 21962 -20501
rect 21916 -20573 21962 -20535
rect 21916 -20607 21922 -20573
rect 21956 -20607 21962 -20573
rect 21916 -20645 21962 -20607
rect 21916 -20679 21922 -20645
rect 21956 -20679 21962 -20645
rect 21916 -20717 21962 -20679
rect 21916 -20751 21922 -20717
rect 21956 -20751 21962 -20717
rect 21916 -20789 21962 -20751
rect 21916 -20823 21922 -20789
rect 21956 -20823 21962 -20789
rect 21916 -20861 21962 -20823
rect 21916 -20895 21922 -20861
rect 21956 -20895 21962 -20861
rect 21916 -20933 21962 -20895
rect 20938 -20967 20952 -20936
rect 21916 -20942 21922 -20933
rect 20168 -21036 20656 -21030
rect 20168 -21070 20215 -21036
rect 20249 -21070 20287 -21036
rect 20321 -21070 20359 -21036
rect 20393 -21070 20431 -21036
rect 20465 -21070 20503 -21036
rect 20537 -21070 20575 -21036
rect 20609 -21070 20656 -21036
rect 20168 -21076 20656 -21070
rect 19868 -21122 19940 -21118
rect 19868 -21174 19878 -21122
rect 19930 -21174 19940 -21122
rect 19868 -21178 19940 -21174
rect 18332 -21332 18404 -21328
rect 18332 -21384 18342 -21332
rect 18394 -21384 18404 -21332
rect 18332 -21388 18404 -21384
rect 20358 -21332 20430 -21328
rect 20358 -21384 20368 -21332
rect 20420 -21384 20430 -21332
rect 20358 -21388 20430 -21384
rect 16156 -21492 16160 -21440
rect 16212 -21492 16216 -21440
rect 16156 -21502 16216 -21492
rect 17830 -21444 17902 -21440
rect 17830 -21496 17840 -21444
rect 17892 -21496 17902 -21444
rect 17830 -21500 17902 -21496
rect 19866 -21444 19938 -21440
rect 19866 -21496 19876 -21444
rect 19928 -21496 19938 -21444
rect 19866 -21500 19938 -21496
rect 16096 -21560 16584 -21554
rect 16096 -21594 16143 -21560
rect 16177 -21594 16215 -21560
rect 16249 -21594 16287 -21560
rect 16321 -21594 16359 -21560
rect 16393 -21594 16431 -21560
rect 16465 -21594 16503 -21560
rect 16537 -21594 16584 -21560
rect 16096 -21600 16584 -21594
rect 17114 -21560 17602 -21554
rect 17114 -21594 17161 -21560
rect 17195 -21594 17233 -21560
rect 17267 -21594 17305 -21560
rect 17339 -21594 17377 -21560
rect 17411 -21594 17449 -21560
rect 17483 -21594 17521 -21560
rect 17555 -21594 17602 -21560
rect 17114 -21600 17602 -21594
rect 15798 -21686 15814 -21663
rect 14790 -21735 14836 -21697
rect 14790 -21769 14796 -21735
rect 14830 -21769 14836 -21735
rect 14790 -21807 14836 -21769
rect 14790 -21841 14796 -21807
rect 14830 -21841 14836 -21807
rect 14790 -21879 14836 -21841
rect 14790 -21913 14796 -21879
rect 14830 -21913 14836 -21879
rect 14790 -21951 14836 -21913
rect 14790 -21985 14796 -21951
rect 14830 -21985 14836 -21951
rect 14790 -22023 14836 -21985
rect 14790 -22057 14796 -22023
rect 14830 -22057 14836 -22023
rect 14790 -22095 14836 -22057
rect 14790 -22129 14796 -22095
rect 14830 -22129 14836 -22095
rect 14790 -22150 14836 -22129
rect 15808 -21697 15814 -21686
rect 15848 -21686 15858 -21663
rect 16826 -21663 16872 -21632
rect 15848 -21697 15854 -21686
rect 15808 -21735 15854 -21697
rect 15808 -21769 15814 -21735
rect 15848 -21769 15854 -21735
rect 15808 -21807 15854 -21769
rect 15808 -21841 15814 -21807
rect 15848 -21841 15854 -21807
rect 15808 -21879 15854 -21841
rect 15808 -21913 15814 -21879
rect 15848 -21913 15854 -21879
rect 15808 -21951 15854 -21913
rect 15808 -21985 15814 -21951
rect 15848 -21985 15854 -21951
rect 15808 -22023 15854 -21985
rect 15808 -22057 15814 -22023
rect 15848 -22057 15854 -22023
rect 15808 -22095 15854 -22057
rect 15808 -22129 15814 -22095
rect 15848 -22129 15854 -22095
rect 13772 -22201 13778 -22167
rect 13812 -22201 13818 -22167
rect 13772 -22232 13818 -22201
rect 14782 -22167 14842 -22150
rect 14782 -22201 14796 -22167
rect 14830 -22201 14842 -22167
rect 13042 -22270 13530 -22264
rect 13042 -22304 13089 -22270
rect 13123 -22304 13161 -22270
rect 13195 -22304 13233 -22270
rect 13267 -22304 13305 -22270
rect 13339 -22304 13377 -22270
rect 13411 -22304 13449 -22270
rect 13483 -22304 13530 -22270
rect 13042 -22310 13530 -22304
rect 14060 -22270 14548 -22264
rect 14060 -22304 14107 -22270
rect 14141 -22304 14179 -22270
rect 14213 -22304 14251 -22270
rect 14285 -22304 14323 -22270
rect 14357 -22304 14395 -22270
rect 14429 -22304 14467 -22270
rect 14501 -22304 14548 -22270
rect 14060 -22310 14548 -22304
rect 12744 -22348 12816 -22344
rect 12744 -22400 12754 -22348
rect 12806 -22400 12816 -22348
rect 12744 -22404 12816 -22400
rect 13266 -22450 13326 -22310
rect 14280 -22450 14340 -22310
rect 14782 -22344 14842 -22201
rect 15808 -22167 15854 -22129
rect 15808 -22201 15814 -22167
rect 15848 -22201 15854 -22167
rect 16826 -21697 16832 -21663
rect 16866 -21697 16872 -21663
rect 17836 -21663 17896 -21500
rect 18132 -21560 18620 -21554
rect 18132 -21594 18179 -21560
rect 18213 -21594 18251 -21560
rect 18285 -21594 18323 -21560
rect 18357 -21594 18395 -21560
rect 18429 -21594 18467 -21560
rect 18501 -21594 18539 -21560
rect 18573 -21594 18620 -21560
rect 18132 -21600 18620 -21594
rect 19150 -21560 19638 -21554
rect 19150 -21594 19197 -21560
rect 19231 -21594 19269 -21560
rect 19303 -21594 19341 -21560
rect 19375 -21594 19413 -21560
rect 19447 -21594 19485 -21560
rect 19519 -21594 19557 -21560
rect 19591 -21594 19638 -21560
rect 19150 -21600 19638 -21594
rect 17836 -21682 17850 -21663
rect 16826 -21735 16872 -21697
rect 16826 -21769 16832 -21735
rect 16866 -21769 16872 -21735
rect 16826 -21807 16872 -21769
rect 16826 -21841 16832 -21807
rect 16866 -21841 16872 -21807
rect 16826 -21879 16872 -21841
rect 16826 -21913 16832 -21879
rect 16866 -21913 16872 -21879
rect 16826 -21951 16872 -21913
rect 16826 -21985 16832 -21951
rect 16866 -21985 16872 -21951
rect 16826 -22023 16872 -21985
rect 16826 -22057 16832 -22023
rect 16866 -22057 16872 -22023
rect 16826 -22095 16872 -22057
rect 16826 -22129 16832 -22095
rect 16866 -22129 16872 -22095
rect 16826 -22167 16872 -22129
rect 16826 -22184 16832 -22167
rect 15808 -22232 15854 -22201
rect 16822 -22201 16832 -22184
rect 16866 -22184 16872 -22167
rect 17844 -21697 17850 -21682
rect 17884 -21682 17896 -21663
rect 18862 -21663 18908 -21632
rect 17884 -21697 17890 -21682
rect 17844 -21735 17890 -21697
rect 17844 -21769 17850 -21735
rect 17884 -21769 17890 -21735
rect 17844 -21807 17890 -21769
rect 17844 -21841 17850 -21807
rect 17884 -21841 17890 -21807
rect 17844 -21879 17890 -21841
rect 17844 -21913 17850 -21879
rect 17884 -21913 17890 -21879
rect 17844 -21951 17890 -21913
rect 17844 -21985 17850 -21951
rect 17884 -21985 17890 -21951
rect 17844 -22023 17890 -21985
rect 17844 -22057 17850 -22023
rect 17884 -22057 17890 -22023
rect 17844 -22095 17890 -22057
rect 17844 -22129 17850 -22095
rect 17884 -22129 17890 -22095
rect 17844 -22167 17890 -22129
rect 17844 -22168 17850 -22167
rect 16866 -22201 16882 -22184
rect 15078 -22270 15566 -22264
rect 15078 -22304 15125 -22270
rect 15159 -22304 15197 -22270
rect 15231 -22304 15269 -22270
rect 15303 -22304 15341 -22270
rect 15375 -22304 15413 -22270
rect 15447 -22304 15485 -22270
rect 15519 -22304 15566 -22270
rect 15078 -22310 15566 -22304
rect 16096 -22270 16584 -22264
rect 16096 -22304 16143 -22270
rect 16177 -22304 16215 -22270
rect 16249 -22304 16287 -22270
rect 16321 -22304 16359 -22270
rect 16393 -22304 16431 -22270
rect 16465 -22304 16503 -22270
rect 16537 -22304 16584 -22270
rect 16096 -22310 16584 -22304
rect 14776 -22348 14848 -22344
rect 14776 -22400 14786 -22348
rect 14838 -22400 14848 -22348
rect 14776 -22404 14848 -22400
rect 15282 -22350 15342 -22310
rect 16308 -22350 16368 -22310
rect 16822 -22344 16882 -22201
rect 17840 -22201 17850 -22168
rect 17884 -22168 17890 -22167
rect 18862 -21697 18868 -21663
rect 18902 -21697 18908 -21663
rect 18862 -21735 18908 -21697
rect 19872 -21663 19932 -21500
rect 20364 -21554 20424 -21388
rect 20168 -21560 20656 -21554
rect 20168 -21594 20215 -21560
rect 20249 -21594 20287 -21560
rect 20321 -21594 20359 -21560
rect 20393 -21594 20431 -21560
rect 20465 -21594 20503 -21560
rect 20537 -21594 20575 -21560
rect 20609 -21594 20656 -21560
rect 20168 -21600 20656 -21594
rect 19872 -21697 19886 -21663
rect 19920 -21697 19932 -21663
rect 20892 -21663 20952 -20967
rect 21908 -20967 21922 -20942
rect 21956 -20942 21962 -20933
rect 22934 -20463 22940 -20429
rect 22974 -20463 22980 -20429
rect 22934 -20501 22980 -20463
rect 22934 -20535 22940 -20501
rect 22974 -20535 22980 -20501
rect 22934 -20573 22980 -20535
rect 22934 -20607 22940 -20573
rect 22974 -20607 22980 -20573
rect 22934 -20645 22980 -20607
rect 22934 -20679 22940 -20645
rect 22974 -20679 22980 -20645
rect 22934 -20717 22980 -20679
rect 22934 -20751 22940 -20717
rect 22974 -20751 22980 -20717
rect 22934 -20789 22980 -20751
rect 22934 -20823 22940 -20789
rect 22974 -20823 22980 -20789
rect 22934 -20861 22980 -20823
rect 22934 -20895 22940 -20861
rect 22974 -20895 22980 -20861
rect 22934 -20933 22980 -20895
rect 21956 -20967 21968 -20942
rect 22934 -20956 22940 -20933
rect 21186 -21036 21674 -21030
rect 21186 -21070 21233 -21036
rect 21267 -21070 21305 -21036
rect 21339 -21070 21377 -21036
rect 21411 -21070 21449 -21036
rect 21483 -21070 21521 -21036
rect 21555 -21070 21593 -21036
rect 21627 -21070 21674 -21036
rect 21186 -21076 21674 -21070
rect 21394 -21328 21454 -21076
rect 21908 -21168 21968 -20967
rect 22924 -20967 22940 -20956
rect 22974 -20956 22980 -20933
rect 22974 -20967 22984 -20956
rect 22204 -21036 22692 -21030
rect 22204 -21070 22251 -21036
rect 22285 -21070 22323 -21036
rect 22357 -21070 22395 -21036
rect 22429 -21070 22467 -21036
rect 22501 -21070 22539 -21036
rect 22573 -21070 22611 -21036
rect 22645 -21070 22692 -21036
rect 22204 -21076 22692 -21070
rect 22414 -21168 22474 -21076
rect 22924 -21168 22984 -20967
rect 21908 -21228 22984 -21168
rect 21388 -21332 21460 -21328
rect 21388 -21384 21398 -21332
rect 21450 -21384 21460 -21332
rect 21388 -21388 21460 -21384
rect 21908 -21440 21968 -21228
rect 21902 -21444 21974 -21440
rect 21902 -21496 21912 -21444
rect 21964 -21496 21974 -21444
rect 21902 -21500 21974 -21496
rect 21186 -21560 21674 -21554
rect 21186 -21594 21233 -21560
rect 21267 -21594 21305 -21560
rect 21339 -21594 21377 -21560
rect 21411 -21594 21449 -21560
rect 21483 -21594 21521 -21560
rect 21555 -21594 21593 -21560
rect 21627 -21594 21674 -21560
rect 21186 -21600 21674 -21594
rect 22204 -21560 22692 -21554
rect 22204 -21594 22251 -21560
rect 22285 -21594 22323 -21560
rect 22357 -21594 22395 -21560
rect 22429 -21594 22467 -21560
rect 22501 -21594 22539 -21560
rect 22573 -21594 22611 -21560
rect 22645 -21594 22692 -21560
rect 22204 -21600 22692 -21594
rect 20892 -21686 20904 -21663
rect 19872 -21702 19932 -21697
rect 20898 -21697 20904 -21686
rect 20938 -21686 20952 -21663
rect 21916 -21663 21962 -21632
rect 20938 -21697 20944 -21686
rect 18862 -21769 18868 -21735
rect 18902 -21769 18908 -21735
rect 18862 -21807 18908 -21769
rect 18862 -21841 18868 -21807
rect 18902 -21841 18908 -21807
rect 18862 -21879 18908 -21841
rect 18862 -21913 18868 -21879
rect 18902 -21913 18908 -21879
rect 18862 -21951 18908 -21913
rect 18862 -21985 18868 -21951
rect 18902 -21985 18908 -21951
rect 18862 -22023 18908 -21985
rect 18862 -22057 18868 -22023
rect 18902 -22057 18908 -22023
rect 18862 -22095 18908 -22057
rect 18862 -22129 18868 -22095
rect 18902 -22129 18908 -22095
rect 18862 -22167 18908 -22129
rect 17884 -22201 17900 -22168
rect 18862 -22176 18868 -22167
rect 17114 -22270 17602 -22264
rect 17114 -22304 17161 -22270
rect 17195 -22304 17233 -22270
rect 17267 -22304 17305 -22270
rect 17339 -22304 17377 -22270
rect 17411 -22304 17449 -22270
rect 17483 -22304 17521 -22270
rect 17555 -22304 17602 -22270
rect 17114 -22310 17602 -22304
rect 15282 -22410 16368 -22350
rect 16816 -22348 16888 -22344
rect 16816 -22400 16826 -22348
rect 16878 -22400 16888 -22348
rect 16816 -22404 16888 -22400
rect 15282 -22450 15342 -22410
rect 12244 -22510 15342 -22450
rect 15794 -22446 15866 -22442
rect 15794 -22498 15804 -22446
rect 15856 -22498 15866 -22446
rect 15794 -22502 15866 -22498
rect 12244 -22614 12304 -22510
rect 12736 -22556 12808 -22552
rect 12736 -22608 12746 -22556
rect 12798 -22608 12808 -22556
rect 12736 -22612 12808 -22608
rect 11230 -22674 12304 -22614
rect 11230 -22786 11290 -22674
rect 12244 -22786 12304 -22674
rect 11006 -22792 11494 -22786
rect 11006 -22826 11053 -22792
rect 11087 -22826 11125 -22792
rect 11159 -22826 11197 -22792
rect 11231 -22826 11269 -22792
rect 11303 -22826 11341 -22792
rect 11375 -22826 11413 -22792
rect 11447 -22826 11494 -22792
rect 11006 -22832 11494 -22826
rect 12024 -22792 12512 -22786
rect 12024 -22826 12071 -22792
rect 12105 -22826 12143 -22792
rect 12177 -22826 12215 -22792
rect 12249 -22826 12287 -22792
rect 12321 -22826 12359 -22792
rect 12393 -22826 12431 -22792
rect 12465 -22826 12512 -22792
rect 12024 -22832 12512 -22826
rect 9740 -22929 9746 -22916
rect 10714 -22920 10724 -22895
rect 7664 -23001 7670 -22967
rect 7704 -23001 7710 -22967
rect 7664 -23039 7710 -23001
rect 7664 -23073 7670 -23039
rect 7704 -23073 7710 -23039
rect 7664 -23111 7710 -23073
rect 7664 -23145 7670 -23111
rect 7704 -23145 7710 -23111
rect 7664 -23183 7710 -23145
rect 7664 -23217 7670 -23183
rect 7704 -23217 7710 -23183
rect 7664 -23255 7710 -23217
rect 7664 -23289 7670 -23255
rect 7704 -23289 7710 -23255
rect 7664 -23327 7710 -23289
rect 7664 -23361 7670 -23327
rect 7704 -23361 7710 -23327
rect 7664 -23398 7710 -23361
rect 8682 -22967 8728 -22936
rect 8682 -23001 8688 -22967
rect 8722 -23001 8728 -22967
rect 8682 -23039 8728 -23001
rect 8682 -23073 8688 -23039
rect 8722 -23073 8728 -23039
rect 8682 -23111 8728 -23073
rect 8682 -23145 8688 -23111
rect 8722 -23145 8728 -23111
rect 8682 -23183 8728 -23145
rect 8682 -23217 8688 -23183
rect 8722 -23217 8728 -23183
rect 8682 -23255 8728 -23217
rect 8682 -23289 8688 -23255
rect 8722 -23289 8728 -23255
rect 8682 -23327 8728 -23289
rect 8682 -23361 8688 -23327
rect 8722 -23361 8728 -23327
rect 5668 -23433 5680 -23410
rect 2862 -23502 3350 -23496
rect 2862 -23536 2909 -23502
rect 2943 -23536 2981 -23502
rect 3015 -23536 3053 -23502
rect 3087 -23536 3125 -23502
rect 3159 -23536 3197 -23502
rect 3231 -23536 3269 -23502
rect 3303 -23536 3350 -23502
rect 2862 -23542 3350 -23536
rect 3880 -23502 4368 -23496
rect 3880 -23536 3927 -23502
rect 3961 -23536 3999 -23502
rect 4033 -23536 4071 -23502
rect 4105 -23536 4143 -23502
rect 4177 -23536 4215 -23502
rect 4249 -23536 4287 -23502
rect 4321 -23536 4368 -23502
rect 3880 -23542 4368 -23536
rect 4898 -23502 5386 -23496
rect 4898 -23536 4945 -23502
rect 4979 -23536 5017 -23502
rect 5051 -23536 5089 -23502
rect 5123 -23536 5161 -23502
rect 5195 -23536 5233 -23502
rect 5267 -23536 5305 -23502
rect 5339 -23536 5386 -23502
rect 4898 -23542 5386 -23536
rect 2330 -23598 2402 -23594
rect 2330 -23650 2340 -23598
rect 2392 -23650 2402 -23598
rect 2330 -23654 2402 -23650
rect 2224 -23724 2296 -23720
rect 2224 -23776 2234 -23724
rect 2286 -23776 2296 -23724
rect 2224 -23780 2296 -23776
rect 2564 -23960 3644 -23900
rect 2564 -24129 2624 -23960
rect 3072 -24020 3132 -23960
rect 2862 -24026 3350 -24020
rect 2862 -24060 2909 -24026
rect 2943 -24060 2981 -24026
rect 3015 -24060 3053 -24026
rect 3087 -24060 3125 -24026
rect 3159 -24060 3197 -24026
rect 3231 -24060 3269 -24026
rect 3303 -24060 3350 -24026
rect 2862 -24066 3350 -24060
rect 2564 -24163 2580 -24129
rect 2614 -24163 2624 -24129
rect 2564 -24166 2624 -24163
rect 3584 -24129 3644 -23960
rect 4082 -24020 4142 -23542
rect 5620 -23720 5680 -23433
rect 6646 -23433 6652 -23399
rect 6686 -23433 6692 -23399
rect 6646 -23464 6692 -23433
rect 7658 -23399 7718 -23398
rect 7658 -23433 7670 -23399
rect 7704 -23433 7718 -23399
rect 5916 -23502 6404 -23496
rect 5916 -23536 5963 -23502
rect 5997 -23536 6035 -23502
rect 6069 -23536 6107 -23502
rect 6141 -23536 6179 -23502
rect 6213 -23536 6251 -23502
rect 6285 -23536 6323 -23502
rect 6357 -23536 6404 -23502
rect 5916 -23542 6256 -23536
rect 6316 -23542 6404 -23536
rect 6934 -23502 7422 -23496
rect 6934 -23536 6981 -23502
rect 7015 -23536 7053 -23502
rect 7087 -23536 7125 -23502
rect 7159 -23536 7197 -23502
rect 7231 -23536 7269 -23502
rect 7303 -23536 7341 -23502
rect 7375 -23536 7422 -23502
rect 6934 -23542 7422 -23536
rect 6140 -23708 6200 -23542
rect 6134 -23712 6206 -23708
rect 5614 -23724 5686 -23720
rect 5614 -23776 5624 -23724
rect 5676 -23776 5686 -23724
rect 6134 -23764 6144 -23712
rect 6196 -23764 6206 -23712
rect 6134 -23768 6206 -23764
rect 5614 -23780 5686 -23776
rect 4596 -23826 4668 -23822
rect 4596 -23878 4606 -23826
rect 4658 -23878 4668 -23826
rect 4596 -23882 4668 -23878
rect 6632 -23826 6704 -23822
rect 6632 -23878 6642 -23826
rect 6694 -23878 6704 -23826
rect 6632 -23882 6704 -23878
rect 3880 -24026 4368 -24020
rect 3880 -24060 3927 -24026
rect 3961 -24060 3999 -24026
rect 4033 -24060 4071 -24026
rect 4105 -24060 4143 -24026
rect 4177 -24060 4215 -24026
rect 4249 -24060 4287 -24026
rect 4321 -24060 4368 -24026
rect 3880 -24066 4368 -24060
rect 3584 -24163 3598 -24129
rect 3632 -24163 3644 -24129
rect 2574 -24201 2620 -24166
rect 2574 -24235 2580 -24201
rect 2614 -24235 2620 -24201
rect 2574 -24273 2620 -24235
rect 2574 -24307 2580 -24273
rect 2614 -24307 2620 -24273
rect 2574 -24345 2620 -24307
rect 2574 -24379 2580 -24345
rect 2614 -24379 2620 -24345
rect 2574 -24417 2620 -24379
rect 2574 -24451 2580 -24417
rect 2614 -24451 2620 -24417
rect 2574 -24489 2620 -24451
rect 2574 -24523 2580 -24489
rect 2614 -24523 2620 -24489
rect 2574 -24561 2620 -24523
rect 2574 -24592 2580 -24561
rect 2614 -24592 2620 -24561
rect 3584 -24201 3644 -24163
rect 4602 -24129 4662 -23882
rect 5614 -23930 5686 -23926
rect 5614 -23982 5624 -23930
rect 5676 -23982 5686 -23930
rect 5614 -23986 5686 -23982
rect 4898 -24026 5386 -24020
rect 4898 -24060 4945 -24026
rect 4979 -24060 5017 -24026
rect 5051 -24060 5089 -24026
rect 5123 -24060 5161 -24026
rect 5195 -24060 5233 -24026
rect 5267 -24060 5305 -24026
rect 5339 -24060 5386 -24026
rect 4898 -24066 5386 -24060
rect 4602 -24163 4616 -24129
rect 4650 -24163 4662 -24129
rect 4602 -24170 4662 -24163
rect 5620 -24129 5680 -23986
rect 5916 -24026 6140 -24020
rect 6200 -24026 6256 -24020
rect 6316 -24026 6404 -24020
rect 5916 -24060 5963 -24026
rect 5997 -24060 6035 -24026
rect 6069 -24060 6107 -24026
rect 6141 -24060 6179 -24026
rect 6213 -24060 6251 -24026
rect 6285 -24060 6323 -24026
rect 6357 -24060 6404 -24026
rect 5916 -24066 6404 -24060
rect 5620 -24163 5634 -24129
rect 5668 -24163 5680 -24129
rect 6638 -24129 6698 -23882
rect 7140 -24020 7200 -23542
rect 7658 -23822 7718 -23433
rect 8682 -23399 8728 -23361
rect 9700 -22967 9746 -22929
rect 9700 -23001 9706 -22967
rect 9740 -23001 9746 -22967
rect 9700 -23039 9746 -23001
rect 9700 -23073 9706 -23039
rect 9740 -23073 9746 -23039
rect 9700 -23111 9746 -23073
rect 9700 -23145 9706 -23111
rect 9740 -23145 9746 -23111
rect 9700 -23183 9746 -23145
rect 9700 -23217 9706 -23183
rect 9740 -23217 9746 -23183
rect 9700 -23255 9746 -23217
rect 9700 -23289 9706 -23255
rect 9740 -23289 9746 -23255
rect 9700 -23327 9746 -23289
rect 9700 -23361 9706 -23327
rect 9740 -23361 9746 -23327
rect 9700 -23386 9746 -23361
rect 10718 -22929 10724 -22920
rect 10758 -22920 10774 -22895
rect 11736 -22895 11782 -22864
rect 10758 -22929 10764 -22920
rect 10718 -22967 10764 -22929
rect 10718 -23001 10724 -22967
rect 10758 -23001 10764 -22967
rect 10718 -23039 10764 -23001
rect 10718 -23073 10724 -23039
rect 10758 -23073 10764 -23039
rect 10718 -23111 10764 -23073
rect 10718 -23145 10724 -23111
rect 10758 -23145 10764 -23111
rect 10718 -23183 10764 -23145
rect 10718 -23217 10724 -23183
rect 10758 -23217 10764 -23183
rect 10718 -23255 10764 -23217
rect 10718 -23289 10724 -23255
rect 10758 -23289 10764 -23255
rect 10718 -23327 10764 -23289
rect 10718 -23361 10724 -23327
rect 10758 -23361 10764 -23327
rect 8682 -23433 8688 -23399
rect 8722 -23433 8728 -23399
rect 8682 -23464 8728 -23433
rect 9694 -23399 9754 -23386
rect 10718 -23394 10764 -23361
rect 11736 -22929 11742 -22895
rect 11776 -22929 11782 -22895
rect 12742 -22895 12802 -22612
rect 13266 -22786 13326 -22510
rect 14280 -22786 14340 -22510
rect 14780 -22556 14852 -22552
rect 14780 -22608 14790 -22556
rect 14842 -22608 14852 -22556
rect 14780 -22612 14852 -22608
rect 13042 -22792 13530 -22786
rect 13042 -22826 13089 -22792
rect 13123 -22826 13161 -22792
rect 13195 -22826 13233 -22792
rect 13267 -22826 13305 -22792
rect 13339 -22826 13377 -22792
rect 13411 -22826 13449 -22792
rect 13483 -22826 13530 -22792
rect 13042 -22832 13530 -22826
rect 14060 -22792 14548 -22786
rect 14060 -22826 14107 -22792
rect 14141 -22826 14179 -22792
rect 14213 -22826 14251 -22792
rect 14285 -22826 14323 -22792
rect 14357 -22826 14395 -22792
rect 14429 -22826 14467 -22792
rect 14501 -22826 14548 -22792
rect 14060 -22832 14548 -22826
rect 12742 -22920 12760 -22895
rect 11736 -22967 11782 -22929
rect 11736 -23001 11742 -22967
rect 11776 -23001 11782 -22967
rect 11736 -23039 11782 -23001
rect 11736 -23073 11742 -23039
rect 11776 -23073 11782 -23039
rect 11736 -23111 11782 -23073
rect 11736 -23145 11742 -23111
rect 11776 -23145 11782 -23111
rect 11736 -23183 11782 -23145
rect 11736 -23217 11742 -23183
rect 11776 -23217 11782 -23183
rect 11736 -23255 11782 -23217
rect 11736 -23289 11742 -23255
rect 11776 -23289 11782 -23255
rect 11736 -23327 11782 -23289
rect 11736 -23361 11742 -23327
rect 11776 -23361 11782 -23327
rect 9694 -23433 9706 -23399
rect 9740 -23433 9754 -23399
rect 7952 -23502 8440 -23496
rect 7952 -23536 7999 -23502
rect 8033 -23536 8071 -23502
rect 8105 -23536 8143 -23502
rect 8177 -23536 8215 -23502
rect 8249 -23536 8287 -23502
rect 8321 -23536 8359 -23502
rect 8393 -23536 8440 -23502
rect 7952 -23542 8440 -23536
rect 8970 -23502 9458 -23496
rect 8970 -23536 9017 -23502
rect 9051 -23536 9089 -23502
rect 9123 -23536 9161 -23502
rect 9195 -23536 9233 -23502
rect 9267 -23536 9305 -23502
rect 9339 -23536 9377 -23502
rect 9411 -23536 9458 -23502
rect 8970 -23542 9458 -23536
rect 7652 -23826 7724 -23822
rect 7652 -23878 7662 -23826
rect 7714 -23878 7724 -23826
rect 7652 -23882 7724 -23878
rect 8162 -24020 8222 -23542
rect 8668 -23826 8740 -23822
rect 8668 -23878 8678 -23826
rect 8730 -23878 8740 -23826
rect 8668 -23882 8740 -23878
rect 6934 -24026 7422 -24020
rect 6934 -24060 6981 -24026
rect 7015 -24060 7053 -24026
rect 7087 -24060 7125 -24026
rect 7159 -24060 7197 -24026
rect 7231 -24060 7269 -24026
rect 7303 -24060 7341 -24026
rect 7375 -24060 7422 -24026
rect 6934 -24066 7422 -24060
rect 7952 -24026 8440 -24020
rect 7952 -24060 7999 -24026
rect 8033 -24060 8071 -24026
rect 8105 -24060 8143 -24026
rect 8177 -24060 8215 -24026
rect 8249 -24060 8287 -24026
rect 8321 -24060 8359 -24026
rect 8393 -24060 8440 -24026
rect 7952 -24066 8440 -24060
rect 6638 -24160 6652 -24129
rect 5620 -24164 5680 -24163
rect 6646 -24163 6652 -24160
rect 6686 -24160 6698 -24129
rect 7664 -24129 7710 -24098
rect 6686 -24163 6692 -24160
rect 3584 -24235 3598 -24201
rect 3632 -24235 3644 -24201
rect 3584 -24273 3644 -24235
rect 3584 -24307 3598 -24273
rect 3632 -24307 3644 -24273
rect 3584 -24345 3644 -24307
rect 3584 -24379 3598 -24345
rect 3632 -24379 3644 -24345
rect 3584 -24417 3644 -24379
rect 3584 -24451 3598 -24417
rect 3632 -24451 3644 -24417
rect 3584 -24489 3644 -24451
rect 3584 -24523 3598 -24489
rect 3632 -24523 3644 -24489
rect 3584 -24561 3644 -24523
rect 2580 -24633 2614 -24595
rect 2580 -24686 2614 -24667
rect 3584 -24595 3598 -24561
rect 3632 -24595 3644 -24561
rect 4610 -24201 4656 -24170
rect 4610 -24235 4616 -24201
rect 4650 -24235 4656 -24201
rect 4610 -24273 4656 -24235
rect 4610 -24307 4616 -24273
rect 4650 -24307 4656 -24273
rect 4610 -24345 4656 -24307
rect 4610 -24379 4616 -24345
rect 4650 -24379 4656 -24345
rect 4610 -24417 4656 -24379
rect 4610 -24451 4616 -24417
rect 4650 -24451 4656 -24417
rect 4610 -24489 4656 -24451
rect 4610 -24523 4616 -24489
rect 4650 -24523 4656 -24489
rect 4610 -24561 4656 -24523
rect 4610 -24592 4616 -24561
rect 3584 -24633 3644 -24595
rect 3584 -24667 3598 -24633
rect 3632 -24667 3644 -24633
rect 4650 -24592 4656 -24561
rect 5628 -24201 5674 -24164
rect 5628 -24235 5634 -24201
rect 5668 -24235 5674 -24201
rect 5628 -24273 5674 -24235
rect 5628 -24307 5634 -24273
rect 5668 -24307 5674 -24273
rect 5628 -24345 5674 -24307
rect 5628 -24379 5634 -24345
rect 5668 -24379 5674 -24345
rect 5628 -24417 5674 -24379
rect 5628 -24451 5634 -24417
rect 5668 -24451 5674 -24417
rect 5628 -24489 5674 -24451
rect 5628 -24523 5634 -24489
rect 5668 -24523 5674 -24489
rect 5628 -24561 5674 -24523
rect 5628 -24592 5634 -24561
rect 4616 -24633 4650 -24595
rect 2874 -24770 2909 -24736
rect 2943 -24770 2981 -24736
rect 3015 -24770 3053 -24736
rect 3087 -24770 3125 -24736
rect 3159 -24770 3197 -24736
rect 3231 -24770 3269 -24736
rect 3303 -24770 3338 -24736
rect 2442 -24828 2514 -24824
rect 2442 -24880 2452 -24828
rect 2504 -24880 2514 -24828
rect 2442 -24884 2514 -24880
rect 2114 -24932 2186 -24928
rect 2114 -24984 2124 -24932
rect 2176 -24984 2186 -24932
rect 2114 -24988 2186 -24984
rect 2448 -25154 2508 -24884
rect 3584 -24928 3644 -24667
rect 4604 -24667 4616 -24650
rect 5668 -24592 5674 -24561
rect 6646 -24201 6692 -24163
rect 6646 -24235 6652 -24201
rect 6686 -24235 6692 -24201
rect 6646 -24273 6692 -24235
rect 6646 -24307 6652 -24273
rect 6686 -24307 6692 -24273
rect 6646 -24345 6692 -24307
rect 6646 -24379 6652 -24345
rect 6686 -24379 6692 -24345
rect 6646 -24417 6692 -24379
rect 6646 -24451 6652 -24417
rect 6686 -24451 6692 -24417
rect 6646 -24489 6692 -24451
rect 6646 -24523 6652 -24489
rect 6686 -24523 6692 -24489
rect 6646 -24561 6692 -24523
rect 6646 -24592 6652 -24561
rect 5634 -24633 5668 -24595
rect 4650 -24667 4664 -24650
rect 3892 -24770 3927 -24736
rect 3961 -24770 3999 -24736
rect 4033 -24770 4071 -24736
rect 4105 -24770 4143 -24736
rect 4177 -24770 4215 -24736
rect 4249 -24770 4287 -24736
rect 4321 -24770 4356 -24736
rect 3578 -24932 3650 -24928
rect 3578 -24984 3588 -24932
rect 3640 -24984 3650 -24932
rect 3578 -24988 3650 -24984
rect 4092 -25034 4152 -24770
rect 4086 -25038 4158 -25034
rect 4086 -25090 4096 -25038
rect 4148 -25090 4158 -25038
rect 4086 -25094 4158 -25090
rect 2448 -25214 3648 -25154
rect 1064 -25992 1136 -25988
rect 1064 -26044 1074 -25992
rect 1126 -26044 1136 -25992
rect 1064 -26048 1136 -26044
rect 2448 -26066 2508 -25214
rect 2568 -25414 2628 -25214
rect 3054 -25298 3114 -25214
rect 3588 -25418 3648 -25214
rect 4092 -25288 4152 -25094
rect 4604 -25144 4664 -24667
rect 5618 -24667 5634 -24646
rect 6686 -24592 6692 -24561
rect 7664 -24163 7670 -24129
rect 7704 -24163 7710 -24129
rect 7664 -24201 7710 -24163
rect 7664 -24235 7670 -24201
rect 7704 -24235 7710 -24201
rect 7664 -24273 7710 -24235
rect 7664 -24307 7670 -24273
rect 7704 -24307 7710 -24273
rect 7664 -24345 7710 -24307
rect 7664 -24379 7670 -24345
rect 7704 -24379 7710 -24345
rect 7664 -24417 7710 -24379
rect 7664 -24451 7670 -24417
rect 7704 -24451 7710 -24417
rect 7664 -24489 7710 -24451
rect 7664 -24523 7670 -24489
rect 7704 -24523 7710 -24489
rect 7664 -24561 7710 -24523
rect 7664 -24592 7670 -24561
rect 6652 -24633 6686 -24595
rect 5668 -24667 5678 -24646
rect 4910 -24770 4945 -24736
rect 4979 -24770 5017 -24736
rect 5051 -24770 5089 -24736
rect 5123 -24770 5161 -24736
rect 5195 -24770 5233 -24736
rect 5267 -24770 5305 -24736
rect 5339 -24770 5374 -24736
rect 5112 -25034 5172 -24770
rect 5618 -24824 5678 -24667
rect 6640 -24667 6652 -24662
rect 7704 -24592 7710 -24561
rect 8674 -24129 8734 -23882
rect 9174 -24020 9234 -23542
rect 9694 -23822 9754 -23433
rect 10706 -23399 10766 -23394
rect 10706 -23433 10724 -23399
rect 10758 -23433 10766 -23399
rect 11736 -23399 11782 -23361
rect 11736 -23400 11742 -23399
rect 9988 -23502 10476 -23496
rect 9988 -23536 10035 -23502
rect 10069 -23536 10107 -23502
rect 10141 -23536 10179 -23502
rect 10213 -23536 10251 -23502
rect 10285 -23536 10323 -23502
rect 10357 -23536 10395 -23502
rect 10429 -23536 10476 -23502
rect 9988 -23542 10476 -23536
rect 9688 -23826 9760 -23822
rect 9688 -23878 9698 -23826
rect 9750 -23878 9760 -23826
rect 9688 -23882 9760 -23878
rect 10204 -24020 10264 -23542
rect 10706 -23654 10766 -23433
rect 11724 -23433 11742 -23400
rect 11776 -23400 11782 -23399
rect 12754 -22929 12760 -22920
rect 12794 -22920 12802 -22895
rect 13772 -22895 13818 -22864
rect 12794 -22929 12800 -22920
rect 12754 -22967 12800 -22929
rect 12754 -23001 12760 -22967
rect 12794 -23001 12800 -22967
rect 12754 -23039 12800 -23001
rect 12754 -23073 12760 -23039
rect 12794 -23073 12800 -23039
rect 12754 -23111 12800 -23073
rect 12754 -23145 12760 -23111
rect 12794 -23145 12800 -23111
rect 12754 -23183 12800 -23145
rect 12754 -23217 12760 -23183
rect 12794 -23217 12800 -23183
rect 12754 -23255 12800 -23217
rect 12754 -23289 12760 -23255
rect 12794 -23289 12800 -23255
rect 12754 -23327 12800 -23289
rect 12754 -23361 12760 -23327
rect 12794 -23361 12800 -23327
rect 12754 -23399 12800 -23361
rect 11776 -23433 11784 -23400
rect 11006 -23502 11494 -23496
rect 11006 -23536 11053 -23502
rect 11087 -23536 11125 -23502
rect 11159 -23536 11197 -23502
rect 11231 -23536 11269 -23502
rect 11303 -23536 11341 -23502
rect 11375 -23536 11413 -23502
rect 11447 -23536 11494 -23502
rect 11006 -23542 11494 -23536
rect 10556 -23714 10766 -23654
rect 11220 -23708 11280 -23542
rect 11724 -23594 11784 -23433
rect 12754 -23433 12760 -23399
rect 12794 -23433 12800 -23399
rect 13772 -22929 13778 -22895
rect 13812 -22929 13818 -22895
rect 14786 -22895 14846 -22612
rect 15282 -22786 15342 -22510
rect 15078 -22792 15566 -22786
rect 15078 -22826 15125 -22792
rect 15159 -22826 15197 -22792
rect 15231 -22826 15269 -22792
rect 15303 -22826 15341 -22792
rect 15375 -22826 15413 -22792
rect 15447 -22826 15485 -22792
rect 15519 -22826 15566 -22792
rect 15078 -22832 15566 -22826
rect 14786 -22924 14796 -22895
rect 13772 -22967 13818 -22929
rect 13772 -23001 13778 -22967
rect 13812 -23001 13818 -22967
rect 13772 -23039 13818 -23001
rect 13772 -23073 13778 -23039
rect 13812 -23073 13818 -23039
rect 13772 -23111 13818 -23073
rect 13772 -23145 13778 -23111
rect 13812 -23145 13818 -23111
rect 13772 -23183 13818 -23145
rect 13772 -23217 13778 -23183
rect 13812 -23217 13818 -23183
rect 13772 -23255 13818 -23217
rect 13772 -23289 13778 -23255
rect 13812 -23289 13818 -23255
rect 13772 -23327 13818 -23289
rect 13772 -23361 13778 -23327
rect 13812 -23361 13818 -23327
rect 13772 -23399 13818 -23361
rect 13772 -23400 13778 -23399
rect 12754 -23464 12800 -23433
rect 13766 -23433 13778 -23400
rect 13812 -23400 13818 -23399
rect 14790 -22929 14796 -22924
rect 14830 -22924 14846 -22895
rect 15800 -22895 15860 -22502
rect 16308 -22786 16368 -22410
rect 16808 -22556 16880 -22552
rect 16808 -22608 16818 -22556
rect 16870 -22608 16880 -22556
rect 16808 -22612 16880 -22608
rect 16096 -22792 16584 -22786
rect 16096 -22826 16143 -22792
rect 16177 -22826 16215 -22792
rect 16249 -22826 16287 -22792
rect 16321 -22826 16359 -22792
rect 16393 -22826 16431 -22792
rect 16465 -22826 16503 -22792
rect 16537 -22826 16584 -22792
rect 16096 -22832 16584 -22826
rect 15800 -22912 15814 -22895
rect 14830 -22929 14836 -22924
rect 14790 -22967 14836 -22929
rect 14790 -23001 14796 -22967
rect 14830 -23001 14836 -22967
rect 14790 -23039 14836 -23001
rect 14790 -23073 14796 -23039
rect 14830 -23073 14836 -23039
rect 14790 -23111 14836 -23073
rect 14790 -23145 14796 -23111
rect 14830 -23145 14836 -23111
rect 14790 -23183 14836 -23145
rect 14790 -23217 14796 -23183
rect 14830 -23217 14836 -23183
rect 14790 -23255 14836 -23217
rect 14790 -23289 14796 -23255
rect 14830 -23289 14836 -23255
rect 14790 -23327 14836 -23289
rect 14790 -23361 14796 -23327
rect 14830 -23361 14836 -23327
rect 14790 -23399 14836 -23361
rect 13812 -23433 13826 -23400
rect 12024 -23502 12512 -23496
rect 12024 -23536 12071 -23502
rect 12105 -23536 12143 -23502
rect 12177 -23536 12215 -23502
rect 12249 -23536 12287 -23502
rect 12321 -23536 12359 -23502
rect 12393 -23536 12431 -23502
rect 12465 -23536 12512 -23502
rect 12024 -23542 12512 -23536
rect 13042 -23502 13530 -23496
rect 13042 -23536 13089 -23502
rect 13123 -23536 13161 -23502
rect 13195 -23536 13233 -23502
rect 13267 -23536 13305 -23502
rect 13339 -23536 13377 -23502
rect 13411 -23536 13449 -23502
rect 13483 -23536 13530 -23502
rect 13042 -23542 13530 -23536
rect 13766 -23594 13826 -23433
rect 14790 -23433 14796 -23399
rect 14830 -23433 14836 -23399
rect 15808 -22929 15814 -22912
rect 15848 -22912 15860 -22895
rect 16814 -22895 16874 -22612
rect 17328 -22786 17388 -22310
rect 17840 -22678 17900 -22201
rect 18852 -22201 18868 -22176
rect 18902 -22176 18908 -22167
rect 19880 -21735 19926 -21702
rect 19880 -21769 19886 -21735
rect 19920 -21769 19926 -21735
rect 19880 -21807 19926 -21769
rect 19880 -21841 19886 -21807
rect 19920 -21841 19926 -21807
rect 19880 -21879 19926 -21841
rect 19880 -21913 19886 -21879
rect 19920 -21913 19926 -21879
rect 19880 -21951 19926 -21913
rect 19880 -21985 19886 -21951
rect 19920 -21985 19926 -21951
rect 19880 -22023 19926 -21985
rect 19880 -22057 19886 -22023
rect 19920 -22057 19926 -22023
rect 19880 -22095 19926 -22057
rect 19880 -22129 19886 -22095
rect 19920 -22129 19926 -22095
rect 19880 -22167 19926 -22129
rect 20898 -21735 20944 -21697
rect 20898 -21769 20904 -21735
rect 20938 -21769 20944 -21735
rect 20898 -21807 20944 -21769
rect 20898 -21841 20904 -21807
rect 20938 -21841 20944 -21807
rect 20898 -21879 20944 -21841
rect 20898 -21913 20904 -21879
rect 20938 -21913 20944 -21879
rect 20898 -21951 20944 -21913
rect 20898 -21985 20904 -21951
rect 20938 -21985 20944 -21951
rect 20898 -22023 20944 -21985
rect 20898 -22057 20904 -22023
rect 20938 -22057 20944 -22023
rect 20898 -22095 20944 -22057
rect 20898 -22129 20904 -22095
rect 20938 -22129 20944 -22095
rect 20898 -22166 20944 -22129
rect 21916 -21697 21922 -21663
rect 21956 -21697 21962 -21663
rect 21916 -21735 21962 -21697
rect 21916 -21769 21922 -21735
rect 21956 -21769 21962 -21735
rect 21916 -21807 21962 -21769
rect 21916 -21841 21922 -21807
rect 21956 -21841 21962 -21807
rect 21916 -21879 21962 -21841
rect 21916 -21913 21922 -21879
rect 21956 -21913 21962 -21879
rect 21916 -21951 21962 -21913
rect 21916 -21985 21922 -21951
rect 21956 -21985 21962 -21951
rect 21916 -22023 21962 -21985
rect 21916 -22057 21922 -22023
rect 21956 -22057 21962 -22023
rect 21916 -22095 21962 -22057
rect 21916 -22129 21922 -22095
rect 21956 -22129 21962 -22095
rect 18902 -22201 18912 -22176
rect 19880 -22180 19886 -22167
rect 18132 -22270 18620 -22264
rect 18132 -22304 18179 -22270
rect 18213 -22304 18251 -22270
rect 18285 -22304 18323 -22270
rect 18357 -22304 18395 -22270
rect 18429 -22304 18467 -22270
rect 18501 -22304 18539 -22270
rect 18573 -22304 18620 -22270
rect 18132 -22310 18620 -22304
rect 17834 -22682 17906 -22678
rect 17834 -22734 17844 -22682
rect 17896 -22734 17906 -22682
rect 17834 -22738 17906 -22734
rect 17114 -22792 17602 -22786
rect 17114 -22826 17161 -22792
rect 17195 -22826 17233 -22792
rect 17267 -22826 17305 -22792
rect 17339 -22826 17377 -22792
rect 17411 -22826 17449 -22792
rect 17483 -22826 17521 -22792
rect 17555 -22826 17602 -22792
rect 17114 -22832 17602 -22826
rect 15848 -22929 15854 -22912
rect 16814 -22924 16832 -22895
rect 15808 -22967 15854 -22929
rect 15808 -23001 15814 -22967
rect 15848 -23001 15854 -22967
rect 15808 -23039 15854 -23001
rect 15808 -23073 15814 -23039
rect 15848 -23073 15854 -23039
rect 15808 -23111 15854 -23073
rect 15808 -23145 15814 -23111
rect 15848 -23145 15854 -23111
rect 15808 -23183 15854 -23145
rect 15808 -23217 15814 -23183
rect 15848 -23217 15854 -23183
rect 15808 -23255 15854 -23217
rect 15808 -23289 15814 -23255
rect 15848 -23289 15854 -23255
rect 15808 -23327 15854 -23289
rect 15808 -23361 15814 -23327
rect 15848 -23361 15854 -23327
rect 15808 -23399 15854 -23361
rect 15808 -23408 15814 -23399
rect 14790 -23464 14836 -23433
rect 15802 -23433 15814 -23408
rect 15848 -23408 15854 -23399
rect 16826 -22929 16832 -22924
rect 16866 -22924 16874 -22895
rect 17840 -22895 17900 -22738
rect 18344 -22786 18404 -22310
rect 18852 -22552 18912 -22201
rect 19870 -22201 19886 -22180
rect 19920 -22180 19926 -22167
rect 20892 -22167 20952 -22166
rect 19920 -22201 19930 -22180
rect 19150 -22270 19638 -22264
rect 19150 -22304 19197 -22270
rect 19231 -22304 19269 -22270
rect 19303 -22304 19341 -22270
rect 19375 -22304 19413 -22270
rect 19447 -22304 19485 -22270
rect 19519 -22304 19557 -22270
rect 19591 -22304 19638 -22270
rect 19150 -22310 19638 -22304
rect 18846 -22556 18918 -22552
rect 18846 -22608 18856 -22556
rect 18908 -22608 18918 -22556
rect 18846 -22612 18918 -22608
rect 19378 -22786 19438 -22310
rect 19870 -22678 19930 -22201
rect 20892 -22201 20904 -22167
rect 20938 -22201 20952 -22167
rect 21916 -22167 21962 -22129
rect 21916 -22174 21922 -22167
rect 20168 -22270 20656 -22264
rect 20168 -22304 20215 -22270
rect 20249 -22304 20287 -22270
rect 20321 -22304 20359 -22270
rect 20393 -22304 20431 -22270
rect 20465 -22304 20503 -22270
rect 20537 -22304 20575 -22270
rect 20609 -22304 20656 -22270
rect 20168 -22310 20656 -22304
rect 19864 -22682 19936 -22678
rect 19864 -22734 19874 -22682
rect 19926 -22734 19936 -22682
rect 19864 -22738 19936 -22734
rect 20396 -22680 20456 -22310
rect 20892 -22552 20952 -22201
rect 21906 -22201 21922 -22174
rect 21956 -22174 21962 -22167
rect 22934 -21663 22980 -21632
rect 22934 -21697 22940 -21663
rect 22974 -21697 22980 -21663
rect 22934 -21735 22980 -21697
rect 22934 -21769 22940 -21735
rect 22974 -21769 22980 -21735
rect 22934 -21807 22980 -21769
rect 22934 -21841 22940 -21807
rect 22974 -21841 22980 -21807
rect 22934 -21879 22980 -21841
rect 22934 -21913 22940 -21879
rect 22974 -21913 22980 -21879
rect 22934 -21951 22980 -21913
rect 22934 -21985 22940 -21951
rect 22974 -21985 22980 -21951
rect 22934 -22023 22980 -21985
rect 22934 -22057 22940 -22023
rect 22974 -22057 22980 -22023
rect 22934 -22095 22980 -22057
rect 22934 -22129 22940 -22095
rect 22974 -22129 22980 -22095
rect 22934 -22167 22980 -22129
rect 21956 -22201 21966 -22174
rect 22934 -22192 22940 -22167
rect 21186 -22270 21674 -22264
rect 21186 -22304 21233 -22270
rect 21267 -22304 21305 -22270
rect 21339 -22304 21377 -22270
rect 21411 -22304 21449 -22270
rect 21483 -22304 21521 -22270
rect 21555 -22304 21593 -22270
rect 21627 -22304 21674 -22270
rect 21186 -22310 21674 -22304
rect 21410 -22548 21470 -22310
rect 21906 -22346 21966 -22201
rect 22926 -22201 22940 -22192
rect 22974 -22192 22980 -22167
rect 22974 -22201 22986 -22192
rect 22204 -22270 22692 -22264
rect 22204 -22304 22251 -22270
rect 22285 -22304 22323 -22270
rect 22357 -22304 22395 -22270
rect 22429 -22304 22467 -22270
rect 22501 -22304 22539 -22270
rect 22573 -22304 22611 -22270
rect 22645 -22304 22692 -22270
rect 22204 -22310 22692 -22304
rect 22412 -22344 22472 -22310
rect 22926 -22344 22986 -22201
rect 22412 -22346 22986 -22344
rect 21906 -22406 22986 -22346
rect 21906 -22442 21966 -22406
rect 21900 -22446 21972 -22442
rect 21900 -22498 21910 -22446
rect 21962 -22498 21972 -22446
rect 21900 -22502 21972 -22498
rect 21404 -22552 21476 -22548
rect 20886 -22556 20958 -22552
rect 20886 -22608 20896 -22556
rect 20948 -22608 20958 -22556
rect 21404 -22604 21414 -22552
rect 21466 -22604 21476 -22552
rect 21404 -22608 21476 -22604
rect 22916 -22552 22988 -22548
rect 22916 -22604 22926 -22552
rect 22978 -22604 22988 -22552
rect 22916 -22608 22988 -22604
rect 20886 -22612 20958 -22608
rect 20396 -22732 20400 -22680
rect 20452 -22732 20456 -22680
rect 18132 -22792 18620 -22786
rect 18132 -22826 18179 -22792
rect 18213 -22826 18251 -22792
rect 18285 -22826 18323 -22792
rect 18357 -22826 18395 -22792
rect 18429 -22826 18467 -22792
rect 18501 -22826 18539 -22792
rect 18573 -22826 18620 -22792
rect 18132 -22832 18620 -22826
rect 19150 -22792 19638 -22786
rect 19150 -22826 19197 -22792
rect 19231 -22826 19269 -22792
rect 19303 -22826 19341 -22792
rect 19375 -22826 19413 -22792
rect 19447 -22826 19485 -22792
rect 19519 -22826 19557 -22792
rect 19591 -22826 19638 -22792
rect 19150 -22832 19638 -22826
rect 17840 -22922 17850 -22895
rect 16866 -22929 16872 -22924
rect 16826 -22967 16872 -22929
rect 16826 -23001 16832 -22967
rect 16866 -23001 16872 -22967
rect 16826 -23039 16872 -23001
rect 16826 -23073 16832 -23039
rect 16866 -23073 16872 -23039
rect 16826 -23111 16872 -23073
rect 16826 -23145 16832 -23111
rect 16866 -23145 16872 -23111
rect 16826 -23183 16872 -23145
rect 16826 -23217 16832 -23183
rect 16866 -23217 16872 -23183
rect 16826 -23255 16872 -23217
rect 16826 -23289 16832 -23255
rect 16866 -23289 16872 -23255
rect 16826 -23327 16872 -23289
rect 16826 -23361 16832 -23327
rect 16866 -23361 16872 -23327
rect 16826 -23399 16872 -23361
rect 17844 -22929 17850 -22922
rect 17884 -22922 17900 -22895
rect 18862 -22895 18908 -22864
rect 17884 -22929 17890 -22922
rect 17844 -22967 17890 -22929
rect 17844 -23001 17850 -22967
rect 17884 -23001 17890 -22967
rect 17844 -23039 17890 -23001
rect 17844 -23073 17850 -23039
rect 17884 -23073 17890 -23039
rect 17844 -23111 17890 -23073
rect 17844 -23145 17850 -23111
rect 17884 -23145 17890 -23111
rect 17844 -23183 17890 -23145
rect 17844 -23217 17850 -23183
rect 17884 -23217 17890 -23183
rect 17844 -23255 17890 -23217
rect 17844 -23289 17850 -23255
rect 17884 -23289 17890 -23255
rect 17844 -23327 17890 -23289
rect 17844 -23361 17850 -23327
rect 17884 -23361 17890 -23327
rect 17844 -23392 17890 -23361
rect 18862 -22929 18868 -22895
rect 18902 -22929 18908 -22895
rect 19870 -22895 19930 -22738
rect 20396 -22786 20456 -22732
rect 21410 -22786 21470 -22608
rect 21904 -22680 21976 -22676
rect 21904 -22732 21914 -22680
rect 21966 -22732 21976 -22680
rect 21904 -22736 21976 -22732
rect 20168 -22792 20656 -22786
rect 20168 -22826 20215 -22792
rect 20249 -22826 20287 -22792
rect 20321 -22826 20359 -22792
rect 20393 -22826 20431 -22792
rect 20465 -22826 20503 -22792
rect 20537 -22826 20575 -22792
rect 20609 -22826 20656 -22792
rect 20168 -22832 20656 -22826
rect 21186 -22792 21674 -22786
rect 21186 -22826 21233 -22792
rect 21267 -22826 21305 -22792
rect 21339 -22826 21377 -22792
rect 21411 -22826 21449 -22792
rect 21483 -22826 21521 -22792
rect 21555 -22826 21593 -22792
rect 21627 -22826 21674 -22792
rect 21186 -22832 21674 -22826
rect 19870 -22922 19886 -22895
rect 18862 -22967 18908 -22929
rect 18862 -23001 18868 -22967
rect 18902 -23001 18908 -22967
rect 18862 -23039 18908 -23001
rect 18862 -23073 18868 -23039
rect 18902 -23073 18908 -23039
rect 18862 -23111 18908 -23073
rect 18862 -23145 18868 -23111
rect 18902 -23145 18908 -23111
rect 18862 -23183 18908 -23145
rect 18862 -23217 18868 -23183
rect 18902 -23217 18908 -23183
rect 18862 -23255 18908 -23217
rect 18862 -23289 18868 -23255
rect 18902 -23289 18908 -23255
rect 18862 -23327 18908 -23289
rect 18862 -23361 18868 -23327
rect 18902 -23361 18908 -23327
rect 15848 -23433 15862 -23408
rect 16826 -23412 16832 -23399
rect 14060 -23502 14548 -23496
rect 14060 -23536 14107 -23502
rect 14141 -23536 14179 -23502
rect 14213 -23536 14251 -23502
rect 14285 -23536 14323 -23502
rect 14357 -23536 14395 -23502
rect 14429 -23536 14467 -23502
rect 14501 -23536 14548 -23502
rect 14060 -23542 14548 -23536
rect 15078 -23502 15566 -23496
rect 15078 -23536 15125 -23502
rect 15159 -23536 15197 -23502
rect 15231 -23536 15269 -23502
rect 15303 -23536 15341 -23502
rect 15375 -23536 15413 -23502
rect 15447 -23536 15485 -23502
rect 15519 -23536 15566 -23502
rect 15078 -23542 15566 -23536
rect 15802 -23594 15862 -23433
rect 16816 -23433 16832 -23412
rect 16866 -23412 16872 -23399
rect 17838 -23399 17898 -23392
rect 16866 -23433 16876 -23412
rect 16096 -23502 16584 -23496
rect 16096 -23536 16143 -23502
rect 16177 -23536 16215 -23502
rect 16249 -23536 16287 -23502
rect 16321 -23536 16359 -23502
rect 16393 -23536 16431 -23502
rect 16465 -23536 16503 -23502
rect 16537 -23536 16584 -23502
rect 16096 -23542 16584 -23536
rect 11718 -23598 11790 -23594
rect 11718 -23650 11728 -23598
rect 11780 -23650 11790 -23598
rect 11718 -23654 11790 -23650
rect 13760 -23598 13832 -23594
rect 13760 -23650 13770 -23598
rect 13822 -23650 13832 -23598
rect 13760 -23654 13832 -23650
rect 15796 -23598 15868 -23594
rect 15796 -23650 15806 -23598
rect 15858 -23650 15868 -23598
rect 15796 -23654 15868 -23650
rect 16308 -23704 16368 -23542
rect 16816 -23602 16876 -23433
rect 17838 -23433 17850 -23399
rect 17884 -23433 17898 -23399
rect 18862 -23399 18908 -23361
rect 18862 -23408 18868 -23399
rect 17114 -23502 17602 -23496
rect 17114 -23536 17161 -23502
rect 17195 -23536 17233 -23502
rect 17267 -23536 17305 -23502
rect 17339 -23536 17377 -23502
rect 17411 -23536 17449 -23502
rect 17483 -23536 17521 -23502
rect 17555 -23536 17602 -23502
rect 17114 -23542 17602 -23536
rect 16816 -23662 17022 -23602
rect 16302 -23708 16374 -23704
rect 11214 -23712 11286 -23708
rect 10556 -23926 10616 -23714
rect 11214 -23764 11224 -23712
rect 11276 -23764 11286 -23712
rect 16302 -23760 16312 -23708
rect 16364 -23760 16374 -23708
rect 16302 -23764 16374 -23760
rect 11214 -23768 11286 -23764
rect 10706 -23826 10778 -23822
rect 10706 -23878 10716 -23826
rect 10768 -23878 10778 -23826
rect 10706 -23882 10778 -23878
rect 12736 -23826 12808 -23822
rect 12736 -23878 12746 -23826
rect 12798 -23878 12808 -23826
rect 12736 -23882 12808 -23878
rect 14774 -23826 14846 -23822
rect 14774 -23878 14784 -23826
rect 14836 -23878 14846 -23826
rect 14774 -23882 14846 -23878
rect 16810 -23826 16882 -23822
rect 16810 -23878 16820 -23826
rect 16872 -23878 16882 -23826
rect 16810 -23882 16882 -23878
rect 10550 -23930 10622 -23926
rect 10550 -23982 10560 -23930
rect 10612 -23982 10622 -23930
rect 10550 -23986 10622 -23982
rect 8970 -24026 9458 -24020
rect 8970 -24060 9017 -24026
rect 9051 -24060 9089 -24026
rect 9123 -24060 9161 -24026
rect 9195 -24060 9233 -24026
rect 9267 -24060 9305 -24026
rect 9339 -24060 9377 -24026
rect 9411 -24060 9458 -24026
rect 8970 -24066 9458 -24060
rect 9988 -24026 10476 -24020
rect 9988 -24060 10035 -24026
rect 10069 -24060 10107 -24026
rect 10141 -24060 10179 -24026
rect 10213 -24060 10251 -24026
rect 10285 -24060 10323 -24026
rect 10357 -24060 10395 -24026
rect 10429 -24060 10476 -24026
rect 9988 -24066 10476 -24060
rect 8674 -24163 8688 -24129
rect 8722 -24163 8734 -24129
rect 8674 -24201 8734 -24163
rect 8674 -24235 8688 -24201
rect 8722 -24235 8734 -24201
rect 8674 -24273 8734 -24235
rect 8674 -24307 8688 -24273
rect 8722 -24307 8734 -24273
rect 8674 -24345 8734 -24307
rect 8674 -24379 8688 -24345
rect 8722 -24379 8734 -24345
rect 8674 -24417 8734 -24379
rect 8674 -24451 8688 -24417
rect 8722 -24451 8734 -24417
rect 8674 -24489 8734 -24451
rect 8674 -24523 8688 -24489
rect 8722 -24523 8734 -24489
rect 8674 -24561 8734 -24523
rect 8674 -24592 8688 -24561
rect 7670 -24633 7704 -24595
rect 6686 -24667 6700 -24662
rect 5928 -24770 5963 -24736
rect 5997 -24770 6035 -24736
rect 6069 -24770 6107 -24736
rect 6141 -24770 6179 -24736
rect 6213 -24770 6251 -24736
rect 6285 -24770 6323 -24736
rect 6357 -24770 6392 -24736
rect 5612 -24828 5684 -24824
rect 5612 -24880 5622 -24828
rect 5674 -24880 5684 -24828
rect 5612 -24884 5684 -24880
rect 5618 -24932 5690 -24928
rect 5618 -24984 5628 -24932
rect 5680 -24984 5690 -24932
rect 5618 -24988 5690 -24984
rect 5106 -25038 5178 -25034
rect 5106 -25090 5116 -25038
rect 5168 -25090 5178 -25038
rect 5106 -25094 5178 -25090
rect 4598 -25148 4670 -25144
rect 4598 -25200 4608 -25148
rect 4660 -25200 4670 -25148
rect 4598 -25204 4670 -25200
rect 3584 -26066 3644 -25870
rect 2442 -26070 2514 -26066
rect 2442 -26122 2452 -26070
rect 2504 -26122 2514 -26070
rect 2442 -26126 2514 -26122
rect 3578 -26070 3650 -26066
rect 3578 -26122 3588 -26070
rect 3640 -26122 3650 -26070
rect 3578 -26126 3650 -26122
rect 4096 -26174 4156 -25970
rect 4090 -26178 4162 -26174
rect 4090 -26230 4100 -26178
rect 4152 -26230 4162 -26178
rect 4090 -26234 4162 -26230
rect 4604 -26430 4664 -25204
rect 5112 -25284 5172 -25094
rect 5624 -25356 5684 -24988
rect 6136 -25034 6196 -24770
rect 6130 -25038 6202 -25034
rect 6130 -25090 6140 -25038
rect 6192 -25090 6202 -25038
rect 6130 -25094 6202 -25090
rect 6136 -25290 6196 -25094
rect 6640 -25144 6700 -24667
rect 8722 -24592 8734 -24561
rect 9700 -24129 9746 -24098
rect 9700 -24163 9706 -24129
rect 9740 -24163 9746 -24129
rect 9700 -24201 9746 -24163
rect 10712 -24129 10772 -23882
rect 11006 -24026 11218 -24020
rect 11278 -24026 11494 -24020
rect 11006 -24060 11053 -24026
rect 11087 -24060 11125 -24026
rect 11159 -24060 11197 -24026
rect 11231 -24060 11269 -24026
rect 11303 -24060 11341 -24026
rect 11375 -24060 11413 -24026
rect 11447 -24060 11494 -24026
rect 11006 -24066 11494 -24060
rect 12024 -24026 12228 -24020
rect 12288 -24026 12512 -24020
rect 12024 -24060 12071 -24026
rect 12105 -24060 12143 -24026
rect 12177 -24060 12215 -24026
rect 12249 -24060 12287 -24026
rect 12321 -24060 12359 -24026
rect 12393 -24060 12431 -24026
rect 12465 -24060 12512 -24026
rect 12024 -24066 12512 -24060
rect 10712 -24163 10724 -24129
rect 10758 -24163 10772 -24129
rect 11730 -24129 11790 -24110
rect 11730 -24146 11742 -24129
rect 10712 -24166 10772 -24163
rect 11736 -24163 11742 -24146
rect 11776 -24146 11790 -24129
rect 12742 -24129 12802 -23882
rect 13042 -24026 13242 -24020
rect 13302 -24026 13530 -24020
rect 13042 -24060 13089 -24026
rect 13123 -24060 13161 -24026
rect 13195 -24060 13233 -24026
rect 13267 -24060 13305 -24026
rect 13339 -24060 13377 -24026
rect 13411 -24060 13449 -24026
rect 13483 -24060 13530 -24026
rect 13042 -24066 13530 -24060
rect 14060 -24026 14270 -24020
rect 14330 -24026 14548 -24020
rect 14060 -24060 14107 -24026
rect 14141 -24060 14179 -24026
rect 14213 -24060 14251 -24026
rect 14285 -24060 14323 -24026
rect 14357 -24060 14395 -24026
rect 14429 -24060 14467 -24026
rect 14501 -24060 14548 -24026
rect 14060 -24066 14548 -24060
rect 11776 -24163 11782 -24146
rect 12742 -24160 12760 -24129
rect 9700 -24235 9706 -24201
rect 9740 -24235 9746 -24201
rect 9700 -24273 9746 -24235
rect 9700 -24307 9706 -24273
rect 9740 -24307 9746 -24273
rect 9700 -24345 9746 -24307
rect 9700 -24379 9706 -24345
rect 9740 -24379 9746 -24345
rect 9700 -24417 9746 -24379
rect 9700 -24451 9706 -24417
rect 9740 -24451 9746 -24417
rect 9700 -24489 9746 -24451
rect 9700 -24523 9706 -24489
rect 9740 -24523 9746 -24489
rect 9700 -24561 9746 -24523
rect 9700 -24592 9706 -24561
rect 8688 -24633 8722 -24595
rect 7670 -24672 7704 -24667
rect 8678 -24667 8688 -24666
rect 9740 -24592 9746 -24561
rect 10718 -24201 10764 -24166
rect 10718 -24235 10724 -24201
rect 10758 -24235 10764 -24201
rect 10718 -24273 10764 -24235
rect 10718 -24307 10724 -24273
rect 10758 -24307 10764 -24273
rect 10718 -24345 10764 -24307
rect 10718 -24379 10724 -24345
rect 10758 -24379 10764 -24345
rect 10718 -24417 10764 -24379
rect 10718 -24451 10724 -24417
rect 10758 -24451 10764 -24417
rect 10718 -24489 10764 -24451
rect 10718 -24523 10724 -24489
rect 10758 -24523 10764 -24489
rect 10718 -24561 10764 -24523
rect 10718 -24592 10724 -24561
rect 9706 -24633 9740 -24595
rect 8722 -24667 8738 -24666
rect 6946 -24770 6981 -24736
rect 7015 -24770 7053 -24736
rect 7087 -24770 7125 -24736
rect 7159 -24770 7197 -24736
rect 7231 -24770 7269 -24736
rect 7303 -24770 7341 -24736
rect 7375 -24770 7410 -24736
rect 7154 -25034 7214 -24770
rect 7654 -24928 7714 -24672
rect 7964 -24770 7999 -24736
rect 8033 -24770 8071 -24736
rect 8105 -24770 8143 -24736
rect 8177 -24770 8215 -24736
rect 8249 -24770 8287 -24736
rect 8321 -24770 8359 -24736
rect 8393 -24770 8428 -24736
rect 7648 -24932 7720 -24928
rect 7648 -24984 7658 -24932
rect 7710 -24984 7720 -24932
rect 7648 -24988 7720 -24984
rect 8168 -25034 8228 -24770
rect 7148 -25038 7220 -25034
rect 7148 -25090 7158 -25038
rect 7210 -25090 7220 -25038
rect 7148 -25094 7220 -25090
rect 8162 -25038 8234 -25034
rect 8162 -25090 8172 -25038
rect 8224 -25090 8234 -25038
rect 8162 -25094 8234 -25090
rect 6634 -25148 6706 -25144
rect 6634 -25200 6644 -25148
rect 6696 -25200 6706 -25148
rect 6634 -25204 6706 -25200
rect 5110 -26178 5170 -25968
rect 5110 -26230 5114 -26178
rect 5166 -26230 5170 -26178
rect 5110 -26240 5170 -26230
rect 6132 -26178 6192 -25968
rect 6132 -26230 6136 -26178
rect 6188 -26230 6192 -26178
rect 6132 -26240 6192 -26230
rect 6640 -26430 6700 -25204
rect 7154 -25294 7214 -25094
rect 8168 -25284 8228 -25094
rect 8678 -25144 8738 -24667
rect 9694 -24667 9706 -24660
rect 10758 -24592 10764 -24561
rect 11736 -24201 11782 -24163
rect 11736 -24235 11742 -24201
rect 11776 -24235 11782 -24201
rect 11736 -24273 11782 -24235
rect 11736 -24307 11742 -24273
rect 11776 -24307 11782 -24273
rect 11736 -24345 11782 -24307
rect 11736 -24379 11742 -24345
rect 11776 -24379 11782 -24345
rect 11736 -24417 11782 -24379
rect 11736 -24451 11742 -24417
rect 11776 -24451 11782 -24417
rect 11736 -24489 11782 -24451
rect 11736 -24523 11742 -24489
rect 11776 -24523 11782 -24489
rect 11736 -24561 11782 -24523
rect 11736 -24592 11742 -24561
rect 10724 -24633 10758 -24595
rect 9740 -24667 9754 -24660
rect 8982 -24770 9017 -24736
rect 9051 -24770 9089 -24736
rect 9123 -24770 9161 -24736
rect 9195 -24770 9233 -24736
rect 9267 -24770 9305 -24736
rect 9339 -24770 9377 -24736
rect 9411 -24770 9446 -24736
rect 9200 -25034 9260 -24770
rect 9694 -24928 9754 -24667
rect 10716 -24667 10724 -24662
rect 11776 -24592 11782 -24561
rect 12754 -24163 12760 -24160
rect 12794 -24160 12802 -24129
rect 13766 -24129 13826 -24110
rect 13766 -24142 13778 -24129
rect 12794 -24163 12800 -24160
rect 12754 -24201 12800 -24163
rect 12754 -24235 12760 -24201
rect 12794 -24235 12800 -24201
rect 12754 -24273 12800 -24235
rect 12754 -24307 12760 -24273
rect 12794 -24307 12800 -24273
rect 12754 -24345 12800 -24307
rect 12754 -24379 12760 -24345
rect 12794 -24379 12800 -24345
rect 12754 -24417 12800 -24379
rect 12754 -24451 12760 -24417
rect 12794 -24451 12800 -24417
rect 12754 -24489 12800 -24451
rect 12754 -24523 12760 -24489
rect 12794 -24523 12800 -24489
rect 12754 -24561 12800 -24523
rect 12754 -24592 12760 -24561
rect 11742 -24633 11776 -24595
rect 10758 -24667 10776 -24662
rect 10212 -24736 10272 -24734
rect 10000 -24770 10035 -24736
rect 10069 -24770 10107 -24736
rect 10141 -24770 10179 -24736
rect 10213 -24770 10251 -24736
rect 10285 -24770 10323 -24736
rect 10357 -24770 10395 -24736
rect 10429 -24770 10464 -24736
rect 9842 -24826 9914 -24822
rect 9842 -24878 9852 -24826
rect 9904 -24878 9914 -24826
rect 9842 -24882 9914 -24878
rect 9688 -24932 9760 -24928
rect 9688 -24984 9698 -24932
rect 9750 -24984 9760 -24932
rect 9688 -24988 9760 -24984
rect 9194 -25038 9266 -25034
rect 9194 -25090 9204 -25038
rect 9256 -25090 9266 -25038
rect 9848 -25066 9908 -24882
rect 10212 -25034 10272 -24770
rect 9194 -25094 9266 -25090
rect 8672 -25148 8744 -25144
rect 8672 -25200 8682 -25148
rect 8734 -25200 8744 -25148
rect 8672 -25204 8744 -25200
rect 7144 -26168 7204 -25964
rect 7654 -26066 7714 -25876
rect 7648 -26070 7720 -26066
rect 7648 -26122 7658 -26070
rect 7710 -26122 7720 -26070
rect 7648 -26126 7720 -26122
rect 8170 -26168 8230 -25964
rect 7144 -26178 7206 -26168
rect 7144 -26180 7150 -26178
rect 7146 -26230 7150 -26180
rect 7202 -26230 7206 -26178
rect 8170 -26178 8232 -26168
rect 8170 -26180 8176 -26178
rect 7146 -26240 7206 -26230
rect 8172 -26230 8176 -26180
rect 8228 -26230 8232 -26178
rect 8172 -26240 8232 -26230
rect 8678 -26430 8738 -25204
rect 9200 -25290 9260 -25094
rect 9692 -25126 9908 -25066
rect 10206 -25038 10278 -25034
rect 10206 -25090 10216 -25038
rect 10268 -25090 10278 -25038
rect 10206 -25094 10278 -25090
rect 9692 -25368 9752 -25126
rect 10212 -25288 10272 -25094
rect 10716 -25144 10776 -24667
rect 11726 -24667 11742 -24634
rect 12794 -24592 12800 -24561
rect 13772 -24163 13778 -24142
rect 13812 -24142 13826 -24129
rect 14780 -24129 14840 -23882
rect 15078 -24026 15566 -24020
rect 15078 -24060 15125 -24026
rect 15159 -24060 15197 -24026
rect 15231 -24060 15269 -24026
rect 15303 -24060 15341 -24026
rect 15375 -24060 15413 -24026
rect 15447 -24060 15485 -24026
rect 15519 -24060 15566 -24026
rect 15078 -24066 15566 -24060
rect 16096 -24026 16584 -24020
rect 16096 -24060 16143 -24026
rect 16177 -24060 16215 -24026
rect 16249 -24060 16287 -24026
rect 16321 -24060 16359 -24026
rect 16393 -24060 16431 -24026
rect 16465 -24060 16503 -24026
rect 16537 -24060 16584 -24026
rect 16096 -24066 16584 -24060
rect 13812 -24163 13818 -24142
rect 14780 -24154 14796 -24129
rect 13772 -24201 13818 -24163
rect 13772 -24235 13778 -24201
rect 13812 -24235 13818 -24201
rect 13772 -24273 13818 -24235
rect 13772 -24307 13778 -24273
rect 13812 -24307 13818 -24273
rect 13772 -24345 13818 -24307
rect 13772 -24379 13778 -24345
rect 13812 -24379 13818 -24345
rect 13772 -24417 13818 -24379
rect 13772 -24451 13778 -24417
rect 13812 -24451 13818 -24417
rect 13772 -24489 13818 -24451
rect 13772 -24523 13778 -24489
rect 13812 -24523 13818 -24489
rect 13772 -24561 13818 -24523
rect 13772 -24592 13778 -24561
rect 12760 -24633 12794 -24595
rect 11776 -24667 11786 -24634
rect 11018 -24770 11053 -24736
rect 11087 -24770 11125 -24736
rect 11159 -24770 11197 -24736
rect 11231 -24770 11269 -24736
rect 11303 -24770 11341 -24736
rect 11375 -24770 11413 -24736
rect 11447 -24770 11482 -24736
rect 11220 -25034 11280 -24770
rect 11726 -24822 11786 -24667
rect 12752 -24667 12760 -24656
rect 13812 -24592 13818 -24561
rect 14790 -24163 14796 -24154
rect 14830 -24154 14840 -24129
rect 15808 -24129 15854 -24098
rect 14830 -24163 14836 -24154
rect 14790 -24201 14836 -24163
rect 14790 -24235 14796 -24201
rect 14830 -24235 14836 -24201
rect 14790 -24273 14836 -24235
rect 14790 -24307 14796 -24273
rect 14830 -24307 14836 -24273
rect 14790 -24345 14836 -24307
rect 14790 -24379 14796 -24345
rect 14830 -24379 14836 -24345
rect 14790 -24417 14836 -24379
rect 14790 -24451 14796 -24417
rect 14830 -24451 14836 -24417
rect 14790 -24489 14836 -24451
rect 14790 -24523 14796 -24489
rect 14830 -24523 14836 -24489
rect 14790 -24561 14836 -24523
rect 14790 -24592 14796 -24561
rect 13778 -24633 13812 -24595
rect 12794 -24667 12812 -24656
rect 12036 -24770 12071 -24736
rect 12105 -24770 12143 -24736
rect 12177 -24770 12215 -24736
rect 12249 -24770 12287 -24736
rect 12321 -24770 12359 -24736
rect 12393 -24770 12431 -24736
rect 12465 -24770 12500 -24736
rect 11720 -24826 11792 -24822
rect 11720 -24878 11730 -24826
rect 11782 -24878 11792 -24826
rect 11720 -24882 11792 -24878
rect 11724 -24932 11796 -24928
rect 11724 -24984 11734 -24932
rect 11786 -24984 11796 -24932
rect 11724 -24988 11796 -24984
rect 11214 -25038 11286 -25034
rect 11214 -25090 11224 -25038
rect 11276 -25090 11286 -25038
rect 11214 -25094 11286 -25090
rect 10710 -25148 10782 -25144
rect 10710 -25200 10720 -25148
rect 10772 -25200 10782 -25148
rect 10710 -25204 10782 -25200
rect 9184 -26178 9244 -25968
rect 9184 -26230 9188 -26178
rect 9240 -26230 9244 -26178
rect 9184 -26240 9244 -26230
rect 10220 -26178 10280 -25972
rect 10220 -26230 10224 -26178
rect 10276 -26230 10280 -26178
rect 10220 -26240 10280 -26230
rect 10716 -26430 10776 -25204
rect 11220 -25290 11280 -25094
rect 11730 -25368 11790 -24988
rect 12238 -25034 12298 -24770
rect 12232 -25038 12304 -25034
rect 12232 -25090 12242 -25038
rect 12294 -25090 12304 -25038
rect 12232 -25094 12304 -25090
rect 12238 -25288 12298 -25094
rect 12752 -25144 12812 -24667
rect 13764 -24667 13778 -24646
rect 14830 -24592 14836 -24561
rect 15808 -24163 15814 -24129
rect 15848 -24163 15854 -24129
rect 16816 -24129 16876 -23882
rect 16962 -23926 17022 -23662
rect 16956 -23930 17028 -23926
rect 16956 -23982 16966 -23930
rect 17018 -23982 17028 -23930
rect 16956 -23986 17028 -23982
rect 17326 -24020 17386 -23542
rect 17838 -23822 17898 -23433
rect 18856 -23433 18868 -23408
rect 18902 -23408 18908 -23399
rect 19880 -22929 19886 -22922
rect 19920 -22922 19930 -22895
rect 20898 -22895 20944 -22864
rect 21910 -22876 21970 -22736
rect 22204 -22792 22410 -22786
rect 22470 -22792 22692 -22786
rect 22204 -22826 22251 -22792
rect 22285 -22826 22323 -22792
rect 22357 -22826 22395 -22792
rect 22429 -22826 22467 -22792
rect 22501 -22826 22539 -22792
rect 22573 -22826 22611 -22792
rect 22645 -22826 22692 -22792
rect 22204 -22832 22692 -22826
rect 19920 -22929 19926 -22922
rect 19880 -22967 19926 -22929
rect 19880 -23001 19886 -22967
rect 19920 -23001 19926 -22967
rect 19880 -23039 19926 -23001
rect 19880 -23073 19886 -23039
rect 19920 -23073 19926 -23039
rect 19880 -23111 19926 -23073
rect 19880 -23145 19886 -23111
rect 19920 -23145 19926 -23111
rect 19880 -23183 19926 -23145
rect 19880 -23217 19886 -23183
rect 19920 -23217 19926 -23183
rect 19880 -23255 19926 -23217
rect 19880 -23289 19886 -23255
rect 19920 -23289 19926 -23255
rect 19880 -23327 19926 -23289
rect 19880 -23361 19886 -23327
rect 19920 -23361 19926 -23327
rect 19880 -23399 19926 -23361
rect 19880 -23404 19886 -23399
rect 18902 -23433 18916 -23408
rect 18132 -23502 18620 -23496
rect 18132 -23536 18179 -23502
rect 18213 -23536 18251 -23502
rect 18285 -23536 18323 -23502
rect 18357 -23536 18395 -23502
rect 18429 -23536 18467 -23502
rect 18501 -23536 18539 -23502
rect 18573 -23536 18620 -23502
rect 18132 -23542 18620 -23536
rect 17832 -23826 17904 -23822
rect 17832 -23878 17842 -23826
rect 17894 -23878 17904 -23826
rect 17832 -23882 17904 -23878
rect 18346 -24020 18406 -23542
rect 18856 -23594 18916 -23433
rect 19872 -23433 19886 -23404
rect 19920 -23404 19926 -23399
rect 20898 -22929 20904 -22895
rect 20938 -22929 20944 -22895
rect 21908 -22895 21970 -22876
rect 21908 -22910 21922 -22895
rect 21910 -22920 21922 -22910
rect 20898 -22967 20944 -22929
rect 20898 -23001 20904 -22967
rect 20938 -23001 20944 -22967
rect 20898 -23039 20944 -23001
rect 20898 -23073 20904 -23039
rect 20938 -23073 20944 -23039
rect 20898 -23111 20944 -23073
rect 20898 -23145 20904 -23111
rect 20938 -23145 20944 -23111
rect 20898 -23183 20944 -23145
rect 20898 -23217 20904 -23183
rect 20938 -23217 20944 -23183
rect 20898 -23255 20944 -23217
rect 20898 -23289 20904 -23255
rect 20938 -23289 20944 -23255
rect 20898 -23327 20944 -23289
rect 20898 -23361 20904 -23327
rect 20938 -23361 20944 -23327
rect 20898 -23399 20944 -23361
rect 19920 -23433 19932 -23404
rect 20898 -23408 20904 -23399
rect 19150 -23502 19638 -23496
rect 19150 -23536 19197 -23502
rect 19231 -23536 19269 -23502
rect 19303 -23536 19341 -23502
rect 19375 -23536 19413 -23502
rect 19447 -23536 19485 -23502
rect 19519 -23536 19557 -23502
rect 19591 -23536 19638 -23502
rect 19150 -23542 19638 -23536
rect 18850 -23598 18922 -23594
rect 18850 -23650 18860 -23598
rect 18912 -23650 18922 -23598
rect 18850 -23654 18922 -23650
rect 18852 -23826 18924 -23822
rect 18852 -23878 18862 -23826
rect 18914 -23878 18924 -23826
rect 18852 -23882 18924 -23878
rect 17114 -24026 17602 -24020
rect 17114 -24060 17161 -24026
rect 17195 -24060 17233 -24026
rect 17267 -24060 17305 -24026
rect 17339 -24060 17377 -24026
rect 17411 -24060 17449 -24026
rect 17483 -24060 17521 -24026
rect 17555 -24060 17602 -24026
rect 17114 -24066 17602 -24060
rect 18132 -24026 18620 -24020
rect 18132 -24060 18179 -24026
rect 18213 -24060 18251 -24026
rect 18285 -24060 18323 -24026
rect 18357 -24060 18395 -24026
rect 18429 -24060 18467 -24026
rect 18501 -24060 18539 -24026
rect 18573 -24060 18620 -24026
rect 18132 -24066 18620 -24060
rect 16816 -24154 16832 -24129
rect 15808 -24201 15854 -24163
rect 15808 -24235 15814 -24201
rect 15848 -24235 15854 -24201
rect 15808 -24273 15854 -24235
rect 15808 -24307 15814 -24273
rect 15848 -24307 15854 -24273
rect 15808 -24345 15854 -24307
rect 15808 -24379 15814 -24345
rect 15848 -24379 15854 -24345
rect 15808 -24417 15854 -24379
rect 15808 -24451 15814 -24417
rect 15848 -24451 15854 -24417
rect 15808 -24489 15854 -24451
rect 15808 -24523 15814 -24489
rect 15848 -24523 15854 -24489
rect 15808 -24561 15854 -24523
rect 15808 -24592 15814 -24561
rect 14796 -24633 14830 -24595
rect 13812 -24667 13824 -24646
rect 13054 -24770 13089 -24736
rect 13123 -24770 13161 -24736
rect 13195 -24770 13233 -24736
rect 13267 -24770 13305 -24736
rect 13339 -24770 13377 -24736
rect 13411 -24770 13449 -24736
rect 13483 -24770 13518 -24736
rect 13264 -25034 13324 -24770
rect 13764 -24822 13824 -24667
rect 14788 -24667 14796 -24662
rect 15848 -24592 15854 -24561
rect 16826 -24163 16832 -24154
rect 16866 -24154 16876 -24129
rect 17844 -24129 17890 -24098
rect 16866 -24163 16872 -24154
rect 16826 -24201 16872 -24163
rect 16826 -24235 16832 -24201
rect 16866 -24235 16872 -24201
rect 16826 -24273 16872 -24235
rect 16826 -24307 16832 -24273
rect 16866 -24307 16872 -24273
rect 16826 -24345 16872 -24307
rect 16826 -24379 16832 -24345
rect 16866 -24379 16872 -24345
rect 16826 -24417 16872 -24379
rect 16826 -24451 16832 -24417
rect 16866 -24451 16872 -24417
rect 16826 -24489 16872 -24451
rect 16826 -24523 16832 -24489
rect 16866 -24523 16872 -24489
rect 16826 -24561 16872 -24523
rect 16826 -24592 16832 -24561
rect 15814 -24633 15848 -24595
rect 14830 -24667 14848 -24662
rect 14072 -24770 14107 -24736
rect 14141 -24770 14179 -24736
rect 14213 -24770 14251 -24736
rect 14285 -24770 14323 -24736
rect 14357 -24770 14395 -24736
rect 14429 -24770 14467 -24736
rect 14501 -24770 14536 -24736
rect 13758 -24826 13830 -24822
rect 13758 -24878 13768 -24826
rect 13820 -24878 13830 -24826
rect 13758 -24882 13830 -24878
rect 13760 -24932 13832 -24928
rect 13760 -24984 13770 -24932
rect 13822 -24984 13832 -24932
rect 13760 -24988 13832 -24984
rect 13258 -25038 13330 -25034
rect 13258 -25090 13268 -25038
rect 13320 -25090 13330 -25038
rect 13258 -25094 13330 -25090
rect 12746 -25148 12818 -25144
rect 12746 -25200 12756 -25148
rect 12808 -25200 12818 -25148
rect 12746 -25204 12818 -25200
rect 11226 -26178 11286 -25972
rect 12240 -26174 12300 -25972
rect 11226 -26230 11230 -26178
rect 11282 -26230 11286 -26178
rect 11226 -26240 11286 -26230
rect 12234 -26178 12306 -26174
rect 12234 -26230 12244 -26178
rect 12296 -26230 12306 -26178
rect 12234 -26234 12306 -26230
rect 12752 -26430 12812 -25204
rect 13264 -25288 13324 -25094
rect 13766 -25378 13826 -24988
rect 14266 -25034 14326 -24770
rect 14260 -25038 14332 -25034
rect 14260 -25090 14270 -25038
rect 14322 -25090 14332 -25038
rect 14260 -25094 14332 -25090
rect 14266 -25290 14326 -25094
rect 14788 -25144 14848 -24667
rect 15800 -24667 15814 -24640
rect 16866 -24592 16872 -24561
rect 17844 -24163 17850 -24129
rect 17884 -24163 17890 -24129
rect 17844 -24201 17890 -24163
rect 18858 -24129 18918 -23882
rect 19360 -24020 19420 -23542
rect 19872 -23822 19932 -23433
rect 20888 -23433 20904 -23408
rect 20938 -23408 20944 -23399
rect 21916 -22929 21922 -22920
rect 21956 -22920 21970 -22895
rect 22922 -22876 22982 -22608
rect 22922 -22895 22986 -22876
rect 21956 -22929 21962 -22920
rect 21916 -22967 21962 -22929
rect 22922 -22929 22940 -22895
rect 22974 -22914 22986 -22895
rect 22974 -22929 22982 -22914
rect 22922 -22930 22982 -22929
rect 21916 -23001 21922 -22967
rect 21956 -23001 21962 -22967
rect 21916 -23039 21962 -23001
rect 21916 -23073 21922 -23039
rect 21956 -23073 21962 -23039
rect 21916 -23111 21962 -23073
rect 21916 -23145 21922 -23111
rect 21956 -23145 21962 -23111
rect 21916 -23183 21962 -23145
rect 21916 -23217 21922 -23183
rect 21956 -23217 21962 -23183
rect 21916 -23255 21962 -23217
rect 21916 -23289 21922 -23255
rect 21956 -23289 21962 -23255
rect 21916 -23327 21962 -23289
rect 21916 -23361 21922 -23327
rect 21956 -23361 21962 -23327
rect 21916 -23399 21962 -23361
rect 20938 -23433 20948 -23408
rect 20168 -23502 20656 -23496
rect 20168 -23536 20215 -23502
rect 20249 -23536 20287 -23502
rect 20321 -23536 20359 -23502
rect 20393 -23536 20431 -23502
rect 20465 -23536 20503 -23502
rect 20537 -23536 20575 -23502
rect 20609 -23536 20656 -23502
rect 20168 -23542 20656 -23536
rect 19866 -23826 19938 -23822
rect 19866 -23878 19876 -23826
rect 19928 -23878 19938 -23826
rect 19866 -23882 19938 -23878
rect 19866 -23930 19938 -23926
rect 19866 -23982 19876 -23930
rect 19928 -23982 19938 -23930
rect 19866 -23986 19938 -23982
rect 19150 -24026 19420 -24020
rect 19428 -24026 19638 -24020
rect 19150 -24060 19197 -24026
rect 19231 -24060 19269 -24026
rect 19303 -24060 19341 -24026
rect 19375 -24060 19413 -24026
rect 19447 -24060 19485 -24026
rect 19519 -24060 19557 -24026
rect 19591 -24060 19638 -24026
rect 19150 -24066 19638 -24060
rect 19368 -24070 19428 -24066
rect 18858 -24163 18868 -24129
rect 18902 -24163 18918 -24129
rect 19872 -24129 19932 -23986
rect 20396 -24020 20456 -23542
rect 20888 -23594 20948 -23433
rect 21916 -23433 21922 -23399
rect 21956 -23433 21962 -23399
rect 21916 -23464 21962 -23433
rect 22934 -22967 22980 -22930
rect 22934 -23001 22940 -22967
rect 22974 -23001 22980 -22967
rect 22934 -23039 22980 -23001
rect 22934 -23073 22940 -23039
rect 22974 -23073 22980 -23039
rect 22934 -23111 22980 -23073
rect 22934 -23145 22940 -23111
rect 22974 -23145 22980 -23111
rect 22934 -23183 22980 -23145
rect 22934 -23217 22940 -23183
rect 22974 -23217 22980 -23183
rect 22934 -23255 22980 -23217
rect 22934 -23289 22940 -23255
rect 22974 -23289 22980 -23255
rect 22934 -23327 22980 -23289
rect 22934 -23361 22940 -23327
rect 22974 -23361 22980 -23327
rect 22934 -23399 22980 -23361
rect 22934 -23433 22940 -23399
rect 22974 -23433 22980 -23399
rect 22934 -23464 22980 -23433
rect 21186 -23502 21674 -23496
rect 21186 -23536 21233 -23502
rect 21267 -23536 21305 -23502
rect 21339 -23536 21377 -23502
rect 21411 -23536 21449 -23502
rect 21483 -23536 21521 -23502
rect 21555 -23536 21593 -23502
rect 21627 -23536 21674 -23502
rect 21186 -23542 21674 -23536
rect 22204 -23502 22692 -23496
rect 22204 -23536 22251 -23502
rect 22285 -23536 22323 -23502
rect 22357 -23536 22395 -23502
rect 22429 -23536 22467 -23502
rect 22501 -23536 22539 -23502
rect 22573 -23536 22611 -23502
rect 22645 -23536 22692 -23502
rect 22204 -23542 22692 -23536
rect 20882 -23598 20954 -23594
rect 20882 -23650 20892 -23598
rect 20944 -23650 20954 -23598
rect 20882 -23654 20954 -23650
rect 21408 -23704 21468 -23542
rect 22416 -23704 22476 -23542
rect 23034 -23594 23094 -17804
rect 23156 -18662 23228 -18658
rect 23156 -18714 23166 -18662
rect 23218 -18714 23228 -18662
rect 23156 -18718 23228 -18714
rect 23162 -20216 23222 -18718
rect 23278 -18982 23338 -17690
rect 23394 -18884 23466 -18880
rect 23394 -18936 23404 -18884
rect 23456 -18936 23466 -18884
rect 23394 -18940 23466 -18936
rect 23272 -18986 23344 -18982
rect 23272 -19038 23282 -18986
rect 23334 -19038 23344 -18986
rect 23272 -19042 23344 -19038
rect 23156 -20220 23228 -20216
rect 23156 -20272 23166 -20220
rect 23218 -20272 23228 -20220
rect 23156 -20276 23228 -20272
rect 23152 -21122 23224 -21118
rect 23152 -21174 23162 -21122
rect 23214 -21174 23224 -21122
rect 23152 -21178 23224 -21174
rect 23158 -22442 23218 -21178
rect 23278 -22344 23338 -19042
rect 23272 -22348 23344 -22344
rect 23272 -22400 23282 -22348
rect 23334 -22400 23344 -22348
rect 23272 -22404 23344 -22400
rect 23152 -22446 23224 -22442
rect 23152 -22498 23162 -22446
rect 23214 -22498 23224 -22446
rect 23152 -22502 23224 -22498
rect 23028 -23598 23100 -23594
rect 23028 -23650 23038 -23598
rect 23090 -23650 23100 -23598
rect 23028 -23654 23100 -23650
rect 21402 -23708 21474 -23704
rect 21402 -23760 21412 -23708
rect 21464 -23760 21474 -23708
rect 21402 -23764 21474 -23760
rect 22410 -23708 22482 -23704
rect 22410 -23760 22420 -23708
rect 22472 -23760 22482 -23708
rect 22410 -23764 22482 -23760
rect 23278 -23820 23338 -22404
rect 23400 -22676 23460 -18940
rect 23528 -20108 23588 -17586
rect 23526 -20118 23588 -20108
rect 23526 -20170 23530 -20118
rect 23582 -20170 23588 -20118
rect 23526 -20180 23588 -20170
rect 23528 -22548 23588 -20180
rect 23522 -22552 23594 -22548
rect 23522 -22604 23532 -22552
rect 23584 -22604 23594 -22552
rect 23522 -22608 23594 -22604
rect 23394 -22680 23466 -22676
rect 23394 -22732 23404 -22680
rect 23456 -22732 23466 -22680
rect 23394 -22736 23466 -22732
rect 23650 -23704 23710 -12776
rect 24816 -12739 24928 -12701
rect 24816 -12773 24855 -12739
rect 24889 -12773 24928 -12739
rect 24816 -12811 24928 -12773
rect 24816 -12845 24855 -12811
rect 24889 -12845 24928 -12811
rect 24816 -12883 24928 -12845
rect 24816 -12917 24855 -12883
rect 24889 -12917 24928 -12883
rect 24816 -12955 24928 -12917
rect 24816 -12989 24855 -12955
rect 24889 -12989 24928 -12955
rect 24816 -13027 24928 -12989
rect 24816 -13061 24855 -13027
rect 24889 -13061 24928 -13027
rect 24816 -13099 24928 -13061
rect 24816 -13133 24855 -13099
rect 24889 -13133 24928 -13099
rect 24816 -13171 24928 -13133
rect 24816 -13205 24855 -13171
rect 24889 -13205 24928 -13171
rect 24816 -13243 24928 -13205
rect 24816 -13277 24855 -13243
rect 24889 -13277 24928 -13243
rect 24816 -13315 24928 -13277
rect 24816 -13349 24855 -13315
rect 24889 -13349 24928 -13315
rect 24816 -13387 24928 -13349
rect 24816 -13421 24855 -13387
rect 24889 -13421 24928 -13387
rect 24816 -13459 24928 -13421
rect 24816 -13493 24855 -13459
rect 24889 -13493 24928 -13459
rect 24816 -13531 24928 -13493
rect 24816 -13565 24855 -13531
rect 24889 -13565 24928 -13531
rect 24816 -13603 24928 -13565
rect 24816 -13637 24855 -13603
rect 24889 -13637 24928 -13603
rect 24816 -13675 24928 -13637
rect 24816 -13709 24855 -13675
rect 24889 -13709 24928 -13675
rect 24816 -13747 24928 -13709
rect 24816 -13781 24855 -13747
rect 24889 -13781 24928 -13747
rect 24816 -13819 24928 -13781
rect 24816 -13853 24855 -13819
rect 24889 -13853 24928 -13819
rect 24816 -13891 24928 -13853
rect 24816 -13925 24855 -13891
rect 24889 -13925 24928 -13891
rect 24816 -13963 24928 -13925
rect 24816 -13997 24855 -13963
rect 24889 -13997 24928 -13963
rect 24816 -14035 24928 -13997
rect 24816 -14069 24855 -14035
rect 24889 -14069 24928 -14035
rect 24816 -14107 24928 -14069
rect 24816 -14141 24855 -14107
rect 24889 -14141 24928 -14107
rect 24816 -14179 24928 -14141
rect 24816 -14213 24855 -14179
rect 24889 -14213 24928 -14179
rect 24816 -14251 24928 -14213
rect 24816 -14285 24855 -14251
rect 24889 -14285 24928 -14251
rect 24816 -14323 24928 -14285
rect 24816 -14357 24855 -14323
rect 24889 -14357 24928 -14323
rect 24816 -14395 24928 -14357
rect 24816 -14429 24855 -14395
rect 24889 -14429 24928 -14395
rect 24816 -14467 24928 -14429
rect 24816 -14501 24855 -14467
rect 24889 -14501 24928 -14467
rect 24816 -14539 24928 -14501
rect 24816 -14573 24855 -14539
rect 24889 -14573 24928 -14539
rect 24816 -14611 24928 -14573
rect 24816 -14645 24855 -14611
rect 24889 -14645 24928 -14611
rect 24816 -14683 24928 -14645
rect 24816 -14717 24855 -14683
rect 24889 -14717 24928 -14683
rect 24816 -14755 24928 -14717
rect 24816 -14789 24855 -14755
rect 24889 -14789 24928 -14755
rect 24816 -14827 24928 -14789
rect 24816 -14861 24855 -14827
rect 24889 -14861 24928 -14827
rect 24816 -14899 24928 -14861
rect 24816 -14933 24855 -14899
rect 24889 -14933 24928 -14899
rect 24816 -14971 24928 -14933
rect 24816 -15005 24855 -14971
rect 24889 -15005 24928 -14971
rect 24816 -15043 24928 -15005
rect 24816 -15077 24855 -15043
rect 24889 -15077 24928 -15043
rect 24816 -15115 24928 -15077
rect 24816 -15149 24855 -15115
rect 24889 -15149 24928 -15115
rect 24816 -15187 24928 -15149
rect 24816 -15221 24855 -15187
rect 24889 -15221 24928 -15187
rect 24816 -15259 24928 -15221
rect 24816 -15293 24855 -15259
rect 24889 -15293 24928 -15259
rect 24816 -15331 24928 -15293
rect 24816 -15365 24855 -15331
rect 24889 -15365 24928 -15331
rect 24816 -15403 24928 -15365
rect 24816 -15437 24855 -15403
rect 24889 -15437 24928 -15403
rect 24816 -15475 24928 -15437
rect 24816 -15509 24855 -15475
rect 24889 -15509 24928 -15475
rect 24816 -15547 24928 -15509
rect 24816 -15581 24855 -15547
rect 24889 -15581 24928 -15547
rect 24816 -15619 24928 -15581
rect 24816 -15653 24855 -15619
rect 24889 -15653 24928 -15619
rect 24816 -15691 24928 -15653
rect 24816 -15725 24855 -15691
rect 24889 -15725 24928 -15691
rect 24816 -15763 24928 -15725
rect 24816 -15797 24855 -15763
rect 24889 -15797 24928 -15763
rect 24816 -15835 24928 -15797
rect 24816 -15869 24855 -15835
rect 24889 -15869 24928 -15835
rect 24816 -15907 24928 -15869
rect 24816 -15941 24855 -15907
rect 24889 -15941 24928 -15907
rect 24816 -15979 24928 -15941
rect 24816 -16013 24855 -15979
rect 24889 -16013 24928 -15979
rect 24816 -16051 24928 -16013
rect 24816 -16085 24855 -16051
rect 24889 -16085 24928 -16051
rect 24816 -16123 24928 -16085
rect 24816 -16157 24855 -16123
rect 24889 -16157 24928 -16123
rect 24816 -16195 24928 -16157
rect 24816 -16229 24855 -16195
rect 24889 -16229 24928 -16195
rect 24816 -16267 24928 -16229
rect 24816 -16301 24855 -16267
rect 24889 -16301 24928 -16267
rect 24816 -16339 24928 -16301
rect 24816 -16373 24855 -16339
rect 24889 -16373 24928 -16339
rect 24816 -16411 24928 -16373
rect 24816 -16445 24855 -16411
rect 24889 -16445 24928 -16411
rect 24816 -16483 24928 -16445
rect 24816 -16517 24855 -16483
rect 24889 -16517 24928 -16483
rect 23756 -16530 23828 -16526
rect 23756 -16582 23766 -16530
rect 23818 -16582 23828 -16530
rect 23756 -16586 23828 -16582
rect 24816 -16555 24928 -16517
rect 23644 -23708 23716 -23704
rect 23644 -23760 23654 -23708
rect 23706 -23760 23716 -23708
rect 23644 -23764 23716 -23760
rect 20888 -23826 20960 -23822
rect 20888 -23878 20898 -23826
rect 20950 -23878 20960 -23826
rect 20888 -23882 20960 -23878
rect 21910 -23880 23338 -23820
rect 20168 -24026 20656 -24020
rect 20168 -24060 20215 -24026
rect 20249 -24060 20287 -24026
rect 20321 -24060 20359 -24026
rect 20393 -24060 20431 -24026
rect 20465 -24060 20503 -24026
rect 20537 -24060 20575 -24026
rect 20609 -24060 20656 -24026
rect 20168 -24066 20656 -24060
rect 19872 -24156 19886 -24129
rect 18858 -24176 18918 -24163
rect 19880 -24163 19886 -24156
rect 19920 -24156 19932 -24129
rect 20894 -24129 20954 -23882
rect 21186 -24026 21408 -24020
rect 21468 -24026 21674 -24020
rect 21186 -24060 21233 -24026
rect 21267 -24060 21305 -24026
rect 21339 -24060 21377 -24026
rect 21411 -24060 21449 -24026
rect 21483 -24060 21521 -24026
rect 21555 -24060 21593 -24026
rect 21627 -24060 21674 -24026
rect 21186 -24066 21674 -24060
rect 19920 -24163 19926 -24156
rect 17844 -24235 17850 -24201
rect 17884 -24235 17890 -24201
rect 17844 -24273 17890 -24235
rect 17844 -24307 17850 -24273
rect 17884 -24307 17890 -24273
rect 17844 -24345 17890 -24307
rect 17844 -24379 17850 -24345
rect 17884 -24379 17890 -24345
rect 17844 -24417 17890 -24379
rect 17844 -24451 17850 -24417
rect 17884 -24451 17890 -24417
rect 17844 -24489 17890 -24451
rect 17844 -24523 17850 -24489
rect 17884 -24523 17890 -24489
rect 17844 -24561 17890 -24523
rect 17844 -24592 17850 -24561
rect 16832 -24633 16866 -24595
rect 15848 -24667 15860 -24640
rect 15090 -24770 15125 -24736
rect 15159 -24770 15197 -24736
rect 15231 -24770 15269 -24736
rect 15303 -24770 15341 -24736
rect 15375 -24770 15413 -24736
rect 15447 -24770 15485 -24736
rect 15519 -24770 15554 -24736
rect 15286 -25034 15346 -24770
rect 15628 -24826 15700 -24822
rect 15628 -24878 15638 -24826
rect 15690 -24878 15700 -24826
rect 15628 -24882 15700 -24878
rect 15280 -25038 15352 -25034
rect 15280 -25090 15290 -25038
rect 15342 -25090 15352 -25038
rect 15280 -25094 15352 -25090
rect 15634 -25074 15694 -24882
rect 15800 -24928 15860 -24667
rect 16820 -24667 16832 -24660
rect 17884 -24592 17890 -24561
rect 18862 -24201 18908 -24176
rect 18862 -24235 18868 -24201
rect 18902 -24235 18908 -24201
rect 18862 -24273 18908 -24235
rect 18862 -24307 18868 -24273
rect 18902 -24307 18908 -24273
rect 18862 -24345 18908 -24307
rect 18862 -24379 18868 -24345
rect 18902 -24379 18908 -24345
rect 18862 -24417 18908 -24379
rect 18862 -24451 18868 -24417
rect 18902 -24451 18908 -24417
rect 18862 -24489 18908 -24451
rect 18862 -24523 18868 -24489
rect 18902 -24523 18908 -24489
rect 18862 -24561 18908 -24523
rect 18862 -24592 18868 -24561
rect 17850 -24633 17884 -24595
rect 16866 -24667 16880 -24660
rect 16108 -24770 16143 -24736
rect 16177 -24770 16215 -24736
rect 16249 -24770 16287 -24736
rect 16321 -24770 16359 -24736
rect 16393 -24770 16431 -24736
rect 16465 -24770 16503 -24736
rect 16537 -24770 16572 -24736
rect 15794 -24932 15866 -24928
rect 15794 -24984 15804 -24932
rect 15856 -24984 15866 -24932
rect 15794 -24988 15866 -24984
rect 16306 -25034 16366 -24770
rect 16300 -25038 16372 -25034
rect 14782 -25148 14854 -25144
rect 14782 -25200 14792 -25148
rect 14844 -25200 14854 -25148
rect 14782 -25204 14854 -25200
rect 13256 -26178 13316 -25968
rect 14266 -26168 14326 -25972
rect 13256 -26230 13260 -26178
rect 13312 -26230 13316 -26178
rect 13256 -26240 13316 -26230
rect 14264 -26178 14326 -26168
rect 14264 -26230 14268 -26178
rect 14320 -26180 14326 -26178
rect 14320 -26230 14324 -26180
rect 14264 -26240 14324 -26230
rect 14788 -26430 14848 -25204
rect 15286 -25288 15346 -25094
rect 15634 -25134 15860 -25074
rect 16300 -25090 16310 -25038
rect 16362 -25090 16372 -25038
rect 16300 -25094 16372 -25090
rect 15800 -25378 15860 -25134
rect 16306 -25288 16366 -25094
rect 16820 -25144 16880 -24667
rect 17840 -24667 17850 -24646
rect 18902 -24592 18908 -24561
rect 19880 -24201 19926 -24163
rect 20894 -24163 20904 -24129
rect 20938 -24163 20954 -24129
rect 20894 -24170 20954 -24163
rect 21910 -24129 21970 -23880
rect 22408 -24020 22468 -23880
rect 22204 -24026 22692 -24020
rect 22204 -24060 22251 -24026
rect 22285 -24060 22323 -24026
rect 22357 -24060 22395 -24026
rect 22429 -24060 22467 -24026
rect 22501 -24060 22539 -24026
rect 22573 -24060 22611 -24026
rect 22645 -24060 22692 -24026
rect 22204 -24066 22692 -24060
rect 21910 -24163 21922 -24129
rect 21956 -24163 21970 -24129
rect 19880 -24235 19886 -24201
rect 19920 -24235 19926 -24201
rect 19880 -24273 19926 -24235
rect 19880 -24307 19886 -24273
rect 19920 -24307 19926 -24273
rect 19880 -24345 19926 -24307
rect 19880 -24379 19886 -24345
rect 19920 -24379 19926 -24345
rect 19880 -24417 19926 -24379
rect 19880 -24451 19886 -24417
rect 19920 -24451 19926 -24417
rect 19880 -24489 19926 -24451
rect 19880 -24523 19886 -24489
rect 19920 -24523 19926 -24489
rect 19880 -24561 19926 -24523
rect 19880 -24592 19886 -24561
rect 18868 -24633 18902 -24595
rect 17884 -24667 17900 -24646
rect 17126 -24770 17161 -24736
rect 17195 -24770 17233 -24736
rect 17267 -24770 17305 -24736
rect 17339 -24770 17377 -24736
rect 17411 -24770 17449 -24736
rect 17483 -24770 17521 -24736
rect 17555 -24770 17590 -24736
rect 17332 -25034 17392 -24770
rect 17840 -24928 17900 -24667
rect 18852 -24667 18868 -24640
rect 19920 -24592 19926 -24561
rect 20898 -24201 20944 -24170
rect 20898 -24235 20904 -24201
rect 20938 -24235 20944 -24201
rect 20898 -24273 20944 -24235
rect 20898 -24307 20904 -24273
rect 20938 -24307 20944 -24273
rect 20898 -24345 20944 -24307
rect 20898 -24379 20904 -24345
rect 20938 -24379 20944 -24345
rect 20898 -24417 20944 -24379
rect 20898 -24451 20904 -24417
rect 20938 -24451 20944 -24417
rect 20898 -24489 20944 -24451
rect 20898 -24523 20904 -24489
rect 20938 -24523 20944 -24489
rect 20898 -24561 20944 -24523
rect 20898 -24592 20904 -24561
rect 19886 -24633 19920 -24595
rect 18902 -24667 18912 -24640
rect 18350 -24736 18410 -24734
rect 18144 -24770 18179 -24736
rect 18213 -24770 18251 -24736
rect 18285 -24770 18323 -24736
rect 18357 -24770 18395 -24736
rect 18429 -24770 18467 -24736
rect 18501 -24770 18539 -24736
rect 18573 -24770 18608 -24736
rect 17834 -24932 17906 -24928
rect 17834 -24984 17844 -24932
rect 17896 -24984 17906 -24932
rect 17834 -24988 17906 -24984
rect 18350 -25034 18410 -24770
rect 17326 -25038 17398 -25034
rect 17326 -25090 17336 -25038
rect 17388 -25090 17398 -25038
rect 17326 -25094 17398 -25090
rect 18344 -25038 18416 -25034
rect 18344 -25090 18354 -25038
rect 18406 -25090 18416 -25038
rect 18344 -25094 18416 -25090
rect 16814 -25148 16886 -25144
rect 16814 -25200 16824 -25148
rect 16876 -25200 16886 -25148
rect 16814 -25204 16886 -25200
rect 15282 -26168 15342 -25972
rect 15280 -26178 15342 -26168
rect 15280 -26230 15284 -26178
rect 15336 -26180 15342 -26178
rect 16304 -26178 16364 -25960
rect 15336 -26230 15340 -26180
rect 15280 -26240 15340 -26230
rect 16304 -26230 16308 -26178
rect 16360 -26230 16364 -26178
rect 16304 -26240 16364 -26230
rect 16820 -26430 16880 -25204
rect 17332 -25294 17392 -25094
rect 18350 -25294 18410 -25094
rect 18852 -25144 18912 -24667
rect 20938 -24592 20944 -24561
rect 21910 -24201 21970 -24163
rect 22924 -24129 22984 -23880
rect 23048 -23930 23120 -23926
rect 23048 -23982 23058 -23930
rect 23110 -23982 23120 -23930
rect 23048 -23986 23120 -23982
rect 22924 -24163 22940 -24129
rect 22974 -24163 22984 -24129
rect 22924 -24164 22984 -24163
rect 21910 -24235 21922 -24201
rect 21956 -24235 21970 -24201
rect 21910 -24273 21970 -24235
rect 21910 -24307 21922 -24273
rect 21956 -24307 21970 -24273
rect 21910 -24345 21970 -24307
rect 21910 -24379 21922 -24345
rect 21956 -24379 21970 -24345
rect 21910 -24417 21970 -24379
rect 21910 -24451 21922 -24417
rect 21956 -24451 21970 -24417
rect 21910 -24489 21970 -24451
rect 21910 -24523 21922 -24489
rect 21956 -24523 21970 -24489
rect 21910 -24561 21970 -24523
rect 20904 -24633 20938 -24595
rect 19886 -24686 19920 -24667
rect 20892 -24667 20904 -24662
rect 21910 -24595 21922 -24561
rect 21956 -24595 21970 -24561
rect 22934 -24201 22980 -24164
rect 22934 -24235 22940 -24201
rect 22974 -24235 22980 -24201
rect 22934 -24273 22980 -24235
rect 22934 -24307 22940 -24273
rect 22974 -24307 22980 -24273
rect 22934 -24345 22980 -24307
rect 22934 -24379 22940 -24345
rect 22974 -24379 22980 -24345
rect 22934 -24417 22980 -24379
rect 22934 -24451 22940 -24417
rect 22974 -24451 22980 -24417
rect 22934 -24489 22980 -24451
rect 22934 -24523 22940 -24489
rect 22974 -24523 22980 -24489
rect 22934 -24561 22980 -24523
rect 22934 -24592 22940 -24561
rect 21910 -24633 21970 -24595
rect 20938 -24667 20952 -24662
rect 19162 -24770 19197 -24736
rect 19231 -24770 19269 -24736
rect 19303 -24770 19341 -24736
rect 19375 -24770 19413 -24736
rect 19447 -24770 19485 -24736
rect 19519 -24770 19557 -24736
rect 19591 -24770 19626 -24736
rect 20180 -24770 20215 -24736
rect 20249 -24770 20287 -24736
rect 20321 -24770 20359 -24736
rect 20393 -24770 20431 -24736
rect 20465 -24770 20503 -24736
rect 20537 -24770 20575 -24736
rect 20609 -24770 20644 -24736
rect 19364 -25034 19424 -24770
rect 19864 -24932 19936 -24928
rect 19864 -24984 19874 -24932
rect 19926 -24984 19936 -24932
rect 19864 -24988 19936 -24984
rect 19358 -25038 19430 -25034
rect 19358 -25090 19368 -25038
rect 19420 -25090 19430 -25038
rect 19358 -25094 19430 -25090
rect 18846 -25148 18918 -25144
rect 18846 -25200 18856 -25148
rect 18908 -25200 18918 -25148
rect 18846 -25204 18918 -25200
rect 17326 -26178 17386 -25964
rect 17834 -26066 17894 -25866
rect 17828 -26070 17900 -26066
rect 17828 -26122 17838 -26070
rect 17890 -26122 17900 -26070
rect 17828 -26126 17900 -26122
rect 17326 -26230 17330 -26178
rect 17382 -26230 17386 -26178
rect 18346 -26168 18406 -25972
rect 18346 -26178 18408 -26168
rect 18346 -26180 18352 -26178
rect 17326 -26240 17386 -26230
rect 18348 -26230 18352 -26180
rect 18404 -26230 18408 -26178
rect 18348 -26240 18408 -26230
rect 18852 -26430 18912 -25204
rect 19364 -25284 19424 -25094
rect 19870 -25386 19930 -24988
rect 20378 -25034 20438 -24770
rect 20372 -25038 20444 -25034
rect 20372 -25090 20382 -25038
rect 20434 -25090 20444 -25038
rect 20372 -25094 20444 -25090
rect 20378 -25284 20438 -25094
rect 20892 -25144 20952 -24667
rect 21910 -24667 21922 -24633
rect 21956 -24667 21970 -24633
rect 21400 -24736 21460 -24734
rect 21198 -24770 21233 -24736
rect 21267 -24770 21305 -24736
rect 21339 -24770 21377 -24736
rect 21411 -24770 21449 -24736
rect 21483 -24770 21521 -24736
rect 21555 -24770 21593 -24736
rect 21627 -24770 21662 -24736
rect 21400 -25034 21460 -24770
rect 21910 -24822 21970 -24667
rect 22974 -24592 22980 -24561
rect 22940 -24633 22974 -24595
rect 22940 -24686 22974 -24667
rect 22216 -24770 22251 -24736
rect 22285 -24770 22323 -24736
rect 22357 -24770 22395 -24736
rect 22429 -24770 22467 -24736
rect 22501 -24770 22539 -24736
rect 22573 -24770 22611 -24736
rect 22645 -24770 22680 -24736
rect 21904 -24826 21976 -24822
rect 21904 -24878 21914 -24826
rect 21966 -24878 21976 -24826
rect 21904 -24882 21976 -24878
rect 21904 -24932 21976 -24928
rect 21904 -24984 21914 -24932
rect 21966 -24984 21976 -24932
rect 21904 -24988 21976 -24984
rect 21394 -25038 21466 -25034
rect 21394 -25090 21404 -25038
rect 21456 -25090 21466 -25038
rect 21394 -25094 21466 -25090
rect 20886 -25148 20958 -25144
rect 20886 -25200 20896 -25148
rect 20948 -25200 20958 -25148
rect 20886 -25204 20958 -25200
rect 19368 -26168 19428 -25960
rect 20382 -26168 20442 -25968
rect 19366 -26178 19428 -26168
rect 19366 -26230 19370 -26178
rect 19422 -26180 19428 -26178
rect 20380 -26178 20442 -26168
rect 19422 -26230 19426 -26180
rect 19366 -26240 19426 -26230
rect 20380 -26230 20384 -26178
rect 20436 -26180 20442 -26178
rect 20436 -26230 20440 -26180
rect 20380 -26240 20440 -26230
rect 20892 -26430 20952 -25204
rect 21400 -25284 21460 -25094
rect 21910 -25144 21970 -24988
rect 21910 -25204 22988 -25144
rect 21910 -25350 21970 -25204
rect 22426 -25294 22486 -25204
rect 22928 -25360 22988 -25204
rect 21402 -26168 21462 -25960
rect 23054 -26066 23114 -23986
rect 23762 -24928 23822 -16586
rect 24816 -16589 24855 -16555
rect 24889 -16589 24928 -16555
rect 24816 -16627 24928 -16589
rect 24816 -16661 24855 -16627
rect 24889 -16661 24928 -16627
rect 24816 -16699 24928 -16661
rect 24816 -16733 24855 -16699
rect 24889 -16733 24928 -16699
rect 24816 -16771 24928 -16733
rect 24816 -16805 24855 -16771
rect 24889 -16805 24928 -16771
rect 24816 -16843 24928 -16805
rect 24816 -16877 24855 -16843
rect 24889 -16877 24928 -16843
rect 24816 -16915 24928 -16877
rect 24816 -16949 24855 -16915
rect 24889 -16949 24928 -16915
rect 24816 -16987 24928 -16949
rect 24816 -17021 24855 -16987
rect 24889 -17021 24928 -16987
rect 24816 -17059 24928 -17021
rect 24816 -17093 24855 -17059
rect 24889 -17093 24928 -17059
rect 24816 -17131 24928 -17093
rect 24816 -17165 24855 -17131
rect 24889 -17165 24928 -17131
rect 24816 -17203 24928 -17165
rect 24816 -17237 24855 -17203
rect 24889 -17237 24928 -17203
rect 24816 -17275 24928 -17237
rect 24816 -17309 24855 -17275
rect 24889 -17309 24928 -17275
rect 24816 -17347 24928 -17309
rect 24816 -17381 24855 -17347
rect 24889 -17381 24928 -17347
rect 24816 -17419 24928 -17381
rect 24816 -17453 24855 -17419
rect 24889 -17453 24928 -17419
rect 24816 -17491 24928 -17453
rect 24816 -17525 24855 -17491
rect 24889 -17525 24928 -17491
rect 24816 -17563 24928 -17525
rect 24816 -17597 24855 -17563
rect 24889 -17597 24928 -17563
rect 24816 -17635 24928 -17597
rect 24816 -17669 24855 -17635
rect 24889 -17669 24928 -17635
rect 24816 -17707 24928 -17669
rect 24816 -17741 24855 -17707
rect 24889 -17741 24928 -17707
rect 24816 -17779 24928 -17741
rect 24816 -17813 24855 -17779
rect 24889 -17813 24928 -17779
rect 24816 -17851 24928 -17813
rect 24816 -17885 24855 -17851
rect 24889 -17885 24928 -17851
rect 24816 -17923 24928 -17885
rect 24816 -17957 24855 -17923
rect 24889 -17957 24928 -17923
rect 24816 -17995 24928 -17957
rect 24816 -18029 24855 -17995
rect 24889 -18029 24928 -17995
rect 24816 -18067 24928 -18029
rect 24816 -18101 24855 -18067
rect 24889 -18101 24928 -18067
rect 24816 -18139 24928 -18101
rect 24816 -18173 24855 -18139
rect 24889 -18173 24928 -18139
rect 24816 -18211 24928 -18173
rect 24816 -18245 24855 -18211
rect 24889 -18245 24928 -18211
rect 24816 -18283 24928 -18245
rect 24816 -18317 24855 -18283
rect 24889 -18317 24928 -18283
rect 24816 -18355 24928 -18317
rect 24816 -18389 24855 -18355
rect 24889 -18389 24928 -18355
rect 24816 -18427 24928 -18389
rect 24816 -18461 24855 -18427
rect 24889 -18461 24928 -18427
rect 24816 -18499 24928 -18461
rect 24816 -18533 24855 -18499
rect 24889 -18533 24928 -18499
rect 24816 -18571 24928 -18533
rect 24816 -18605 24855 -18571
rect 24889 -18605 24928 -18571
rect 24816 -18643 24928 -18605
rect 24816 -18677 24855 -18643
rect 24889 -18677 24928 -18643
rect 24816 -18715 24928 -18677
rect 24816 -18749 24855 -18715
rect 24889 -18749 24928 -18715
rect 24816 -18787 24928 -18749
rect 24816 -18821 24855 -18787
rect 24889 -18821 24928 -18787
rect 24816 -18859 24928 -18821
rect 24816 -18893 24855 -18859
rect 24889 -18893 24928 -18859
rect 24816 -18931 24928 -18893
rect 24816 -18965 24855 -18931
rect 24889 -18965 24928 -18931
rect 24816 -19003 24928 -18965
rect 24816 -19037 24855 -19003
rect 24889 -19037 24928 -19003
rect 24816 -19075 24928 -19037
rect 24816 -19109 24855 -19075
rect 24889 -19109 24928 -19075
rect 24816 -19147 24928 -19109
rect 24816 -19181 24855 -19147
rect 24889 -19181 24928 -19147
rect 24816 -19219 24928 -19181
rect 24816 -19253 24855 -19219
rect 24889 -19253 24928 -19219
rect 24816 -19291 24928 -19253
rect 24816 -19325 24855 -19291
rect 24889 -19325 24928 -19291
rect 24816 -19363 24928 -19325
rect 24816 -19397 24855 -19363
rect 24889 -19397 24928 -19363
rect 24816 -19435 24928 -19397
rect 24816 -19469 24855 -19435
rect 24889 -19469 24928 -19435
rect 24816 -19507 24928 -19469
rect 24816 -19541 24855 -19507
rect 24889 -19541 24928 -19507
rect 24816 -19579 24928 -19541
rect 24816 -19613 24855 -19579
rect 24889 -19613 24928 -19579
rect 24816 -19651 24928 -19613
rect 24816 -19685 24855 -19651
rect 24889 -19685 24928 -19651
rect 24816 -19723 24928 -19685
rect 24816 -19757 24855 -19723
rect 24889 -19757 24928 -19723
rect 24816 -19795 24928 -19757
rect 24816 -19829 24855 -19795
rect 24889 -19829 24928 -19795
rect 24816 -19867 24928 -19829
rect 24816 -19901 24855 -19867
rect 24889 -19901 24928 -19867
rect 24816 -19939 24928 -19901
rect 24816 -19973 24855 -19939
rect 24889 -19973 24928 -19939
rect 24816 -20011 24928 -19973
rect 24816 -20045 24855 -20011
rect 24889 -20045 24928 -20011
rect 24816 -20083 24928 -20045
rect 24816 -20117 24855 -20083
rect 24889 -20117 24928 -20083
rect 24816 -20155 24928 -20117
rect 24816 -20189 24855 -20155
rect 24889 -20189 24928 -20155
rect 24816 -20227 24928 -20189
rect 24816 -20261 24855 -20227
rect 24889 -20261 24928 -20227
rect 24816 -20299 24928 -20261
rect 24816 -20333 24855 -20299
rect 24889 -20333 24928 -20299
rect 24816 -20371 24928 -20333
rect 24816 -20405 24855 -20371
rect 24889 -20405 24928 -20371
rect 24816 -20443 24928 -20405
rect 24816 -20477 24855 -20443
rect 24889 -20477 24928 -20443
rect 24816 -20515 24928 -20477
rect 24816 -20549 24855 -20515
rect 24889 -20549 24928 -20515
rect 24816 -20587 24928 -20549
rect 24816 -20621 24855 -20587
rect 24889 -20621 24928 -20587
rect 24816 -20659 24928 -20621
rect 24816 -20693 24855 -20659
rect 24889 -20693 24928 -20659
rect 24816 -20731 24928 -20693
rect 24816 -20765 24855 -20731
rect 24889 -20765 24928 -20731
rect 24816 -20803 24928 -20765
rect 24816 -20837 24855 -20803
rect 24889 -20837 24928 -20803
rect 24816 -20875 24928 -20837
rect 24816 -20909 24855 -20875
rect 24889 -20909 24928 -20875
rect 24816 -20947 24928 -20909
rect 24816 -20981 24855 -20947
rect 24889 -20981 24928 -20947
rect 24816 -21019 24928 -20981
rect 24816 -21053 24855 -21019
rect 24889 -21053 24928 -21019
rect 24816 -21091 24928 -21053
rect 24816 -21125 24855 -21091
rect 24889 -21125 24928 -21091
rect 24816 -21163 24928 -21125
rect 24816 -21197 24855 -21163
rect 24889 -21197 24928 -21163
rect 24816 -21235 24928 -21197
rect 24816 -21269 24855 -21235
rect 24889 -21269 24928 -21235
rect 24816 -21307 24928 -21269
rect 24816 -21341 24855 -21307
rect 24889 -21341 24928 -21307
rect 24816 -21379 24928 -21341
rect 24816 -21413 24855 -21379
rect 24889 -21413 24928 -21379
rect 24816 -21451 24928 -21413
rect 24816 -21485 24855 -21451
rect 24889 -21485 24928 -21451
rect 24816 -21523 24928 -21485
rect 24816 -21557 24855 -21523
rect 24889 -21557 24928 -21523
rect 24816 -21595 24928 -21557
rect 24816 -21629 24855 -21595
rect 24889 -21629 24928 -21595
rect 24816 -21667 24928 -21629
rect 24816 -21701 24855 -21667
rect 24889 -21701 24928 -21667
rect 24816 -21739 24928 -21701
rect 24816 -21773 24855 -21739
rect 24889 -21773 24928 -21739
rect 24816 -21811 24928 -21773
rect 24816 -21845 24855 -21811
rect 24889 -21845 24928 -21811
rect 24816 -21883 24928 -21845
rect 24816 -21917 24855 -21883
rect 24889 -21917 24928 -21883
rect 24816 -21955 24928 -21917
rect 24816 -21989 24855 -21955
rect 24889 -21989 24928 -21955
rect 24816 -22027 24928 -21989
rect 24816 -22061 24855 -22027
rect 24889 -22061 24928 -22027
rect 24816 -22099 24928 -22061
rect 24816 -22133 24855 -22099
rect 24889 -22133 24928 -22099
rect 24816 -22171 24928 -22133
rect 24816 -22205 24855 -22171
rect 24889 -22205 24928 -22171
rect 24816 -22243 24928 -22205
rect 24816 -22277 24855 -22243
rect 24889 -22277 24928 -22243
rect 24816 -22315 24928 -22277
rect 24816 -22349 24855 -22315
rect 24889 -22349 24928 -22315
rect 24816 -22387 24928 -22349
rect 24816 -22421 24855 -22387
rect 24889 -22421 24928 -22387
rect 24816 -22459 24928 -22421
rect 24816 -22493 24855 -22459
rect 24889 -22493 24928 -22459
rect 24816 -22531 24928 -22493
rect 24816 -22565 24855 -22531
rect 24889 -22565 24928 -22531
rect 24816 -22603 24928 -22565
rect 24816 -22637 24855 -22603
rect 24889 -22637 24928 -22603
rect 24816 -22675 24928 -22637
rect 24816 -22709 24855 -22675
rect 24889 -22709 24928 -22675
rect 24816 -22747 24928 -22709
rect 24816 -22781 24855 -22747
rect 24889 -22781 24928 -22747
rect 24816 -22819 24928 -22781
rect 24816 -22853 24855 -22819
rect 24889 -22853 24928 -22819
rect 24816 -22891 24928 -22853
rect 24816 -22925 24855 -22891
rect 24889 -22925 24928 -22891
rect 24816 -22963 24928 -22925
rect 24816 -22997 24855 -22963
rect 24889 -22997 24928 -22963
rect 24816 -23035 24928 -22997
rect 24816 -23069 24855 -23035
rect 24889 -23069 24928 -23035
rect 24816 -23107 24928 -23069
rect 24816 -23141 24855 -23107
rect 24889 -23141 24928 -23107
rect 24816 -23179 24928 -23141
rect 24816 -23213 24855 -23179
rect 24889 -23213 24928 -23179
rect 24816 -23251 24928 -23213
rect 24816 -23285 24855 -23251
rect 24889 -23285 24928 -23251
rect 24816 -23323 24928 -23285
rect 24816 -23357 24855 -23323
rect 24889 -23357 24928 -23323
rect 24816 -23395 24928 -23357
rect 24816 -23429 24855 -23395
rect 24889 -23429 24928 -23395
rect 24816 -23467 24928 -23429
rect 24816 -23501 24855 -23467
rect 24889 -23501 24928 -23467
rect 24816 -23539 24928 -23501
rect 24816 -23573 24855 -23539
rect 24889 -23573 24928 -23539
rect 24816 -23611 24928 -23573
rect 24816 -23645 24855 -23611
rect 24889 -23645 24928 -23611
rect 24816 -23683 24928 -23645
rect 24816 -23717 24855 -23683
rect 24889 -23717 24928 -23683
rect 24816 -23755 24928 -23717
rect 24816 -23789 24855 -23755
rect 24889 -23789 24928 -23755
rect 24816 -23827 24928 -23789
rect 24816 -23861 24855 -23827
rect 24889 -23861 24928 -23827
rect 24816 -23899 24928 -23861
rect 24816 -23933 24855 -23899
rect 24889 -23933 24928 -23899
rect 24816 -23971 24928 -23933
rect 24816 -24005 24855 -23971
rect 24889 -24005 24928 -23971
rect 24816 -24043 24928 -24005
rect 24816 -24077 24855 -24043
rect 24889 -24077 24928 -24043
rect 24816 -24115 24928 -24077
rect 24816 -24149 24855 -24115
rect 24889 -24149 24928 -24115
rect 24816 -24187 24928 -24149
rect 24816 -24221 24855 -24187
rect 24889 -24221 24928 -24187
rect 24816 -24259 24928 -24221
rect 24816 -24293 24855 -24259
rect 24889 -24293 24928 -24259
rect 24816 -24331 24928 -24293
rect 24816 -24365 24855 -24331
rect 24889 -24365 24928 -24331
rect 24816 -24403 24928 -24365
rect 24816 -24437 24855 -24403
rect 24889 -24437 24928 -24403
rect 24816 -24475 24928 -24437
rect 24816 -24509 24855 -24475
rect 24889 -24509 24928 -24475
rect 24816 -24547 24928 -24509
rect 24816 -24581 24855 -24547
rect 24889 -24581 24928 -24547
rect 24816 -24619 24928 -24581
rect 24816 -24653 24855 -24619
rect 24889 -24653 24928 -24619
rect 24816 -24691 24928 -24653
rect 24816 -24725 24855 -24691
rect 24889 -24725 24928 -24691
rect 24816 -24763 24928 -24725
rect 24816 -24797 24855 -24763
rect 24889 -24797 24928 -24763
rect 24816 -24835 24928 -24797
rect 24816 -24869 24855 -24835
rect 24889 -24869 24928 -24835
rect 24816 -24907 24928 -24869
rect 23756 -24932 23828 -24928
rect 23756 -24984 23766 -24932
rect 23818 -24984 23828 -24932
rect 23756 -24988 23828 -24984
rect 24816 -24941 24855 -24907
rect 24889 -24941 24928 -24907
rect 24816 -24979 24928 -24941
rect 24816 -25013 24855 -24979
rect 24889 -25013 24928 -24979
rect 24816 -25051 24928 -25013
rect 24816 -25085 24855 -25051
rect 24889 -25085 24928 -25051
rect 24816 -25123 24928 -25085
rect 24816 -25157 24855 -25123
rect 24889 -25157 24928 -25123
rect 24816 -25195 24928 -25157
rect 24816 -25229 24855 -25195
rect 24889 -25229 24928 -25195
rect 24816 -25267 24928 -25229
rect 24816 -25301 24855 -25267
rect 24889 -25301 24928 -25267
rect 24816 -25339 24928 -25301
rect 24816 -25373 24855 -25339
rect 24889 -25373 24928 -25339
rect 24816 -25411 24928 -25373
rect 24816 -25445 24855 -25411
rect 24889 -25445 24928 -25411
rect 24816 -25483 24928 -25445
rect 24816 -25517 24855 -25483
rect 24889 -25517 24928 -25483
rect 24816 -25555 24928 -25517
rect 24816 -25589 24855 -25555
rect 24889 -25589 24928 -25555
rect 24816 -25627 24928 -25589
rect 24816 -25661 24855 -25627
rect 24889 -25661 24928 -25627
rect 24816 -25699 24928 -25661
rect 24816 -25733 24855 -25699
rect 24889 -25733 24928 -25699
rect 24816 -25771 24928 -25733
rect 24816 -25805 24855 -25771
rect 24889 -25805 24928 -25771
rect 24816 -25843 24928 -25805
rect 24816 -25877 24855 -25843
rect 24889 -25877 24928 -25843
rect 24816 -25915 24928 -25877
rect 24816 -25949 24855 -25915
rect 24889 -25949 24928 -25915
rect 24816 -25987 24928 -25949
rect 24816 -26021 24855 -25987
rect 24889 -26021 24928 -25987
rect 24816 -26059 24928 -26021
rect 23048 -26070 23120 -26066
rect 23048 -26122 23058 -26070
rect 23110 -26122 23120 -26070
rect 23048 -26126 23120 -26122
rect 24816 -26093 24855 -26059
rect 24889 -26093 24928 -26059
rect 24816 -26131 24928 -26093
rect 24816 -26165 24855 -26131
rect 24889 -26165 24928 -26131
rect 21402 -26178 21464 -26168
rect 21402 -26180 21408 -26178
rect 21404 -26230 21408 -26180
rect 21460 -26230 21464 -26178
rect 21404 -26240 21464 -26230
rect 24816 -26203 24928 -26165
rect 24816 -26237 24855 -26203
rect 24889 -26237 24928 -26203
rect 24816 -26275 24928 -26237
rect 24816 -26309 24855 -26275
rect 24889 -26309 24928 -26275
rect -8118 -26476 -7968 -26430
rect -7922 -26476 -4748 -26430
rect -4688 -26476 1704 -26430
rect 1764 -26476 23806 -26430
rect 23866 -26476 23968 -26430
rect -8118 -26495 23968 -26476
rect -8118 -26611 -8066 -26495
rect 23922 -26611 23968 -26495
rect -8118 -26676 23968 -26611
rect 24816 -26816 24928 -26309
rect -12328 -26844 -11606 -26816
rect -12328 -27088 -12198 -26844
rect -11634 -27088 -11606 -26844
rect -12328 -27116 -11606 -27088
rect 24206 -26844 24928 -26816
rect 24206 -27088 24234 -26844
rect 24798 -27088 24928 -26844
rect 24206 -27116 24928 -27088
rect -12328 -27155 24928 -27116
rect -12328 -27189 -12221 -27155
rect -12187 -27189 -12149 -27155
rect -12115 -27189 -12077 -27155
rect -12043 -27189 -12005 -27155
rect -11971 -27189 -11933 -27155
rect -11899 -27189 -11861 -27155
rect -11827 -27189 -11789 -27155
rect -11755 -27189 -11717 -27155
rect -11683 -27189 -11645 -27155
rect -11611 -27189 -11573 -27155
rect -11539 -27189 -11501 -27155
rect -11467 -27189 -11429 -27155
rect -11395 -27189 -11357 -27155
rect -11323 -27189 -11285 -27155
rect -11251 -27189 -11213 -27155
rect -11179 -27189 -11141 -27155
rect -11107 -27189 -11069 -27155
rect -11035 -27189 -10997 -27155
rect -10963 -27189 -10925 -27155
rect -10891 -27189 -10853 -27155
rect -10819 -27189 -10781 -27155
rect -10747 -27189 -10709 -27155
rect -10675 -27189 -10637 -27155
rect -10603 -27189 -10565 -27155
rect -10531 -27189 -10493 -27155
rect -10459 -27189 -10421 -27155
rect -10387 -27189 -10349 -27155
rect -10315 -27189 -10277 -27155
rect -10243 -27189 -10205 -27155
rect -10171 -27189 -10133 -27155
rect -10099 -27189 -10061 -27155
rect -10027 -27189 -9989 -27155
rect -9955 -27189 -9917 -27155
rect -9883 -27189 -9845 -27155
rect -9811 -27189 -9773 -27155
rect -9739 -27189 -9701 -27155
rect -9667 -27189 -9629 -27155
rect -9595 -27189 -9557 -27155
rect -9523 -27189 -9485 -27155
rect -9451 -27189 -9413 -27155
rect -9379 -27189 -9341 -27155
rect -9307 -27189 -9269 -27155
rect -9235 -27189 -9197 -27155
rect -9163 -27189 -9125 -27155
rect -9091 -27189 -9053 -27155
rect -9019 -27189 -8981 -27155
rect -8947 -27189 -8909 -27155
rect -8875 -27189 -8837 -27155
rect -8803 -27189 -8765 -27155
rect -8731 -27189 -8693 -27155
rect -8659 -27189 -8621 -27155
rect -8587 -27189 -8549 -27155
rect -8515 -27189 -8477 -27155
rect -8443 -27189 -8405 -27155
rect -8371 -27189 -8333 -27155
rect -8299 -27189 -8261 -27155
rect -8227 -27189 -8189 -27155
rect -8155 -27189 -8117 -27155
rect -8083 -27189 -8045 -27155
rect -8011 -27189 -7973 -27155
rect -7939 -27189 -7901 -27155
rect -7867 -27189 -7829 -27155
rect -7795 -27189 -7757 -27155
rect -7723 -27189 -7685 -27155
rect -7651 -27189 -7613 -27155
rect -7579 -27189 -7541 -27155
rect -7507 -27189 -7469 -27155
rect -7435 -27189 -7397 -27155
rect -7363 -27189 -7325 -27155
rect -7291 -27189 -7253 -27155
rect -7219 -27189 -7181 -27155
rect -7147 -27189 -7109 -27155
rect -7075 -27189 -7037 -27155
rect -7003 -27189 -6965 -27155
rect -6931 -27189 -6893 -27155
rect -6859 -27189 -6821 -27155
rect -6787 -27189 -6749 -27155
rect -6715 -27189 -6677 -27155
rect -6643 -27189 -6605 -27155
rect -6571 -27189 -6533 -27155
rect -6499 -27189 -6461 -27155
rect -6427 -27189 -6389 -27155
rect -6355 -27189 -6317 -27155
rect -6283 -27189 -6245 -27155
rect -6211 -27189 -6173 -27155
rect -6139 -27189 -6101 -27155
rect -6067 -27189 -6029 -27155
rect -5995 -27189 -5957 -27155
rect -5923 -27189 -5885 -27155
rect -5851 -27189 -5813 -27155
rect -5779 -27189 -5741 -27155
rect -5707 -27189 -5669 -27155
rect -5635 -27189 -5597 -27155
rect -5563 -27189 -5525 -27155
rect -5491 -27189 -5453 -27155
rect -5419 -27189 -5381 -27155
rect -5347 -27189 -5309 -27155
rect -5275 -27189 -5237 -27155
rect -5203 -27189 -5165 -27155
rect -5131 -27189 -5093 -27155
rect -5059 -27189 -5021 -27155
rect -4987 -27189 -4949 -27155
rect -4915 -27189 -4877 -27155
rect -4843 -27189 -4805 -27155
rect -4771 -27189 -4733 -27155
rect -4699 -27189 -4661 -27155
rect -4627 -27189 -4589 -27155
rect -4555 -27189 -4517 -27155
rect -4483 -27189 -4445 -27155
rect -4411 -27189 -4373 -27155
rect -4339 -27189 -4301 -27155
rect -4267 -27189 -4229 -27155
rect -4195 -27189 -4157 -27155
rect -4123 -27189 -4085 -27155
rect -4051 -27189 -4013 -27155
rect -3979 -27189 -3941 -27155
rect -3907 -27189 -3869 -27155
rect -3835 -27189 -3797 -27155
rect -3763 -27189 -3725 -27155
rect -3691 -27189 -3653 -27155
rect -3619 -27189 -3581 -27155
rect -3547 -27189 -3509 -27155
rect -3475 -27189 -3437 -27155
rect -3403 -27189 -3365 -27155
rect -3331 -27189 -3293 -27155
rect -3259 -27189 -3221 -27155
rect -3187 -27189 -3149 -27155
rect -3115 -27189 -3077 -27155
rect -3043 -27189 -3005 -27155
rect -2971 -27189 -2933 -27155
rect -2899 -27189 -2861 -27155
rect -2827 -27189 -2789 -27155
rect -2755 -27189 -2717 -27155
rect -2683 -27189 -2645 -27155
rect -2611 -27189 -2573 -27155
rect -2539 -27189 -2501 -27155
rect -2467 -27189 -2429 -27155
rect -2395 -27189 -2357 -27155
rect -2323 -27189 -2285 -27155
rect -2251 -27189 -2213 -27155
rect -2179 -27189 -2141 -27155
rect -2107 -27189 -2069 -27155
rect -2035 -27189 -1997 -27155
rect -1963 -27189 -1925 -27155
rect -1891 -27189 -1853 -27155
rect -1819 -27189 -1781 -27155
rect -1747 -27189 -1709 -27155
rect -1675 -27189 -1637 -27155
rect -1603 -27189 -1565 -27155
rect -1531 -27189 -1493 -27155
rect -1459 -27189 -1421 -27155
rect -1387 -27189 -1349 -27155
rect -1315 -27189 -1277 -27155
rect -1243 -27189 -1205 -27155
rect -1171 -27189 -1133 -27155
rect -1099 -27189 -1061 -27155
rect -1027 -27189 -989 -27155
rect -955 -27189 -917 -27155
rect -883 -27189 -845 -27155
rect -811 -27189 -773 -27155
rect -739 -27189 -701 -27155
rect -667 -27189 -629 -27155
rect -595 -27189 -557 -27155
rect -523 -27189 -485 -27155
rect -451 -27189 -413 -27155
rect -379 -27189 -341 -27155
rect -307 -27189 -269 -27155
rect -235 -27189 -197 -27155
rect -163 -27189 -125 -27155
rect -91 -27189 -53 -27155
rect -19 -27189 19 -27155
rect 53 -27189 91 -27155
rect 125 -27189 163 -27155
rect 197 -27189 235 -27155
rect 269 -27189 307 -27155
rect 341 -27189 379 -27155
rect 413 -27189 451 -27155
rect 485 -27189 523 -27155
rect 557 -27189 595 -27155
rect 629 -27189 667 -27155
rect 701 -27189 739 -27155
rect 773 -27189 811 -27155
rect 845 -27189 883 -27155
rect 917 -27189 955 -27155
rect 989 -27189 1027 -27155
rect 1061 -27189 1099 -27155
rect 1133 -27189 1171 -27155
rect 1205 -27189 1243 -27155
rect 1277 -27189 1315 -27155
rect 1349 -27189 1387 -27155
rect 1421 -27189 1459 -27155
rect 1493 -27189 1531 -27155
rect 1565 -27189 1603 -27155
rect 1637 -27189 1675 -27155
rect 1709 -27189 1747 -27155
rect 1781 -27189 1819 -27155
rect 1853 -27189 1891 -27155
rect 1925 -27189 1963 -27155
rect 1997 -27189 2035 -27155
rect 2069 -27189 2107 -27155
rect 2141 -27189 2179 -27155
rect 2213 -27189 2251 -27155
rect 2285 -27189 2323 -27155
rect 2357 -27189 2395 -27155
rect 2429 -27189 2467 -27155
rect 2501 -27189 2539 -27155
rect 2573 -27189 2611 -27155
rect 2645 -27189 2683 -27155
rect 2717 -27189 2755 -27155
rect 2789 -27189 2827 -27155
rect 2861 -27189 2899 -27155
rect 2933 -27189 2971 -27155
rect 3005 -27189 3043 -27155
rect 3077 -27189 3115 -27155
rect 3149 -27189 3187 -27155
rect 3221 -27189 3259 -27155
rect 3293 -27189 3331 -27155
rect 3365 -27189 3403 -27155
rect 3437 -27189 3475 -27155
rect 3509 -27189 3547 -27155
rect 3581 -27189 3619 -27155
rect 3653 -27189 3691 -27155
rect 3725 -27189 3763 -27155
rect 3797 -27189 3835 -27155
rect 3869 -27189 3907 -27155
rect 3941 -27189 3979 -27155
rect 4013 -27189 4051 -27155
rect 4085 -27189 4123 -27155
rect 4157 -27189 4195 -27155
rect 4229 -27189 4267 -27155
rect 4301 -27189 4339 -27155
rect 4373 -27189 4411 -27155
rect 4445 -27189 4483 -27155
rect 4517 -27189 4555 -27155
rect 4589 -27189 4627 -27155
rect 4661 -27189 4699 -27155
rect 4733 -27189 4771 -27155
rect 4805 -27189 4843 -27155
rect 4877 -27189 4915 -27155
rect 4949 -27189 4987 -27155
rect 5021 -27189 5059 -27155
rect 5093 -27189 5131 -27155
rect 5165 -27189 5203 -27155
rect 5237 -27189 5275 -27155
rect 5309 -27189 5347 -27155
rect 5381 -27189 5419 -27155
rect 5453 -27189 5491 -27155
rect 5525 -27189 5563 -27155
rect 5597 -27189 5635 -27155
rect 5669 -27189 5707 -27155
rect 5741 -27189 5779 -27155
rect 5813 -27189 5851 -27155
rect 5885 -27189 5923 -27155
rect 5957 -27189 5995 -27155
rect 6029 -27189 6067 -27155
rect 6101 -27189 6139 -27155
rect 6173 -27189 6211 -27155
rect 6245 -27189 6283 -27155
rect 6317 -27189 6355 -27155
rect 6389 -27189 6427 -27155
rect 6461 -27189 6499 -27155
rect 6533 -27189 6571 -27155
rect 6605 -27189 6643 -27155
rect 6677 -27189 6715 -27155
rect 6749 -27189 6787 -27155
rect 6821 -27189 6859 -27155
rect 6893 -27189 6931 -27155
rect 6965 -27189 7003 -27155
rect 7037 -27189 7075 -27155
rect 7109 -27189 7147 -27155
rect 7181 -27189 7219 -27155
rect 7253 -27189 7291 -27155
rect 7325 -27189 7363 -27155
rect 7397 -27189 7435 -27155
rect 7469 -27189 7507 -27155
rect 7541 -27189 7579 -27155
rect 7613 -27189 7651 -27155
rect 7685 -27189 7723 -27155
rect 7757 -27189 7795 -27155
rect 7829 -27189 7867 -27155
rect 7901 -27189 7939 -27155
rect 7973 -27189 8011 -27155
rect 8045 -27189 8083 -27155
rect 8117 -27189 8155 -27155
rect 8189 -27189 8227 -27155
rect 8261 -27189 8299 -27155
rect 8333 -27189 8371 -27155
rect 8405 -27189 8443 -27155
rect 8477 -27189 8515 -27155
rect 8549 -27189 8587 -27155
rect 8621 -27189 8659 -27155
rect 8693 -27189 8731 -27155
rect 8765 -27189 8803 -27155
rect 8837 -27189 8875 -27155
rect 8909 -27189 8947 -27155
rect 8981 -27189 9019 -27155
rect 9053 -27189 9091 -27155
rect 9125 -27189 9163 -27155
rect 9197 -27189 9235 -27155
rect 9269 -27189 9307 -27155
rect 9341 -27189 9379 -27155
rect 9413 -27189 9451 -27155
rect 9485 -27189 9523 -27155
rect 9557 -27189 9595 -27155
rect 9629 -27189 9667 -27155
rect 9701 -27189 9739 -27155
rect 9773 -27189 9811 -27155
rect 9845 -27189 9883 -27155
rect 9917 -27189 9955 -27155
rect 9989 -27189 10027 -27155
rect 10061 -27189 10099 -27155
rect 10133 -27189 10171 -27155
rect 10205 -27189 10243 -27155
rect 10277 -27189 10315 -27155
rect 10349 -27189 10387 -27155
rect 10421 -27189 10459 -27155
rect 10493 -27189 10531 -27155
rect 10565 -27189 10603 -27155
rect 10637 -27189 10675 -27155
rect 10709 -27189 10747 -27155
rect 10781 -27189 10819 -27155
rect 10853 -27189 10891 -27155
rect 10925 -27189 10963 -27155
rect 10997 -27189 11035 -27155
rect 11069 -27189 11107 -27155
rect 11141 -27189 11179 -27155
rect 11213 -27189 11251 -27155
rect 11285 -27189 11323 -27155
rect 11357 -27189 11395 -27155
rect 11429 -27189 11467 -27155
rect 11501 -27189 11539 -27155
rect 11573 -27189 11611 -27155
rect 11645 -27189 11683 -27155
rect 11717 -27189 11755 -27155
rect 11789 -27189 11827 -27155
rect 11861 -27189 11899 -27155
rect 11933 -27189 11971 -27155
rect 12005 -27189 12043 -27155
rect 12077 -27189 12115 -27155
rect 12149 -27189 12187 -27155
rect 12221 -27189 12259 -27155
rect 12293 -27189 12331 -27155
rect 12365 -27189 12403 -27155
rect 12437 -27189 12475 -27155
rect 12509 -27189 12547 -27155
rect 12581 -27189 12619 -27155
rect 12653 -27189 12691 -27155
rect 12725 -27189 12763 -27155
rect 12797 -27189 12835 -27155
rect 12869 -27189 12907 -27155
rect 12941 -27189 12979 -27155
rect 13013 -27189 13051 -27155
rect 13085 -27189 13123 -27155
rect 13157 -27189 13195 -27155
rect 13229 -27189 13267 -27155
rect 13301 -27189 13339 -27155
rect 13373 -27189 13411 -27155
rect 13445 -27189 13483 -27155
rect 13517 -27189 13555 -27155
rect 13589 -27189 13627 -27155
rect 13661 -27189 13699 -27155
rect 13733 -27189 13771 -27155
rect 13805 -27189 13843 -27155
rect 13877 -27189 13915 -27155
rect 13949 -27189 13987 -27155
rect 14021 -27189 14059 -27155
rect 14093 -27189 14131 -27155
rect 14165 -27189 14203 -27155
rect 14237 -27189 14275 -27155
rect 14309 -27189 14347 -27155
rect 14381 -27189 14419 -27155
rect 14453 -27189 14491 -27155
rect 14525 -27189 14563 -27155
rect 14597 -27189 14635 -27155
rect 14669 -27189 14707 -27155
rect 14741 -27189 14779 -27155
rect 14813 -27189 14851 -27155
rect 14885 -27189 14923 -27155
rect 14957 -27189 14995 -27155
rect 15029 -27189 15067 -27155
rect 15101 -27189 15139 -27155
rect 15173 -27189 15211 -27155
rect 15245 -27189 15283 -27155
rect 15317 -27189 15355 -27155
rect 15389 -27189 15427 -27155
rect 15461 -27189 15499 -27155
rect 15533 -27189 15571 -27155
rect 15605 -27189 15643 -27155
rect 15677 -27189 15715 -27155
rect 15749 -27189 15787 -27155
rect 15821 -27189 15859 -27155
rect 15893 -27189 15931 -27155
rect 15965 -27189 16003 -27155
rect 16037 -27189 16075 -27155
rect 16109 -27189 16147 -27155
rect 16181 -27189 16219 -27155
rect 16253 -27189 16291 -27155
rect 16325 -27189 16363 -27155
rect 16397 -27189 16435 -27155
rect 16469 -27189 16507 -27155
rect 16541 -27189 16579 -27155
rect 16613 -27189 16651 -27155
rect 16685 -27189 16723 -27155
rect 16757 -27189 16795 -27155
rect 16829 -27189 16867 -27155
rect 16901 -27189 16939 -27155
rect 16973 -27189 17011 -27155
rect 17045 -27189 17083 -27155
rect 17117 -27189 17155 -27155
rect 17189 -27189 17227 -27155
rect 17261 -27189 17299 -27155
rect 17333 -27189 17371 -27155
rect 17405 -27189 17443 -27155
rect 17477 -27189 17515 -27155
rect 17549 -27189 17587 -27155
rect 17621 -27189 17659 -27155
rect 17693 -27189 17731 -27155
rect 17765 -27189 17803 -27155
rect 17837 -27189 17875 -27155
rect 17909 -27189 17947 -27155
rect 17981 -27189 18019 -27155
rect 18053 -27189 18091 -27155
rect 18125 -27189 18163 -27155
rect 18197 -27189 18235 -27155
rect 18269 -27189 18307 -27155
rect 18341 -27189 18379 -27155
rect 18413 -27189 18451 -27155
rect 18485 -27189 18523 -27155
rect 18557 -27189 18595 -27155
rect 18629 -27189 18667 -27155
rect 18701 -27189 18739 -27155
rect 18773 -27189 18811 -27155
rect 18845 -27189 18883 -27155
rect 18917 -27189 18955 -27155
rect 18989 -27189 19027 -27155
rect 19061 -27189 19099 -27155
rect 19133 -27189 19171 -27155
rect 19205 -27189 19243 -27155
rect 19277 -27189 19315 -27155
rect 19349 -27189 19387 -27155
rect 19421 -27189 19459 -27155
rect 19493 -27189 19531 -27155
rect 19565 -27189 19603 -27155
rect 19637 -27189 19675 -27155
rect 19709 -27189 19747 -27155
rect 19781 -27189 19819 -27155
rect 19853 -27189 19891 -27155
rect 19925 -27189 19963 -27155
rect 19997 -27189 20035 -27155
rect 20069 -27189 20107 -27155
rect 20141 -27189 20179 -27155
rect 20213 -27189 20251 -27155
rect 20285 -27189 20323 -27155
rect 20357 -27189 20395 -27155
rect 20429 -27189 20467 -27155
rect 20501 -27189 20539 -27155
rect 20573 -27189 20611 -27155
rect 20645 -27189 20683 -27155
rect 20717 -27189 20755 -27155
rect 20789 -27189 20827 -27155
rect 20861 -27189 20899 -27155
rect 20933 -27189 20971 -27155
rect 21005 -27189 21043 -27155
rect 21077 -27189 21115 -27155
rect 21149 -27189 21187 -27155
rect 21221 -27189 21259 -27155
rect 21293 -27189 21331 -27155
rect 21365 -27189 21403 -27155
rect 21437 -27189 21475 -27155
rect 21509 -27189 21547 -27155
rect 21581 -27189 21619 -27155
rect 21653 -27189 21691 -27155
rect 21725 -27189 21763 -27155
rect 21797 -27189 21835 -27155
rect 21869 -27189 21907 -27155
rect 21941 -27189 21979 -27155
rect 22013 -27189 22051 -27155
rect 22085 -27189 22123 -27155
rect 22157 -27189 22195 -27155
rect 22229 -27189 22267 -27155
rect 22301 -27189 22339 -27155
rect 22373 -27189 22411 -27155
rect 22445 -27189 22483 -27155
rect 22517 -27189 22555 -27155
rect 22589 -27189 22627 -27155
rect 22661 -27189 22699 -27155
rect 22733 -27189 22771 -27155
rect 22805 -27189 22843 -27155
rect 22877 -27189 22915 -27155
rect 22949 -27189 22987 -27155
rect 23021 -27189 23059 -27155
rect 23093 -27189 23131 -27155
rect 23165 -27189 23203 -27155
rect 23237 -27189 23275 -27155
rect 23309 -27189 23347 -27155
rect 23381 -27189 23419 -27155
rect 23453 -27189 23491 -27155
rect 23525 -27189 23563 -27155
rect 23597 -27189 23635 -27155
rect 23669 -27189 23707 -27155
rect 23741 -27189 23779 -27155
rect 23813 -27189 23851 -27155
rect 23885 -27189 23923 -27155
rect 23957 -27189 23995 -27155
rect 24029 -27189 24067 -27155
rect 24101 -27189 24139 -27155
rect 24173 -27189 24211 -27155
rect 24245 -27189 24283 -27155
rect 24317 -27189 24355 -27155
rect 24389 -27189 24427 -27155
rect 24461 -27189 24499 -27155
rect 24533 -27189 24571 -27155
rect 24605 -27189 24643 -27155
rect 24677 -27189 24715 -27155
rect 24749 -27189 24787 -27155
rect 24821 -27189 24928 -27155
rect -12328 -27228 24928 -27189
<< via1 >>
rect 502 3944 1066 4188
rect 24134 3944 24698 4188
rect 4075 3637 20831 3817
rect 7990 1862 8042 1914
rect 9072 1862 9124 1914
rect 10030 1862 10082 1914
rect 8516 1616 8568 1668
rect 10552 1616 10604 1668
rect 13094 1862 13146 1914
rect 14112 1862 14164 1914
rect 12590 1618 12642 1670
rect 15136 1862 15188 1914
rect 16148 1862 16200 1914
rect 14620 1618 14672 1670
rect 16662 1620 16714 1672
rect 17672 1620 17724 1672
rect 19206 1862 19258 1914
rect 20218 1862 20270 1914
rect 18694 1620 18746 1672
rect 21236 1862 21288 1914
rect 20730 1620 20782 1672
rect 6334 684 6386 736
rect 7498 684 7550 736
rect 6204 480 6256 532
rect 4196 -1704 4248 -1652
rect 3680 -5962 3732 -5910
rect 3788 -6074 3840 -6022
rect 2018 -6996 2070 -6944
rect 3178 -7106 3230 -7054
rect 1892 -8084 1944 -8032
rect 3694 -8030 3746 -7978
rect 3800 -8130 3852 -8078
rect 7498 480 7550 532
rect 9534 580 9586 632
rect 11570 580 11622 632
rect 13608 684 13660 736
rect 13604 480 13656 532
rect 15642 684 15694 736
rect 15640 480 15692 532
rect 16142 480 16194 532
rect 17676 580 17728 632
rect 17162 480 17214 532
rect 19710 580 19762 632
rect 18188 480 18240 532
rect 18694 476 18746 528
rect 19208 476 19260 528
rect 19712 476 19764 528
rect 20218 476 20270 528
rect 20738 476 20790 528
rect 21750 684 21802 736
rect 23000 684 23052 736
rect 7984 -670 8036 -618
rect 10040 -454 10092 -402
rect 10550 -454 10602 -402
rect 9534 -554 9586 -502
rect 9022 -670 9074 -618
rect 10034 -670 10086 -618
rect 11410 -554 11462 -502
rect 12584 -454 12636 -402
rect 11044 -662 11096 -610
rect 12068 -662 12120 -610
rect 13096 -662 13148 -610
rect 14622 -456 14674 -404
rect 15642 -554 15694 -502
rect 16658 -456 16710 -404
rect 17158 -456 17210 -404
rect 17672 -456 17724 -404
rect 18196 -456 18248 -404
rect 18694 -456 18746 -404
rect 19196 -456 19248 -404
rect 19710 -458 19762 -406
rect 20218 -458 20270 -406
rect 20728 -458 20780 -406
rect 19200 -670 19252 -618
rect 20212 -670 20264 -618
rect 21750 -554 21802 -502
rect 21214 -670 21266 -618
rect 6334 -1990 6386 -1938
rect 6690 -4398 6742 -4346
rect 6564 -5008 6616 -4956
rect 4702 -5962 4754 -5910
rect 4572 -6074 4624 -6022
rect 5212 -6996 5264 -6944
rect 6364 -7106 6416 -7054
rect 4704 -8030 4756 -7978
rect 6556 -7234 6608 -7182
rect 4586 -8130 4638 -8078
rect 1406 -9140 1458 -9088
rect 1546 -9316 1598 -9264
rect 2446 -9490 2498 -9438
rect 6806 -5008 6858 -4956
rect 7494 -1842 7546 -1790
rect 7316 -1990 7368 -1938
rect 8514 -1592 8566 -1540
rect 9532 -1704 9584 -1652
rect 10550 -1592 10602 -1540
rect 11072 -1592 11124 -1540
rect 11570 -1592 11622 -1540
rect 12044 -1596 12096 -1544
rect 7432 -2096 7484 -2044
rect 7994 -2096 8046 -2044
rect 9036 -2096 9088 -2044
rect 10036 -2096 10088 -2044
rect 12568 -1593 12620 -1541
rect 13044 -1592 13096 -1540
rect 13604 -1846 13656 -1794
rect 14088 -1590 14140 -1538
rect 13198 -2096 13250 -2044
rect 14620 -1592 14672 -1540
rect 16132 -1590 16184 -1538
rect 15640 -1988 15692 -1936
rect 14208 -2096 14260 -2044
rect 15150 -2096 15202 -2044
rect 16642 -1595 16694 -1543
rect 17154 -1600 17206 -1548
rect 17659 -1597 17711 -1545
rect 18154 -1600 18206 -1548
rect 18694 -1596 18746 -1544
rect 20728 -1596 20780 -1544
rect 19712 -1704 19764 -1652
rect 22998 -1842 23050 -1790
rect 21744 -1990 21796 -1938
rect 7546 -2298 7598 -2246
rect 8690 -3234 8742 -3182
rect 9194 -3342 9246 -3290
rect 8686 -4266 8738 -4214
rect 9192 -4400 9244 -4348
rect 10724 -2298 10776 -2246
rect 10724 -3234 10776 -3182
rect 10216 -3342 10268 -3290
rect 11234 -3342 11286 -3290
rect 10206 -4404 10258 -4352
rect 11238 -4396 11290 -4344
rect 12766 -3234 12818 -3182
rect 12258 -3342 12310 -3290
rect 13272 -3342 13324 -3290
rect 12766 -4266 12818 -4214
rect 12236 -4396 12288 -4344
rect 13280 -4396 13332 -4344
rect 14792 -2298 14844 -2246
rect 14792 -3234 14844 -3182
rect 14290 -3342 14342 -3290
rect 15300 -3342 15352 -3290
rect 14284 -4400 14336 -4348
rect 15300 -4400 15352 -4348
rect 14084 -4608 14136 -4556
rect 7316 -4926 7368 -4874
rect 8482 -4926 8534 -4874
rect 7048 -5972 7100 -5920
rect 6806 -7130 6858 -7078
rect 6802 -7344 6854 -7292
rect 6690 -8386 6742 -8334
rect 1286 -9640 1338 -9588
rect 7184 -6070 7236 -6018
rect 7048 -9644 7100 -9592
rect 10518 -4926 10570 -4874
rect 11028 -4928 11080 -4876
rect 9500 -5874 9552 -5822
rect 11536 -5874 11588 -5822
rect 11878 -5872 11930 -5820
rect 18868 -2298 18920 -2246
rect 16834 -3234 16886 -3182
rect 16322 -3342 16374 -3290
rect 17336 -3342 17388 -3290
rect 16834 -4266 16886 -4214
rect 16304 -4400 16356 -4348
rect 17336 -4396 17388 -4344
rect 15820 -4608 15872 -4556
rect 15102 -4806 15154 -4754
rect 18870 -3234 18922 -3182
rect 18368 -3342 18420 -3290
rect 19378 -3342 19430 -3290
rect 18352 -4400 18404 -4348
rect 19380 -4400 19432 -4348
rect 22064 -2298 22116 -2246
rect 20906 -3234 20958 -3182
rect 20400 -3342 20452 -3290
rect 20902 -4266 20954 -4214
rect 20400 -4400 20452 -4348
rect 22858 -4398 22910 -4346
rect 21718 -4624 21770 -4572
rect 19166 -4806 19218 -4754
rect 20190 -4806 20242 -4754
rect 21202 -4806 21254 -4754
rect 15104 -4928 15156 -4876
rect 14592 -5872 14644 -5820
rect 9500 -6070 9552 -6018
rect 10520 -6068 10572 -6016
rect 8486 -6180 8538 -6128
rect 10520 -6180 10572 -6128
rect 18664 -4926 18716 -4874
rect 20698 -4926 20750 -4874
rect 15610 -6068 15662 -6016
rect 13576 -6182 13628 -6130
rect 15610 -6182 15662 -6130
rect 18666 -6182 18718 -6130
rect 19680 -5874 19732 -5822
rect 20700 -6182 20752 -6130
rect 21716 -5874 21768 -5822
rect 7468 -7344 7520 -7292
rect 9502 -7234 9554 -7182
rect 9502 -7438 9554 -7386
rect 13572 -7130 13624 -7078
rect 11538 -7234 11590 -7182
rect 11536 -7336 11588 -7284
rect 11536 -7438 11588 -7386
rect 14592 -7130 14644 -7078
rect 14592 -7436 14644 -7384
rect 15610 -7436 15662 -7384
rect 16628 -7130 16680 -7078
rect 16626 -7436 16678 -7384
rect 18662 -7234 18714 -7182
rect 19530 -7116 19582 -7064
rect 19678 -7226 19730 -7174
rect 19530 -7436 19582 -7384
rect 19682 -7434 19734 -7382
rect 20698 -7336 20750 -7284
rect 23294 -4266 23346 -4214
rect 23000 -4626 23052 -4574
rect 23142 -4926 23194 -4874
rect 22982 -6068 23034 -6016
rect 21718 -7226 21770 -7174
rect 22858 -7226 22910 -7174
rect 21716 -7434 21768 -7382
rect 8484 -8386 8536 -8334
rect 7316 -8594 7368 -8542
rect 9498 -8696 9550 -8644
rect 10520 -8386 10572 -8334
rect 10520 -8494 10572 -8442
rect 11538 -8378 11590 -8326
rect 13340 -8378 13392 -8326
rect 11532 -8696 11584 -8644
rect 11736 -8708 11788 -8656
rect 13574 -8384 13626 -8332
rect 15610 -8384 15662 -8332
rect 15608 -8494 15660 -8442
rect 15098 -8708 15150 -8656
rect 18664 -8382 18716 -8330
rect 16114 -8708 16166 -8656
rect 19174 -8708 19226 -8656
rect 19686 -8696 19738 -8644
rect 20700 -8382 20752 -8330
rect 22982 -7434 23034 -7382
rect 22858 -8494 22910 -8442
rect 21720 -8696 21772 -8644
rect 8480 -9644 8532 -9592
rect 10516 -9644 10568 -9592
rect 7184 -9774 7236 -9722
rect 2340 -9902 2392 -9850
rect 2220 -10020 2272 -9968
rect 18668 -9644 18720 -9592
rect 20704 -9644 20756 -9592
rect 11538 -9914 11590 -9862
rect 23294 -6182 23346 -6130
rect 23142 -9914 23194 -9862
rect 1774 -10138 1826 -10086
rect -13618 -10646 -2878 -10402
rect 1892 -11414 1944 -11362
rect 2220 -11404 2272 -11352
rect 1286 -11550 1338 -11498
rect 1406 -11548 1458 -11496
rect 1546 -11530 1598 -11478
rect 1774 -11514 1826 -11462
rect 1154 -11678 1206 -11626
rect -1558 -12276 -1506 -12224
rect -32 -12410 20 -12358
rect 1154 -18878 1206 -18826
rect -3394 -19804 -3342 -19752
rect -9504 -19950 -9452 -19898
rect -10658 -20078 -10606 -20026
rect -5424 -19950 -5372 -19898
rect -7980 -20078 -7928 -20026
rect -6948 -20078 -6896 -20026
rect -3888 -20078 -3836 -20026
rect -9000 -21040 -8948 -20988
rect -9500 -21144 -9448 -21092
rect -10658 -22310 -10606 -22258
rect -7976 -21040 -7924 -20988
rect -8482 -21248 -8430 -21196
rect -9008 -22310 -8956 -22258
rect -6944 -21040 -6892 -20988
rect -7464 -21144 -7412 -21092
rect -5944 -21040 -5892 -20988
rect -4924 -21040 -4872 -20988
rect -5428 -21144 -5376 -21092
rect -6446 -21248 -6394 -21196
rect -7470 -22190 -7418 -22138
rect -8482 -23254 -8430 -23202
rect -9496 -23362 -9444 -23310
rect -9002 -23474 -8950 -23422
rect -7460 -23362 -7408 -23310
rect -7978 -23474 -7926 -23422
rect -5938 -22310 -5886 -22258
rect -3904 -21040 -3852 -20988
rect -4414 -21248 -4362 -21196
rect -4930 -22310 -4878 -22258
rect -6446 -23254 -6394 -23202
rect -6946 -23474 -6894 -23422
rect -1364 -19950 -1312 -19898
rect 820 -19950 872 -19898
rect -2892 -20078 -2840 -20026
rect -2894 -21040 -2842 -20988
rect -3394 -21144 -3342 -21092
rect -1880 -21040 -1828 -20988
rect -862 -21040 -810 -20988
rect -1358 -21144 -1306 -21092
rect -2380 -21248 -2328 -21196
rect -3394 -22190 -3342 -22138
rect -4414 -23254 -4362 -23202
rect -5424 -23362 -5372 -23310
rect -5946 -23474 -5894 -23422
rect -4926 -23474 -4874 -23422
rect -3390 -23362 -3338 -23310
rect -3906 -23474 -3854 -23422
rect -2896 -23474 -2844 -23422
rect -1868 -22310 -1816 -22258
rect -336 -21248 -284 -21196
rect 940 -21040 992 -20988
rect 820 -22190 872 -22138
rect -842 -22310 -790 -22258
rect -2380 -23254 -2328 -23202
rect -336 -23254 -284 -23202
rect -1354 -23362 -1302 -23310
rect -1882 -23474 -1830 -23422
rect -864 -23474 -812 -23422
rect -10658 -24436 -10606 -24384
rect -7988 -24436 -7936 -24384
rect -6956 -24436 -6904 -24384
rect -3896 -24436 -3844 -24384
rect -2900 -24436 -2848 -24384
rect 940 -23474 992 -23422
rect -9502 -24566 -9450 -24514
rect -5422 -24566 -5370 -24514
rect -1362 -24566 -1310 -24514
rect 820 -24566 872 -24514
rect -8024 -25932 -7972 -25880
rect -5986 -25932 -5934 -25880
rect -3950 -25932 -3898 -25880
rect -7006 -26044 -6954 -25992
rect -1914 -25932 -1862 -25880
rect -2932 -26044 -2880 -25992
rect 1286 -19950 1338 -19898
rect 1406 -20078 1458 -20026
rect 1664 -11668 1716 -11616
rect 1774 -12410 1826 -12358
rect 2340 -11412 2392 -11360
rect 2220 -12276 2272 -12224
rect 2016 -13634 2068 -13582
rect 1890 -15336 1942 -15284
rect 1664 -17796 1716 -17744
rect 1546 -21040 1598 -20988
rect 2228 -13970 2280 -13918
rect 2124 -15230 2176 -15178
rect 2016 -16330 2068 -16278
rect 2446 -11548 2498 -11496
rect 13258 -11898 13310 -11846
rect 18362 -11898 18414 -11846
rect 22422 -11904 22474 -11852
rect 3590 -13634 3642 -13582
rect 4604 -13850 4656 -13798
rect 6644 -13850 6696 -13798
rect 8684 -13850 8736 -13798
rect 10714 -13850 10766 -13798
rect 12754 -13850 12806 -13798
rect 14786 -13850 14838 -13798
rect 16826 -13850 16878 -13798
rect 18862 -13850 18914 -13798
rect 20896 -13850 20948 -13798
rect 2572 -13970 2624 -13918
rect 4096 -13976 4148 -13924
rect 2446 -14092 2498 -14040
rect 5110 -13976 5162 -13924
rect 6132 -13976 6184 -13924
rect 7146 -13976 7198 -13924
rect 8172 -13976 8224 -13924
rect 7660 -14092 7712 -14040
rect 9184 -13976 9236 -13924
rect 10220 -13976 10272 -13924
rect 11226 -13976 11278 -13924
rect 12240 -13976 12292 -13924
rect 13256 -13976 13308 -13924
rect 14264 -13976 14316 -13924
rect 15280 -13976 15332 -13924
rect 16304 -13976 16356 -13924
rect 4608 -15014 4660 -14962
rect 4100 -15124 4152 -15072
rect 3590 -15230 3642 -15178
rect 2576 -15336 2628 -15284
rect 3074 -15336 3126 -15284
rect 3586 -15336 3638 -15284
rect 5122 -15124 5174 -15072
rect 6648 -15014 6700 -14962
rect 6136 -15124 6188 -15072
rect 5630 -15230 5682 -15178
rect 8680 -15014 8732 -14962
rect 7150 -15124 7202 -15072
rect 8168 -15124 8220 -15072
rect 7660 -15230 7712 -15178
rect 17326 -13976 17378 -13924
rect 18348 -13976 18400 -13924
rect 17848 -14092 17900 -14040
rect 9194 -15124 9246 -15072
rect 19366 -13976 19418 -13924
rect 20380 -13976 20432 -13924
rect 21404 -13976 21456 -13924
rect 21920 -14092 21972 -14040
rect 23052 -14092 23104 -14040
rect 10712 -15014 10764 -14962
rect 9700 -15230 9752 -15178
rect 10214 -15124 10266 -15072
rect 9866 -15336 9918 -15284
rect 2446 -16226 2498 -16174
rect 2570 -16330 2622 -16278
rect 4090 -16330 4142 -16278
rect 4602 -16330 4654 -16278
rect 2340 -16452 2392 -16400
rect 2228 -16566 2280 -16514
rect 3076 -16566 3128 -16514
rect 4608 -16564 4660 -16512
rect 5624 -16226 5676 -16174
rect 5626 -16330 5678 -16278
rect 11234 -15124 11286 -15072
rect 12748 -15014 12800 -14962
rect 12236 -15124 12288 -15072
rect 11734 -15230 11786 -15178
rect 11734 -15336 11786 -15284
rect 13262 -15124 13314 -15072
rect 14784 -15014 14836 -14962
rect 14280 -15124 14332 -15072
rect 13770 -15230 13822 -15178
rect 13772 -15336 13824 -15284
rect 6638 -16330 6690 -16278
rect 6644 -16564 6696 -16512
rect 7658 -16330 7710 -16278
rect 8680 -16226 8732 -16174
rect 2452 -17494 2504 -17442
rect 3590 -17494 3642 -17442
rect 2340 -17694 2392 -17642
rect 2234 -17796 2286 -17744
rect 2124 -21248 2176 -21196
rect 2340 -18930 2392 -18878
rect 1892 -21398 1944 -21346
rect 2234 -21286 2286 -21234
rect 3588 -17694 3640 -17642
rect 4606 -17574 4658 -17522
rect 15288 -15124 15340 -15072
rect 16822 -15014 16874 -14962
rect 16300 -15124 16352 -15072
rect 15806 -15230 15858 -15178
rect 15652 -15336 15704 -15284
rect 18860 -15014 18912 -14962
rect 17332 -15124 17384 -15072
rect 18346 -15124 18398 -15072
rect 17846 -15230 17898 -15178
rect 19364 -15124 19416 -15072
rect 20896 -15014 20948 -14962
rect 20388 -15124 20440 -15072
rect 19876 -15230 19928 -15178
rect 19876 -15334 19928 -15282
rect 21408 -15124 21460 -15072
rect 21916 -15230 21968 -15178
rect 14786 -16226 14838 -16174
rect 10716 -16330 10768 -16278
rect 12754 -16330 12806 -16278
rect 9700 -16452 9752 -16400
rect 11734 -16452 11786 -16400
rect 13764 -16452 13816 -16400
rect 5624 -17470 5676 -17418
rect 5120 -17688 5172 -17636
rect 6646 -17574 6698 -17522
rect 6124 -17688 6176 -17636
rect 7660 -17470 7712 -17418
rect 7136 -17688 7188 -17636
rect 3588 -18726 3640 -18674
rect 4094 -18828 4146 -18776
rect 8678 -17574 8730 -17522
rect 15804 -16330 15856 -16278
rect 8156 -17688 8208 -17636
rect 8678 -17686 8730 -17634
rect 10712 -17574 10764 -17522
rect 9696 -17796 9748 -17744
rect 10714 -17686 10766 -17634
rect 11730 -17796 11782 -17744
rect 5626 -18726 5678 -18674
rect 5624 -18930 5676 -18878
rect 23052 -15334 23104 -15282
rect 16822 -16330 16874 -16278
rect 17842 -16330 17894 -16278
rect 12752 -17574 12804 -17522
rect 19880 -16226 19932 -16174
rect 18858 -16330 18910 -16278
rect 20894 -16330 20946 -16278
rect 12750 -17686 12802 -17634
rect 14786 -17574 14838 -17522
rect 14982 -17578 15034 -17526
rect 13770 -17796 13822 -17744
rect 14786 -17686 14838 -17634
rect 15804 -17470 15856 -17418
rect 14982 -17796 15034 -17744
rect 15276 -17794 15328 -17742
rect 16820 -17686 16872 -17634
rect 16304 -17794 16356 -17742
rect 16822 -17800 16874 -17748
rect 7662 -18726 7714 -18674
rect 4608 -19030 4660 -18978
rect 6132 -18936 6184 -18884
rect 7154 -18936 7206 -18884
rect 6642 -19030 6694 -18978
rect 9694 -18726 9746 -18674
rect 9186 -18828 9238 -18776
rect 8168 -18936 8220 -18884
rect 9186 -18936 9238 -18884
rect 8678 -19030 8730 -18978
rect 4090 -19954 4142 -19902
rect 5000 -19954 5052 -19902
rect 4090 -20170 4142 -20118
rect 2454 -20274 2506 -20222
rect 6002 -19954 6054 -19902
rect 5128 -20170 5180 -20118
rect 7154 -19954 7206 -19902
rect 6642 -20056 6694 -20004
rect 6142 -20170 6194 -20118
rect 10206 -18936 10258 -18884
rect 17840 -17470 17892 -17418
rect 18858 -17686 18910 -17634
rect 23038 -16564 23090 -16512
rect 19874 -17578 19926 -17526
rect 20378 -17582 20430 -17530
rect 20898 -17686 20950 -17634
rect 18858 -17800 18910 -17748
rect 20896 -17800 20948 -17748
rect 14276 -18714 14328 -18662
rect 13770 -18842 13822 -18790
rect 15806 -19040 15858 -18988
rect 8164 -19954 8216 -19902
rect 9170 -19954 9222 -19902
rect 10214 -19954 10266 -19902
rect 10714 -19948 10766 -19896
rect 9168 -20170 9220 -20118
rect 10208 -20170 10260 -20118
rect 9692 -20274 9744 -20222
rect 4088 -21182 4140 -21130
rect 3590 -21286 3642 -21234
rect 3586 -21496 3638 -21444
rect 5096 -21182 5148 -21130
rect 4606 -21398 4658 -21346
rect 6110 -21182 6162 -21130
rect 11222 -20170 11274 -20118
rect 12750 -19948 12802 -19896
rect 12230 -20170 12282 -20118
rect 13274 -20170 13326 -20118
rect 11734 -20274 11786 -20222
rect 21914 -17470 21966 -17418
rect 22932 -17452 22984 -17400
rect 23166 -16582 23218 -16530
rect 23532 -17582 23584 -17530
rect 23282 -17686 23334 -17634
rect 17318 -18936 17370 -18884
rect 19370 -18714 19422 -18662
rect 19508 -18710 19560 -18658
rect 23038 -17800 23090 -17748
rect 20390 -18710 20442 -18658
rect 21396 -18710 21448 -18658
rect 21914 -18714 21966 -18662
rect 18348 -18936 18400 -18884
rect 19508 -18936 19560 -18884
rect 19876 -18936 19928 -18884
rect 19876 -19040 19928 -18988
rect 21914 -18842 21966 -18790
rect 20892 -19038 20944 -18986
rect 14786 -19948 14838 -19896
rect 14264 -20170 14316 -20118
rect 15282 -20170 15334 -20118
rect 13772 -20274 13824 -20222
rect 7148 -21182 7200 -21130
rect 6644 -21398 6696 -21346
rect 5624 -21496 5676 -21444
rect 8166 -21182 8218 -21130
rect 8682 -21176 8734 -21124
rect 16824 -19948 16876 -19896
rect 16816 -20056 16868 -20004
rect 16316 -20170 16368 -20118
rect 15806 -20274 15858 -20222
rect 16318 -20278 16370 -20226
rect 17340 -20278 17392 -20226
rect 17840 -20272 17892 -20220
rect 18860 -19948 18912 -19896
rect 18856 -20056 18908 -20004
rect 19348 -20170 19400 -20118
rect 20898 -19948 20950 -19896
rect 20894 -20056 20946 -20004
rect 20386 -20170 20438 -20118
rect 19874 -20272 19926 -20220
rect 21412 -20170 21464 -20118
rect 21916 -20272 21968 -20220
rect 10718 -21176 10770 -21124
rect 7664 -21496 7716 -21444
rect 2452 -22518 2504 -22466
rect 3592 -22734 3644 -22682
rect 12750 -21176 12802 -21124
rect 14784 -21176 14836 -21124
rect 11734 -21286 11786 -21234
rect 13770 -21286 13822 -21234
rect 10716 -21398 10768 -21346
rect 9700 -21496 9752 -21444
rect 4606 -22420 4658 -22368
rect 4610 -22614 4662 -22562
rect 5624 -22518 5676 -22466
rect 6642 -22420 6694 -22368
rect 7148 -22518 7200 -22466
rect 6646 -22614 6698 -22562
rect 8680 -22420 8732 -22368
rect 8170 -22518 8222 -22466
rect 7660 -22734 7712 -22682
rect 9192 -22518 9244 -22466
rect 8674 -22614 8726 -22562
rect 15806 -21174 15858 -21122
rect 16160 -21174 16212 -21122
rect 15802 -21286 15854 -21234
rect 15312 -21384 15364 -21332
rect 10542 -22400 10594 -22348
rect 10196 -22518 10248 -22466
rect 9694 -22734 9746 -22682
rect 10712 -22400 10764 -22348
rect 10542 -22614 10594 -22562
rect 10718 -22608 10770 -22556
rect 16350 -21384 16402 -21332
rect 17326 -21384 17378 -21332
rect 19878 -21174 19930 -21122
rect 18342 -21384 18394 -21332
rect 20368 -21384 20420 -21332
rect 16160 -21492 16212 -21440
rect 17840 -21496 17892 -21444
rect 19876 -21496 19928 -21444
rect 12754 -22400 12806 -22348
rect 14786 -22400 14838 -22348
rect 21398 -21384 21450 -21332
rect 21912 -21496 21964 -21444
rect 16826 -22400 16878 -22348
rect 15804 -22498 15856 -22446
rect 12746 -22608 12798 -22556
rect 2340 -23650 2392 -23598
rect 2234 -23776 2286 -23724
rect 5624 -23776 5676 -23724
rect 6144 -23764 6196 -23712
rect 4606 -23878 4658 -23826
rect 6642 -23878 6694 -23826
rect 5624 -23982 5676 -23930
rect 14790 -22608 14842 -22556
rect 7662 -23878 7714 -23826
rect 8678 -23878 8730 -23826
rect 2452 -24880 2504 -24828
rect 2124 -24984 2176 -24932
rect 3588 -24984 3640 -24932
rect 4096 -25090 4148 -25038
rect 1074 -26044 1126 -25992
rect 9698 -23878 9750 -23826
rect 16818 -22608 16870 -22556
rect 17844 -22734 17896 -22682
rect 18856 -22608 18908 -22556
rect 19874 -22734 19926 -22682
rect 21910 -22498 21962 -22446
rect 20896 -22608 20948 -22556
rect 21414 -22604 21466 -22552
rect 22926 -22604 22978 -22552
rect 20400 -22732 20452 -22680
rect 21914 -22732 21966 -22680
rect 11728 -23650 11780 -23598
rect 13770 -23650 13822 -23598
rect 15806 -23650 15858 -23598
rect 11224 -23764 11276 -23712
rect 16312 -23760 16364 -23708
rect 10716 -23878 10768 -23826
rect 12746 -23878 12798 -23826
rect 14784 -23878 14836 -23826
rect 16820 -23878 16872 -23826
rect 10560 -23982 10612 -23930
rect 5622 -24880 5674 -24828
rect 5628 -24984 5680 -24932
rect 5116 -25090 5168 -25038
rect 4608 -25200 4660 -25148
rect 2452 -26122 2504 -26070
rect 3588 -26122 3640 -26070
rect 4100 -26230 4152 -26178
rect 6140 -25090 6192 -25038
rect 7658 -24984 7710 -24932
rect 7158 -25090 7210 -25038
rect 8172 -25090 8224 -25038
rect 6644 -25200 6696 -25148
rect 5114 -26230 5166 -26178
rect 6136 -26230 6188 -26178
rect 9852 -24878 9904 -24826
rect 9698 -24984 9750 -24932
rect 9204 -25090 9256 -25038
rect 8682 -25200 8734 -25148
rect 7658 -26122 7710 -26070
rect 7150 -26230 7202 -26178
rect 8176 -26230 8228 -26178
rect 10216 -25090 10268 -25038
rect 11730 -24878 11782 -24826
rect 11734 -24984 11786 -24932
rect 11224 -25090 11276 -25038
rect 10720 -25200 10772 -25148
rect 9188 -26230 9240 -26178
rect 10224 -26230 10276 -26178
rect 12242 -25090 12294 -25038
rect 16966 -23982 17018 -23930
rect 17842 -23878 17894 -23826
rect 18860 -23650 18912 -23598
rect 18862 -23878 18914 -23826
rect 13768 -24878 13820 -24826
rect 13770 -24984 13822 -24932
rect 13268 -25090 13320 -25038
rect 12756 -25200 12808 -25148
rect 11230 -26230 11282 -26178
rect 12244 -26230 12296 -26178
rect 14270 -25090 14322 -25038
rect 19876 -23878 19928 -23826
rect 19876 -23982 19928 -23930
rect 20892 -23650 20944 -23598
rect 23166 -18714 23218 -18662
rect 23404 -18936 23456 -18884
rect 23282 -19038 23334 -18986
rect 23166 -20272 23218 -20220
rect 23162 -21174 23214 -21122
rect 23282 -22400 23334 -22348
rect 23162 -22498 23214 -22446
rect 23038 -23650 23090 -23598
rect 21412 -23760 21464 -23708
rect 22420 -23760 22472 -23708
rect 23530 -20170 23582 -20118
rect 23532 -22604 23584 -22552
rect 23404 -22732 23456 -22680
rect 23766 -16582 23818 -16530
rect 23654 -23760 23706 -23708
rect 20898 -23878 20950 -23826
rect 15638 -24878 15690 -24826
rect 15290 -25090 15342 -25038
rect 15804 -24984 15856 -24932
rect 14792 -25200 14844 -25148
rect 13260 -26230 13312 -26178
rect 14268 -26230 14320 -26178
rect 16310 -25090 16362 -25038
rect 17844 -24984 17896 -24932
rect 17336 -25090 17388 -25038
rect 18354 -25090 18406 -25038
rect 16824 -25200 16876 -25148
rect 15284 -26230 15336 -26178
rect 16308 -26230 16360 -26178
rect 23058 -23982 23110 -23930
rect 19874 -24984 19926 -24932
rect 19368 -25090 19420 -25038
rect 18856 -25200 18908 -25148
rect 17838 -26122 17890 -26070
rect 17330 -26230 17382 -26178
rect 18352 -26230 18404 -26178
rect 20382 -25090 20434 -25038
rect 21914 -24878 21966 -24826
rect 21914 -24984 21966 -24932
rect 21404 -25090 21456 -25038
rect 20896 -25200 20948 -25148
rect 19370 -26230 19422 -26178
rect 20384 -26230 20436 -26178
rect 23766 -24984 23818 -24932
rect 23058 -26122 23110 -26070
rect 21408 -26230 21460 -26178
rect -8066 -26611 23922 -26495
rect -12198 -27088 -11634 -26844
rect 24234 -27088 24798 -26844
<< metal2 >>
rect 484 4214 1084 4226
rect 484 4188 516 4214
rect 1052 4188 1084 4214
rect 484 3944 502 4188
rect 1066 3944 1084 4188
rect 484 3918 516 3944
rect 1052 3918 1084 3944
rect 484 3906 1084 3918
rect 24116 4214 24716 4226
rect 24116 4188 24148 4214
rect 24684 4188 24716 4214
rect 24116 3944 24134 4188
rect 24698 3944 24716 4188
rect 24116 3918 24148 3944
rect 24684 3918 24716 3944
rect 24116 3906 24716 3918
rect 3998 3817 20878 3866
rect 3998 3795 4075 3817
rect 20831 3795 20878 3817
rect 3998 3659 4065 3795
rect 20841 3659 20878 3795
rect 3998 3637 4075 3659
rect 20831 3637 20878 3659
rect 3998 3600 20878 3637
rect 3998 3598 8352 3600
rect 7986 1918 8046 1924
rect 9068 1918 9128 1924
rect 10026 1918 10086 1924
rect 13090 1918 13150 1924
rect 14108 1918 14168 1924
rect 15132 1918 15192 1924
rect 16144 1918 16204 1924
rect 19202 1918 19262 1924
rect 20214 1918 20274 1924
rect 21232 1918 21292 1924
rect 7986 1914 21292 1918
rect 7986 1862 7990 1914
rect 8042 1862 9072 1914
rect 9124 1862 10030 1914
rect 10082 1862 13094 1914
rect 13146 1862 14112 1914
rect 14164 1862 15136 1914
rect 15188 1862 16148 1914
rect 16200 1862 19206 1914
rect 19258 1862 20218 1914
rect 20270 1862 21236 1914
rect 21288 1862 21292 1914
rect 7986 1858 21292 1862
rect 7986 1852 8046 1858
rect 9068 1852 9128 1858
rect 10026 1852 10086 1858
rect 13090 1852 13150 1858
rect 14108 1852 14168 1858
rect 15132 1852 15192 1858
rect 16144 1852 16204 1858
rect 19202 1852 19262 1858
rect 20214 1852 20274 1858
rect 21232 1852 21292 1858
rect 8512 1672 8572 1678
rect 10548 1672 10608 1678
rect 12586 1674 12646 1680
rect 14616 1674 14676 1680
rect 16658 1676 16718 1682
rect 17668 1676 17728 1682
rect 18690 1676 18750 1682
rect 20726 1676 20786 1682
rect 16658 1674 20786 1676
rect 12586 1672 20786 1674
rect 8512 1670 16662 1672
rect 8512 1668 12590 1670
rect 8512 1616 8516 1668
rect 8568 1616 10552 1668
rect 10604 1618 12590 1668
rect 12642 1618 14620 1670
rect 14672 1620 16662 1670
rect 16714 1620 17672 1672
rect 17724 1620 18694 1672
rect 18746 1620 20730 1672
rect 20782 1620 20786 1672
rect 14672 1618 20786 1620
rect 10604 1616 20786 1618
rect 8512 1614 16856 1616
rect 8512 1612 12768 1614
rect 8512 1606 8572 1612
rect 10548 1606 10608 1612
rect 12586 1608 12646 1612
rect 14616 1608 14676 1614
rect 16658 1610 16718 1614
rect 17668 1610 17728 1616
rect 18690 1610 18750 1616
rect 20726 1610 20786 1616
rect 6330 740 6390 746
rect 7494 740 7554 746
rect 13604 740 13664 746
rect 6330 736 13664 740
rect 6330 684 6334 736
rect 6386 684 7498 736
rect 7550 684 13608 736
rect 13660 684 13664 736
rect 6330 680 13664 684
rect 6330 674 6390 680
rect 7494 674 7554 680
rect 13604 674 13664 680
rect 15638 740 15698 746
rect 21746 740 21806 746
rect 22996 740 23056 746
rect 15638 736 23056 740
rect 15638 684 15642 736
rect 15694 684 21750 736
rect 21802 684 23000 736
rect 23052 684 23056 736
rect 15638 680 23056 684
rect 15638 674 15698 680
rect 21746 674 21806 680
rect 22996 674 23056 680
rect 9530 636 9590 642
rect 11566 636 11626 642
rect 17672 636 17732 642
rect 19706 636 19766 642
rect 9530 632 12044 636
rect 9530 580 9534 632
rect 9586 580 11570 632
rect 11622 628 12044 632
rect 12260 632 19766 636
rect 12260 628 17676 632
rect 11622 582 17676 628
rect 11622 580 14060 582
rect 9530 578 14060 580
rect 9530 576 13034 578
rect 13272 576 14060 578
rect 14276 580 17676 582
rect 17728 580 19710 632
rect 19762 580 19766 632
rect 14276 576 19766 580
rect 9530 570 9590 576
rect 11566 570 11626 576
rect 17672 570 17732 576
rect 19706 570 19766 576
rect 6200 536 6260 542
rect 7494 536 7554 542
rect 13600 536 13660 542
rect 15636 536 15696 542
rect 6200 532 15696 536
rect 6200 480 6204 532
rect 6256 480 7498 532
rect 7550 480 13604 532
rect 13656 480 15640 532
rect 15692 480 15696 532
rect 6200 476 15696 480
rect 6200 470 6260 476
rect 7494 470 7554 476
rect 13600 470 13660 476
rect 15636 470 15696 476
rect 16138 536 16198 542
rect 17158 536 17218 542
rect 18184 536 18244 542
rect 16138 532 18244 536
rect 16138 480 16142 532
rect 16194 480 17162 532
rect 17214 480 18188 532
rect 18240 480 18244 532
rect 16138 476 18244 480
rect 16138 470 16198 476
rect 17158 470 17218 476
rect 18184 470 18244 476
rect 18690 532 18750 538
rect 19204 532 19264 538
rect 19708 532 19768 538
rect 20214 532 20274 538
rect 18690 528 20800 532
rect 18690 476 18694 528
rect 18746 476 19208 528
rect 19260 476 19712 528
rect 19764 476 20218 528
rect 20270 476 20738 528
rect 20790 476 20800 528
rect 18690 472 20800 476
rect 18690 466 18750 472
rect 19204 466 19264 472
rect 19708 466 19768 472
rect 20214 466 20274 472
rect 10546 -398 10606 -392
rect 12580 -398 12640 -392
rect 14618 -398 14678 -394
rect 10030 -400 14822 -398
rect 16654 -400 16714 -394
rect 17154 -400 17214 -394
rect 17668 -400 17728 -394
rect 18192 -400 18252 -394
rect 18690 -400 18750 -394
rect 19192 -400 19252 -394
rect 10030 -402 19560 -400
rect 19706 -402 19766 -396
rect 20214 -402 20274 -396
rect 20724 -402 20784 -396
rect 10030 -454 10040 -402
rect 10092 -454 10550 -402
rect 10602 -454 12584 -402
rect 12636 -404 20784 -402
rect 12636 -454 14622 -404
rect 10030 -456 14622 -454
rect 14674 -456 16658 -404
rect 16710 -456 17158 -404
rect 17210 -456 17672 -404
rect 17724 -456 18196 -404
rect 18248 -456 18694 -404
rect 18746 -456 19196 -404
rect 19248 -406 20784 -404
rect 19248 -456 19710 -406
rect 10030 -458 19710 -456
rect 19762 -458 20218 -406
rect 20270 -458 20728 -406
rect 20780 -458 20784 -406
rect 10546 -464 10606 -458
rect 12580 -464 12640 -458
rect 14618 -460 20784 -458
rect 14618 -466 14678 -460
rect 16654 -466 16714 -460
rect 17154 -466 17214 -460
rect 17668 -466 17728 -460
rect 18192 -466 18252 -460
rect 18589 -462 19104 -460
rect 18690 -466 18750 -462
rect 19192 -466 19252 -460
rect 19354 -462 20784 -460
rect 19706 -468 19766 -462
rect 20214 -468 20274 -462
rect 20724 -468 20784 -462
rect 9528 -496 9592 -490
rect 11404 -496 11468 -490
rect 9528 -502 11468 -496
rect 9528 -554 9534 -502
rect 9586 -554 11410 -502
rect 11462 -554 11468 -502
rect 9528 -560 11468 -554
rect 9528 -566 9592 -560
rect 11404 -566 11468 -560
rect 15638 -498 15698 -492
rect 21746 -498 21806 -492
rect 15638 -502 21806 -498
rect 15638 -554 15642 -502
rect 15694 -554 21750 -502
rect 21802 -554 21806 -502
rect 15638 -558 21806 -554
rect 15638 -564 15698 -558
rect 21746 -564 21806 -558
rect 11040 -606 11100 -600
rect 12064 -606 12124 -600
rect 13092 -606 13152 -600
rect 9018 -614 9078 -608
rect 10030 -614 10090 -608
rect 7974 -618 10090 -614
rect 7974 -670 7984 -618
rect 8036 -670 9022 -618
rect 9074 -670 10034 -618
rect 10086 -670 10090 -618
rect 7974 -674 10090 -670
rect 11040 -610 13152 -606
rect 11040 -662 11044 -610
rect 11096 -662 12068 -610
rect 12120 -662 13096 -610
rect 13148 -662 13152 -610
rect 11040 -666 13152 -662
rect 11040 -672 11100 -666
rect 12064 -672 12124 -666
rect 13092 -672 13152 -666
rect 19196 -614 19256 -608
rect 20208 -614 20268 -608
rect 21210 -614 21270 -608
rect 19196 -618 21270 -614
rect 19196 -670 19200 -618
rect 19252 -670 20212 -618
rect 20264 -670 21214 -618
rect 21266 -670 21270 -618
rect 9018 -680 9078 -674
rect 10030 -680 10090 -674
rect 19196 -674 21270 -670
rect 19196 -680 19256 -674
rect 20208 -680 20268 -674
rect 21210 -680 21270 -674
rect 8510 -1536 8570 -1530
rect 10546 -1536 10606 -1530
rect 11068 -1536 11128 -1530
rect 11566 -1536 11626 -1530
rect 12580 -1536 12640 -1530
rect 13040 -1536 13100 -1530
rect 14078 -1536 14150 -1534
rect 14616 -1536 14676 -1530
rect 16122 -1536 16194 -1534
rect 8510 -1538 16500 -1536
rect 16654 -1538 16714 -1532
rect 18690 -1538 18750 -1534
rect 8510 -1540 14088 -1538
rect 8510 -1592 8514 -1540
rect 8566 -1592 10550 -1540
rect 10602 -1592 11072 -1540
rect 11124 -1592 11570 -1540
rect 11622 -1541 13044 -1540
rect 11622 -1544 12568 -1541
rect 11622 -1592 12044 -1544
rect 8510 -1596 12044 -1592
rect 12096 -1593 12568 -1544
rect 12620 -1592 13044 -1541
rect 13096 -1590 14088 -1540
rect 14140 -1540 16132 -1538
rect 14140 -1590 14620 -1540
rect 13096 -1592 14620 -1590
rect 14672 -1590 16132 -1540
rect 16184 -1540 18878 -1538
rect 20724 -1540 20784 -1534
rect 16184 -1543 20784 -1540
rect 16184 -1590 16642 -1543
rect 14672 -1592 16642 -1590
rect 12620 -1593 16642 -1592
rect 12096 -1595 16642 -1593
rect 16694 -1544 20784 -1543
rect 16694 -1545 18694 -1544
rect 16694 -1548 17659 -1545
rect 16694 -1595 17154 -1548
rect 12096 -1596 17154 -1595
rect 8510 -1602 8570 -1596
rect 10546 -1602 10606 -1596
rect 11068 -1602 11128 -1596
rect 11566 -1602 11626 -1596
rect 12034 -1600 12106 -1596
rect 12542 -1598 12640 -1596
rect 12580 -1602 12640 -1598
rect 13040 -1602 13100 -1596
rect 14616 -1602 14676 -1596
rect 14760 -1598 16086 -1596
rect 16292 -1598 17154 -1596
rect 16616 -1600 16714 -1598
rect 16654 -1604 16714 -1600
rect 17144 -1600 17154 -1598
rect 17206 -1597 17659 -1548
rect 17711 -1548 18694 -1545
rect 17711 -1597 18154 -1548
rect 17206 -1598 18154 -1597
rect 17206 -1600 17216 -1598
rect 17632 -1600 17738 -1598
rect 17144 -1604 17216 -1600
rect 17666 -1602 17738 -1600
rect 18144 -1600 18154 -1598
rect 18206 -1596 18694 -1548
rect 18746 -1596 20728 -1544
rect 20780 -1596 20784 -1544
rect 18206 -1598 20784 -1596
rect 18206 -1600 18216 -1598
rect 18144 -1604 18216 -1600
rect 18690 -1600 20784 -1598
rect 18690 -1606 18750 -1600
rect 20724 -1606 20784 -1600
rect 4192 -1646 4252 -1642
rect 9526 -1646 9590 -1640
rect 19706 -1646 19770 -1640
rect 4190 -1652 19770 -1646
rect 4190 -1704 4196 -1652
rect 4248 -1704 9532 -1652
rect 9584 -1704 19712 -1652
rect 19764 -1704 19770 -1652
rect 4190 -1710 19770 -1704
rect 4192 -1714 4252 -1710
rect 9526 -1716 9590 -1710
rect 19706 -1716 19770 -1710
rect 7488 -1784 7552 -1778
rect 7488 -1790 23062 -1784
rect 7488 -1842 7494 -1790
rect 7546 -1794 22998 -1790
rect 7546 -1842 13604 -1794
rect 7488 -1846 13604 -1842
rect 13656 -1842 22998 -1794
rect 23050 -1842 23062 -1790
rect 13656 -1846 23062 -1842
rect 7488 -1848 23062 -1846
rect 7488 -1854 7552 -1848
rect 13592 -1852 13668 -1848
rect 6330 -1934 6390 -1928
rect 15634 -1934 15698 -1924
rect 21740 -1934 21800 -1928
rect 6330 -1936 21800 -1934
rect 6330 -1938 15640 -1936
rect 6330 -1990 6334 -1938
rect 6386 -1990 7316 -1938
rect 7368 -1988 15640 -1938
rect 15692 -1938 21800 -1936
rect 15692 -1988 21744 -1938
rect 7368 -1990 21744 -1988
rect 21796 -1990 21800 -1938
rect 6330 -1994 21800 -1990
rect 6330 -2000 6390 -1994
rect 15634 -2000 15698 -1994
rect 21740 -2000 21800 -1994
rect 7428 -2040 7488 -2034
rect 7990 -2040 8050 -2034
rect 9032 -2040 9092 -2034
rect 10032 -2040 10092 -2034
rect 13194 -2040 13254 -2034
rect 14204 -2040 14264 -2034
rect 15146 -2040 15206 -2034
rect 7428 -2044 15206 -2040
rect 7428 -2096 7432 -2044
rect 7484 -2096 7994 -2044
rect 8046 -2096 9036 -2044
rect 9088 -2096 10036 -2044
rect 10088 -2096 13198 -2044
rect 13250 -2096 14208 -2044
rect 14260 -2096 15150 -2044
rect 15202 -2096 15206 -2044
rect 7428 -2100 15206 -2096
rect 7428 -2106 7488 -2100
rect 7990 -2106 8050 -2100
rect 9032 -2106 9092 -2100
rect 10032 -2106 10092 -2100
rect 13194 -2106 13254 -2100
rect 14204 -2106 14264 -2100
rect 15146 -2106 15206 -2100
rect 7542 -2242 7602 -2236
rect 10720 -2242 10780 -2236
rect 14788 -2242 14848 -2236
rect 18864 -2242 18924 -2236
rect 22060 -2242 22120 -2236
rect 7542 -2246 22120 -2242
rect 7542 -2298 7546 -2246
rect 7598 -2298 10724 -2246
rect 10776 -2298 14792 -2246
rect 14844 -2298 18868 -2246
rect 18920 -2298 22064 -2246
rect 22116 -2298 22120 -2246
rect 7542 -2302 22120 -2298
rect 7542 -2308 7602 -2302
rect 10720 -2308 10780 -2302
rect 14788 -2308 14848 -2302
rect 18864 -2308 18924 -2302
rect 22060 -2308 22120 -2302
rect 8686 -3178 8746 -3172
rect 10720 -3178 10780 -3172
rect 12762 -3178 12822 -3172
rect 14788 -3178 14848 -3172
rect 16830 -3178 16890 -3172
rect 18866 -3178 18926 -3172
rect 20902 -3178 20962 -3172
rect 8686 -3182 20962 -3178
rect 8686 -3234 8690 -3182
rect 8742 -3234 10724 -3182
rect 10776 -3234 12766 -3182
rect 12818 -3234 14792 -3182
rect 14844 -3234 16834 -3182
rect 16886 -3234 18870 -3182
rect 18922 -3234 20906 -3182
rect 20958 -3234 20962 -3182
rect 8686 -3238 20962 -3234
rect 8686 -3244 8746 -3238
rect 10720 -3244 10780 -3238
rect 12762 -3244 12822 -3238
rect 14788 -3244 14848 -3238
rect 16830 -3244 16890 -3238
rect 18866 -3244 18926 -3238
rect 20902 -3244 20962 -3238
rect 9190 -3286 9250 -3280
rect 9190 -3290 20462 -3286
rect 9190 -3342 9194 -3290
rect 9246 -3342 10216 -3290
rect 10268 -3342 11234 -3290
rect 11286 -3342 12258 -3290
rect 12310 -3342 13272 -3290
rect 13324 -3342 14290 -3290
rect 14342 -3342 15300 -3290
rect 15352 -3342 16322 -3290
rect 16374 -3342 17336 -3290
rect 17388 -3342 18368 -3290
rect 18420 -3342 19378 -3290
rect 19430 -3342 20400 -3290
rect 20452 -3342 20462 -3290
rect 9190 -3346 20462 -3342
rect 9190 -3352 9250 -3346
rect 8682 -4210 8742 -4204
rect 12762 -4210 12822 -4204
rect 16830 -4210 16890 -4204
rect 20898 -4210 20958 -4204
rect 23290 -4210 23350 -4204
rect 1150 -4214 23350 -4210
rect 1150 -4266 8686 -4214
rect 8738 -4266 12766 -4214
rect 12818 -4266 16834 -4214
rect 16886 -4266 20902 -4214
rect 20954 -4266 23294 -4214
rect 23346 -4266 23350 -4214
rect 1150 -4270 23350 -4266
rect -13992 -10402 -2722 -10122
rect -13992 -10646 -13618 -10402
rect -2878 -10646 -2722 -10402
rect -13992 -10978 -2722 -10646
rect -13992 -11300 -1640 -10978
rect 1150 -11626 1210 -4270
rect 8682 -4276 8742 -4270
rect 12762 -4276 12822 -4270
rect 16830 -4276 16890 -4270
rect 20898 -4276 20958 -4270
rect 23290 -4276 23350 -4270
rect 6686 -4342 6746 -4336
rect 11228 -4342 11300 -4340
rect 12226 -4342 12298 -4340
rect 13270 -4342 13342 -4340
rect 17326 -4342 17398 -4340
rect 22854 -4342 22914 -4336
rect 6686 -4344 22914 -4342
rect 6686 -4346 11238 -4344
rect 6686 -4398 6690 -4346
rect 6742 -4348 11238 -4346
rect 6742 -4398 9192 -4348
rect 6686 -4400 9192 -4398
rect 9244 -4352 11238 -4348
rect 9244 -4400 10206 -4352
rect 6686 -4402 10206 -4400
rect 6686 -4408 6746 -4402
rect 9182 -4404 9254 -4402
rect 10196 -4404 10206 -4402
rect 10258 -4396 11238 -4352
rect 11290 -4396 12236 -4344
rect 12288 -4396 13280 -4344
rect 13332 -4348 17336 -4344
rect 13332 -4396 14284 -4348
rect 10258 -4400 14284 -4396
rect 14336 -4400 15300 -4348
rect 15352 -4400 16304 -4348
rect 16356 -4396 17336 -4348
rect 17388 -4346 22914 -4344
rect 17388 -4348 22858 -4346
rect 17388 -4396 18352 -4348
rect 16356 -4400 18352 -4396
rect 18404 -4400 19380 -4348
rect 19432 -4400 20400 -4348
rect 20452 -4398 22858 -4348
rect 22910 -4398 22914 -4346
rect 20452 -4400 22914 -4398
rect 10258 -4402 22914 -4400
rect 10258 -4404 10268 -4402
rect 14274 -4404 14346 -4402
rect 15290 -4404 15362 -4402
rect 16294 -4404 16366 -4402
rect 18342 -4404 18414 -4402
rect 19370 -4404 19442 -4402
rect 20390 -4404 20462 -4402
rect 10196 -4408 10268 -4404
rect 22854 -4408 22914 -4402
rect 14080 -4552 14140 -4546
rect 14080 -4556 15882 -4552
rect 14080 -4608 14084 -4556
rect 14136 -4608 15820 -4556
rect 15872 -4608 15882 -4556
rect 21714 -4566 21774 -4562
rect 14080 -4612 15882 -4608
rect 21712 -4570 23056 -4566
rect 21712 -4572 23062 -4570
rect 14080 -4618 14140 -4612
rect 21712 -4624 21718 -4572
rect 21770 -4574 23062 -4572
rect 21770 -4624 23000 -4574
rect 21712 -4626 23000 -4624
rect 23052 -4626 23062 -4574
rect 21712 -4630 23062 -4626
rect 21714 -4634 21774 -4630
rect 15096 -4748 15160 -4742
rect 19160 -4748 19224 -4742
rect 20184 -4748 20248 -4742
rect 21196 -4748 21260 -4742
rect 15096 -4754 21260 -4748
rect 15096 -4806 15102 -4754
rect 15154 -4806 19166 -4754
rect 19218 -4806 20190 -4754
rect 20242 -4806 21202 -4754
rect 21254 -4806 21260 -4754
rect 15096 -4812 21260 -4806
rect 15096 -4818 15160 -4812
rect 19160 -4818 19224 -4812
rect 20184 -4818 20248 -4812
rect 21196 -4818 21260 -4812
rect 7312 -4870 7372 -4864
rect 8478 -4870 8538 -4864
rect 10514 -4870 10574 -4864
rect 7312 -4874 10574 -4870
rect 7312 -4926 7316 -4874
rect 7368 -4926 8482 -4874
rect 8534 -4926 10518 -4874
rect 10570 -4926 10574 -4874
rect 7312 -4930 10574 -4926
rect 7312 -4936 7372 -4930
rect 8478 -4936 8538 -4930
rect 10514 -4936 10574 -4930
rect 11022 -4870 11086 -4864
rect 15098 -4870 15162 -4864
rect 11022 -4876 15162 -4870
rect 11022 -4928 11028 -4876
rect 11080 -4928 15104 -4876
rect 15156 -4928 15162 -4876
rect 11022 -4934 15162 -4928
rect 11022 -4940 11086 -4934
rect 15098 -4940 15162 -4934
rect 18660 -4870 18720 -4864
rect 20694 -4870 20754 -4864
rect 23138 -4870 23198 -4864
rect 18660 -4874 23198 -4870
rect 18660 -4926 18664 -4874
rect 18716 -4926 20698 -4874
rect 20750 -4926 23142 -4874
rect 23194 -4926 23198 -4874
rect 18660 -4930 23198 -4926
rect 18660 -4936 18720 -4930
rect 20694 -4936 20754 -4930
rect 23138 -4936 23198 -4930
rect 6560 -4952 6620 -4946
rect 6802 -4952 6862 -4946
rect 6560 -4956 6862 -4952
rect 6560 -5008 6564 -4956
rect 6616 -5008 6806 -4956
rect 6858 -5008 6862 -4956
rect 6560 -5012 6862 -5008
rect 6560 -5018 6620 -5012
rect 6802 -5018 6862 -5012
rect 9496 -5818 9556 -5812
rect 11532 -5818 11592 -5812
rect 9496 -5822 11592 -5818
rect 9496 -5874 9500 -5822
rect 9552 -5874 11536 -5822
rect 11588 -5874 11592 -5822
rect 9496 -5878 11592 -5874
rect 9496 -5884 9556 -5878
rect 11532 -5884 11592 -5878
rect 11874 -5816 11934 -5810
rect 14588 -5816 14648 -5810
rect 11874 -5820 14648 -5816
rect 11874 -5872 11878 -5820
rect 11930 -5872 14592 -5820
rect 14644 -5872 14648 -5820
rect 11874 -5876 14648 -5872
rect 11874 -5882 11934 -5876
rect 14588 -5882 14648 -5876
rect 19676 -5818 19736 -5812
rect 21712 -5818 21772 -5812
rect 19676 -5822 21772 -5818
rect 19676 -5874 19680 -5822
rect 19732 -5874 21716 -5822
rect 21768 -5874 21772 -5822
rect 19676 -5878 21772 -5874
rect 19676 -5884 19736 -5878
rect 3676 -5906 3736 -5900
rect 4698 -5906 4758 -5900
rect 3676 -5910 4758 -5906
rect 3676 -5962 3680 -5910
rect 3732 -5962 4702 -5910
rect 4754 -5962 4758 -5910
rect 3676 -5966 4758 -5962
rect 3676 -5972 3736 -5966
rect 4698 -5972 4758 -5966
rect 7044 -5916 7104 -5910
rect 19784 -5916 19844 -5878
rect 21712 -5884 21772 -5878
rect 7044 -5920 19844 -5916
rect 7044 -5972 7048 -5920
rect 7100 -5972 19844 -5920
rect 7044 -5976 19844 -5972
rect 7044 -5982 7104 -5976
rect 3784 -6018 3844 -6012
rect 4568 -6018 4628 -6012
rect 3784 -6022 4628 -6018
rect 3784 -6074 3788 -6022
rect 3840 -6074 4572 -6022
rect 4624 -6074 4628 -6022
rect 3784 -6078 4628 -6074
rect 3784 -6084 3844 -6078
rect 4568 -6084 4628 -6078
rect 7180 -6014 7240 -6008
rect 9496 -6014 9556 -6008
rect 7180 -6018 9556 -6014
rect 7180 -6070 7184 -6018
rect 7236 -6070 9500 -6018
rect 9552 -6070 9556 -6018
rect 7180 -6074 9556 -6070
rect 7180 -6080 7240 -6074
rect 9496 -6080 9556 -6074
rect 10516 -6012 10576 -6006
rect 15606 -6012 15666 -6006
rect 22978 -6012 23038 -6006
rect 10516 -6016 23038 -6012
rect 10516 -6068 10520 -6016
rect 10572 -6068 15610 -6016
rect 15662 -6068 22982 -6016
rect 23034 -6068 23038 -6016
rect 10516 -6072 23038 -6068
rect 10516 -6078 10576 -6072
rect 15606 -6078 15666 -6072
rect 22978 -6078 23038 -6072
rect 8482 -6124 8542 -6118
rect 10516 -6124 10576 -6118
rect 8482 -6128 10576 -6124
rect 8482 -6180 8486 -6128
rect 8538 -6180 10520 -6128
rect 10572 -6180 10576 -6128
rect 8482 -6184 10576 -6180
rect 8482 -6190 8542 -6184
rect 10516 -6190 10576 -6184
rect 13572 -6126 13632 -6120
rect 15606 -6126 15666 -6120
rect 13572 -6130 15666 -6126
rect 13572 -6182 13576 -6130
rect 13628 -6182 15610 -6130
rect 15662 -6182 15666 -6130
rect 13572 -6186 15666 -6182
rect 13572 -6192 13632 -6186
rect 15606 -6192 15666 -6186
rect 18662 -6126 18722 -6120
rect 20696 -6124 20756 -6120
rect 20628 -6126 20756 -6124
rect 23290 -6126 23350 -6120
rect 18662 -6130 23350 -6126
rect 18662 -6182 18666 -6130
rect 18718 -6182 20700 -6130
rect 20752 -6182 23294 -6130
rect 23346 -6182 23350 -6130
rect 18662 -6186 23350 -6182
rect 18662 -6192 18722 -6186
rect 20628 -6188 20756 -6186
rect 20696 -6192 20756 -6188
rect 23290 -6192 23350 -6186
rect 2014 -6940 2074 -6934
rect 5208 -6940 5268 -6934
rect 2014 -6944 5268 -6940
rect 2014 -6996 2018 -6944
rect 2070 -6996 5212 -6944
rect 5264 -6996 5268 -6944
rect 2014 -7000 5268 -6996
rect 2014 -7006 2074 -7000
rect 5208 -7006 5268 -7000
rect 3174 -7050 3234 -7044
rect 6360 -7050 6420 -7044
rect 3174 -7054 6420 -7050
rect 3174 -7106 3178 -7054
rect 3230 -7106 6364 -7054
rect 6416 -7106 6420 -7054
rect 19526 -7060 19586 -7054
rect 19526 -7064 23948 -7060
rect 3174 -7110 6420 -7106
rect 3174 -7116 3234 -7110
rect 6360 -7116 6420 -7110
rect 6802 -7074 6862 -7068
rect 13568 -7074 13628 -7068
rect 14588 -7074 14648 -7068
rect 16624 -7074 16684 -7068
rect 6802 -7078 16684 -7074
rect 6802 -7130 6806 -7078
rect 6858 -7130 13572 -7078
rect 13624 -7130 14592 -7078
rect 14644 -7130 16628 -7078
rect 16680 -7130 16684 -7078
rect 19526 -7116 19530 -7064
rect 19582 -7116 23948 -7064
rect 19526 -7120 23948 -7116
rect 19526 -7126 19586 -7120
rect 6802 -7134 16684 -7130
rect 6802 -7140 6862 -7134
rect 13568 -7140 13628 -7134
rect 14588 -7140 14648 -7134
rect 16624 -7140 16684 -7134
rect 19674 -7170 19734 -7164
rect 21714 -7170 21774 -7164
rect 22854 -7170 22914 -7164
rect 6552 -7178 6612 -7172
rect 11534 -7178 11594 -7172
rect 18658 -7178 18718 -7172
rect 6552 -7182 18718 -7178
rect 6552 -7234 6556 -7182
rect 6608 -7234 9502 -7182
rect 9554 -7234 11538 -7182
rect 11590 -7234 18662 -7182
rect 18714 -7234 18718 -7182
rect 6552 -7238 18718 -7234
rect 19674 -7174 22914 -7170
rect 19674 -7226 19678 -7174
rect 19730 -7226 21718 -7174
rect 21770 -7226 22858 -7174
rect 22910 -7226 22914 -7174
rect 19674 -7230 22914 -7226
rect 19674 -7236 19734 -7230
rect 21714 -7236 21774 -7230
rect 22854 -7236 22914 -7230
rect 6552 -7244 6612 -7238
rect 11534 -7244 11594 -7238
rect 18658 -7244 18718 -7238
rect 11532 -7280 11592 -7274
rect 20694 -7280 20754 -7274
rect 6798 -7288 6858 -7282
rect 7464 -7288 7524 -7282
rect 6798 -7292 7524 -7288
rect 6798 -7344 6802 -7292
rect 6854 -7344 7468 -7292
rect 7520 -7344 7524 -7292
rect 6798 -7348 7524 -7344
rect 11532 -7284 20754 -7280
rect 11532 -7336 11536 -7284
rect 11588 -7336 20698 -7284
rect 20750 -7336 20754 -7284
rect 11532 -7340 20754 -7336
rect 11532 -7346 11592 -7340
rect 20694 -7346 20754 -7340
rect 6798 -7354 6858 -7348
rect 7464 -7354 7524 -7348
rect 9498 -7382 9558 -7376
rect 11532 -7382 11592 -7376
rect 9498 -7386 11592 -7382
rect 9498 -7438 9502 -7386
rect 9554 -7438 11536 -7386
rect 11588 -7438 11592 -7386
rect 9498 -7442 11592 -7438
rect 9498 -7448 9558 -7442
rect 11532 -7448 11592 -7442
rect 14588 -7380 14648 -7374
rect 15606 -7380 15666 -7374
rect 16622 -7380 16682 -7374
rect 19526 -7380 19586 -7374
rect 14588 -7384 19586 -7380
rect 14588 -7436 14592 -7384
rect 14644 -7436 15610 -7384
rect 15662 -7436 16626 -7384
rect 16678 -7436 19530 -7384
rect 19582 -7436 19586 -7384
rect 14588 -7440 19586 -7436
rect 14588 -7446 14648 -7440
rect 15606 -7446 15666 -7440
rect 16622 -7446 16682 -7440
rect 19526 -7446 19586 -7440
rect 19678 -7378 19738 -7372
rect 21712 -7378 21772 -7372
rect 22978 -7378 23038 -7372
rect 19678 -7382 23820 -7378
rect 19678 -7434 19682 -7382
rect 19734 -7434 21716 -7382
rect 21768 -7434 22982 -7382
rect 23034 -7434 23820 -7382
rect 19678 -7438 23820 -7434
rect 19678 -7444 19738 -7438
rect 21712 -7444 21772 -7438
rect 22978 -7444 23038 -7438
rect 3690 -7974 3750 -7968
rect 4700 -7974 4760 -7968
rect 3690 -7978 4760 -7974
rect 1882 -8032 1954 -8028
rect 1882 -8084 1892 -8032
rect 1944 -8084 1954 -8032
rect 3690 -8030 3694 -7978
rect 3746 -8030 4704 -7978
rect 4756 -8030 4760 -7978
rect 3690 -8034 4760 -8030
rect 3690 -8040 3750 -8034
rect 4700 -8040 4760 -8034
rect 1882 -8088 1954 -8084
rect 3796 -8074 3856 -8068
rect 4582 -8074 4642 -8068
rect 3796 -8078 4642 -8074
rect 1396 -9088 1468 -9084
rect 1396 -9140 1406 -9088
rect 1458 -9140 1468 -9088
rect 1396 -9144 1468 -9140
rect 1276 -9588 1348 -9584
rect 1276 -9640 1286 -9588
rect 1338 -9640 1348 -9588
rect 1276 -9644 1348 -9640
rect 1282 -11498 1342 -9644
rect 1282 -11550 1286 -11498
rect 1338 -11550 1342 -11498
rect 1282 -11560 1342 -11550
rect 1402 -11496 1462 -9144
rect 1536 -9264 1608 -9260
rect 1536 -9316 1546 -9264
rect 1598 -9316 1608 -9264
rect 1536 -9320 1608 -9316
rect 1402 -11548 1406 -11496
rect 1458 -11548 1462 -11496
rect 1542 -11478 1602 -9320
rect 1764 -10086 1836 -10082
rect 1764 -10138 1774 -10086
rect 1826 -10138 1836 -10086
rect 1764 -10142 1836 -10138
rect 1542 -11530 1546 -11478
rect 1598 -11530 1602 -11478
rect 1770 -11462 1830 -10142
rect 1888 -11358 1948 -8088
rect 3796 -8130 3800 -8078
rect 3852 -8130 4586 -8078
rect 4638 -8130 4642 -8078
rect 3796 -8134 4642 -8130
rect 3796 -8140 3856 -8134
rect 4582 -8140 4642 -8134
rect 11534 -8322 11594 -8316
rect 13336 -8322 13396 -8316
rect 6686 -8330 6746 -8324
rect 8480 -8330 8540 -8324
rect 10516 -8330 10576 -8324
rect 6686 -8334 10576 -8330
rect 6686 -8386 6690 -8334
rect 6742 -8386 8484 -8334
rect 8536 -8386 10520 -8334
rect 10572 -8386 10576 -8334
rect 6686 -8390 10576 -8386
rect 11534 -8326 13396 -8322
rect 11534 -8378 11538 -8326
rect 11590 -8378 13340 -8326
rect 13392 -8378 13396 -8326
rect 11534 -8382 13396 -8378
rect 11534 -8388 11594 -8382
rect 13336 -8388 13396 -8382
rect 13570 -8328 13630 -8322
rect 15606 -8328 15666 -8322
rect 13570 -8332 15666 -8328
rect 13570 -8384 13574 -8332
rect 13626 -8384 15610 -8332
rect 15662 -8384 15666 -8332
rect 13570 -8388 15666 -8384
rect 6686 -8396 6746 -8390
rect 2436 -9438 2508 -9434
rect 2436 -9490 2446 -9438
rect 2498 -9490 2508 -9438
rect 2436 -9494 2508 -9490
rect 2330 -9850 2402 -9846
rect 2330 -9902 2340 -9850
rect 2392 -9902 2402 -9850
rect 2330 -9906 2402 -9902
rect 2210 -9968 2282 -9964
rect 2210 -10020 2220 -9968
rect 2272 -10020 2282 -9968
rect 2210 -10024 2282 -10020
rect 2216 -11352 2276 -10024
rect 2336 -10940 2396 -9906
rect 2319 -10966 2409 -10940
rect 2319 -11022 2336 -10966
rect 2392 -11022 2409 -10966
rect 2319 -11048 2409 -11022
rect 1882 -11362 1954 -11358
rect 1882 -11414 1892 -11362
rect 1944 -11414 1954 -11362
rect 2216 -11404 2220 -11352
rect 2272 -11404 2276 -11352
rect 2336 -11356 2396 -11048
rect 2216 -11414 2276 -11404
rect 2330 -11360 2402 -11356
rect 2330 -11412 2340 -11360
rect 2392 -11412 2402 -11360
rect 1882 -11418 1954 -11414
rect 2330 -11416 2402 -11412
rect 1770 -11514 1774 -11462
rect 1826 -11514 1830 -11462
rect 2442 -11492 2502 -9494
rect 1770 -11524 1830 -11514
rect 2436 -11496 2508 -11492
rect 1542 -11540 1602 -11530
rect 1402 -11558 1462 -11548
rect 2436 -11548 2446 -11496
rect 2498 -11548 2508 -11496
rect 2436 -11552 2508 -11548
rect 1150 -11678 1154 -11626
rect 1206 -11678 1210 -11626
rect 1660 -11612 1720 -11606
rect 6914 -11612 6974 -8390
rect 8480 -8396 8540 -8390
rect 10516 -8396 10576 -8390
rect 13570 -8394 13630 -8388
rect 15606 -8394 15666 -8388
rect 18660 -8326 18720 -8320
rect 20696 -8326 20756 -8320
rect 18660 -8330 20756 -8326
rect 18660 -8382 18664 -8330
rect 18716 -8382 20700 -8330
rect 20752 -8382 20756 -8330
rect 18660 -8386 20756 -8382
rect 18660 -8392 18720 -8386
rect 20696 -8392 20756 -8386
rect 10516 -8438 10576 -8432
rect 15604 -8438 15664 -8432
rect 22854 -8438 22914 -8432
rect 10516 -8442 22914 -8438
rect 10516 -8494 10520 -8442
rect 10572 -8494 15608 -8442
rect 15660 -8494 22858 -8442
rect 22910 -8494 22914 -8442
rect 10516 -8498 22914 -8494
rect 10516 -8504 10576 -8498
rect 15604 -8504 15664 -8498
rect 22854 -8504 22914 -8498
rect 7312 -8538 7372 -8532
rect 7312 -8542 19896 -8538
rect 7312 -8594 7316 -8542
rect 7368 -8594 19896 -8542
rect 7312 -8598 19896 -8594
rect 7312 -8604 7372 -8598
rect 9494 -8640 9554 -8634
rect 11528 -8640 11588 -8634
rect 9494 -8644 11588 -8640
rect 9494 -8696 9498 -8644
rect 9550 -8696 11532 -8644
rect 11584 -8696 11588 -8644
rect 19682 -8640 19742 -8634
rect 19836 -8640 19896 -8598
rect 21716 -8640 21776 -8634
rect 19682 -8644 21776 -8640
rect 9494 -8700 11588 -8696
rect 9494 -8706 9554 -8700
rect 11528 -8706 11588 -8700
rect 11732 -8652 11792 -8646
rect 11732 -8656 19236 -8652
rect 11732 -8708 11736 -8656
rect 11788 -8708 15098 -8656
rect 15150 -8708 16114 -8656
rect 16166 -8708 19174 -8656
rect 19226 -8708 19236 -8656
rect 19682 -8696 19686 -8644
rect 19738 -8696 21720 -8644
rect 21772 -8696 21776 -8644
rect 19682 -8700 21776 -8696
rect 19682 -8706 19742 -8700
rect 21716 -8706 21776 -8700
rect 11732 -8712 19236 -8708
rect 11732 -8718 11792 -8712
rect 7044 -9588 7104 -9582
rect 8476 -9588 8536 -9582
rect 10512 -9588 10572 -9582
rect 7044 -9592 10572 -9588
rect 7044 -9644 7048 -9592
rect 7100 -9644 8480 -9592
rect 8532 -9644 10516 -9592
rect 10568 -9644 10572 -9592
rect 7044 -9648 10572 -9644
rect 7044 -9654 7104 -9648
rect 8476 -9654 8536 -9648
rect 10512 -9654 10572 -9648
rect 18664 -9588 18724 -9582
rect 20700 -9588 20760 -9582
rect 18664 -9592 20760 -9588
rect 18664 -9644 18668 -9592
rect 18720 -9644 20704 -9592
rect 20756 -9644 20760 -9592
rect 18664 -9648 20760 -9644
rect 18664 -9654 18724 -9648
rect 7180 -9718 7240 -9712
rect 18794 -9718 18854 -9648
rect 20700 -9654 20760 -9648
rect 7180 -9722 18854 -9718
rect 7180 -9774 7184 -9722
rect 7236 -9774 18854 -9722
rect 7180 -9778 18854 -9774
rect 7180 -9784 7240 -9778
rect 11534 -9858 11594 -9852
rect 23138 -9858 23198 -9852
rect 11534 -9862 23198 -9858
rect 11534 -9914 11538 -9862
rect 11590 -9914 23142 -9862
rect 23194 -9914 23198 -9862
rect 11534 -9918 23198 -9914
rect 11534 -9924 11594 -9918
rect 1660 -11616 6974 -11612
rect 1660 -11668 1664 -11616
rect 1716 -11668 6974 -11616
rect 1660 -11672 6974 -11668
rect 1660 -11678 1720 -11672
rect 1150 -11688 1210 -11678
rect 13254 -11846 13314 -9918
rect 13254 -11898 13258 -11846
rect 13310 -11898 13314 -11846
rect 13254 -11908 13314 -11898
rect 18358 -11846 18418 -9918
rect 18358 -11898 18362 -11846
rect 18414 -11898 18418 -11846
rect 22418 -11848 22478 -9918
rect 23138 -9924 23198 -9918
rect 18358 -11908 18418 -11898
rect 22412 -11852 22484 -11848
rect 22412 -11904 22422 -11852
rect 22474 -11904 22484 -11852
rect 22412 -11908 22484 -11904
rect -1562 -12220 -1502 -12214
rect 2216 -12220 2276 -12214
rect -1562 -12224 2276 -12220
rect -1562 -12276 -1558 -12224
rect -1506 -12276 2220 -12224
rect 2272 -12276 2276 -12224
rect -1562 -12280 2276 -12276
rect -1562 -12286 -1502 -12280
rect 2216 -12286 2276 -12280
rect -36 -12354 24 -12348
rect 1770 -12354 1830 -12348
rect -36 -12358 1830 -12354
rect -36 -12410 -32 -12358
rect 20 -12410 1774 -12358
rect 1826 -12410 1830 -12358
rect -36 -12414 1830 -12410
rect -36 -12420 24 -12414
rect 1770 -12420 1830 -12414
rect 2012 -13578 2072 -13572
rect 2012 -13582 3652 -13578
rect 2012 -13634 2016 -13582
rect 2068 -13634 3590 -13582
rect 3642 -13634 3652 -13582
rect 2012 -13638 3652 -13634
rect 2012 -13644 2072 -13638
rect 4600 -13794 4660 -13788
rect 6640 -13794 6700 -13788
rect 8680 -13794 8740 -13788
rect 10710 -13794 10770 -13788
rect 12750 -13794 12810 -13788
rect 14782 -13794 14842 -13788
rect 16822 -13794 16882 -13788
rect 18858 -13794 18918 -13788
rect 20892 -13794 20952 -13788
rect 4600 -13798 20952 -13794
rect 4600 -13850 4604 -13798
rect 4656 -13850 6644 -13798
rect 6696 -13850 8684 -13798
rect 8736 -13850 10714 -13798
rect 10766 -13850 12754 -13798
rect 12806 -13850 14786 -13798
rect 14838 -13850 16826 -13798
rect 16878 -13850 18862 -13798
rect 18914 -13850 20896 -13798
rect 20948 -13850 20952 -13798
rect 4600 -13854 20952 -13850
rect 4600 -13860 4660 -13854
rect 6640 -13860 6700 -13854
rect 8680 -13860 8740 -13854
rect 10710 -13860 10770 -13854
rect 12750 -13860 12810 -13854
rect 14782 -13860 14842 -13854
rect 16822 -13860 16882 -13854
rect 18858 -13860 18918 -13854
rect 20892 -13860 20952 -13854
rect 2224 -13914 2284 -13908
rect 2568 -13914 2628 -13908
rect 2224 -13918 2628 -13914
rect 2224 -13970 2228 -13918
rect 2280 -13970 2572 -13918
rect 2624 -13970 2628 -13918
rect 2224 -13974 2628 -13970
rect 2224 -13980 2284 -13974
rect 2568 -13980 2628 -13974
rect 4092 -13920 4152 -13914
rect 12236 -13920 12296 -13914
rect 4092 -13924 21466 -13920
rect 4092 -13976 4096 -13924
rect 4148 -13976 5110 -13924
rect 5162 -13976 6132 -13924
rect 6184 -13976 7146 -13924
rect 7198 -13976 8172 -13924
rect 8224 -13976 9184 -13924
rect 9236 -13976 10220 -13924
rect 10272 -13976 11226 -13924
rect 11278 -13976 12240 -13924
rect 12292 -13976 13256 -13924
rect 13308 -13976 14264 -13924
rect 14316 -13976 15280 -13924
rect 15332 -13976 16304 -13924
rect 16356 -13976 17326 -13924
rect 17378 -13976 18348 -13924
rect 18400 -13976 19366 -13924
rect 19418 -13976 20380 -13924
rect 20432 -13976 21404 -13924
rect 21456 -13976 21466 -13924
rect 4092 -13980 21466 -13976
rect 4092 -13986 4152 -13980
rect 12236 -13986 12296 -13980
rect 2442 -14036 2502 -14030
rect 7656 -14036 7716 -14030
rect 17844 -14036 17904 -14030
rect 21916 -14036 21976 -14030
rect 23048 -14036 23108 -14030
rect 2442 -14040 23108 -14036
rect 2442 -14092 2446 -14040
rect 2498 -14092 7660 -14040
rect 7712 -14092 17848 -14040
rect 17900 -14092 21920 -14040
rect 21972 -14092 23052 -14040
rect 23104 -14092 23108 -14040
rect 2442 -14096 23108 -14092
rect 2442 -14102 2502 -14096
rect 7656 -14102 7716 -14096
rect 17844 -14102 17904 -14096
rect 21916 -14102 21976 -14096
rect 23048 -14102 23108 -14096
rect 4604 -14958 4664 -14952
rect 6644 -14958 6704 -14952
rect 8676 -14958 8736 -14952
rect 10708 -14958 10768 -14952
rect 12744 -14958 12804 -14952
rect 14780 -14958 14840 -14952
rect 16818 -14958 16878 -14952
rect 18856 -14958 18916 -14952
rect 20892 -14958 20952 -14952
rect 4604 -14962 20952 -14958
rect 4604 -15014 4608 -14962
rect 4660 -15014 6648 -14962
rect 6700 -15014 8680 -14962
rect 8732 -15014 10712 -14962
rect 10764 -15014 12748 -14962
rect 12800 -15014 14784 -14962
rect 14836 -15014 16822 -14962
rect 16874 -15014 18860 -14962
rect 18912 -15014 20896 -14962
rect 20948 -15014 20952 -14962
rect 4604 -15018 20952 -15014
rect 4604 -15024 4664 -15018
rect 6644 -15024 6704 -15018
rect 8676 -15024 8736 -15018
rect 10708 -15024 10768 -15018
rect 12744 -15024 12804 -15018
rect 14780 -15024 14840 -15018
rect 16818 -15024 16878 -15018
rect 18856 -15024 18916 -15018
rect 20892 -15024 20952 -15018
rect 4096 -15068 4156 -15062
rect 5118 -15068 5178 -15062
rect 6132 -15068 6192 -15062
rect 7146 -15068 7206 -15062
rect 8164 -15068 8224 -15062
rect 9190 -15068 9250 -15062
rect 10210 -15068 10270 -15062
rect 11230 -15068 11290 -15062
rect 12232 -15068 12292 -15062
rect 13258 -15068 13318 -15062
rect 14276 -15068 14336 -15062
rect 15284 -15068 15344 -15062
rect 16296 -15068 16356 -15062
rect 17328 -15068 17388 -15062
rect 18342 -15068 18402 -15062
rect 19360 -15068 19420 -15062
rect 20384 -15068 20444 -15062
rect 21404 -15068 21464 -15062
rect 4096 -15072 21464 -15068
rect 4096 -15124 4100 -15072
rect 4152 -15124 5122 -15072
rect 5174 -15124 6136 -15072
rect 6188 -15124 7150 -15072
rect 7202 -15124 8168 -15072
rect 8220 -15124 9194 -15072
rect 9246 -15124 10214 -15072
rect 10266 -15124 11234 -15072
rect 11286 -15124 12236 -15072
rect 12288 -15124 13262 -15072
rect 13314 -15124 14280 -15072
rect 14332 -15124 15288 -15072
rect 15340 -15124 16300 -15072
rect 16352 -15124 17332 -15072
rect 17384 -15124 18346 -15072
rect 18398 -15124 19364 -15072
rect 19416 -15124 20388 -15072
rect 20440 -15124 21408 -15072
rect 21460 -15124 21464 -15072
rect 4096 -15128 21464 -15124
rect 4096 -15134 4156 -15128
rect 5118 -15134 5178 -15128
rect 6132 -15134 6192 -15128
rect 7146 -15134 7206 -15128
rect 8164 -15134 8224 -15128
rect 9190 -15134 9250 -15128
rect 10210 -15134 10270 -15128
rect 11230 -15134 11290 -15128
rect 12232 -15134 12292 -15128
rect 13258 -15134 13318 -15128
rect 14276 -15134 14336 -15128
rect 15284 -15134 15344 -15128
rect 16296 -15134 16356 -15128
rect 17328 -15134 17388 -15128
rect 18342 -15134 18402 -15128
rect 19360 -15134 19420 -15128
rect 20384 -15134 20444 -15128
rect 21404 -15134 21464 -15128
rect 2120 -15174 2180 -15168
rect 3586 -15174 3646 -15168
rect 5626 -15174 5686 -15168
rect 7656 -15174 7716 -15168
rect 9696 -15174 9756 -15168
rect 11730 -15174 11790 -15168
rect 13766 -15174 13826 -15168
rect 15802 -15174 15862 -15168
rect 17842 -15174 17902 -15168
rect 19872 -15174 19932 -15168
rect 21912 -15174 21972 -15168
rect 2120 -15178 21972 -15174
rect 2120 -15230 2124 -15178
rect 2176 -15230 3590 -15178
rect 3642 -15230 5630 -15178
rect 5682 -15230 7660 -15178
rect 7712 -15230 9700 -15178
rect 9752 -15230 11734 -15178
rect 11786 -15230 13770 -15178
rect 13822 -15230 15806 -15178
rect 15858 -15230 17846 -15178
rect 17898 -15230 19876 -15178
rect 19928 -15230 21916 -15178
rect 21968 -15230 21972 -15178
rect 2120 -15234 21972 -15230
rect 2120 -15240 2180 -15234
rect 3586 -15240 3646 -15234
rect 5626 -15240 5686 -15234
rect 7656 -15240 7716 -15234
rect 9696 -15240 9756 -15234
rect 11730 -15240 11790 -15234
rect 13766 -15240 13826 -15234
rect 15802 -15240 15862 -15234
rect 17842 -15240 17902 -15234
rect 19872 -15240 19932 -15234
rect 21912 -15240 21972 -15234
rect 2572 -15280 2632 -15274
rect 3070 -15280 3130 -15274
rect 3582 -15280 3642 -15274
rect 9862 -15280 9922 -15274
rect 11730 -15280 11790 -15274
rect 13768 -15280 13828 -15274
rect 15648 -15280 15708 -15274
rect 1880 -15284 15708 -15280
rect 1880 -15336 1890 -15284
rect 1942 -15336 2576 -15284
rect 2628 -15336 3074 -15284
rect 3126 -15336 3586 -15284
rect 3638 -15336 9866 -15284
rect 9918 -15336 11734 -15284
rect 11786 -15336 13772 -15284
rect 13824 -15336 15652 -15284
rect 15704 -15336 15708 -15284
rect 1880 -15340 15708 -15336
rect 2572 -15346 2632 -15340
rect 3070 -15346 3130 -15340
rect 3582 -15346 3642 -15340
rect 9862 -15346 9922 -15340
rect 11730 -15346 11790 -15340
rect 13768 -15346 13828 -15340
rect 15648 -15346 15708 -15340
rect 19872 -15278 19932 -15272
rect 23048 -15278 23108 -15272
rect 19872 -15282 23108 -15278
rect 19872 -15334 19876 -15282
rect 19928 -15334 23052 -15282
rect 23104 -15334 23108 -15282
rect 19872 -15338 23108 -15334
rect 19872 -15344 19932 -15338
rect 23048 -15344 23108 -15338
rect 2442 -16170 2502 -16164
rect 5620 -16170 5680 -16164
rect 8676 -16170 8736 -16164
rect 14782 -16170 14842 -16164
rect 19876 -16170 19936 -16164
rect 2442 -16174 19936 -16170
rect 2442 -16226 2446 -16174
rect 2498 -16226 5624 -16174
rect 5676 -16226 8680 -16174
rect 8732 -16226 14786 -16174
rect 14838 -16226 19880 -16174
rect 19932 -16226 19936 -16174
rect 2442 -16230 19936 -16226
rect 2442 -16236 2502 -16230
rect 5620 -16236 5680 -16230
rect 8676 -16236 8736 -16230
rect 14782 -16236 14842 -16230
rect 19876 -16236 19936 -16230
rect 2012 -16274 2072 -16268
rect 2566 -16274 2626 -16268
rect 4086 -16274 4146 -16268
rect 2012 -16278 4146 -16274
rect 2012 -16330 2016 -16278
rect 2068 -16330 2570 -16278
rect 2622 -16330 4090 -16278
rect 4142 -16330 4146 -16278
rect 2012 -16334 4146 -16330
rect 2012 -16340 2072 -16334
rect 2566 -16340 2626 -16334
rect 4086 -16340 4146 -16334
rect 4598 -16274 4658 -16268
rect 5622 -16274 5682 -16268
rect 6634 -16274 6694 -16268
rect 7654 -16274 7714 -16268
rect 10712 -16274 10772 -16268
rect 12750 -16274 12810 -16268
rect 15800 -16274 15860 -16268
rect 16818 -16274 16878 -16268
rect 17838 -16274 17898 -16268
rect 18854 -16274 18914 -16268
rect 20890 -16274 20950 -16268
rect 4598 -16278 20950 -16274
rect 4598 -16330 4602 -16278
rect 4654 -16330 5626 -16278
rect 5678 -16330 6638 -16278
rect 6690 -16330 7658 -16278
rect 7710 -16330 10716 -16278
rect 10768 -16330 12754 -16278
rect 12806 -16330 15804 -16278
rect 15856 -16330 16822 -16278
rect 16874 -16330 17842 -16278
rect 17894 -16330 18858 -16278
rect 18910 -16330 20894 -16278
rect 20946 -16330 20950 -16278
rect 4598 -16334 20950 -16330
rect 4598 -16340 4658 -16334
rect 5622 -16340 5682 -16334
rect 6634 -16340 6694 -16334
rect 7654 -16340 7714 -16334
rect 10712 -16340 10772 -16334
rect 12750 -16340 12810 -16334
rect 15800 -16340 15860 -16334
rect 16818 -16340 16878 -16334
rect 17838 -16340 17898 -16334
rect 18854 -16340 18914 -16334
rect 20890 -16340 20950 -16334
rect 2336 -16396 2396 -16390
rect 9696 -16396 9756 -16390
rect 11730 -16396 11790 -16390
rect 13760 -16396 13820 -16390
rect 23760 -16396 23820 -7438
rect 2336 -16400 23820 -16396
rect 2336 -16452 2340 -16400
rect 2392 -16452 9700 -16400
rect 9752 -16452 11734 -16400
rect 11786 -16452 13764 -16400
rect 13816 -16452 23820 -16400
rect 2336 -16456 23820 -16452
rect 2336 -16462 2396 -16456
rect 9696 -16462 9756 -16456
rect 11730 -16462 11790 -16456
rect 13760 -16462 13820 -16456
rect 2224 -16510 2284 -16504
rect 3072 -16510 3132 -16504
rect 2224 -16514 3132 -16510
rect 2224 -16566 2228 -16514
rect 2280 -16566 3076 -16514
rect 3128 -16566 3132 -16514
rect 2224 -16570 3132 -16566
rect 2224 -16576 2284 -16570
rect 3072 -16576 3132 -16570
rect 4604 -16508 4664 -16502
rect 6640 -16508 6700 -16502
rect 23034 -16508 23094 -16502
rect 4604 -16512 23094 -16508
rect 4604 -16564 4608 -16512
rect 4660 -16564 6644 -16512
rect 6696 -16564 23038 -16512
rect 23090 -16564 23094 -16512
rect 4604 -16568 23094 -16564
rect 4604 -16574 4664 -16568
rect 6640 -16574 6700 -16568
rect 23034 -16574 23094 -16568
rect 23162 -16526 23222 -16520
rect 23762 -16526 23822 -16520
rect 23162 -16530 23822 -16526
rect 23162 -16582 23166 -16530
rect 23218 -16582 23766 -16530
rect 23818 -16582 23822 -16530
rect 23162 -16586 23822 -16582
rect 23162 -16592 23222 -16586
rect 23762 -16592 23822 -16586
rect 22928 -17396 22988 -17390
rect 23888 -17396 23948 -7120
rect 22928 -17400 23948 -17396
rect 5620 -17414 5680 -17408
rect 7656 -17414 7716 -17408
rect 15800 -17414 15860 -17408
rect 17836 -17414 17896 -17408
rect 21910 -17414 21970 -17408
rect 5620 -17418 21970 -17414
rect 2448 -17438 2508 -17432
rect 3586 -17438 3646 -17432
rect 2448 -17442 4468 -17438
rect 2448 -17494 2452 -17442
rect 2504 -17494 3590 -17442
rect 3642 -17494 4468 -17442
rect 5620 -17470 5624 -17418
rect 5676 -17470 7660 -17418
rect 7712 -17470 15804 -17418
rect 15856 -17470 17840 -17418
rect 17892 -17470 21914 -17418
rect 21966 -17470 21970 -17418
rect 22928 -17452 22932 -17400
rect 22984 -17452 23948 -17400
rect 22928 -17456 23948 -17452
rect 22928 -17462 22988 -17456
rect 5620 -17474 21970 -17470
rect 5620 -17480 5680 -17474
rect 7656 -17480 7716 -17474
rect 15800 -17480 15860 -17474
rect 17836 -17480 17896 -17474
rect 21910 -17480 21970 -17474
rect 2448 -17498 4468 -17494
rect 2448 -17504 2508 -17498
rect 3586 -17504 3646 -17498
rect 2336 -17638 2396 -17632
rect 3584 -17638 3644 -17632
rect 2336 -17642 3644 -17638
rect 2336 -17694 2340 -17642
rect 2392 -17694 3588 -17642
rect 3640 -17694 3644 -17642
rect 4408 -17634 4468 -17498
rect 4602 -17518 4662 -17512
rect 6642 -17518 6702 -17512
rect 8674 -17518 8734 -17512
rect 10708 -17518 10768 -17512
rect 12748 -17518 12808 -17512
rect 14782 -17518 14842 -17512
rect 4602 -17522 14842 -17518
rect 4602 -17574 4606 -17522
rect 4658 -17574 6646 -17522
rect 6698 -17574 8678 -17522
rect 8730 -17574 10712 -17522
rect 10764 -17574 12752 -17522
rect 12804 -17574 14786 -17522
rect 14838 -17574 14842 -17522
rect 4602 -17578 14842 -17574
rect 4602 -17584 4662 -17578
rect 6642 -17584 6702 -17578
rect 8674 -17584 8734 -17578
rect 10708 -17584 10768 -17578
rect 12748 -17584 12808 -17578
rect 14782 -17584 14842 -17578
rect 14978 -17522 15038 -17516
rect 19870 -17522 19930 -17516
rect 14978 -17526 19930 -17522
rect 23528 -17526 23588 -17520
rect 14978 -17578 14982 -17526
rect 15034 -17578 19874 -17526
rect 19926 -17578 19930 -17526
rect 14978 -17582 19930 -17578
rect 14978 -17588 15038 -17582
rect 19870 -17588 19930 -17582
rect 20368 -17530 23588 -17526
rect 20368 -17582 20378 -17530
rect 20430 -17582 23532 -17530
rect 23584 -17582 23588 -17530
rect 20368 -17586 23588 -17582
rect 23528 -17592 23588 -17586
rect 5116 -17632 5176 -17626
rect 8674 -17630 8734 -17624
rect 10710 -17630 10770 -17624
rect 12746 -17630 12806 -17624
rect 14782 -17630 14842 -17624
rect 16816 -17630 16876 -17624
rect 18854 -17630 18914 -17624
rect 20894 -17630 20954 -17624
rect 23278 -17630 23338 -17624
rect 5116 -17634 8218 -17632
rect 4408 -17636 8218 -17634
rect 4408 -17688 5120 -17636
rect 5172 -17688 6124 -17636
rect 6176 -17688 7136 -17636
rect 7188 -17688 8156 -17636
rect 8208 -17688 8218 -17636
rect 4408 -17692 8218 -17688
rect 8674 -17634 23338 -17630
rect 8674 -17686 8678 -17634
rect 8730 -17686 10714 -17634
rect 10766 -17686 12750 -17634
rect 12802 -17686 14786 -17634
rect 14838 -17686 16820 -17634
rect 16872 -17686 18858 -17634
rect 18910 -17686 20898 -17634
rect 20950 -17686 23282 -17634
rect 23334 -17686 23338 -17634
rect 8674 -17690 23338 -17686
rect 4408 -17694 5458 -17692
rect 2336 -17698 3644 -17694
rect 5116 -17698 5176 -17694
rect 8674 -17696 8734 -17690
rect 10710 -17696 10770 -17690
rect 12746 -17696 12806 -17690
rect 14782 -17696 14842 -17690
rect 16816 -17696 16876 -17690
rect 18854 -17696 18914 -17690
rect 20894 -17696 20954 -17690
rect 23278 -17696 23338 -17690
rect 2336 -17704 2396 -17698
rect 3584 -17704 3644 -17698
rect 1660 -17740 1720 -17734
rect 2230 -17740 2290 -17734
rect 9692 -17740 9752 -17734
rect 11726 -17740 11786 -17734
rect 13766 -17740 13826 -17734
rect 14978 -17740 15038 -17734
rect 1660 -17744 15038 -17740
rect 1660 -17796 1664 -17744
rect 1716 -17796 2234 -17744
rect 2286 -17796 9696 -17744
rect 9748 -17796 11730 -17744
rect 11782 -17796 13770 -17744
rect 13822 -17796 14982 -17744
rect 15034 -17796 15038 -17744
rect 1660 -17800 15038 -17796
rect 1660 -17806 1720 -17800
rect 2230 -17806 2290 -17800
rect 9692 -17806 9752 -17800
rect 11726 -17806 11786 -17800
rect 13766 -17806 13826 -17800
rect 14978 -17806 15038 -17800
rect 15272 -17738 15332 -17732
rect 15272 -17742 16366 -17738
rect 15272 -17794 15276 -17742
rect 15328 -17794 16304 -17742
rect 16356 -17794 16366 -17742
rect 15272 -17798 16366 -17794
rect 16818 -17744 16878 -17738
rect 18854 -17744 18914 -17738
rect 20892 -17744 20952 -17738
rect 23034 -17744 23094 -17738
rect 16818 -17748 23094 -17744
rect 15272 -17804 15332 -17798
rect 16818 -17800 16822 -17748
rect 16874 -17800 18858 -17748
rect 18910 -17800 20896 -17748
rect 20948 -17800 23038 -17748
rect 23090 -17800 23094 -17748
rect 16818 -17804 23094 -17800
rect 16818 -17810 16878 -17804
rect 18854 -17810 18914 -17804
rect 20892 -17810 20952 -17804
rect 23034 -17810 23094 -17804
rect 19366 -18658 19426 -18652
rect 14266 -18662 19426 -18658
rect 3584 -18670 3644 -18664
rect 5622 -18670 5682 -18664
rect 7658 -18670 7718 -18664
rect 9690 -18670 9750 -18664
rect 3584 -18674 9750 -18670
rect 3584 -18726 3588 -18674
rect 3640 -18726 5626 -18674
rect 5678 -18726 7662 -18674
rect 7714 -18726 9694 -18674
rect 9746 -18726 9750 -18674
rect 14266 -18714 14276 -18662
rect 14328 -18714 19370 -18662
rect 19422 -18714 19426 -18662
rect 14266 -18718 19426 -18714
rect 19366 -18724 19426 -18718
rect 19504 -18654 19564 -18648
rect 20386 -18654 20446 -18648
rect 21392 -18654 21452 -18648
rect 19504 -18658 21452 -18654
rect 19504 -18710 19508 -18658
rect 19560 -18710 20390 -18658
rect 20442 -18710 21396 -18658
rect 21448 -18710 21452 -18658
rect 19504 -18714 21452 -18710
rect 19504 -18720 19564 -18714
rect 20386 -18720 20446 -18714
rect 21392 -18720 21452 -18714
rect 21910 -18658 21970 -18652
rect 23162 -18658 23222 -18652
rect 21910 -18662 23222 -18658
rect 21910 -18714 21914 -18662
rect 21966 -18714 23166 -18662
rect 23218 -18714 23222 -18662
rect 21910 -18718 23222 -18714
rect 21910 -18724 21970 -18718
rect 23162 -18724 23222 -18718
rect 3584 -18730 9750 -18726
rect 3584 -18736 3644 -18730
rect 5622 -18736 5682 -18730
rect 7658 -18736 7718 -18730
rect 9690 -18736 9750 -18730
rect 4090 -18772 4150 -18766
rect 9182 -18772 9242 -18766
rect 4090 -18776 9242 -18772
rect 1150 -18826 1210 -18816
rect 1150 -18878 1154 -18826
rect 1206 -18878 1210 -18826
rect 4090 -18828 4094 -18776
rect 4146 -18828 9186 -18776
rect 9238 -18828 9242 -18776
rect 4090 -18832 9242 -18828
rect 4090 -18838 4150 -18832
rect 9182 -18838 9242 -18832
rect 13766 -18786 13826 -18780
rect 21910 -18786 21970 -18780
rect 13766 -18790 21970 -18786
rect 13766 -18842 13770 -18790
rect 13822 -18842 21914 -18790
rect 21966 -18842 21970 -18790
rect 13766 -18846 21970 -18842
rect 13766 -18852 13826 -18846
rect 21910 -18852 21970 -18846
rect -3398 -19748 -3338 -19742
rect 1150 -19748 1210 -18878
rect 2336 -18874 2396 -18868
rect 5620 -18874 5680 -18868
rect 2336 -18878 5680 -18874
rect 2336 -18930 2340 -18878
rect 2392 -18930 5624 -18878
rect 5676 -18930 5680 -18878
rect 2336 -18934 5680 -18930
rect 2336 -18940 2396 -18934
rect 5620 -18940 5680 -18934
rect 6128 -18880 6188 -18874
rect 7150 -18880 7210 -18874
rect 8164 -18880 8224 -18874
rect 9182 -18880 9242 -18874
rect 10202 -18880 10262 -18874
rect 17314 -18880 17374 -18874
rect 18344 -18880 18404 -18874
rect 19504 -18880 19564 -18874
rect 6128 -18884 19564 -18880
rect 6128 -18936 6132 -18884
rect 6184 -18936 7154 -18884
rect 7206 -18936 8168 -18884
rect 8220 -18936 9186 -18884
rect 9238 -18936 10206 -18884
rect 10258 -18936 17318 -18884
rect 17370 -18936 18348 -18884
rect 18400 -18936 19508 -18884
rect 19560 -18936 19564 -18884
rect 6128 -18940 19564 -18936
rect 6128 -18946 6188 -18940
rect 7150 -18946 7210 -18940
rect 8164 -18946 8224 -18940
rect 9182 -18946 9242 -18940
rect 10202 -18946 10262 -18940
rect 17314 -18946 17374 -18940
rect 18344 -18946 18404 -18940
rect 19504 -18946 19564 -18940
rect 19872 -18880 19932 -18874
rect 23400 -18880 23460 -18874
rect 19872 -18884 23460 -18880
rect 19872 -18936 19876 -18884
rect 19928 -18936 23404 -18884
rect 23456 -18936 23460 -18884
rect 19872 -18940 23460 -18936
rect 19872 -18946 19932 -18940
rect 23400 -18946 23460 -18940
rect 4604 -18974 4664 -18968
rect 6638 -18974 6698 -18968
rect 8674 -18974 8734 -18968
rect 4604 -18978 8734 -18974
rect 4604 -19030 4608 -18978
rect 4660 -19030 6642 -18978
rect 6694 -19030 8678 -18978
rect 8730 -19030 8734 -18978
rect 4604 -19034 8734 -19030
rect 4604 -19040 4664 -19034
rect 6638 -19040 6698 -19034
rect 8674 -19040 8734 -19034
rect 15802 -18984 15862 -18978
rect 19872 -18984 19932 -18978
rect 15802 -18988 19932 -18984
rect 15802 -19040 15806 -18988
rect 15858 -19040 19876 -18988
rect 19928 -19040 19932 -18988
rect 15802 -19044 19932 -19040
rect 15802 -19050 15862 -19044
rect 19872 -19050 19932 -19044
rect 20888 -18982 20948 -18976
rect 23278 -18982 23338 -18976
rect 20888 -18986 23338 -18982
rect 20888 -19038 20892 -18986
rect 20944 -19038 23282 -18986
rect 23334 -19038 23338 -18986
rect 20888 -19042 23338 -19038
rect 20888 -19048 20948 -19042
rect 23278 -19048 23338 -19042
rect -3398 -19752 1210 -19748
rect -3398 -19804 -3394 -19752
rect -3342 -19804 1210 -19752
rect -3398 -19808 1210 -19804
rect -3398 -19814 -3338 -19808
rect -5428 -19894 -5368 -19888
rect -1368 -19894 -1308 -19888
rect 816 -19894 876 -19888
rect 1282 -19894 1342 -19888
rect 10710 -19892 10770 -19886
rect 12746 -19892 12806 -19886
rect 14782 -19892 14842 -19886
rect 16820 -19892 16880 -19886
rect -9514 -19898 1342 -19894
rect -9514 -19950 -9504 -19898
rect -9452 -19950 -5424 -19898
rect -5372 -19950 -1364 -19898
rect -1312 -19950 820 -19898
rect 872 -19950 1286 -19898
rect 1338 -19950 1342 -19898
rect -9514 -19954 1342 -19950
rect -5428 -19960 -5368 -19954
rect -1368 -19960 -1308 -19954
rect 816 -19960 876 -19954
rect 1282 -19960 1342 -19954
rect 4086 -19898 4146 -19892
rect 4996 -19898 5056 -19892
rect 5998 -19898 6058 -19892
rect 7150 -19898 7210 -19892
rect 8160 -19898 8220 -19892
rect 9166 -19898 9226 -19892
rect 10210 -19898 10270 -19892
rect 4086 -19902 10270 -19898
rect 4086 -19954 4090 -19902
rect 4142 -19954 5000 -19902
rect 5052 -19954 6002 -19902
rect 6054 -19954 7154 -19902
rect 7206 -19954 8164 -19902
rect 8216 -19954 9170 -19902
rect 9222 -19954 10214 -19902
rect 10266 -19954 10270 -19902
rect 4086 -19958 10270 -19954
rect 10710 -19896 16880 -19892
rect 10710 -19948 10714 -19896
rect 10766 -19948 12750 -19896
rect 12802 -19948 14786 -19896
rect 14838 -19948 16824 -19896
rect 16876 -19948 16880 -19896
rect 10710 -19952 16880 -19948
rect 10710 -19958 10770 -19952
rect 12746 -19958 12806 -19952
rect 14782 -19958 14842 -19952
rect 16820 -19958 16880 -19952
rect 18856 -19892 18916 -19886
rect 20894 -19892 20954 -19886
rect 18856 -19896 20954 -19892
rect 18856 -19948 18860 -19896
rect 18912 -19948 20898 -19896
rect 20950 -19948 20954 -19896
rect 18856 -19952 20954 -19948
rect 18856 -19958 18916 -19952
rect 20894 -19958 20954 -19952
rect 4086 -19964 4146 -19958
rect 4996 -19964 5056 -19958
rect 5998 -19964 6058 -19958
rect 7150 -19964 7210 -19958
rect 8160 -19964 8220 -19958
rect 9166 -19964 9226 -19958
rect 10210 -19964 10270 -19958
rect 6638 -20000 6698 -19994
rect 16812 -20000 16872 -19994
rect 18852 -20000 18912 -19994
rect 20890 -20000 20950 -19994
rect 6638 -20004 20950 -20000
rect -10662 -20022 -10602 -20016
rect -7984 -20022 -7924 -20016
rect -6952 -20022 -6892 -20016
rect -3892 -20022 -3832 -20016
rect -2896 -20022 -2836 -20016
rect 1402 -20022 1462 -20016
rect -10662 -20026 1462 -20022
rect -10662 -20078 -10658 -20026
rect -10606 -20078 -7980 -20026
rect -7928 -20078 -6948 -20026
rect -6896 -20078 -3888 -20026
rect -3836 -20078 -2892 -20026
rect -2840 -20078 1406 -20026
rect 1458 -20078 1462 -20026
rect 6638 -20056 6642 -20004
rect 6694 -20056 16816 -20004
rect 16868 -20056 18856 -20004
rect 18908 -20056 20894 -20004
rect 20946 -20056 20950 -20004
rect 6638 -20060 20950 -20056
rect 6638 -20066 6698 -20060
rect 16812 -20066 16872 -20060
rect 18852 -20066 18912 -20060
rect 20890 -20066 20950 -20060
rect -10662 -20082 1462 -20078
rect -10662 -20088 -10602 -20082
rect -7984 -20088 -7924 -20082
rect -6952 -20088 -6892 -20082
rect -3892 -20088 -3832 -20082
rect -2896 -20088 -2836 -20082
rect 1402 -20088 1462 -20082
rect 4086 -20114 4146 -20108
rect 6138 -20114 6198 -20108
rect 9164 -20114 9224 -20108
rect 10204 -20114 10264 -20108
rect 11218 -20114 11278 -20108
rect 12226 -20114 12286 -20108
rect 13270 -20114 13330 -20108
rect 14260 -20114 14320 -20108
rect 15278 -20114 15338 -20108
rect 16312 -20114 16372 -20108
rect 19344 -20114 19404 -20108
rect 20382 -20114 20442 -20108
rect 21408 -20114 21468 -20108
rect 4086 -20118 23592 -20114
rect 4086 -20170 4090 -20118
rect 4142 -20170 5128 -20118
rect 5180 -20170 6142 -20118
rect 6194 -20170 9168 -20118
rect 9220 -20170 10208 -20118
rect 10260 -20170 11222 -20118
rect 11274 -20170 12230 -20118
rect 12282 -20170 13274 -20118
rect 13326 -20170 14264 -20118
rect 14316 -20170 15282 -20118
rect 15334 -20170 16316 -20118
rect 16368 -20170 19348 -20118
rect 19400 -20170 20386 -20118
rect 20438 -20170 21412 -20118
rect 21464 -20170 23530 -20118
rect 23582 -20170 23592 -20118
rect 4086 -20174 23592 -20170
rect 4086 -20180 4146 -20174
rect 6138 -20180 6198 -20174
rect 9164 -20180 9224 -20174
rect 10204 -20180 10264 -20174
rect 11218 -20180 11278 -20174
rect 12226 -20180 12286 -20174
rect 13270 -20180 13330 -20174
rect 14260 -20180 14320 -20174
rect 15278 -20180 15338 -20174
rect 16312 -20180 16372 -20174
rect 19344 -20180 19404 -20174
rect 20382 -20180 20442 -20174
rect 21408 -20180 21468 -20174
rect 9688 -20218 9748 -20212
rect 11730 -20218 11790 -20212
rect 13768 -20218 13828 -20212
rect 15802 -20218 15862 -20212
rect 17836 -20216 17896 -20210
rect 19870 -20216 19930 -20210
rect 21912 -20216 21972 -20210
rect 23162 -20216 23222 -20210
rect 2444 -20222 15862 -20218
rect 2444 -20274 2454 -20222
rect 2506 -20274 9692 -20222
rect 9744 -20274 11734 -20222
rect 11786 -20274 13772 -20222
rect 13824 -20274 15806 -20222
rect 15858 -20274 15862 -20222
rect 2444 -20278 15862 -20274
rect 9688 -20284 9748 -20278
rect 11730 -20284 11790 -20278
rect 13768 -20284 13828 -20278
rect 15802 -20284 15862 -20278
rect 16314 -20222 16374 -20216
rect 17336 -20222 17396 -20216
rect 16314 -20226 17396 -20222
rect 16314 -20278 16318 -20226
rect 16370 -20278 17340 -20226
rect 17392 -20278 17396 -20226
rect 16314 -20282 17396 -20278
rect 17836 -20220 23222 -20216
rect 17836 -20272 17840 -20220
rect 17892 -20272 19874 -20220
rect 19926 -20272 21916 -20220
rect 21968 -20272 23166 -20220
rect 23218 -20272 23222 -20220
rect 17836 -20276 23222 -20272
rect 17836 -20282 17896 -20276
rect 19870 -20282 19930 -20276
rect 21912 -20282 21972 -20276
rect 23162 -20282 23222 -20276
rect 16314 -20288 16374 -20282
rect 17336 -20288 17396 -20282
rect -9004 -20984 -8944 -20978
rect -7980 -20984 -7920 -20978
rect -6948 -20984 -6888 -20978
rect -5948 -20984 -5888 -20978
rect -4928 -20984 -4868 -20978
rect -3908 -20984 -3848 -20978
rect -1884 -20984 -1824 -20978
rect 936 -20984 996 -20978
rect 1542 -20984 1602 -20978
rect -9004 -20988 1602 -20984
rect -9004 -21040 -9000 -20988
rect -8948 -21040 -7976 -20988
rect -7924 -21040 -6944 -20988
rect -6892 -21040 -5944 -20988
rect -5892 -21040 -4924 -20988
rect -4872 -21040 -3904 -20988
rect -3852 -21040 -2894 -20988
rect -2842 -21040 -1880 -20988
rect -1828 -21040 -862 -20988
rect -810 -21040 940 -20988
rect 992 -21040 1546 -20988
rect 1598 -21040 1602 -20988
rect -9004 -21044 1602 -21040
rect -9004 -21050 -8944 -21044
rect -7980 -21050 -7920 -21044
rect -6948 -21050 -6888 -21044
rect -5948 -21050 -5888 -21044
rect -4928 -21050 -4868 -21044
rect -3908 -21050 -3848 -21044
rect -1884 -21050 -1824 -21044
rect 936 -21050 996 -21044
rect 1542 -21050 1602 -21044
rect -9504 -21088 -9444 -21082
rect -7468 -21088 -7408 -21082
rect -5432 -21088 -5372 -21082
rect -3398 -21088 -3338 -21082
rect -1362 -21088 -1302 -21082
rect -9504 -21092 -1302 -21088
rect -9504 -21144 -9500 -21092
rect -9448 -21144 -7464 -21092
rect -7412 -21144 -5428 -21092
rect -5376 -21144 -3394 -21092
rect -3342 -21144 -1358 -21092
rect -1306 -21144 -1302 -21092
rect 8678 -21120 8738 -21114
rect 12746 -21120 12806 -21114
rect 14780 -21120 14840 -21114
rect -9504 -21148 -1302 -21144
rect -9504 -21154 -9444 -21148
rect -7468 -21154 -7408 -21148
rect -5432 -21154 -5372 -21148
rect -3398 -21154 -3338 -21148
rect -1362 -21154 -1302 -21148
rect 4084 -21126 4144 -21120
rect 5092 -21126 5152 -21120
rect 6106 -21126 6166 -21120
rect 7144 -21126 7204 -21120
rect 8162 -21126 8222 -21120
rect 4084 -21130 8222 -21126
rect 4084 -21182 4088 -21130
rect 4140 -21182 5096 -21130
rect 5148 -21182 6110 -21130
rect 6162 -21182 7148 -21130
rect 7200 -21182 8166 -21130
rect 8218 -21182 8222 -21130
rect 4084 -21186 8222 -21182
rect 8678 -21124 14840 -21120
rect 8678 -21176 8682 -21124
rect 8734 -21176 10718 -21124
rect 10770 -21176 12750 -21124
rect 12802 -21176 14784 -21124
rect 14836 -21176 14840 -21124
rect 8678 -21180 14840 -21176
rect 8678 -21186 8738 -21180
rect 12746 -21186 12806 -21180
rect 14780 -21186 14840 -21180
rect 15802 -21118 15862 -21112
rect 16156 -21118 16216 -21112
rect 15802 -21122 16216 -21118
rect 15802 -21174 15806 -21122
rect 15858 -21174 16160 -21122
rect 16212 -21174 16216 -21122
rect 15802 -21178 16216 -21174
rect 15802 -21184 15862 -21178
rect 16156 -21184 16216 -21178
rect 19874 -21118 19934 -21112
rect 23158 -21118 23218 -21112
rect 19874 -21122 23218 -21118
rect 19874 -21174 19878 -21122
rect 19930 -21174 23162 -21122
rect 23214 -21174 23218 -21122
rect 19874 -21178 23218 -21174
rect 19874 -21184 19934 -21178
rect 23158 -21184 23218 -21178
rect -4418 -21192 -4358 -21186
rect 2120 -21192 2180 -21186
rect 4084 -21192 4144 -21186
rect 5092 -21192 5152 -21186
rect 6106 -21192 6166 -21186
rect 7144 -21192 7204 -21186
rect 8162 -21192 8222 -21186
rect -8492 -21196 2180 -21192
rect -8492 -21248 -8482 -21196
rect -8430 -21248 -6446 -21196
rect -6394 -21248 -4414 -21196
rect -4362 -21248 -2380 -21196
rect -2328 -21248 -336 -21196
rect -284 -21248 2124 -21196
rect 2176 -21248 2180 -21196
rect -8492 -21252 2180 -21248
rect -4418 -21258 -4358 -21252
rect 2120 -21258 2180 -21252
rect 2230 -21230 2290 -21224
rect 3586 -21230 3646 -21224
rect 11730 -21230 11790 -21224
rect 13766 -21230 13826 -21224
rect 15798 -21230 15858 -21224
rect 2230 -21234 15858 -21230
rect 2230 -21286 2234 -21234
rect 2286 -21286 3590 -21234
rect 3642 -21286 11734 -21234
rect 11786 -21286 13770 -21234
rect 13822 -21286 15802 -21234
rect 15854 -21286 15858 -21234
rect 2230 -21290 15858 -21286
rect 2230 -21296 2290 -21290
rect 3586 -21296 3646 -21290
rect 11730 -21296 11790 -21290
rect 13766 -21296 13826 -21290
rect 15798 -21296 15858 -21290
rect 15308 -21328 15368 -21322
rect 16346 -21328 16406 -21322
rect 17322 -21328 17382 -21322
rect 18338 -21328 18398 -21322
rect 20364 -21328 20424 -21322
rect 21394 -21328 21454 -21322
rect 15308 -21332 21454 -21328
rect 1888 -21342 1948 -21336
rect 4602 -21342 4662 -21336
rect 6640 -21342 6700 -21336
rect 10712 -21342 10772 -21336
rect 1888 -21346 10772 -21342
rect 1888 -21398 1892 -21346
rect 1944 -21398 4606 -21346
rect 4658 -21398 6644 -21346
rect 6696 -21398 10716 -21346
rect 10768 -21398 10772 -21346
rect 15308 -21384 15312 -21332
rect 15364 -21384 16350 -21332
rect 16402 -21384 17326 -21332
rect 17378 -21384 18342 -21332
rect 18394 -21384 20368 -21332
rect 20420 -21384 21398 -21332
rect 21450 -21384 21454 -21332
rect 15308 -21388 21454 -21384
rect 15308 -21394 15368 -21388
rect 16346 -21394 16406 -21388
rect 17322 -21394 17382 -21388
rect 18338 -21394 18398 -21388
rect 20364 -21394 20424 -21388
rect 21394 -21394 21454 -21388
rect 1888 -21402 10772 -21398
rect 1888 -21408 1948 -21402
rect 4602 -21408 4662 -21402
rect 6640 -21408 6700 -21402
rect 10712 -21408 10772 -21402
rect 3582 -21440 3642 -21434
rect 5620 -21440 5680 -21434
rect 7660 -21440 7720 -21434
rect 9696 -21440 9756 -21434
rect 15800 -21440 15860 -21434
rect 16150 -21440 16222 -21436
rect 17836 -21440 17896 -21434
rect 19872 -21440 19932 -21434
rect 21908 -21440 21968 -21434
rect 3582 -21444 16160 -21440
rect 3582 -21496 3586 -21444
rect 3638 -21496 5624 -21444
rect 5676 -21496 7664 -21444
rect 7716 -21496 9700 -21444
rect 9752 -21492 16160 -21444
rect 16212 -21444 21968 -21440
rect 16212 -21492 17840 -21444
rect 9752 -21496 17840 -21492
rect 17892 -21496 19876 -21444
rect 19928 -21496 21912 -21444
rect 21964 -21496 21968 -21444
rect 3582 -21500 21968 -21496
rect 3582 -21506 3642 -21500
rect 5620 -21506 5680 -21500
rect 7660 -21506 7720 -21500
rect 9696 -21506 9756 -21500
rect 15800 -21506 15860 -21500
rect 17836 -21506 17896 -21500
rect 19872 -21506 19932 -21500
rect 21908 -21506 21968 -21500
rect -7474 -22134 -7414 -22128
rect -3398 -22134 -3338 -22128
rect 816 -22134 876 -22128
rect -7474 -22138 876 -22134
rect -7474 -22190 -7470 -22138
rect -7418 -22190 -3394 -22138
rect -3342 -22190 820 -22138
rect 872 -22190 876 -22138
rect -7474 -22194 876 -22190
rect -7474 -22200 -7414 -22194
rect -3398 -22200 -3338 -22194
rect 816 -22200 876 -22194
rect -10662 -22254 -10602 -22248
rect -9012 -22254 -8952 -22248
rect -5942 -22254 -5882 -22248
rect -4934 -22254 -4874 -22248
rect -1872 -22254 -1812 -22248
rect -846 -22254 -786 -22248
rect -10662 -22258 -786 -22254
rect -10662 -22310 -10658 -22258
rect -10606 -22310 -9008 -22258
rect -8956 -22310 -5938 -22258
rect -5886 -22310 -4930 -22258
rect -4878 -22310 -1868 -22258
rect -1816 -22310 -842 -22258
rect -790 -22310 -786 -22258
rect -10662 -22314 -786 -22310
rect -10662 -22320 -10602 -22314
rect -9012 -22320 -8952 -22314
rect -5942 -22320 -5882 -22314
rect -4934 -22320 -4874 -22314
rect -1872 -22320 -1812 -22314
rect -846 -22320 -786 -22314
rect 10708 -22344 10768 -22338
rect 12750 -22344 12810 -22338
rect 14782 -22344 14842 -22338
rect 16822 -22344 16882 -22338
rect 23278 -22344 23338 -22338
rect 10532 -22348 23338 -22344
rect 4602 -22364 4662 -22358
rect 6638 -22364 6698 -22358
rect 8676 -22364 8736 -22358
rect 4602 -22368 8736 -22364
rect 4602 -22420 4606 -22368
rect 4658 -22420 6642 -22368
rect 6694 -22420 8680 -22368
rect 8732 -22420 8736 -22368
rect 10532 -22400 10542 -22348
rect 10594 -22400 10712 -22348
rect 10764 -22400 12754 -22348
rect 12806 -22400 14786 -22348
rect 14838 -22400 16826 -22348
rect 16878 -22400 23282 -22348
rect 23334 -22400 23338 -22348
rect 10532 -22404 23338 -22400
rect 10708 -22410 10768 -22404
rect 12750 -22410 12810 -22404
rect 14782 -22410 14842 -22404
rect 16822 -22410 16882 -22404
rect 23278 -22410 23338 -22404
rect 4602 -22424 8736 -22420
rect 4602 -22430 4662 -22424
rect 6638 -22430 6698 -22424
rect 8676 -22430 8736 -22424
rect 15800 -22442 15860 -22436
rect 21906 -22442 21966 -22436
rect 23158 -22442 23218 -22436
rect 15800 -22446 23218 -22442
rect 2448 -22462 2508 -22456
rect 5620 -22462 5680 -22456
rect 2448 -22466 5680 -22462
rect 2448 -22518 2452 -22466
rect 2504 -22518 5624 -22466
rect 5676 -22518 5680 -22466
rect 2448 -22522 5680 -22518
rect 2448 -22528 2508 -22522
rect 5620 -22528 5680 -22522
rect 7144 -22462 7204 -22456
rect 10192 -22462 10252 -22456
rect 7144 -22466 10252 -22462
rect 7144 -22518 7148 -22466
rect 7200 -22518 8170 -22466
rect 8222 -22518 9192 -22466
rect 9244 -22518 10196 -22466
rect 10248 -22518 10252 -22466
rect 15800 -22498 15804 -22446
rect 15856 -22498 21910 -22446
rect 21962 -22498 23162 -22446
rect 23214 -22498 23218 -22446
rect 15800 -22502 23218 -22498
rect 15800 -22508 15860 -22502
rect 21906 -22508 21966 -22502
rect 23158 -22508 23218 -22502
rect 7144 -22522 10252 -22518
rect 7144 -22528 7204 -22522
rect 10192 -22528 10252 -22522
rect 10714 -22552 10774 -22546
rect 12742 -22552 12802 -22546
rect 14786 -22552 14846 -22546
rect 16814 -22552 16874 -22546
rect 18852 -22552 18912 -22546
rect 20892 -22552 20952 -22546
rect 4606 -22558 4666 -22552
rect 6642 -22558 6702 -22552
rect 8670 -22558 8730 -22552
rect 10538 -22558 10598 -22552
rect 4606 -22562 10598 -22558
rect 4606 -22614 4610 -22562
rect 4662 -22614 6646 -22562
rect 6698 -22614 8674 -22562
rect 8726 -22614 10542 -22562
rect 10594 -22614 10598 -22562
rect 4606 -22618 10598 -22614
rect 10714 -22556 20952 -22552
rect 10714 -22608 10718 -22556
rect 10770 -22608 12746 -22556
rect 12798 -22608 14790 -22556
rect 14842 -22608 16818 -22556
rect 16870 -22608 18856 -22556
rect 18908 -22608 20896 -22556
rect 20948 -22608 20952 -22556
rect 10714 -22612 20952 -22608
rect 10714 -22618 10774 -22612
rect 12742 -22618 12802 -22612
rect 14786 -22618 14846 -22612
rect 16814 -22618 16874 -22612
rect 18852 -22618 18912 -22612
rect 20892 -22618 20952 -22612
rect 21410 -22548 21470 -22542
rect 22922 -22548 22982 -22542
rect 23528 -22548 23588 -22542
rect 21410 -22552 23588 -22548
rect 21410 -22604 21414 -22552
rect 21466 -22604 22926 -22552
rect 22978 -22604 23532 -22552
rect 23584 -22604 23588 -22552
rect 21410 -22608 23588 -22604
rect 21410 -22614 21470 -22608
rect 22922 -22614 22982 -22608
rect 23528 -22614 23588 -22608
rect 4606 -22624 4666 -22618
rect 6642 -22624 6702 -22618
rect 8670 -22624 8730 -22618
rect 10538 -22624 10598 -22618
rect 3588 -22678 3648 -22672
rect 7656 -22678 7716 -22672
rect 9690 -22678 9750 -22672
rect 17840 -22678 17900 -22672
rect 19870 -22678 19930 -22672
rect 21910 -22676 21970 -22670
rect 23400 -22676 23460 -22670
rect 3588 -22682 19930 -22678
rect 3588 -22734 3592 -22682
rect 3644 -22734 7660 -22682
rect 7712 -22734 9694 -22682
rect 9746 -22734 17844 -22682
rect 17896 -22734 19874 -22682
rect 19926 -22734 19930 -22682
rect 3588 -22738 19930 -22734
rect 20390 -22680 23460 -22676
rect 20390 -22732 20400 -22680
rect 20452 -22732 21914 -22680
rect 21966 -22732 23404 -22680
rect 23456 -22732 23460 -22680
rect 20390 -22736 23460 -22732
rect 3588 -22744 3648 -22738
rect 7656 -22744 7716 -22738
rect 9690 -22744 9750 -22738
rect 17840 -22744 17900 -22738
rect 19870 -22744 19930 -22738
rect 21910 -22742 21970 -22736
rect 23400 -22742 23460 -22736
rect -340 -23198 -280 -23192
rect -8492 -23202 -280 -23198
rect -8492 -23254 -8482 -23202
rect -8430 -23254 -6446 -23202
rect -6394 -23254 -4414 -23202
rect -4362 -23254 -2380 -23202
rect -2328 -23254 -336 -23202
rect -284 -23254 -280 -23202
rect -8492 -23258 -280 -23254
rect -340 -23264 -280 -23258
rect -9500 -23306 -9440 -23300
rect -7464 -23306 -7404 -23300
rect -5428 -23306 -5368 -23300
rect -3394 -23306 -3334 -23300
rect -1358 -23306 -1298 -23300
rect -9500 -23310 -1298 -23306
rect -9500 -23362 -9496 -23310
rect -9444 -23362 -7460 -23310
rect -7408 -23362 -5424 -23310
rect -5372 -23362 -3390 -23310
rect -3338 -23362 -1354 -23310
rect -1302 -23362 -1298 -23310
rect -9500 -23366 -1298 -23362
rect -9500 -23372 -9440 -23366
rect -7464 -23372 -7404 -23366
rect -5428 -23372 -5368 -23366
rect -3394 -23372 -3334 -23366
rect -1358 -23372 -1298 -23366
rect -9006 -23418 -8946 -23412
rect -7982 -23418 -7922 -23412
rect -6950 -23418 -6890 -23412
rect -5950 -23418 -5890 -23412
rect -4930 -23418 -4870 -23412
rect -3910 -23418 -3850 -23412
rect -1886 -23418 -1826 -23412
rect 936 -23418 996 -23412
rect -9006 -23422 996 -23418
rect -9006 -23474 -9002 -23422
rect -8950 -23474 -7978 -23422
rect -7926 -23474 -6946 -23422
rect -6894 -23474 -5946 -23422
rect -5894 -23474 -4926 -23422
rect -4874 -23474 -3906 -23422
rect -3854 -23474 -2896 -23422
rect -2844 -23474 -1882 -23422
rect -1830 -23474 -864 -23422
rect -812 -23474 940 -23422
rect 992 -23474 996 -23422
rect -9006 -23478 996 -23474
rect -9006 -23484 -8946 -23478
rect -7982 -23484 -7922 -23478
rect -6950 -23484 -6890 -23478
rect -5950 -23484 -5890 -23478
rect -4930 -23484 -4870 -23478
rect -3910 -23484 -3850 -23478
rect -1886 -23484 -1826 -23478
rect 936 -23484 996 -23478
rect 2336 -23594 2396 -23588
rect 11724 -23594 11784 -23588
rect 13766 -23594 13826 -23588
rect 15802 -23594 15862 -23588
rect 2336 -23598 15862 -23594
rect 2336 -23650 2340 -23598
rect 2392 -23650 11728 -23598
rect 11780 -23650 13770 -23598
rect 13822 -23650 15806 -23598
rect 15858 -23650 15862 -23598
rect 2336 -23654 15862 -23650
rect 2336 -23660 2396 -23654
rect 11724 -23660 11784 -23654
rect 13766 -23660 13826 -23654
rect 15802 -23660 15862 -23654
rect 18856 -23594 18916 -23588
rect 20888 -23594 20948 -23588
rect 23034 -23594 23094 -23588
rect 18856 -23598 23094 -23594
rect 18856 -23650 18860 -23598
rect 18912 -23650 20892 -23598
rect 20944 -23650 23038 -23598
rect 23090 -23650 23094 -23598
rect 18856 -23654 23094 -23650
rect 18856 -23660 18916 -23654
rect 20888 -23660 20948 -23654
rect 23034 -23660 23094 -23654
rect 6140 -23708 6200 -23702
rect 11220 -23708 11280 -23702
rect 6140 -23712 11280 -23708
rect 2230 -23720 2290 -23714
rect 5620 -23720 5680 -23714
rect 2230 -23724 5680 -23720
rect 2230 -23776 2234 -23724
rect 2286 -23776 5624 -23724
rect 5676 -23776 5680 -23724
rect 6140 -23764 6144 -23712
rect 6196 -23764 11224 -23712
rect 11276 -23764 11280 -23712
rect 6140 -23768 11280 -23764
rect 6140 -23774 6200 -23768
rect 11220 -23774 11280 -23768
rect 16308 -23704 16368 -23698
rect 21408 -23704 21468 -23698
rect 16308 -23708 21468 -23704
rect 16308 -23760 16312 -23708
rect 16364 -23760 21412 -23708
rect 21464 -23760 21468 -23708
rect 16308 -23764 21468 -23760
rect 16308 -23770 16368 -23764
rect 21408 -23770 21468 -23764
rect 22416 -23704 22476 -23698
rect 23650 -23704 23710 -23698
rect 22416 -23708 23710 -23704
rect 22416 -23760 22420 -23708
rect 22472 -23760 23654 -23708
rect 23706 -23760 23710 -23708
rect 22416 -23764 23710 -23760
rect 22416 -23770 22476 -23764
rect 23650 -23770 23710 -23764
rect 2230 -23780 5680 -23776
rect 2230 -23786 2290 -23780
rect 5620 -23786 5680 -23780
rect 4602 -23822 4662 -23816
rect 6638 -23822 6698 -23816
rect 7658 -23822 7718 -23816
rect 8674 -23822 8734 -23816
rect 9694 -23822 9754 -23816
rect 10712 -23822 10772 -23816
rect 12742 -23822 12802 -23816
rect 14780 -23822 14840 -23816
rect 16816 -23822 16876 -23816
rect 17838 -23822 17898 -23816
rect 18858 -23822 18918 -23816
rect 19872 -23822 19932 -23816
rect 20894 -23822 20954 -23816
rect 4602 -23826 20954 -23822
rect 4602 -23878 4606 -23826
rect 4658 -23878 6642 -23826
rect 6694 -23878 7662 -23826
rect 7714 -23878 8678 -23826
rect 8730 -23878 9698 -23826
rect 9750 -23878 10716 -23826
rect 10768 -23878 12746 -23826
rect 12798 -23878 14784 -23826
rect 14836 -23878 16820 -23826
rect 16872 -23878 17842 -23826
rect 17894 -23878 18862 -23826
rect 18914 -23878 19876 -23826
rect 19928 -23878 20898 -23826
rect 20950 -23878 20954 -23826
rect 4602 -23882 20954 -23878
rect 4602 -23888 4662 -23882
rect 6638 -23888 6698 -23882
rect 7658 -23888 7718 -23882
rect 8674 -23888 8734 -23882
rect 9694 -23888 9754 -23882
rect 10712 -23888 10772 -23882
rect 12742 -23888 12802 -23882
rect 14780 -23888 14840 -23882
rect 16816 -23888 16876 -23882
rect 17838 -23888 17898 -23882
rect 18858 -23888 18918 -23882
rect 19872 -23888 19932 -23882
rect 20894 -23888 20954 -23882
rect 5620 -23926 5680 -23920
rect 10556 -23926 10616 -23920
rect 16962 -23926 17022 -23920
rect 19872 -23926 19932 -23920
rect 23054 -23926 23114 -23920
rect 5620 -23930 23114 -23926
rect 5620 -23982 5624 -23930
rect 5676 -23982 10560 -23930
rect 10612 -23982 16966 -23930
rect 17018 -23982 19876 -23930
rect 19928 -23982 23058 -23930
rect 23110 -23982 23114 -23930
rect 5620 -23986 23114 -23982
rect 5620 -23992 5680 -23986
rect 10556 -23992 10616 -23986
rect 16962 -23992 17022 -23986
rect 19872 -23992 19932 -23986
rect 23054 -23992 23114 -23986
rect -10662 -24380 -10602 -24374
rect -7992 -24380 -7932 -24374
rect -6960 -24380 -6900 -24374
rect -3900 -24380 -3840 -24374
rect -2904 -24380 -2844 -24374
rect -10662 -24384 -2844 -24380
rect -10662 -24436 -10658 -24384
rect -10606 -24436 -7988 -24384
rect -7936 -24436 -6956 -24384
rect -6904 -24436 -3896 -24384
rect -3844 -24436 -2900 -24384
rect -2848 -24436 -2844 -24384
rect -10662 -24440 -2844 -24436
rect -10662 -24446 -10602 -24440
rect -7992 -24446 -7932 -24440
rect -6960 -24446 -6900 -24440
rect -3900 -24446 -3840 -24440
rect -2904 -24446 -2844 -24440
rect -5426 -24510 -5366 -24504
rect -1366 -24510 -1306 -24504
rect 816 -24510 876 -24504
rect -9512 -24514 876 -24510
rect -9512 -24566 -9502 -24514
rect -9450 -24566 -5422 -24514
rect -5370 -24566 -1362 -24514
rect -1310 -24566 820 -24514
rect 872 -24566 876 -24514
rect -9512 -24570 876 -24566
rect -5426 -24576 -5366 -24570
rect -1366 -24576 -1306 -24570
rect 816 -24576 876 -24570
rect 2448 -24824 2508 -24818
rect 5618 -24824 5678 -24818
rect 2448 -24828 5678 -24824
rect 2448 -24880 2452 -24828
rect 2504 -24880 5622 -24828
rect 5674 -24880 5678 -24828
rect 2448 -24884 5678 -24880
rect 2448 -24890 2508 -24884
rect 5618 -24890 5678 -24884
rect 9848 -24822 9908 -24816
rect 11726 -24822 11786 -24816
rect 13764 -24822 13824 -24816
rect 15634 -24822 15694 -24816
rect 21910 -24822 21970 -24816
rect 9848 -24826 21970 -24822
rect 9848 -24878 9852 -24826
rect 9904 -24878 11730 -24826
rect 11782 -24878 13768 -24826
rect 13820 -24878 15638 -24826
rect 15690 -24878 21914 -24826
rect 21966 -24878 21970 -24826
rect 9848 -24882 21970 -24878
rect 9848 -24888 9908 -24882
rect 11726 -24888 11786 -24882
rect 13764 -24888 13824 -24882
rect 15634 -24888 15694 -24882
rect 21910 -24888 21970 -24882
rect 2120 -24928 2180 -24922
rect 3584 -24928 3644 -24922
rect 5624 -24928 5684 -24922
rect 7654 -24928 7714 -24922
rect 9694 -24928 9754 -24922
rect 11730 -24928 11790 -24922
rect 13766 -24928 13826 -24922
rect 15800 -24928 15860 -24922
rect 17840 -24928 17900 -24922
rect 19870 -24928 19930 -24922
rect 21910 -24928 21970 -24922
rect 23762 -24928 23822 -24922
rect 2120 -24932 23822 -24928
rect 2120 -24984 2124 -24932
rect 2176 -24984 3588 -24932
rect 3640 -24984 5628 -24932
rect 5680 -24984 7658 -24932
rect 7710 -24984 9698 -24932
rect 9750 -24984 11734 -24932
rect 11786 -24984 13770 -24932
rect 13822 -24984 15804 -24932
rect 15856 -24984 17844 -24932
rect 17896 -24984 19874 -24932
rect 19926 -24984 21914 -24932
rect 21966 -24984 23766 -24932
rect 23818 -24984 23822 -24932
rect 2120 -24988 23822 -24984
rect 2120 -24994 2180 -24988
rect 3584 -24994 3644 -24988
rect 5624 -24994 5684 -24988
rect 7654 -24994 7714 -24988
rect 9694 -24994 9754 -24988
rect 11730 -24994 11790 -24988
rect 13766 -24994 13826 -24988
rect 15800 -24994 15860 -24988
rect 17840 -24994 17900 -24988
rect 19870 -24994 19930 -24988
rect 21910 -24994 21970 -24988
rect 23762 -24994 23822 -24988
rect 4092 -25034 4152 -25028
rect 5112 -25034 5172 -25028
rect 6136 -25034 6196 -25028
rect 7154 -25034 7214 -25028
rect 8168 -25034 8228 -25028
rect 9200 -25034 9260 -25028
rect 10212 -25034 10272 -25028
rect 11220 -25034 11280 -25028
rect 12238 -25034 12298 -25028
rect 13264 -25034 13324 -25028
rect 14266 -25034 14326 -25028
rect 15286 -25034 15346 -25028
rect 16306 -25034 16366 -25028
rect 17332 -25034 17392 -25028
rect 18350 -25034 18410 -25028
rect 19364 -25034 19424 -25028
rect 20378 -25034 20438 -25028
rect 21400 -25034 21460 -25028
rect 4092 -25038 21460 -25034
rect 4092 -25090 4096 -25038
rect 4148 -25090 5116 -25038
rect 5168 -25090 6140 -25038
rect 6192 -25090 7158 -25038
rect 7210 -25090 8172 -25038
rect 8224 -25090 9204 -25038
rect 9256 -25090 10216 -25038
rect 10268 -25090 11224 -25038
rect 11276 -25090 12242 -25038
rect 12294 -25090 13268 -25038
rect 13320 -25090 14270 -25038
rect 14322 -25090 15290 -25038
rect 15342 -25090 16310 -25038
rect 16362 -25090 17336 -25038
rect 17388 -25090 18354 -25038
rect 18406 -25090 19368 -25038
rect 19420 -25090 20382 -25038
rect 20434 -25090 21404 -25038
rect 21456 -25090 21460 -25038
rect 4092 -25094 21460 -25090
rect 4092 -25100 4152 -25094
rect 5112 -25100 5172 -25094
rect 6136 -25100 6196 -25094
rect 7154 -25100 7214 -25094
rect 8168 -25100 8228 -25094
rect 9200 -25100 9260 -25094
rect 10212 -25100 10272 -25094
rect 11220 -25100 11280 -25094
rect 12238 -25100 12298 -25094
rect 13264 -25100 13324 -25094
rect 14266 -25100 14326 -25094
rect 15286 -25100 15346 -25094
rect 16306 -25100 16366 -25094
rect 17332 -25100 17392 -25094
rect 18350 -25100 18410 -25094
rect 19364 -25100 19424 -25094
rect 20378 -25100 20438 -25094
rect 21400 -25100 21460 -25094
rect 4604 -25144 4664 -25138
rect 6640 -25144 6700 -25138
rect 8678 -25144 8738 -25138
rect 10716 -25144 10776 -25138
rect 12752 -25144 12812 -25138
rect 14788 -25144 14848 -25138
rect 16820 -25144 16880 -25138
rect 18852 -25144 18912 -25138
rect 20892 -25144 20952 -25138
rect 4604 -25148 20952 -25144
rect 4604 -25200 4608 -25148
rect 4660 -25200 6644 -25148
rect 6696 -25200 8682 -25148
rect 8734 -25200 10720 -25148
rect 10772 -25200 12756 -25148
rect 12808 -25200 14792 -25148
rect 14844 -25200 16824 -25148
rect 16876 -25200 18856 -25148
rect 18908 -25200 20896 -25148
rect 20948 -25200 20952 -25148
rect 4604 -25204 20952 -25200
rect 4604 -25210 4664 -25204
rect 6640 -25210 6700 -25204
rect 8678 -25210 8738 -25204
rect 10716 -25210 10776 -25204
rect 12752 -25210 12812 -25204
rect 14788 -25210 14848 -25204
rect 16820 -25210 16880 -25204
rect 18852 -25210 18912 -25204
rect 20892 -25210 20952 -25204
rect -8028 -25876 -7968 -25870
rect -5990 -25876 -5930 -25870
rect -3954 -25876 -3894 -25870
rect -1918 -25876 -1858 -25870
rect -8028 -25880 -1858 -25876
rect -8028 -25932 -8024 -25880
rect -7972 -25932 -5986 -25880
rect -5934 -25932 -3950 -25880
rect -3898 -25932 -1914 -25880
rect -1862 -25932 -1858 -25880
rect -8028 -25936 -1858 -25932
rect -8028 -25942 -7968 -25936
rect -5990 -25942 -5930 -25936
rect -3954 -25942 -3894 -25936
rect -1918 -25942 -1858 -25936
rect -7010 -25988 -6950 -25982
rect -2936 -25988 -2876 -25982
rect 1070 -25988 1130 -25982
rect -7010 -25992 1130 -25988
rect -7010 -26044 -7006 -25992
rect -6954 -26044 -2932 -25992
rect -2880 -26044 1074 -25992
rect 1126 -26044 1130 -25992
rect -7010 -26048 1130 -26044
rect -7010 -26054 -6950 -26048
rect -2936 -26054 -2876 -26048
rect 1070 -26054 1130 -26048
rect 2448 -26066 2508 -26060
rect 3584 -26066 3644 -26060
rect 7654 -26066 7714 -26060
rect 17834 -26066 17894 -26060
rect 23054 -26066 23114 -26060
rect 2448 -26070 23114 -26066
rect 2448 -26122 2452 -26070
rect 2504 -26122 3588 -26070
rect 3640 -26122 7658 -26070
rect 7710 -26122 17838 -26070
rect 17890 -26122 23058 -26070
rect 23110 -26122 23114 -26070
rect 2448 -26126 23114 -26122
rect 2448 -26132 2508 -26126
rect 3584 -26132 3644 -26126
rect 7654 -26132 7714 -26126
rect 17834 -26132 17894 -26126
rect 23054 -26132 23114 -26126
rect 4096 -26174 4156 -26168
rect 12240 -26174 12300 -26168
rect 4096 -26178 21470 -26174
rect 4096 -26230 4100 -26178
rect 4152 -26230 5114 -26178
rect 5166 -26230 6136 -26178
rect 6188 -26230 7150 -26178
rect 7202 -26230 8176 -26178
rect 8228 -26230 9188 -26178
rect 9240 -26230 10224 -26178
rect 10276 -26230 11230 -26178
rect 11282 -26230 12244 -26178
rect 12296 -26230 13260 -26178
rect 13312 -26230 14268 -26178
rect 14320 -26230 15284 -26178
rect 15336 -26230 16308 -26178
rect 16360 -26230 17330 -26178
rect 17382 -26230 18352 -26178
rect 18404 -26230 19370 -26178
rect 19422 -26230 20384 -26178
rect 20436 -26230 21408 -26178
rect 21460 -26230 21470 -26178
rect 4096 -26234 21470 -26230
rect 4096 -26240 4156 -26234
rect 12240 -26240 12300 -26234
rect -8118 -26485 23968 -26430
rect -8118 -26495 -8060 -26485
rect 23916 -26495 23968 -26485
rect -8118 -26611 -8066 -26495
rect 23922 -26611 23968 -26495
rect -8118 -26621 -8060 -26611
rect 23916 -26621 23968 -26611
rect -8118 -26676 23968 -26621
rect -12216 -26818 -11616 -26806
rect -12216 -26844 -12184 -26818
rect -11648 -26844 -11616 -26818
rect -12216 -27088 -12198 -26844
rect -11634 -27088 -11616 -26844
rect -12216 -27114 -12184 -27088
rect -11648 -27114 -11616 -27088
rect -12216 -27126 -11616 -27114
rect 24216 -26818 24816 -26806
rect 24216 -26844 24248 -26818
rect 24784 -26844 24816 -26818
rect 24216 -27088 24234 -26844
rect 24798 -27088 24816 -26844
rect 24216 -27114 24248 -27088
rect 24784 -27114 24816 -27088
rect 24216 -27126 24816 -27114
<< via2 >>
rect 516 4188 1052 4214
rect 516 3944 1052 4188
rect 516 3918 1052 3944
rect 24148 4188 24684 4214
rect 24148 3944 24684 4188
rect 24148 3918 24684 3944
rect 4065 3659 4075 3795
rect 4075 3659 20831 3795
rect 20831 3659 20841 3795
rect -13597 -10632 -2901 -10416
rect 2336 -11022 2392 -10966
rect -8060 -26495 23916 -26485
rect -8060 -26611 23916 -26495
rect -8060 -26621 23916 -26611
rect -12184 -26844 -11648 -26818
rect -12184 -27088 -11648 -26844
rect -12184 -27114 -11648 -27088
rect 24248 -26844 24784 -26818
rect 24248 -27088 24784 -26844
rect 24248 -27114 24784 -27088
<< metal3 >>
rect 474 4214 1094 4221
rect 474 4178 516 4214
rect 1052 4178 1094 4214
rect 474 3954 512 4178
rect 1056 3954 1094 4178
rect 474 3918 516 3954
rect 1052 3918 1094 3954
rect 474 3911 1094 3918
rect 24106 4214 24726 4221
rect 24106 4178 24148 4214
rect 24684 4178 24726 4214
rect 24106 3954 24144 4178
rect 24688 3954 24726 4178
rect 24106 3918 24148 3954
rect 24684 3918 24726 3954
rect 24106 3911 24726 3918
rect 3998 3799 20878 3866
rect 3998 3655 4061 3799
rect 20845 3655 20878 3799
rect 3998 3600 20878 3655
rect 3998 3598 8352 3600
rect -15168 2903 -128 3086
rect -15168 2897 -941 2903
rect -15168 2273 -14980 2897
rect -14356 2279 -941 2897
rect -317 2279 -128 2903
rect -14356 2273 -128 2279
rect -15168 -10416 -128 2273
rect -15168 -10632 -13597 -10416
rect -2901 -10632 -128 -10416
rect -15168 -10978 -128 -10632
rect 2315 -10944 2413 -10939
rect 2314 -10962 2414 -10944
rect -15168 -11472 -1378 -10978
rect 2314 -11026 2332 -10962
rect 2396 -11026 2414 -10962
rect 2314 -11044 2414 -11026
rect 2315 -11049 2413 -11044
rect -15168 -11916 -1376 -11472
rect -1714 -11918 -1376 -11916
rect -8118 -26481 23968 -26430
rect -8118 -26625 -8064 -26481
rect 23920 -26625 23968 -26481
rect -8118 -26676 23968 -26625
rect -12226 -26818 -11606 -26811
rect -12226 -26854 -12184 -26818
rect -11648 -26854 -11606 -26818
rect -12226 -27078 -12188 -26854
rect -11644 -27078 -11606 -26854
rect -12226 -27114 -12184 -27078
rect -11648 -27114 -11606 -27078
rect -12226 -27121 -11606 -27114
rect 24206 -26818 24826 -26811
rect 24206 -26854 24248 -26818
rect 24784 -26854 24826 -26818
rect 24206 -27078 24244 -26854
rect 24788 -27078 24826 -26854
rect 24206 -27114 24248 -27078
rect 24784 -27114 24826 -27078
rect 24206 -27121 24826 -27114
<< via3 >>
rect 512 3954 516 4178
rect 516 3954 1052 4178
rect 1052 3954 1056 4178
rect 24144 3954 24148 4178
rect 24148 3954 24684 4178
rect 24684 3954 24688 4178
rect 4061 3795 20845 3799
rect 4061 3659 4065 3795
rect 4065 3659 20841 3795
rect 20841 3659 20845 3795
rect 4061 3655 20845 3659
rect -14980 2273 -14356 2897
rect -941 2279 -317 2903
rect 2332 -10966 2396 -10962
rect 2332 -11022 2336 -10966
rect 2336 -11022 2392 -10966
rect 2392 -11022 2396 -10966
rect 2332 -11026 2396 -11022
rect -8064 -26485 23920 -26481
rect -8064 -26621 -8060 -26485
rect -8060 -26621 23916 -26485
rect 23916 -26621 23920 -26485
rect -8064 -26625 23920 -26621
rect -12188 -27078 -12184 -26854
rect -12184 -27078 -11648 -26854
rect -11648 -27078 -11644 -26854
rect 24244 -27078 24248 -26854
rect 24248 -27078 24784 -26854
rect 24784 -27078 24788 -26854
<< mimcap >>
rect -13982 2898 -7782 2986
rect -13982 2674 -8094 2898
rect -7870 2674 -7782 2898
rect -13982 2586 -7782 2674
rect -7582 2898 -1382 2986
rect -7582 2674 -1694 2898
rect -1470 2674 -1382 2898
rect -7582 2586 -1382 2674
rect -15068 1836 -14268 1904
rect -15068 -3828 -14580 1836
rect -14356 -3828 -14268 1836
rect -1024 1836 -224 1904
rect -13128 898 -7928 986
rect -13128 -3726 -8240 898
rect -8016 -3726 -7928 898
rect -13128 -3814 -7928 -3726
rect -7528 898 -2328 986
rect -7528 -3726 -2640 898
rect -2416 -3726 -2328 898
rect -7528 -3814 -2328 -3726
rect -15068 -3896 -14268 -3828
rect -1024 -3828 -536 1836
rect -312 -3828 -224 1836
rect -1024 -3896 -224 -3828
rect -15068 -4656 -14268 -4588
rect -15068 -10320 -14580 -4656
rect -14356 -10320 -14268 -4656
rect -13128 -4702 -7928 -4614
rect -13128 -9326 -8240 -4702
rect -8016 -9326 -7928 -4702
rect -13128 -9414 -7928 -9326
rect -7528 -4702 -2328 -4614
rect -7528 -9326 -2640 -4702
rect -2416 -9326 -2328 -4702
rect -7528 -9414 -2328 -9326
rect -1024 -4656 -224 -4588
rect -15068 -10388 -14268 -10320
rect -1024 -10320 -536 -4656
rect -312 -10320 -224 -4656
rect -1024 -10388 -224 -10320
rect -14482 -11102 -8282 -11014
rect -14482 -11326 -8594 -11102
rect -8370 -11326 -8282 -11102
rect -14482 -11414 -8282 -11326
rect -8082 -11102 -1882 -11014
rect -8082 -11326 -2194 -11102
rect -1970 -11326 -1882 -11102
rect -8082 -11414 -1882 -11326
<< mimcapcontact >>
rect -8094 2674 -7870 2898
rect -1694 2674 -1470 2898
rect -14580 -3828 -14356 1836
rect -8240 -3726 -8016 898
rect -2640 -3726 -2416 898
rect -536 -3828 -312 1836
rect -14580 -10320 -14356 -4656
rect -8240 -9326 -8016 -4702
rect -2640 -9326 -2416 -4702
rect -536 -10320 -312 -4656
rect -8594 -11326 -8370 -11102
rect -2194 -11326 -1970 -11102
<< metal4 >>
rect -15168 4178 25000 4400
rect -15168 3954 512 4178
rect 1056 3954 24144 4178
rect 24688 3954 25000 4178
rect -15168 3799 25000 3954
rect -15168 3655 4061 3799
rect 20845 3655 25000 3799
rect -15168 3600 25000 3655
rect -15168 2903 -128 3086
rect -15168 2898 -941 2903
rect -15168 2897 -8094 2898
rect -15168 2273 -14980 2897
rect -14356 2674 -8094 2897
rect -7870 2674 -1694 2898
rect -1470 2674 -941 2898
rect -14356 2279 -941 2674
rect -317 2279 -128 2903
rect -14356 2273 -128 2279
rect -15168 1910 -128 2273
rect -15168 1836 -13986 1910
rect -15168 -3828 -14580 1836
rect -14356 -3828 -13986 1836
rect -1428 1836 -128 1910
rect -15168 -4656 -13986 -3828
rect -15168 -10320 -14580 -4656
rect -14356 -10320 -13986 -4656
rect -13228 898 -2228 1086
rect -13228 -3726 -8240 898
rect -8016 -3726 -2640 898
rect -2416 -3726 -2228 898
rect -13228 -4702 -2228 -3726
rect -13228 -9326 -8240 -4702
rect -8016 -9326 -2640 -4702
rect -2416 -9326 -2228 -4702
rect -13228 -9816 -2228 -9326
rect -1428 -3828 -536 1836
rect -312 -3828 -128 1836
rect -1428 -4656 -128 -3828
rect -1428 -9436 -536 -4656
rect -13228 -9913 -1327 -9816
rect -13228 -9914 -2228 -9913
rect -15168 -10752 -13986 -10320
rect -15168 -10838 -2722 -10752
rect -15166 -10978 -2722 -10838
rect -15166 -11102 -1722 -10978
rect -15166 -11326 -8594 -11102
rect -8370 -11326 -2194 -11102
rect -1970 -11326 -1722 -11102
rect -15166 -11916 -1722 -11326
rect -1424 -11400 -1327 -9913
rect -1058 -10320 -536 -9436
rect -312 -10320 -128 -4656
rect -1058 -10848 -128 -10320
rect 226 -10962 2414 -10944
rect 226 -11026 2332 -10962
rect 2396 -11026 2414 -10962
rect 226 -11044 2414 -11026
rect 226 -11400 326 -11044
rect -1424 -11500 326 -11400
rect -15168 -26481 25000 -26400
rect -15168 -26625 -8064 -26481
rect 23920 -26625 25000 -26481
rect -15168 -26854 25000 -26625
rect -15168 -27078 -12188 -26854
rect -11644 -27078 24244 -26854
rect 24788 -27078 25000 -26854
rect -15168 -27200 25000 -27078
<< via4 >>
rect -14946 2307 -14390 2863
rect -907 2313 -351 2869
<< mimcap2 >>
rect -13982 2504 -8182 2986
rect -13982 2268 -13920 2504
rect -8244 2268 -8182 2504
rect -13982 2186 -8182 2268
rect -7582 2504 -1782 2986
rect -7582 2268 -7520 2504
rect -1844 2268 -1782 2504
rect -7582 2186 -1782 2268
rect -15068 -3978 -14668 1904
rect -15068 -4214 -14986 -3978
rect -14750 -4214 -14668 -3978
rect -13128 -3896 -8328 986
rect -13128 -4132 -12926 -3896
rect -8530 -4132 -8328 -3896
rect -13128 -4214 -8328 -4132
rect -7528 -3896 -2728 986
rect -7528 -4132 -7326 -3896
rect -2930 -4132 -2728 -3896
rect -7528 -4214 -2728 -4132
rect -1024 -3978 -624 1904
rect -1024 -4214 -942 -3978
rect -706 -4214 -624 -3978
rect -15068 -4296 -14668 -4214
rect -1024 -4296 -624 -4214
rect -15068 -10470 -14668 -4588
rect -13128 -9496 -8328 -4614
rect -13128 -9732 -12926 -9496
rect -8530 -9732 -8328 -9496
rect -13128 -9814 -8328 -9732
rect -7528 -9496 -2728 -4614
rect -7528 -9732 -7326 -9496
rect -2930 -9732 -2728 -9496
rect -7528 -9814 -2728 -9732
rect -15068 -10706 -14986 -10470
rect -14750 -10706 -14668 -10470
rect -15068 -10788 -14668 -10706
rect -1024 -10463 -624 -4588
rect -1024 -10699 -942 -10463
rect -706 -10699 -624 -10463
rect -1024 -10788 -624 -10699
rect -14482 -11496 -8682 -11014
rect -14482 -11732 -14420 -11496
rect -8744 -11732 -8682 -11496
rect -14482 -11814 -8682 -11732
rect -8082 -11496 -2282 -11014
rect -8082 -11732 -8020 -11496
rect -2344 -11732 -2282 -11496
rect -8082 -11814 -2282 -11732
<< mimcap2contact >>
rect -13920 2268 -8244 2504
rect -7520 2268 -1844 2504
rect -14986 -4214 -14750 -3978
rect -12926 -4132 -8530 -3896
rect -7326 -4132 -2930 -3896
rect -942 -4214 -706 -3978
rect -12926 -9732 -8530 -9496
rect -7326 -9732 -2930 -9496
rect -14986 -10706 -14750 -10470
rect -942 -10699 -706 -10463
rect -14420 -11732 -8744 -11496
rect -8020 -11732 -2344 -11496
<< metal5 >>
rect -15168 2869 -128 3086
rect -15168 2863 -907 2869
rect -15168 2307 -14946 2863
rect -14390 2504 -907 2863
rect -14390 2307 -13920 2504
rect -15168 2268 -13920 2307
rect -8244 2268 -7520 2504
rect -1844 2313 -907 2504
rect -351 2313 -128 2869
rect -1844 2268 -128 2313
rect -15168 -3896 -128 2268
rect -15168 -3978 -12926 -3896
rect -15168 -4214 -14986 -3978
rect -14750 -4132 -12926 -3978
rect -8530 -4132 -7326 -3896
rect -2930 -3978 -128 -3896
rect -2930 -4132 -942 -3978
rect -14750 -4214 -942 -4132
rect -706 -4214 -128 -3978
rect -15168 -9496 -128 -4214
rect -15168 -9732 -12926 -9496
rect -8530 -9732 -7326 -9496
rect -2930 -9732 -128 -9496
rect -15168 -10463 -128 -9732
rect -15168 -10470 -942 -10463
rect -15168 -10706 -14986 -10470
rect -14750 -10699 -942 -10470
rect -706 -10699 -128 -10463
rect -14750 -10706 -128 -10699
rect -15168 -10764 -128 -10706
rect -15168 -11496 -130 -10764
rect -15168 -11732 -14420 -11496
rect -8744 -11732 -8020 -11496
rect -2344 -11732 -130 -11496
rect -15168 -11916 -130 -11732
use ptap  ptap_395
timestamp 1626486988
transform 1 0 -10304 0 1 -26298
box 62 116 196 250
use ptap  ptap_394
timestamp 1626486988
transform 1 0 -9286 0 1 -26298
box 62 116 196 250
use ptap  ptap_392
timestamp 1626486988
transform 1 0 -8268 0 1 -26298
box 62 116 196 250
use ptap  ptap_391
timestamp 1626486988
transform 1 0 -6232 0 1 -26298
box 62 116 196 250
use ptap  ptap_393
timestamp 1626486988
transform 1 0 -7250 0 1 -26298
box 62 116 196 250
use ptap  ptap_390
timestamp 1626486988
transform 1 0 -5214 0 1 -26298
box 62 116 196 250
use ptap  ptap_389
timestamp 1626486988
transform 1 0 -4196 0 1 -26298
box 62 116 196 250
use ptap  ptap_388
timestamp 1626486988
transform 1 0 -3178 0 1 -26298
box 62 116 196 250
use ptap  ptap_387
timestamp 1626486988
transform 1 0 -2160 0 1 -26298
box 62 116 196 250
use ptap  ptap_386
timestamp 1626486988
transform 1 0 -1142 0 1 -26298
box 62 116 196 250
use ptap  ptap_385
timestamp 1626486988
transform 1 0 -124 0 1 -26298
box 62 116 196 250
use ptap  ptap_384
timestamp 1626486988
transform 1 0 2986 0 1 -26380
box 62 116 196 250
use ptap  ptap_382
timestamp 1626486988
transform 1 0 4004 0 1 -26380
box 62 116 196 250
use ptap  ptap_383
timestamp 1626486988
transform 1 0 5022 0 1 -26380
box 62 116 196 250
use ptap  ptap_381
timestamp 1626486988
transform 1 0 6040 0 1 -26380
box 62 116 196 250
use sky130_fd_pr__nfet_01v8_FYXD5N  sky130_fd_pr__nfet_01v8_FYXD5N_0
timestamp 1626486988
transform 1 0 -4943 0 1 -25440
box -5145 -388 5145 388
use ptap  ptap_380
timestamp 1626486988
transform 1 0 7058 0 1 -26380
box 62 116 196 250
use ptap  ptap_379
timestamp 1626486988
transform 1 0 8076 0 1 -26380
box 62 116 196 250
use ptap  ptap_378
timestamp 1626486988
transform 1 0 9094 0 1 -26380
box 62 116 196 250
use ptap  ptap_377
timestamp 1626486988
transform 1 0 10112 0 1 -26380
box 62 116 196 250
use ptap  ptap_376
timestamp 1626486988
transform 1 0 11130 0 1 -26380
box 62 116 196 250
use ptap  ptap_375
timestamp 1626486988
transform 1 0 12148 0 1 -26380
box 62 116 196 250
use ptap  ptap_374
timestamp 1626486988
transform 1 0 13166 0 1 -26380
box 62 116 196 250
use ptap  ptap_373
timestamp 1626486988
transform 1 0 14184 0 1 -26380
box 62 116 196 250
use ptap  ptap_372
timestamp 1626486988
transform 1 0 15202 0 1 -26380
box 62 116 196 250
use ptap  ptap_371
timestamp 1626486988
transform 1 0 16220 0 1 -26380
box 62 116 196 250
use ptap  ptap_370
timestamp 1626486988
transform 1 0 17238 0 1 -26380
box 62 116 196 250
use ptap  ptap_369
timestamp 1626486988
transform 1 0 18256 0 1 -26380
box 62 116 196 250
use ptap  ptap_368
timestamp 1626486988
transform 1 0 19274 0 1 -26380
box 62 116 196 250
use ptap  ptap_367
timestamp 1626486988
transform 1 0 20292 0 1 -26380
box 62 116 196 250
use ptap  ptap_366
timestamp 1626486988
transform 1 0 21310 0 1 -26380
box 62 116 196 250
use ptap  ptap_365
timestamp 1626486988
transform 1 0 22328 0 1 -26380
box 62 116 196 250
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_9
timestamp 1626486988
transform -1 0 12777 0 -1 -25630
box -10235 -388 10235 388
use ptap  ptap_364
timestamp 1626486988
transform 1 0 -10114 0 1 -24852
box 62 116 196 250
use ptap  ptap_363
timestamp 1626486988
transform 1 0 -9096 0 1 -24852
box 62 116 196 250
use ptap  ptap_362
timestamp 1626486988
transform 1 0 -8078 0 1 -24852
box 62 116 196 250
use ptap  ptap_361
timestamp 1626486988
transform 1 0 -7060 0 1 -24852
box 62 116 196 250
use ptap  ptap_360
timestamp 1626486988
transform 1 0 -6042 0 1 -24852
box 62 116 196 250
use ptap  ptap_359
timestamp 1626486988
transform 1 0 -5024 0 1 -24852
box 62 116 196 250
use ptap  ptap_358
timestamp 1626486988
transform 1 0 -4006 0 1 -24852
box 62 116 196 250
use ptap  ptap_357
timestamp 1626486988
transform 1 0 -2988 0 1 -24852
box 62 116 196 250
use ptap  ptap_356
timestamp 1626486988
transform 1 0 -1970 0 1 -24852
box 62 116 196 250
use ptap  ptap_355
timestamp 1626486988
transform 1 0 -952 0 1 -24852
box 62 116 196 250
use ptap  ptap_354
timestamp 1626486988
transform 1 0 66 0 1 -24852
box 62 116 196 250
use ptap  ptap_353
timestamp 1626486988
transform 1 0 2998 0 1 -25202
box 62 116 196 250
use ptap  ptap_352
timestamp 1626486988
transform 1 0 4016 0 1 -25202
box 62 116 196 250
use ptap  ptap_351
timestamp 1626486988
transform 1 0 5034 0 1 -25202
box 62 116 196 250
use ptap  ptap_350
timestamp 1626486988
transform 1 0 6052 0 1 -25202
box 62 116 196 250
use ptap  ptap_349
timestamp 1626486988
transform 1 0 7070 0 1 -25202
box 62 116 196 250
use ptap  ptap_348
timestamp 1626486988
transform 1 0 8088 0 1 -25202
box 62 116 196 250
use ptap  ptap_347
timestamp 1626486988
transform 1 0 9106 0 1 -25202
box 62 116 196 250
use ptap  ptap_346
timestamp 1626486988
transform 1 0 10124 0 1 -25202
box 62 116 196 250
use ptap  ptap_345
timestamp 1626486988
transform 1 0 11142 0 1 -25202
box 62 116 196 250
use ptap  ptap_344
timestamp 1626486988
transform 1 0 12160 0 1 -25202
box 62 116 196 250
use ptap  ptap_343
timestamp 1626486988
transform 1 0 13178 0 1 -25202
box 62 116 196 250
use ptap  ptap_342
timestamp 1626486988
transform 1 0 14196 0 1 -25202
box 62 116 196 250
use ptap  ptap_341
timestamp 1626486988
transform 1 0 15214 0 1 -25202
box 62 116 196 250
use ptap  ptap_340
timestamp 1626486988
transform 1 0 16232 0 1 -25202
box 62 116 196 250
use ptap  ptap_339
timestamp 1626486988
transform 1 0 17250 0 1 -25202
box 62 116 196 250
use ptap  ptap_338
timestamp 1626486988
transform 1 0 18268 0 1 -25202
box 62 116 196 250
use ptap  ptap_337
timestamp 1626486988
transform 1 0 19286 0 1 -25202
box 62 116 196 250
use ptap  ptap_336
timestamp 1626486988
transform 1 0 20304 0 1 -25202
box 62 116 196 250
use ptap  ptap_335
timestamp 1626486988
transform 1 0 21322 0 1 -25202
box 62 116 196 250
use ptap  ptap_334
timestamp 1626486988
transform 1 0 22340 0 1 -25202
box 62 116 196 250
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_8
timestamp 1626486988
transform 1 0 12777 0 1 -24398
box -10235 -388 10235 388
use sky130_fd_pr__nfet_01v8_lvt_ZYX5GY  sky130_fd_pr__nfet_01v8_lvt_ZYX5GY_3
timestamp 1626486988
transform 1 0 -4892 0 1 -23898
box -5654 -388 5654 388
use ptap  ptap_333
timestamp 1626486988
transform 1 0 2986 0 1 -23956
box 62 116 196 250
use ptap  ptap_332
timestamp 1626486988
transform 1 0 4004 0 1 -23956
box 62 116 196 250
use ptap  ptap_331
timestamp 1626486988
transform 1 0 5022 0 1 -23956
box 62 116 196 250
use ptap  ptap_330
timestamp 1626486988
transform 1 0 6040 0 1 -23956
box 62 116 196 250
use ptap  ptap_328
timestamp 1626486988
transform 1 0 -9096 0 1 -23510
box 62 116 196 250
use ptap  ptap_329
timestamp 1626486988
transform 1 0 -10114 0 1 -23510
box 62 116 196 250
use ptap  ptap_327
timestamp 1626486988
transform 1 0 -8078 0 1 -23510
box 62 116 196 250
use ptap  ptap_325
timestamp 1626486988
transform 1 0 -7060 0 1 -23510
box 62 116 196 250
use ptap  ptap_326
timestamp 1626486988
transform 1 0 -6042 0 1 -23510
box 62 116 196 250
use ptap  ptap_324
timestamp 1626486988
transform 1 0 -5024 0 1 -23510
box 62 116 196 250
use ptap  ptap_322
timestamp 1626486988
transform 1 0 -2988 0 1 -23510
box 62 116 196 250
use ptap  ptap_323
timestamp 1626486988
transform 1 0 -4006 0 1 -23510
box 62 116 196 250
use ptap  ptap_321
timestamp 1626486988
transform 1 0 -1970 0 1 -23510
box 62 116 196 250
use ptap  ptap_319
timestamp 1626486988
transform 1 0 -952 0 1 -23510
box 62 116 196 250
use ptap  ptap_320
timestamp 1626486988
transform 1 0 66 0 1 -23510
box 62 116 196 250
use sky130_fd_pr__nfet_01v8_lvt_ZYX5GY  sky130_fd_pr__nfet_01v8_lvt_ZYX5GY_2
timestamp 1626486988
transform 1 0 -4892 0 1 -22786
box -5654 -388 5654 388
use ptap  ptap_318
timestamp 1626486988
transform 1 0 7058 0 1 -23956
box 62 116 196 250
use ptap  ptap_317
timestamp 1626486988
transform 1 0 8076 0 1 -23956
box 62 116 196 250
use ptap  ptap_316
timestamp 1626486988
transform 1 0 9094 0 1 -23956
box 62 116 196 250
use ptap  ptap_315
timestamp 1626486988
transform 1 0 10112 0 1 -23956
box 62 116 196 250
use ptap  ptap_314
timestamp 1626486988
transform 1 0 11130 0 1 -23956
box 62 116 196 250
use ptap  ptap_313
timestamp 1626486988
transform 1 0 12148 0 1 -23956
box 62 116 196 250
use ptap  ptap_312
timestamp 1626486988
transform 1 0 13166 0 1 -23956
box 62 116 196 250
use ptap  ptap_311
timestamp 1626486988
transform 1 0 14184 0 1 -23956
box 62 116 196 250
use ptap  ptap_310
timestamp 1626486988
transform 1 0 15202 0 1 -23956
box 62 116 196 250
use ptap  ptap_309
timestamp 1626486988
transform 1 0 16220 0 1 -23956
box 62 116 196 250
use ptap  ptap_308
timestamp 1626486988
transform 1 0 17238 0 1 -23956
box 62 116 196 250
use ptap  ptap_307
timestamp 1626486988
transform 1 0 18256 0 1 -23956
box 62 116 196 250
use ptap  ptap_306
timestamp 1626486988
transform 1 0 19274 0 1 -23956
box 62 116 196 250
use ptap  ptap_305
timestamp 1626486988
transform 1 0 20292 0 1 -23956
box 62 116 196 250
use ptap  ptap_304
timestamp 1626486988
transform 1 0 21310 0 1 -23956
box 62 116 196 250
use ptap  ptap_303
timestamp 1626486988
transform 1 0 22328 0 1 -23956
box 62 116 196 250
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_7
timestamp 1626486988
transform 1 0 12777 0 1 -23164
box -10235 -388 10235 388
use ptap  ptap_302
timestamp 1626486988
transform 1 0 -10114 0 1 -22404
box 62 116 196 250
use ptap  ptap_301
timestamp 1626486988
transform 1 0 -9096 0 1 -22404
box 62 116 196 250
use ptap  ptap_300
timestamp 1626486988
transform 1 0 -8078 0 1 -22404
box 62 116 196 250
use ptap  ptap_299
timestamp 1626486988
transform 1 0 -7060 0 1 -22404
box 62 116 196 250
use ptap  ptap_298
timestamp 1626486988
transform 1 0 -6042 0 1 -22404
box 62 116 196 250
use ptap  ptap_297
timestamp 1626486988
transform 1 0 -5024 0 1 -22404
box 62 116 196 250
use ptap  ptap_296
timestamp 1626486988
transform 1 0 -4006 0 1 -22404
box 62 116 196 250
use ptap  ptap_295
timestamp 1626486988
transform 1 0 -2988 0 1 -22404
box 62 116 196 250
use ptap  ptap_294
timestamp 1626486988
transform 1 0 -1970 0 1 -22404
box 62 116 196 250
use ptap  ptap_293
timestamp 1626486988
transform 1 0 -952 0 1 -22404
box 62 116 196 250
use ptap  ptap_292
timestamp 1626486988
transform 1 0 66 0 1 -22404
box 62 116 196 250
use ptap  ptap_291
timestamp 1626486988
transform 1 0 2986 0 1 -22720
box 62 116 196 250
use ptap  ptap_290
timestamp 1626486988
transform 1 0 4004 0 1 -22720
box 62 116 196 250
use ptap  ptap_289
timestamp 1626486988
transform 1 0 5022 0 1 -22720
box 62 116 196 250
use ptap  ptap_288
timestamp 1626486988
transform 1 0 6040 0 1 -22720
box 62 116 196 250
use ptap  ptap_287
timestamp 1626486988
transform 1 0 7058 0 1 -22720
box 62 116 196 250
use ptap  ptap_286
timestamp 1626486988
transform 1 0 8076 0 1 -22720
box 62 116 196 250
use ptap  ptap_285
timestamp 1626486988
transform 1 0 9094 0 1 -22720
box 62 116 196 250
use ptap  ptap_284
timestamp 1626486988
transform 1 0 10112 0 1 -22720
box 62 116 196 250
use ptap  ptap_283
timestamp 1626486988
transform 1 0 11130 0 1 -22720
box 62 116 196 250
use ptap  ptap_282
timestamp 1626486988
transform 1 0 12148 0 1 -22720
box 62 116 196 250
use ptap  ptap_281
timestamp 1626486988
transform 1 0 13166 0 1 -22720
box 62 116 196 250
use ptap  ptap_280
timestamp 1626486988
transform 1 0 14184 0 1 -22720
box 62 116 196 250
use ptap  ptap_279
timestamp 1626486988
transform 1 0 15202 0 1 -22720
box 62 116 196 250
use ptap  ptap_278
timestamp 1626486988
transform 1 0 16220 0 1 -22720
box 62 116 196 250
use ptap  ptap_277
timestamp 1626486988
transform 1 0 17238 0 1 -22720
box 62 116 196 250
use ptap  ptap_276
timestamp 1626486988
transform 1 0 18256 0 1 -22720
box 62 116 196 250
use ptap  ptap_275
timestamp 1626486988
transform 1 0 19274 0 1 -22720
box 62 116 196 250
use ptap  ptap_274
timestamp 1626486988
transform 1 0 20292 0 1 -22720
box 62 116 196 250
use ptap  ptap_273
timestamp 1626486988
transform 1 0 21310 0 1 -22720
box 62 116 196 250
use ptap  ptap_272
timestamp 1626486988
transform 1 0 22328 0 1 -22720
box 62 116 196 250
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_6
timestamp 1626486988
transform 1 0 12777 0 1 -21932
box -10235 -388 10235 388
use sky130_fd_pr__nfet_01v8_lvt_ZYX5GY  sky130_fd_pr__nfet_01v8_lvt_ZYX5GY_1
timestamp 1626486988
transform 1 0 -4892 0 1 -21674
box -5654 -388 5654 388
use ptap  ptap_271
timestamp 1626486988
transform 1 0 -10092 0 1 -21296
box 62 116 196 250
use ptap  ptap_270
timestamp 1626486988
transform 1 0 -9074 0 1 -21296
box 62 116 196 250
use ptap  ptap_269
timestamp 1626486988
transform 1 0 -8056 0 1 -21296
box 62 116 196 250
use ptap  ptap_268
timestamp 1626486988
transform 1 0 -7038 0 1 -21296
box 62 116 196 250
use ptap  ptap_267
timestamp 1626486988
transform 1 0 -6020 0 1 -21296
box 62 116 196 250
use ptap  ptap_265
timestamp 1626486988
transform 1 0 -5002 0 1 -21296
box 62 116 196 250
use ptap  ptap_266
timestamp 1626486988
transform 1 0 -3984 0 1 -21296
box 62 116 196 250
use ptap  ptap_264
timestamp 1626486988
transform 1 0 -2966 0 1 -21296
box 62 116 196 250
use ptap  ptap_263
timestamp 1626486988
transform 1 0 -1948 0 1 -21296
box 62 116 196 250
use ptap  ptap_262
timestamp 1626486988
transform 1 0 -930 0 1 -21296
box 62 116 196 250
use ptap  ptap_261
timestamp 1626486988
transform 1 0 88 0 1 -21296
box 62 116 196 250
use ptap  ptap_260
timestamp 1626486988
transform 1 0 2974 0 1 -21496
box 62 116 196 250
use ptap  ptap_258
timestamp 1626486988
transform 1 0 3992 0 1 -21496
box 62 116 196 250
use ptap  ptap_259
timestamp 1626486988
transform 1 0 5010 0 1 -21496
box 62 116 196 250
use ptap  ptap_257
timestamp 1626486988
transform 1 0 6028 0 1 -21496
box 62 116 196 250
use sky130_fd_pr__nfet_01v8_lvt_ZYX5GY  sky130_fd_pr__nfet_01v8_lvt_ZYX5GY_0
timestamp 1626486988
transform 1 0 -4892 0 1 -20562
box -5654 -388 5654 388
use ptap  ptap_256
timestamp 1626486988
transform 1 0 7046 0 1 -21496
box 62 116 196 250
use ptap  ptap_255
timestamp 1626486988
transform 1 0 8064 0 1 -21496
box 62 116 196 250
use ptap  ptap_254
timestamp 1626486988
transform 1 0 9082 0 1 -21496
box 62 116 196 250
use ptap  ptap_253
timestamp 1626486988
transform 1 0 10100 0 1 -21496
box 62 116 196 250
use ptap  ptap_252
timestamp 1626486988
transform 1 0 11118 0 1 -21496
box 62 116 196 250
use ptap  ptap_251
timestamp 1626486988
transform 1 0 12136 0 1 -21496
box 62 116 196 250
use ptap  ptap_250
timestamp 1626486988
transform 1 0 13154 0 1 -21496
box 62 116 196 250
use ptap  ptap_249
timestamp 1626486988
transform 1 0 14172 0 1 -21496
box 62 116 196 250
use ptap  ptap_248
timestamp 1626486988
transform 1 0 15190 0 1 -21496
box 62 116 196 250
use ptap  ptap_247
timestamp 1626486988
transform 1 0 16208 0 1 -21496
box 62 116 196 250
use ptap  ptap_246
timestamp 1626486988
transform 1 0 17226 0 1 -21496
box 62 116 196 250
use ptap  ptap_245
timestamp 1626486988
transform 1 0 18244 0 1 -21496
box 62 116 196 250
use ptap  ptap_244
timestamp 1626486988
transform 1 0 19262 0 1 -21496
box 62 116 196 250
use ptap  ptap_243
timestamp 1626486988
transform 1 0 20280 0 1 -21496
box 62 116 196 250
use ptap  ptap_242
timestamp 1626486988
transform 1 0 21298 0 1 -21496
box 62 116 196 250
use ptap  ptap_241
timestamp 1626486988
transform 1 0 22316 0 1 -21496
box 62 116 196 250
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_5
timestamp 1626486988
transform 1 0 12777 0 1 -20698
box -10235 -388 10235 388
use ptap  ptap_240
timestamp 1626486988
transform 1 0 -10104 0 1 -20154
box 62 116 196 250
use ptap  ptap_239
timestamp 1626486988
transform 1 0 -9086 0 1 -20154
box 62 116 196 250
use ptap  ptap_238
timestamp 1626486988
transform 1 0 -8068 0 1 -20154
box 62 116 196 250
use ptap  ptap_237
timestamp 1626486988
transform 1 0 -7050 0 1 -20154
box 62 116 196 250
use ptap  ptap_236
timestamp 1626486988
transform 1 0 -6032 0 1 -20154
box 62 116 196 250
use ptap  ptap_235
timestamp 1626486988
transform 1 0 -5014 0 1 -20154
box 62 116 196 250
use ptap  ptap_234
timestamp 1626486988
transform 1 0 -3996 0 1 -20154
box 62 116 196 250
use ptap  ptap_232
timestamp 1626486988
transform 1 0 -2978 0 1 -20154
box 62 116 196 250
use ptap  ptap_233
timestamp 1626486988
transform 1 0 -1960 0 1 -20154
box 62 116 196 250
use ptap  ptap_231
timestamp 1626486988
transform 1 0 -942 0 1 -20154
box 62 116 196 250
use ptap  ptap_230
timestamp 1626486988
transform 1 0 76 0 1 -20154
box 62 116 196 250
use ptap  ptap_229
timestamp 1626486988
transform 1 0 2998 0 1 -20260
box 62 116 196 250
use ptap  ptap_228
timestamp 1626486988
transform 1 0 4016 0 1 -20260
box 62 116 196 250
use ptap  ptap_227
timestamp 1626486988
transform 1 0 5034 0 1 -20260
box 62 116 196 250
use ptap  ptap_226
timestamp 1626486988
transform 1 0 6052 0 1 -20260
box 62 116 196 250
use ptap  ptap_225
timestamp 1626486988
transform 1 0 7070 0 1 -20260
box 62 116 196 250
use ptap  ptap_224
timestamp 1626486988
transform 1 0 8088 0 1 -20260
box 62 116 196 250
use ptap  ptap_223
timestamp 1626486988
transform 1 0 9106 0 1 -20260
box 62 116 196 250
use ptap  ptap_222
timestamp 1626486988
transform 1 0 10124 0 1 -20260
box 62 116 196 250
use ptap  ptap_221
timestamp 1626486988
transform 1 0 11142 0 1 -20260
box 62 116 196 250
use ptap  ptap_219
timestamp 1626486988
transform 1 0 12160 0 1 -20260
box 62 116 196 250
use ptap  ptap_220
timestamp 1626486988
transform 1 0 13178 0 1 -20260
box 62 116 196 250
use ptap  ptap_218
timestamp 1626486988
transform 1 0 14196 0 1 -20260
box 62 116 196 250
use ptap  ptap_217
timestamp 1626486988
transform 1 0 15214 0 1 -20260
box 62 116 196 250
use ptap  ptap_216
timestamp 1626486988
transform 1 0 16232 0 1 -20260
box 62 116 196 250
use ptap  ptap_215
timestamp 1626486988
transform 1 0 17250 0 1 -20260
box 62 116 196 250
use ptap  ptap_214
timestamp 1626486988
transform 1 0 18268 0 1 -20260
box 62 116 196 250
use ptap  ptap_213
timestamp 1626486988
transform 1 0 19286 0 1 -20260
box 62 116 196 250
use ptap  ptap_212
timestamp 1626486988
transform 1 0 20304 0 1 -20260
box 62 116 196 250
use ptap  ptap_211
timestamp 1626486988
transform 1 0 21322 0 1 -20260
box 62 116 196 250
use ptap  ptap_210
timestamp 1626486988
transform 1 0 22340 0 1 -20260
box 62 116 196 250
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_4
timestamp 1626486988
transform 1 0 12777 0 1 -19464
box -10235 -388 10235 388
use ptap  ptap_209
timestamp 1626486988
transform 1 0 -9308 0 1 -19206
box 62 116 196 250
use ptap  ptap_208
timestamp 1626486988
transform 1 0 -7272 0 1 -19206
box 62 116 196 250
use ptap  ptap_207
timestamp 1626486988
transform 1 0 -8290 0 1 -19206
box 62 116 196 250
use ptap  ptap_206
timestamp 1626486988
transform 1 0 -4218 0 1 -19206
box 62 116 196 250
use ptap  ptap_205
timestamp 1626486988
transform 1 0 -6254 0 1 -19206
box 62 116 196 250
use ptap  ptap_204
timestamp 1626486988
transform 1 0 -5236 0 1 -19206
box 62 116 196 250
use ptap  ptap_203
timestamp 1626486988
transform 1 0 -2182 0 1 -19206
box 62 116 196 250
use ptap  ptap_202
timestamp 1626486988
transform 1 0 -1164 0 1 -19206
box 62 116 196 250
use ptap  ptap_201
timestamp 1626486988
transform 1 0 -3200 0 1 -19206
box 62 116 196 250
use ptap  ptap_200
timestamp 1626486988
transform 1 0 -136 0 1 -19206
box 62 116 196 250
use ptap  ptap_198
timestamp 1626486988
transform 1 0 2998 0 1 -19012
box 62 116 196 250
use ptap  ptap_199
timestamp 1626486988
transform 1 0 4016 0 1 -19012
box 62 116 196 250
use ptap  ptap_196
timestamp 1626486988
transform 1 0 5034 0 1 -19012
box 62 116 196 250
use ptap  ptap_197
timestamp 1626486988
transform 1 0 6052 0 1 -19012
box 62 116 196 250
use ptap  ptap_195
timestamp 1626486988
transform 1 0 7070 0 1 -19012
box 62 116 196 250
use ptap  ptap_193
timestamp 1626486988
transform 1 0 9106 0 1 -19012
box 62 116 196 250
use ptap  ptap_194
timestamp 1626486988
transform 1 0 8088 0 1 -19012
box 62 116 196 250
use ptap  ptap_191
timestamp 1626486988
transform 1 0 10124 0 1 -19012
box 62 116 196 250
use ptap  ptap_192
timestamp 1626486988
transform 1 0 11142 0 1 -19012
box 62 116 196 250
use ptap  ptap_190
timestamp 1626486988
transform 1 0 12160 0 1 -19012
box 62 116 196 250
use ptap  ptap_188
timestamp 1626486988
transform 1 0 13178 0 1 -19012
box 62 116 196 250
use ptap  ptap_189
timestamp 1626486988
transform 1 0 14196 0 1 -19012
box 62 116 196 250
use ptap  ptap_185
timestamp 1626486988
transform 1 0 16232 0 1 -19012
box 62 116 196 250
use ptap  ptap_187
timestamp 1626486988
transform 1 0 15214 0 1 -19012
box 62 116 196 250
use ptap  ptap_186
timestamp 1626486988
transform 1 0 17250 0 1 -19012
box 62 116 196 250
use ptap  ptap_183
timestamp 1626486988
transform 1 0 18268 0 1 -19012
box 62 116 196 250
use ptap  ptap_184
timestamp 1626486988
transform 1 0 19286 0 1 -19012
box 62 116 196 250
use ptap  ptap_182
timestamp 1626486988
transform 1 0 20304 0 1 -19012
box 62 116 196 250
use ptap  ptap_180
timestamp 1626486988
transform 1 0 21322 0 1 -19012
box 62 116 196 250
use ptap  ptap_181
timestamp 1626486988
transform 1 0 22340 0 1 -19012
box 62 116 196 250
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_3
timestamp 1626486988
transform 1 0 12777 0 1 -18232
box -10235 -388 10235 388
use ptap  ptap_179
timestamp 1626486988
transform 1 0 -9296 0 1 -18312
box 62 116 196 250
use ptap  ptap_178
timestamp 1626486988
transform 1 0 -7260 0 1 -18312
box 62 116 196 250
use ptap  ptap_177
timestamp 1626486988
transform 1 0 -8278 0 1 -18312
box 62 116 196 250
use ptap  ptap_176
timestamp 1626486988
transform 1 0 -6242 0 1 -18312
box 62 116 196 250
use ptap  ptap_175
timestamp 1626486988
transform 1 0 -5224 0 1 -18312
box 62 116 196 250
use ptap  ptap_174
timestamp 1626486988
transform 1 0 -4206 0 1 -18312
box 62 116 196 250
use ptap  ptap_173
timestamp 1626486988
transform 1 0 -3188 0 1 -18312
box 62 116 196 250
use ptap  ptap_172
timestamp 1626486988
transform 1 0 -2170 0 1 -18312
box 62 116 196 250
use ptap  ptap_171
timestamp 1626486988
transform 1 0 -1152 0 1 -18312
box 62 116 196 250
use ptap  ptap_170
timestamp 1626486988
transform 1 0 -124 0 1 -18312
box 62 116 196 250
use ptap  ptap_169
timestamp 1626486988
transform 1 0 4004 0 1 -17776
box 62 116 196 250
use ptap  ptap_168
timestamp 1626486988
transform 1 0 2986 0 1 -17776
box 62 116 196 250
use ptap  ptap_167
timestamp 1626486988
transform 1 0 6040 0 1 -17776
box 62 116 196 250
use ptap  ptap_166
timestamp 1626486988
transform 1 0 5022 0 1 -17776
box 62 116 196 250
use ptap  ptap_165
timestamp 1626486988
transform 1 0 7058 0 1 -17776
box 62 116 196 250
use ptap  ptap_164
timestamp 1626486988
transform 1 0 8076 0 1 -17776
box 62 116 196 250
use ptap  ptap_163
timestamp 1626486988
transform 1 0 9094 0 1 -17776
box 62 116 196 250
use ptap  ptap_162
timestamp 1626486988
transform 1 0 11130 0 1 -17776
box 62 116 196 250
use ptap  ptap_161
timestamp 1626486988
transform 1 0 10112 0 1 -17776
box 62 116 196 250
use ptap  ptap_160
timestamp 1626486988
transform 1 0 12148 0 1 -17776
box 62 116 196 250
use ptap  ptap_159
timestamp 1626486988
transform 1 0 13166 0 1 -17776
box 62 116 196 250
use ptap  ptap_158
timestamp 1626486988
transform 1 0 14184 0 1 -17776
box 62 116 196 250
use ptap  ptap_157
timestamp 1626486988
transform 1 0 15202 0 1 -17776
box 62 116 196 250
use ptap  ptap_155
timestamp 1626486988
transform 1 0 16220 0 1 -17776
box 62 116 196 250
use ptap  ptap_156
timestamp 1626486988
transform 1 0 17238 0 1 -17776
box 62 116 196 250
use ptap  ptap_154
timestamp 1626486988
transform 1 0 18256 0 1 -17776
box 62 116 196 250
use ptap  ptap_153
timestamp 1626486988
transform 1 0 19274 0 1 -17776
box 62 116 196 250
use ptap  ptap_152
timestamp 1626486988
transform 1 0 20292 0 1 -17776
box 62 116 196 250
use ptap  ptap_151
timestamp 1626486988
transform 1 0 22328 0 1 -17776
box 62 116 196 250
use ptap  ptap_150
timestamp 1626486988
transform 1 0 21310 0 1 -17776
box 62 116 196 250
use ptap  ptap_147
timestamp 1626486988
transform 1 0 -9296 0 1 -17494
box 62 116 196 250
use ptap  ptap_148
timestamp 1626486988
transform 1 0 -7260 0 1 -17494
box 62 116 196 250
use ptap  ptap_149
timestamp 1626486988
transform 1 0 -8278 0 1 -17494
box 62 116 196 250
use ptap  ptap_144
timestamp 1626486988
transform 1 0 -5224 0 1 -17494
box 62 116 196 250
use ptap  ptap_145
timestamp 1626486988
transform 1 0 -6242 0 1 -17494
box 62 116 196 250
use ptap  ptap_146
timestamp 1626486988
transform 1 0 -4206 0 1 -17494
box 62 116 196 250
use ptap  ptap_141
timestamp 1626486988
transform 1 0 -2170 0 1 -17494
box 62 116 196 250
use ptap  ptap_142
timestamp 1626486988
transform 1 0 -3188 0 1 -17494
box 62 116 196 250
use ptap  ptap_143
timestamp 1626486988
transform 1 0 -1152 0 1 -17494
box 62 116 196 250
use ptap  ptap_140
timestamp 1626486988
transform 1 0 -124 0 1 -17494
box 62 116 196 250
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_2
timestamp 1626486988
transform 1 0 12777 0 1 -16998
box -10235 -388 10235 388
use sky130_fd_pr__nfet_01v8_lvt_XH9Q8F  sky130_fd_pr__nfet_01v8_lvt_XH9Q8F_1
timestamp 1626486988
transform 1 0 -4586 0 1 -17311
box -4636 -1615 4636 1615
use ptap  ptap_139
timestamp 1626486988
transform 1 0 -9296 0 1 -16676
box 62 116 196 250
use ptap  ptap_137
timestamp 1626486988
transform 1 0 -7260 0 1 -16676
box 62 116 196 250
use ptap  ptap_138
timestamp 1626486988
transform 1 0 -8278 0 1 -16676
box 62 116 196 250
use ptap  ptap_136
timestamp 1626486988
transform 1 0 -6242 0 1 -16676
box 62 116 196 250
use ptap  ptap_135
timestamp 1626486988
transform 1 0 -5224 0 1 -16676
box 62 116 196 250
use ptap  ptap_134
timestamp 1626486988
transform 1 0 -4206 0 1 -16676
box 62 116 196 250
use ptap  ptap_133
timestamp 1626486988
transform 1 0 -3188 0 1 -16676
box 62 116 196 250
use ptap  ptap_132
timestamp 1626486988
transform 1 0 -2170 0 1 -16676
box 62 116 196 250
use ptap  ptap_131
timestamp 1626486988
transform 1 0 -1152 0 1 -16676
box 62 116 196 250
use ptap  ptap_130
timestamp 1626486988
transform 1 0 -124 0 1 -16676
box 62 116 196 250
use ptap  ptap_129
timestamp 1626486988
transform 1 0 2986 0 1 -16552
box 62 116 196 250
use ptap  ptap_127
timestamp 1626486988
transform 1 0 4004 0 1 -16552
box 62 116 196 250
use ptap  ptap_128
timestamp 1626486988
transform 1 0 5022 0 1 -16552
box 62 116 196 250
use ptap  ptap_126
timestamp 1626486988
transform 1 0 6040 0 1 -16552
box 62 116 196 250
use ptap  ptap_125
timestamp 1626486988
transform 1 0 7058 0 1 -16552
box 62 116 196 250
use ptap  ptap_124
timestamp 1626486988
transform 1 0 8076 0 1 -16552
box 62 116 196 250
use ptap  ptap_123
timestamp 1626486988
transform 1 0 9094 0 1 -16552
box 62 116 196 250
use ptap  ptap_122
timestamp 1626486988
transform 1 0 10112 0 1 -16552
box 62 116 196 250
use ptap  ptap_121
timestamp 1626486988
transform 1 0 11130 0 1 -16552
box 62 116 196 250
use ptap  ptap_120
timestamp 1626486988
transform 1 0 12148 0 1 -16552
box 62 116 196 250
use ptap  ptap_119
timestamp 1626486988
transform 1 0 13166 0 1 -16552
box 62 116 196 250
use ptap  ptap_118
timestamp 1626486988
transform 1 0 14184 0 1 -16552
box 62 116 196 250
use ptap  ptap_116
timestamp 1626486988
transform 1 0 16220 0 1 -16552
box 62 116 196 250
use ptap  ptap_117
timestamp 1626486988
transform 1 0 15202 0 1 -16552
box 62 116 196 250
use ptap  ptap_115
timestamp 1626486988
transform 1 0 17238 0 1 -16552
box 62 116 196 250
use ptap  ptap_114
timestamp 1626486988
transform 1 0 18256 0 1 -16552
box 62 116 196 250
use ptap  ptap_113
timestamp 1626486988
transform 1 0 19274 0 1 -16552
box 62 116 196 250
use ptap  ptap_112
timestamp 1626486988
transform 1 0 20292 0 1 -16552
box 62 116 196 250
use ptap  ptap_111
timestamp 1626486988
transform 1 0 21310 0 1 -16552
box 62 116 196 250
use ptap  ptap_110
timestamp 1626486988
transform 1 0 22328 0 1 -16552
box 62 116 196 250
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_1
timestamp 1626486988
transform 1 0 12779 0 1 -15764
box -10235 -388 10235 388
use ptap  ptap_109
timestamp 1626486988
transform 1 0 -9296 0 1 -15858
box 62 116 196 250
use ptap  ptap_108
timestamp 1626486988
transform 1 0 -7260 0 1 -15858
box 62 116 196 250
use ptap  ptap_107
timestamp 1626486988
transform 1 0 -8278 0 1 -15858
box 62 116 196 250
use ptap  ptap_106
timestamp 1626486988
transform 1 0 -6242 0 1 -15858
box 62 116 196 250
use ptap  ptap_105
timestamp 1626486988
transform 1 0 -5224 0 1 -15858
box 62 116 196 250
use ptap  ptap_104
timestamp 1626486988
transform 1 0 -4206 0 1 -15858
box 62 116 196 250
use ptap  ptap_103
timestamp 1626486988
transform 1 0 -3188 0 1 -15858
box 62 116 196 250
use ptap  ptap_102
timestamp 1626486988
transform 1 0 -2170 0 1 -15858
box 62 116 196 250
use ptap  ptap_101
timestamp 1626486988
transform 1 0 -1152 0 1 -15858
box 62 116 196 250
use ptap  ptap_100
timestamp 1626486988
transform 1 0 -124 0 1 -15858
box 62 116 196 250
use ptap  ptap_99
timestamp 1626486988
transform 1 0 2998 0 1 -15316
box 62 116 196 250
use ptap  ptap_98
timestamp 1626486988
transform 1 0 4016 0 1 -15316
box 62 116 196 250
use ptap  ptap_97
timestamp 1626486988
transform 1 0 5034 0 1 -15316
box 62 116 196 250
use ptap  ptap_96
timestamp 1626486988
transform 1 0 6052 0 1 -15316
box 62 116 196 250
use ptap  ptap_95
timestamp 1626486988
transform 1 0 7070 0 1 -15316
box 62 116 196 250
use ptap  ptap_94
timestamp 1626486988
transform 1 0 8088 0 1 -15316
box 62 116 196 250
use ptap  ptap_93
timestamp 1626486988
transform 1 0 9106 0 1 -15316
box 62 116 196 250
use ptap  ptap_92
timestamp 1626486988
transform 1 0 10124 0 1 -15316
box 62 116 196 250
use ptap  ptap_91
timestamp 1626486988
transform 1 0 11142 0 1 -15316
box 62 116 196 250
use ptap  ptap_90
timestamp 1626486988
transform 1 0 12160 0 1 -15316
box 62 116 196 250
use ptap  ptap_89
timestamp 1626486988
transform 1 0 13178 0 1 -15316
box 62 116 196 250
use ptap  ptap_88
timestamp 1626486988
transform 1 0 14196 0 1 -15316
box 62 116 196 250
use ptap  ptap_87
timestamp 1626486988
transform 1 0 15214 0 1 -15316
box 62 116 196 250
use ptap  ptap_86
timestamp 1626486988
transform 1 0 16232 0 1 -15316
box 62 116 196 250
use ptap  ptap_85
timestamp 1626486988
transform 1 0 17250 0 1 -15316
box 62 116 196 250
use ptap  ptap_84
timestamp 1626486988
transform 1 0 18268 0 1 -15316
box 62 116 196 250
use ptap  ptap_83
timestamp 1626486988
transform 1 0 19286 0 1 -15316
box 62 116 196 250
use ptap  ptap_82
timestamp 1626486988
transform 1 0 20304 0 1 -15316
box 62 116 196 250
use ptap  ptap_81
timestamp 1626486988
transform 1 0 21322 0 1 -15316
box 62 116 196 250
use ptap  ptap_80
timestamp 1626486988
transform 1 0 22340 0 1 -15316
box 62 116 196 250
use ptap  ptap_77
timestamp 1626486988
transform 1 0 -9296 0 1 -15040
box 62 116 196 250
use ptap  ptap_78
timestamp 1626486988
transform 1 0 -8278 0 1 -15040
box 62 116 196 250
use ptap  ptap_79
timestamp 1626486988
transform 1 0 -7260 0 1 -15040
box 62 116 196 250
use ptap  ptap_74
timestamp 1626486988
transform 1 0 -5224 0 1 -15040
box 62 116 196 250
use ptap  ptap_75
timestamp 1626486988
transform 1 0 -6242 0 1 -15040
box 62 116 196 250
use ptap  ptap_76
timestamp 1626486988
transform 1 0 -4206 0 1 -15040
box 62 116 196 250
use ptap  ptap_71
timestamp 1626486988
transform 1 0 -2170 0 1 -15040
box 62 116 196 250
use ptap  ptap_72
timestamp 1626486988
transform 1 0 -3188 0 1 -15040
box 62 116 196 250
use ptap  ptap_73
timestamp 1626486988
transform 1 0 -1152 0 1 -15040
box 62 116 196 250
use ptap  ptap_70
timestamp 1626486988
transform 1 0 -124 0 1 -15040
box 62 116 196 250
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_0
timestamp 1626486988
transform 1 0 12779 0 1 -14532
box -10235 -388 10235 388
use ptap  ptap_69
timestamp 1626486988
transform 1 0 -9296 0 1 -14222
box 62 116 196 250
use ptap  ptap_68
timestamp 1626486988
transform 1 0 -8278 0 1 -14222
box 62 116 196 250
use ptap  ptap_67
timestamp 1626486988
transform 1 0 -7260 0 1 -14222
box 62 116 196 250
use ptap  ptap_66
timestamp 1626486988
transform 1 0 -6242 0 1 -14222
box 62 116 196 250
use ptap  ptap_65
timestamp 1626486988
transform 1 0 -5224 0 1 -14222
box 62 116 196 250
use ptap  ptap_64
timestamp 1626486988
transform 1 0 -4206 0 1 -14222
box 62 116 196 250
use ptap  ptap_63
timestamp 1626486988
transform 1 0 -3188 0 1 -14222
box 62 116 196 250
use ptap  ptap_62
timestamp 1626486988
transform 1 0 -2170 0 1 -14222
box 62 116 196 250
use ptap  ptap_61
timestamp 1626486988
transform 1 0 -1152 0 1 -14222
box 62 116 196 250
use ptap  ptap_60
timestamp 1626486988
transform 1 0 -124 0 1 -14222
box 62 116 196 250
use ptap  ptap_59
timestamp 1626486988
transform 1 0 3010 0 1 -14010
box 62 116 196 250
use ptap  ptap_58
timestamp 1626486988
transform 1 0 4028 0 1 -14010
box 62 116 196 250
use ptap  ptap_57
timestamp 1626486988
transform 1 0 5046 0 1 -14010
box 62 116 196 250
use ptap  ptap_56
timestamp 1626486988
transform 1 0 6064 0 1 -14010
box 62 116 196 250
use ptap  ptap_55
timestamp 1626486988
transform 1 0 7082 0 1 -14010
box 62 116 196 250
use ptap  ptap_54
timestamp 1626486988
transform 1 0 8100 0 1 -14010
box 62 116 196 250
use ptap  ptap_53
timestamp 1626486988
transform 1 0 9118 0 1 -14010
box 62 116 196 250
use ptap  ptap_52
timestamp 1626486988
transform 1 0 10136 0 1 -14010
box 62 116 196 250
use ptap  ptap_51
timestamp 1626486988
transform 1 0 11154 0 1 -14010
box 62 116 196 250
use ptap  ptap_50
timestamp 1626486988
transform 1 0 12172 0 1 -14010
box 62 116 196 250
use ptap  ptap_49
timestamp 1626486988
transform 1 0 13190 0 1 -14010
box 62 116 196 250
use ptap  ptap_48
timestamp 1626486988
transform 1 0 14208 0 1 -14010
box 62 116 196 250
use ptap  ptap_47
timestamp 1626486988
transform 1 0 15226 0 1 -14010
box 62 116 196 250
use ptap  ptap_46
timestamp 1626486988
transform 1 0 16244 0 1 -14010
box 62 116 196 250
use ptap  ptap_45
timestamp 1626486988
transform 1 0 17262 0 1 -14010
box 62 116 196 250
use ptap  ptap_44
timestamp 1626486988
transform 1 0 18280 0 1 -14010
box 62 116 196 250
use ptap  ptap_43
timestamp 1626486988
transform 1 0 19298 0 1 -14010
box 62 116 196 250
use ptap  ptap_42
timestamp 1626486988
transform 1 0 20316 0 1 -14010
box 62 116 196 250
use ptap  ptap_41
timestamp 1626486988
transform 1 0 21334 0 1 -14010
box 62 116 196 250
use ptap  ptap_40
timestamp 1626486988
transform 1 0 22352 0 1 -14010
box 62 116 196 250
use sky130_fd_pr__nfet_01v8_J5YDRX  sky130_fd_pr__nfet_01v8_J5YDRX_0
timestamp 1626486988
transform -1 0 12779 0 -1 -12745
box -10235 -797 10235 797
use sky130_fd_pr__nfet_01v8_lvt_XH9Q8F  sky130_fd_pr__nfet_01v8_lvt_XH9Q8F_0
timestamp 1626486988
transform 1 0 -4586 0 1 -14039
box -4636 -1615 4636 1615
use ptap  ptap_39
timestamp 1626486988
transform 1 0 -9296 0 1 -12586
box 62 116 196 250
use ptap  ptap_38
timestamp 1626486988
transform 1 0 -9296 0 1 -13404
box 62 116 196 250
use ptap  ptap_37
timestamp 1626486988
transform 1 0 -8278 0 1 -13404
box 62 116 196 250
use ptap  ptap_36
timestamp 1626486988
transform 1 0 -8278 0 1 -12586
box 62 116 196 250
use ptap  ptap_35
timestamp 1626486988
transform 1 0 -7260 0 1 -13404
box 62 116 196 250
use ptap  ptap_34
timestamp 1626486988
transform 1 0 -7260 0 1 -12586
box 62 116 196 250
use ptap  ptap_33
timestamp 1626486988
transform 1 0 -6242 0 1 -13404
box 62 116 196 250
use ptap  ptap_32
timestamp 1626486988
transform 1 0 -6242 0 1 -12586
box 62 116 196 250
use ptap  ptap_31
timestamp 1626486988
transform 1 0 -5224 0 1 -13404
box 62 116 196 250
use ptap  ptap_30
timestamp 1626486988
transform 1 0 -5224 0 1 -12586
box 62 116 196 250
use ptap  ptap_29
timestamp 1626486988
transform 1 0 -4206 0 1 -13404
box 62 116 196 250
use ptap  ptap_28
timestamp 1626486988
transform 1 0 -4206 0 1 -12586
box 62 116 196 250
use ptap  ptap_27
timestamp 1626486988
transform 1 0 -3188 0 1 -13404
box 62 116 196 250
use ptap  ptap_26
timestamp 1626486988
transform 1 0 -3188 0 1 -12586
box 62 116 196 250
use ptap  ptap_25
timestamp 1626486988
transform 1 0 -2170 0 1 -13404
box 62 116 196 250
use ptap  ptap_24
timestamp 1626486988
transform 1 0 -2170 0 1 -12586
box 62 116 196 250
use ptap  ptap_23
timestamp 1626486988
transform 1 0 -1152 0 1 -13404
box 62 116 196 250
use ptap  ptap_22
timestamp 1626486988
transform 1 0 -1152 0 1 -12586
box 62 116 196 250
use ptap  ptap_21
timestamp 1626486988
transform 1 0 -124 0 1 -13404
box 62 116 196 250
use ptap  ptap_20
timestamp 1626486988
transform 1 0 -124 0 1 -12586
box 62 116 196 250
use ptap  ptap_19
timestamp 1626486988
transform 1 0 2998 0 1 -11984
box 62 116 196 250
use ptap  ptap_18
timestamp 1626486988
transform 1 0 4016 0 1 -11984
box 62 116 196 250
use ptap  ptap_17
timestamp 1626486988
transform 1 0 5034 0 1 -11984
box 62 116 196 250
use ptap  ptap_16
timestamp 1626486988
transform 1 0 6052 0 1 -11984
box 62 116 196 250
use ptap  ptap_15
timestamp 1626486988
transform 1 0 7070 0 1 -11984
box 62 116 196 250
use ptap  ptap_14
timestamp 1626486988
transform 1 0 8088 0 1 -11984
box 62 116 196 250
use ptap  ptap_13
timestamp 1626486988
transform 1 0 9106 0 1 -11984
box 62 116 196 250
use ptap  ptap_12
timestamp 1626486988
transform 1 0 10124 0 1 -11984
box 62 116 196 250
use ptap  ptap_11
timestamp 1626486988
transform 1 0 11142 0 1 -11984
box 62 116 196 250
use ptap  ptap_10
timestamp 1626486988
transform 1 0 12160 0 1 -11984
box 62 116 196 250
use ptap  ptap_9
timestamp 1626486988
transform 1 0 13178 0 1 -11984
box 62 116 196 250
use ptap  ptap_8
timestamp 1626486988
transform 1 0 14196 0 1 -11984
box 62 116 196 250
use ptap  ptap_7
timestamp 1626486988
transform 1 0 15214 0 1 -11984
box 62 116 196 250
use ptap  ptap_6
timestamp 1626486988
transform 1 0 16232 0 1 -11984
box 62 116 196 250
use ptap  ptap_5
timestamp 1626486988
transform 1 0 17250 0 1 -11984
box 62 116 196 250
use ptap  ptap_4
timestamp 1626486988
transform 1 0 18268 0 1 -11984
box 62 116 196 250
use ptap  ptap_3
timestamp 1626486988
transform 1 0 19286 0 1 -11984
box 62 116 196 250
use ptap  ptap_2
timestamp 1626486988
transform 1 0 20304 0 1 -11984
box 62 116 196 250
use ptap  ptap_1
timestamp 1626486988
transform 1 0 21322 0 1 -11984
box 62 116 196 250
use ptap  ptap_0
timestamp 1626486988
transform 1 0 22340 0 1 -11984
box 62 116 196 250
use ntap  ntap_162
timestamp 1626486988
transform 1 0 4384 0 1 -9532
box 250 218 480 436
use ntap  ntap_161
timestamp 1626486988
transform 1 0 3366 0 1 -9532
box 250 218 480 436
use ntap  ntap_160
timestamp 1626486988
transform 1 0 2348 0 1 -9532
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_MSJKJ2  sky130_fd_pr__pfet_01v8_MSJKJ2_3
timestamp 1626486988
transform 1 0 15126 0 1 -9140
box -7700 -400 7700 400
use ntap  ntap_159
timestamp 1626486988
transform 1 0 5402 0 1 -9532
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_lvt_DHLX6D  sky130_fd_pr__pfet_01v8_lvt_DHLX6D_3
timestamp 1626486988
transform 1 0 4223 0 1 -8572
box -2101 -400 2101 400
use ntap  ntap_158
timestamp 1626486988
transform 1 0 6924 0 1 -8820
box 250 218 480 436
use ntap  ntap_157
timestamp 1626486988
transform 1 0 7942 0 1 -8820
box 250 218 480 436
use ntap  ntap_156
timestamp 1626486988
transform 1 0 8960 0 1 -8820
box 250 218 480 436
use ntap  ntap_155
timestamp 1626486988
transform 1 0 9978 0 1 -8820
box 250 218 480 436
use ntap  ntap_154
timestamp 1626486988
transform 1 0 10996 0 1 -8820
box 250 218 480 436
use ntap  ntap_153
timestamp 1626486988
transform 1 0 12014 0 1 -8820
box 250 218 480 436
use ntap  ntap_151
timestamp 1626486988
transform 1 0 14050 0 1 -8820
box 250 218 480 436
use ntap  ntap_152
timestamp 1626486988
transform 1 0 13032 0 1 -8820
box 250 218 480 436
use ntap  ntap_150
timestamp 1626486988
transform 1 0 15068 0 1 -8820
box 250 218 480 436
use ntap  ntap_149
timestamp 1626486988
transform 1 0 16086 0 1 -8820
box 250 218 480 436
use ntap  ntap_148
timestamp 1626486988
transform 1 0 17104 0 1 -8820
box 250 218 480 436
use ntap  ntap_147
timestamp 1626486988
transform 1 0 18122 0 1 -8820
box 250 218 480 436
use ntap  ntap_146
timestamp 1626486988
transform 1 0 19140 0 1 -8820
box 250 218 480 436
use ntap  ntap_145
timestamp 1626486988
transform 1 0 22194 0 1 -8820
box 250 218 480 436
use ntap  ntap_144
timestamp 1626486988
transform 1 0 21176 0 1 -8820
box 250 218 480 436
use ntap  ntap_143
timestamp 1626486988
transform 1 0 20158 0 1 -8820
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_lvt_DHLX6D  sky130_fd_pr__pfet_01v8_lvt_DHLX6D_2
timestamp 1626486988
transform 1 0 4223 0 1 -7540
box -2101 -400 2101 400
use ntap  ntap_142
timestamp 1626486988
transform 1 0 1824 0 1 -8380
box 250 218 480 436
use ntap  ntap_141
timestamp 1626486988
transform 1 0 2842 0 1 -8380
box 250 218 480 436
use ntap  ntap_140
timestamp 1626486988
transform 1 0 3860 0 1 -8380
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_MSJKJ2  sky130_fd_pr__pfet_01v8_MSJKJ2_2
timestamp 1626486988
transform 1 0 15126 0 1 -7884
box -7700 -400 7700 400
use ntap  ntap_139
timestamp 1626486988
transform 1 0 4878 0 1 -8380
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_lvt_DHLX6D  sky130_fd_pr__pfet_01v8_lvt_DHLX6D_1
timestamp 1626486988
transform 1 0 4223 0 1 -6508
box -2101 -400 2101 400
use ntap  ntap_138
timestamp 1626486988
transform 1 0 3870 0 1 -7352
box 250 218 480 436
use ntap  ntap_137
timestamp 1626486988
transform 1 0 2852 0 1 -7352
box 250 218 480 436
use ntap  ntap_136
timestamp 1626486988
transform 1 0 1834 0 1 -7352
box 250 218 480 436
use ntap  ntap_135
timestamp 1626486988
transform 1 0 8078 0 1 -7576
box 250 218 480 436
use ntap  ntap_134
timestamp 1626486988
transform 1 0 7060 0 1 -7576
box 250 218 480 436
use ntap  ntap_133
timestamp 1626486988
transform 1 0 9096 0 1 -7576
box 250 218 480 436
use ntap  ntap_132
timestamp 1626486988
transform 1 0 10114 0 1 -7576
box 250 218 480 436
use ntap  ntap_131
timestamp 1626486988
transform 1 0 11132 0 1 -7576
box 250 218 480 436
use ntap  ntap_130
timestamp 1626486988
transform 1 0 12150 0 1 -7576
box 250 218 480 436
use ntap  ntap_129
timestamp 1626486988
transform 1 0 13168 0 1 -7576
box 250 218 480 436
use ntap  ntap_128
timestamp 1626486988
transform 1 0 15204 0 1 -7576
box 250 218 480 436
use ntap  ntap_127
timestamp 1626486988
transform 1 0 14186 0 1 -7576
box 250 218 480 436
use ntap  ntap_126
timestamp 1626486988
transform 1 0 16222 0 1 -7576
box 250 218 480 436
use ntap  ntap_125
timestamp 1626486988
transform 1 0 17240 0 1 -7576
box 250 218 480 436
use ntap  ntap_124
timestamp 1626486988
transform 1 0 18258 0 1 -7576
box 250 218 480 436
use ntap  ntap_123
timestamp 1626486988
transform 1 0 19276 0 1 -7576
box 250 218 480 436
use ntap  ntap_122
timestamp 1626486988
transform 1 0 4888 0 1 -7352
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_MSJKJ2  sky130_fd_pr__pfet_01v8_MSJKJ2_1
timestamp 1626486988
transform 1 0 15126 0 1 -6628
box -7700 -400 7700 400
use ntap  ntap_121
timestamp 1626486988
transform 1 0 22330 0 1 -7576
box 250 218 480 436
use ntap  ntap_120
timestamp 1626486988
transform 1 0 21312 0 1 -7576
box 250 218 480 436
use ntap  ntap_119
timestamp 1626486988
transform 1 0 20294 0 1 -7576
box 250 218 480 436
use ntap  ntap_118
timestamp 1626486988
transform 1 0 3860 0 1 -6324
box 250 218 480 436
use ntap  ntap_117
timestamp 1626486988
transform 1 0 1824 0 1 -6324
box 250 218 480 436
use ntap  ntap_116
timestamp 1626486988
transform 1 0 2842 0 1 -6324
box 250 218 480 436
use ntap  ntap_115
timestamp 1626486988
transform 1 0 4878 0 1 -6324
box 250 218 480 436
use ntap  ntap_114
timestamp 1626486988
transform 1 0 7036 0 1 -6308
box 250 218 480 436
use ntap  ntap_113
timestamp 1626486988
transform 1 0 8054 0 1 -6308
box 250 218 480 436
use ntap  ntap_111
timestamp 1626486988
transform 1 0 10090 0 1 -6308
box 250 218 480 436
use ntap  ntap_112
timestamp 1626486988
transform 1 0 9072 0 1 -6308
box 250 218 480 436
use ntap  ntap_110
timestamp 1626486988
transform 1 0 11108 0 1 -6308
box 250 218 480 436
use ntap  ntap_109
timestamp 1626486988
transform 1 0 12126 0 1 -6308
box 250 218 480 436
use ntap  ntap_108
timestamp 1626486988
transform 1 0 13144 0 1 -6308
box 250 218 480 436
use ntap  ntap_107
timestamp 1626486988
transform 1 0 14162 0 1 -6308
box 250 218 480 436
use ntap  ntap_106
timestamp 1626486988
transform 1 0 15180 0 1 -6308
box 250 218 480 436
use ntap  ntap_105
timestamp 1626486988
transform 1 0 16198 0 1 -6308
box 250 218 480 436
use ntap  ntap_104
timestamp 1626486988
transform 1 0 17216 0 1 -6308
box 250 218 480 436
use ntap  ntap_103
timestamp 1626486988
transform 1 0 18234 0 1 -6308
box 250 218 480 436
use ntap  ntap_102
timestamp 1626486988
transform 1 0 19252 0 1 -6308
box 250 218 480 436
use ntap  ntap_101
timestamp 1626486988
transform 1 0 21288 0 1 -6308
box 250 218 480 436
use ntap  ntap_100
timestamp 1626486988
transform 1 0 22306 0 1 -6308
box 250 218 480 436
use ntap  ntap_99
timestamp 1626486988
transform 1 0 20270 0 1 -6308
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_lvt_DHLX6D  sky130_fd_pr__pfet_01v8_lvt_DHLX6D_0
timestamp 1626486988
transform 1 0 4223 0 1 -5476
box -2101 -400 2101 400
use sky130_fd_pr__pfet_01v8_MSJKJ2  sky130_fd_pr__pfet_01v8_MSJKJ2_0
timestamp 1626486988
transform 1 0 15126 0 1 -5372
box -7700 -400 7700 400
use ntap  ntap_98
timestamp 1626486988
transform 1 0 4384 0 1 -5170
box 250 218 480 436
use ntap  ntap_97
timestamp 1626486988
transform 1 0 3366 0 1 -5170
box 250 218 480 436
use ntap  ntap_96
timestamp 1626486988
transform 1 0 2348 0 1 -5170
box 250 218 480 436
use ntap  ntap_95
timestamp 1626486988
transform 1 0 5402 0 1 -5170
box 250 218 480 436
use ntap  ntap_94
timestamp 1626486988
transform 1 0 6946 0 1 -4860
box 250 218 480 436
use ntap  ntap_92
timestamp 1626486988
transform 1 0 7964 0 1 -4860
box 250 218 480 436
use ntap  ntap_93
timestamp 1626486988
transform 1 0 8982 0 1 -4860
box 250 218 480 436
use ntap  ntap_91
timestamp 1626486988
transform 1 0 10000 0 1 -4860
box 250 218 480 436
use ntap  ntap_90
timestamp 1626486988
transform 1 0 11018 0 1 -4860
box 250 218 480 436
use ntap  ntap_89
timestamp 1626486988
transform 1 0 12036 0 1 -4860
box 250 218 480 436
use ntap  ntap_88
timestamp 1626486988
transform 1 0 13054 0 1 -4860
box 250 218 480 436
use ntap  ntap_87
timestamp 1626486988
transform 1 0 14072 0 1 -4860
box 250 218 480 436
use ntap  ntap_86
timestamp 1626486988
transform 1 0 15090 0 1 -4860
box 250 218 480 436
use ntap  ntap_85
timestamp 1626486988
transform 1 0 16108 0 1 -4860
box 250 218 480 436
use ntap  ntap_84
timestamp 1626486988
transform 1 0 17126 0 1 -4860
box 250 218 480 436
use ntap  ntap_83
timestamp 1626486988
transform 1 0 18144 0 1 -4860
box 250 218 480 436
use ntap  ntap_82
timestamp 1626486988
transform 1 0 19162 0 1 -4860
box 250 218 480 436
use ntap  ntap_81
timestamp 1626486988
transform 1 0 22216 0 1 -4860
box 250 218 480 436
use ntap  ntap_80
timestamp 1626486988
transform 1 0 21198 0 1 -4860
box 250 218 480 436
use ntap  ntap_79
timestamp 1626486988
transform 1 0 20180 0 1 -4860
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_lvt_SH2KEA  sky130_fd_pr__pfet_01v8_lvt_SH2KEA_1
timestamp 1626486988
transform 1 0 14825 0 1 -3768
box -7191 -400 7191 400
use ntap  ntap_78
timestamp 1626486988
transform 1 0 7340 0 1 -3582
box 250 218 480 436
use ntap  ntap_77
timestamp 1626486988
transform 1 0 8358 0 1 -3582
box 250 218 480 436
use ntap  ntap_76
timestamp 1626486988
transform 1 0 9376 0 1 -3582
box 250 218 480 436
use ntap  ntap_75
timestamp 1626486988
transform 1 0 10394 0 1 -3582
box 250 218 480 436
use ntap  ntap_74
timestamp 1626486988
transform 1 0 11412 0 1 -3582
box 250 218 480 436
use ntap  ntap_73
timestamp 1626486988
transform 1 0 12430 0 1 -3582
box 250 218 480 436
use ntap  ntap_72
timestamp 1626486988
transform 1 0 13448 0 1 -3582
box 250 218 480 436
use ntap  ntap_70
timestamp 1626486988
transform 1 0 14466 0 1 -3582
box 250 218 480 436
use ntap  ntap_71
timestamp 1626486988
transform 1 0 15484 0 1 -3582
box 250 218 480 436
use ntap  ntap_69
timestamp 1626486988
transform 1 0 16502 0 1 -3582
box 250 218 480 436
use ntap  ntap_68
timestamp 1626486988
transform 1 0 17520 0 1 -3582
box 250 218 480 436
use ntap  ntap_67
timestamp 1626486988
transform 1 0 18538 0 1 -3582
box 250 218 480 436
use ntap  ntap_66
timestamp 1626486988
transform 1 0 19556 0 1 -3582
box 250 218 480 436
use ntap  ntap_65
timestamp 1626486988
transform 1 0 20574 0 1 -3582
box 250 218 480 436
use ntap  ntap_64
timestamp 1626486988
transform 1 0 21592 0 1 -3582
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_lvt_SH2KEA  sky130_fd_pr__pfet_01v8_lvt_SH2KEA_0
timestamp 1626486988
transform 1 0 14825 0 1 -2736
box -7191 -400 7191 400
use ntap  ntap_63
timestamp 1626486988
transform 1 0 6652 0 1 -2234
box 250 218 480 436
use ntap  ntap_62
timestamp 1626486988
transform 1 0 7670 0 1 -2234
box 250 218 480 436
use ntap  ntap_61
timestamp 1626486988
transform 1 0 8688 0 1 -2234
box 250 218 480 436
use ntap  ntap_60
timestamp 1626486988
transform 1 0 9706 0 1 -2234
box 250 218 480 436
use ntap  ntap_59
timestamp 1626486988
transform 1 0 10724 0 1 -2234
box 250 218 480 436
use ntap  ntap_58
timestamp 1626486988
transform 1 0 11742 0 1 -2234
box 250 218 480 436
use ntap  ntap_57
timestamp 1626486988
transform 1 0 12760 0 1 -2234
box 250 218 480 436
use ntap  ntap_56
timestamp 1626486988
transform 1 0 13778 0 1 -2234
box 250 218 480 436
use ntap  ntap_55
timestamp 1626486988
transform 1 0 14796 0 1 -2234
box 250 218 480 436
use ntap  ntap_54
timestamp 1626486988
transform 1 0 15814 0 1 -2234
box 250 218 480 436
use ntap  ntap_53
timestamp 1626486988
transform 1 0 16832 0 1 -2234
box 250 218 480 436
use ntap  ntap_52
timestamp 1626486988
transform 1 0 17850 0 1 -2234
box 250 218 480 436
use ntap  ntap_51
timestamp 1626486988
transform 1 0 18868 0 1 -2234
box 250 218 480 436
use ntap  ntap_50
timestamp 1626486988
transform 1 0 19886 0 1 -2234
box 250 218 480 436
use ntap  ntap_49
timestamp 1626486988
transform 1 0 20904 0 1 -2234
box 250 218 480 436
use ntap  ntap_48
timestamp 1626486988
transform 1 0 21922 0 1 -2234
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_lvt_V2JKJ2  sky130_fd_pr__pfet_01v8_lvt_V2JKJ2_2
timestamp 1626486988
transform 1 0 14649 0 1 -1098
box -8209 -400 8209 400
use ntap  ntap_46
timestamp 1626486988
transform 1 0 7670 0 1 -852
box 250 218 480 436
use ntap  ntap_47
timestamp 1626486988
transform 1 0 6652 0 1 -852
box 250 218 480 436
use ntap  ntap_45
timestamp 1626486988
transform 1 0 8688 0 1 -852
box 250 218 480 436
use ntap  ntap_44
timestamp 1626486988
transform 1 0 9706 0 1 -852
box 250 218 480 436
use ntap  ntap_43
timestamp 1626486988
transform 1 0 10724 0 1 -852
box 250 218 480 436
use ntap  ntap_42
timestamp 1626486988
transform 1 0 11742 0 1 -852
box 250 218 480 436
use ntap  ntap_41
timestamp 1626486988
transform 1 0 12760 0 1 -852
box 250 218 480 436
use ntap  ntap_40
timestamp 1626486988
transform 1 0 13778 0 1 -852
box 250 218 480 436
use ntap  ntap_39
timestamp 1626486988
transform 1 0 14796 0 1 -852
box 250 218 480 436
use ntap  ntap_38
timestamp 1626486988
transform 1 0 15814 0 1 -852
box 250 218 480 436
use ntap  ntap_37
timestamp 1626486988
transform 1 0 16832 0 1 -852
box 250 218 480 436
use ntap  ntap_36
timestamp 1626486988
transform 1 0 17850 0 1 -852
box 250 218 480 436
use ntap  ntap_35
timestamp 1626486988
transform 1 0 18868 0 1 -852
box 250 218 480 436
use ntap  ntap_34
timestamp 1626486988
transform 1 0 19886 0 1 -852
box 250 218 480 436
use ntap  ntap_33
timestamp 1626486988
transform 1 0 20904 0 1 -852
box 250 218 480 436
use ntap  ntap_32
timestamp 1626486988
transform 1 0 21922 0 1 -852
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_lvt_V2JKJ2  sky130_fd_pr__pfet_01v8_lvt_V2JKJ2_1
timestamp 1626486988
transform 1 0 14649 0 1 38
box -8209 -400 8209 400
use ntap  ntap_31
timestamp 1626486988
transform 1 0 6674 0 1 280
box 250 218 480 436
use ntap  ntap_30
timestamp 1626486988
transform 1 0 7692 0 1 280
box 250 218 480 436
use ntap  ntap_29
timestamp 1626486988
transform 1 0 8710 0 1 280
box 250 218 480 436
use ntap  ntap_28
timestamp 1626486988
transform 1 0 9728 0 1 280
box 250 218 480 436
use ntap  ntap_27
timestamp 1626486988
transform 1 0 10746 0 1 280
box 250 218 480 436
use ntap  ntap_26
timestamp 1626486988
transform 1 0 11764 0 1 280
box 250 218 480 436
use ntap  ntap_25
timestamp 1626486988
transform 1 0 12782 0 1 280
box 250 218 480 436
use ntap  ntap_24
timestamp 1626486988
transform 1 0 13800 0 1 280
box 250 218 480 436
use ntap  ntap_23
timestamp 1626486988
transform 1 0 14818 0 1 280
box 250 218 480 436
use ntap  ntap_22
timestamp 1626486988
transform 1 0 15836 0 1 280
box 250 218 480 436
use ntap  ntap_21
timestamp 1626486988
transform 1 0 16854 0 1 280
box 250 218 480 436
use ntap  ntap_20
timestamp 1626486988
transform 1 0 17872 0 1 280
box 250 218 480 436
use ntap  ntap_19
timestamp 1626486988
transform 1 0 18890 0 1 280
box 250 218 480 436
use ntap  ntap_18
timestamp 1626486988
transform 1 0 19908 0 1 280
box 250 218 480 436
use ntap  ntap_17
timestamp 1626486988
transform 1 0 20926 0 1 280
box 250 218 480 436
use ntap  ntap_16
timestamp 1626486988
transform 1 0 21944 0 1 280
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_lvt_V2JKJ2  sky130_fd_pr__pfet_01v8_lvt_V2JKJ2_0
timestamp 1626486988
transform 1 0 14649 0 1 1174
box -8209 -400 8209 400
use ntap  ntap_14
timestamp 1626486988
transform 1 0 7670 0 1 1434
box 250 218 480 436
use ntap  ntap_15
timestamp 1626486988
transform 1 0 6652 0 1 1434
box 250 218 480 436
use ntap  ntap_13
timestamp 1626486988
transform 1 0 8688 0 1 1434
box 250 218 480 436
use ntap  ntap_12
timestamp 1626486988
transform 1 0 9706 0 1 1434
box 250 218 480 436
use ntap  ntap_11
timestamp 1626486988
transform 1 0 10724 0 1 1434
box 250 218 480 436
use ntap  ntap_10
timestamp 1626486988
transform 1 0 11742 0 1 1434
box 250 218 480 436
use ntap  ntap_9
timestamp 1626486988
transform 1 0 12760 0 1 1434
box 250 218 480 436
use ntap  ntap_8
timestamp 1626486988
transform 1 0 13778 0 1 1434
box 250 218 480 436
use ntap  ntap_7
timestamp 1626486988
transform 1 0 14796 0 1 1434
box 250 218 480 436
use ntap  ntap_6
timestamp 1626486988
transform 1 0 15814 0 1 1434
box 250 218 480 436
use ntap  ntap_5
timestamp 1626486988
transform 1 0 16832 0 1 1434
box 250 218 480 436
use ntap  ntap_4
timestamp 1626486988
transform 1 0 17850 0 1 1434
box 250 218 480 436
use ntap  ntap_3
timestamp 1626486988
transform 1 0 18868 0 1 1434
box 250 218 480 436
use ntap  ntap_2
timestamp 1626486988
transform 1 0 19886 0 1 1434
box 250 218 480 436
use ntap  ntap_1
timestamp 1626486988
transform 1 0 20904 0 1 1434
box 250 218 480 436
use ntap  ntap_0
timestamp 1626486988
transform 1 0 21922 0 1 1434
box 250 218 480 436
<< labels >>
flabel metal1 s -8078 -12352 -8078 -12352 1 FreeSans 600 0 0 0 vbias1
flabel metal1 s -6206 -19026 -6206 -19026 1 FreeSans 600 0 0 0 vbias2
flabel metal1 s 23180 -19318 23204 -19288 1 FreeSans 600 0 0 0 VSS
flabel metal1 s 23556 -18470 23556 -18470 1 FreeSans 600 0 0 0 vbias3
flabel metal1 s 23300 -18264 23300 -18264 1 FreeSans 600 0 0 0 vcascnm
flabel metal1 s 23436 -22496 23436 -22496 1 FreeSans 600 0 0 0 vbias4
flabel metal1 s 2138 -18102 2166 -18072 1 FreeSans 600 0 0 0 vtail_cascn
flabel metal1 s 2456 -14760 2488 -14720 1 FreeSans 600 0 0 0 vcascnp
flabel metal1 s 3322 -11898 3412 -11868 1 FreeSans 600 0 0 0 M8d
flabel metal1 s 2244 -18362 2282 -18326 1 FreeSans 600 0 0 0 vmirror
flabel metal1 s 22938 -16630 22974 -16600 1 FreeSans 600 0 0 0 M16d
flabel metal1 s -10646 -21540 -10618 -21496 1 FreeSans 600 0 0 0 vip
flabel metal1 s 954 -21536 986 -21498 1 FreeSans 600 0 0 0 vim
flabel metal1 s -5202 -24966 -5106 -24930 1 FreeSans 600 0 0 0 ibiasn
flabel metal1 s -52 -22240 -4 -22216 1 FreeSans 600 0 0 0 vtail_cascn
flabel metal4 s -10920 -26744 -10894 -26722 1 FreeSans 4000 0 0 0 VSS
flabel metal2 s -6564 -19934 -6516 -19918 1 FreeSans 600 0 0 0 vcascpp
flabel metal1 s -9488 -22168 -9456 -22140 1 FreeSans 600 0 0 0 vcascpm
flabel metal4 s -11704 3910 -11678 4004 1 FreeSans 4000 0 0 0 VDD
flabel metal4 s 594 -11002 614 -10982 1 FreeSans 600 0 0 0 vo
flabel metal1 s 22608 -8372 22614 -8354 1 FreeSans 600 0 0 0 vo
flabel metal1 s 7498 -1550 7530 -1518 1 FreeSans 600 0 0 0 M9d
flabel metal1 s 2932 -5008 3004 -4978 1 FreeSans 600 0 0 0 vcascnm
flabel metal1 s 5656 -5000 5698 -4978 1 FreeSans 600 0 0 0 vcascnp
flabel metal1 s 4210 -5038 4236 -5000 1 FreeSans 600 0 0 0 vtail_cascp
flabel metal1 s 3698 -9046 3728 -9020 1 FreeSans 600 0 0 0 vip
flabel metal1 s 4706 -9050 4736 -9016 1 FreeSans 600 0 0 0 vim
flabel metal2 s 20172 -4390 20234 -4362 1 FreeSans 600 0 0 0 vmirror
flabel metal1 s 16210 -2186 16262 -2160 1 FreeSans 600 0 0 0 VDD
flabel metal2 s 10446 -3228 10514 -3198 1 FreeSans 600 0 0 0 vcascpp
flabel metal2 s 10670 -4260 10722 -4226 1 FreeSans 600 0 0 0 vcascpm
flabel metal2 s 8324 1884 8324 1884 1 FreeSans 600 0 0 0 vbias1
flabel metal2 s 9302 1622 9332 1650 1 FreeSans 600 0 0 0 VDD
flabel metal1 s 6346 610 6380 632 1 FreeSans 600 0 0 0 M7d
flabel metal2 s 7734 486 7792 522 1 FreeSans 600 0 0 0 M13d
flabel metal2 s 9760 -1694 9838 -1660 1 FreeSans 600 0 0 0 vtail_cascp
flabel metal1 s 17510 -5860 17546 -5832 1 FreeSans 600 0 0 0 VDD
flabel metal2 s 11866 -9908 11920 -9874 1 FreeSans 600 0 0 0 M8d
flabel metal2 s 12290 -4920 12372 -4888 1 FreeSans 600 0 0 0 vbias2
flabel metal2 s 16840 -7430 16902 -7400 1 FreeSans 600 0 0 0 M16d
flabel metal2 s 16432 -7118 16496 -7086 1 FreeSans 600 0 0 0 M13d
flabel metal1 s 7324 -5080 7364 -5046 1 FreeSans 600 0 0 0 M7d
flabel metal2 s 22394 -7218 22456 -7186 1 FreeSans 600 0 0 0 vmirror
flabel metal2 s 20508 -7328 20558 -7292 1 FreeSans 600 0 0 0 vcascpm
flabel metal2 s 20560 -8376 20652 -8344 1 FreeSans 600 0 0 0 vcascpp
flabel metal2 s 7618 -6048 7618 -6048 1 FreeSans 600 0 0 0 vbias1
flabel metal2 s 7488 -9634 7544 -9600 1 FreeSans 600 0 0 0 M9d
<< properties >>
string FIXED_BBOX -10872 -26372 24872 -10428
<< end >>
