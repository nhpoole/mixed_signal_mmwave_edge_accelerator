magic
tech sky130A
magscale 1 2
timestamp 1623984492
<< metal1 >>
rect -300 60 300 117
rect -300 -117 300 -60
<< rmetal1 >>
rect -300 -60 300 60
<< properties >>
string gencell sky130_fd_pr__res_generic_m1
string parameters w 3 l 0.6 m 1 nx 1 wmin 0.14 lmin 0.14 rho 0.125 val 24.999m dummy 0 dw 0.0 term 0.0 roverlap 0
string library sky130
<< end >>
