magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -1610 -2560 1609 2560
<< metal3 >>
rect -350 1272 349 1300
rect -350 1208 265 1272
rect 329 1208 349 1272
rect -350 1192 349 1208
rect -350 1128 265 1192
rect 329 1128 349 1192
rect -350 1112 349 1128
rect -350 1048 265 1112
rect 329 1048 349 1112
rect -350 1032 349 1048
rect -350 968 265 1032
rect 329 968 349 1032
rect -350 952 349 968
rect -350 888 265 952
rect 329 888 349 952
rect -350 872 349 888
rect -350 808 265 872
rect 329 808 349 872
rect -350 792 349 808
rect -350 728 265 792
rect 329 728 349 792
rect -350 712 349 728
rect -350 648 265 712
rect 329 648 349 712
rect -350 632 349 648
rect -350 568 265 632
rect 329 568 349 632
rect -350 552 349 568
rect -350 488 265 552
rect 329 488 349 552
rect -350 472 349 488
rect -350 408 265 472
rect 329 408 349 472
rect -350 392 349 408
rect -350 328 265 392
rect 329 328 349 392
rect -350 312 349 328
rect -350 248 265 312
rect 329 248 349 312
rect -350 232 349 248
rect -350 168 265 232
rect 329 168 349 232
rect -350 152 349 168
rect -350 88 265 152
rect 329 88 349 152
rect -350 72 349 88
rect -350 8 265 72
rect 329 8 349 72
rect -350 -8 349 8
rect -350 -72 265 -8
rect 329 -72 349 -8
rect -350 -88 349 -72
rect -350 -152 265 -88
rect 329 -152 349 -88
rect -350 -168 349 -152
rect -350 -232 265 -168
rect 329 -232 349 -168
rect -350 -248 349 -232
rect -350 -312 265 -248
rect 329 -312 349 -248
rect -350 -328 349 -312
rect -350 -392 265 -328
rect 329 -392 349 -328
rect -350 -408 349 -392
rect -350 -472 265 -408
rect 329 -472 349 -408
rect -350 -488 349 -472
rect -350 -552 265 -488
rect 329 -552 349 -488
rect -350 -568 349 -552
rect -350 -632 265 -568
rect 329 -632 349 -568
rect -350 -648 349 -632
rect -350 -712 265 -648
rect 329 -712 349 -648
rect -350 -728 349 -712
rect -350 -792 265 -728
rect 329 -792 349 -728
rect -350 -808 349 -792
rect -350 -872 265 -808
rect 329 -872 349 -808
rect -350 -888 349 -872
rect -350 -952 265 -888
rect 329 -952 349 -888
rect -350 -968 349 -952
rect -350 -1032 265 -968
rect 329 -1032 349 -968
rect -350 -1048 349 -1032
rect -350 -1112 265 -1048
rect 329 -1112 349 -1048
rect -350 -1128 349 -1112
rect -350 -1192 265 -1128
rect 329 -1192 349 -1128
rect -350 -1208 349 -1192
rect -350 -1272 265 -1208
rect 329 -1272 349 -1208
rect -350 -1300 349 -1272
<< via3 >>
rect 265 1208 329 1272
rect 265 1128 329 1192
rect 265 1048 329 1112
rect 265 968 329 1032
rect 265 888 329 952
rect 265 808 329 872
rect 265 728 329 792
rect 265 648 329 712
rect 265 568 329 632
rect 265 488 329 552
rect 265 408 329 472
rect 265 328 329 392
rect 265 248 329 312
rect 265 168 329 232
rect 265 88 329 152
rect 265 8 329 72
rect 265 -72 329 -8
rect 265 -152 329 -88
rect 265 -232 329 -168
rect 265 -312 329 -248
rect 265 -392 329 -328
rect 265 -472 329 -408
rect 265 -552 329 -488
rect 265 -632 329 -568
rect 265 -712 329 -648
rect 265 -792 329 -728
rect 265 -872 329 -808
rect 265 -952 329 -888
rect 265 -1032 329 -968
rect 265 -1112 329 -1048
rect 265 -1192 329 -1128
rect 265 -1272 329 -1208
<< mimcap >>
rect -250 1152 150 1200
rect -250 -1152 -202 1152
rect 102 -1152 150 1152
rect -250 -1200 150 -1152
<< mimcapcontact >>
rect -202 -1152 102 1152
<< metal4 >>
rect 249 1272 345 1288
rect 249 1208 265 1272
rect 329 1208 345 1272
rect 249 1192 345 1208
rect -211 1152 111 1161
rect -211 -1152 -202 1152
rect 102 -1152 111 1152
rect -211 -1161 111 -1152
rect 249 1128 265 1192
rect 329 1128 345 1192
rect 249 1112 345 1128
rect 249 1048 265 1112
rect 329 1048 345 1112
rect 249 1032 345 1048
rect 249 968 265 1032
rect 329 968 345 1032
rect 249 952 345 968
rect 249 888 265 952
rect 329 888 345 952
rect 249 872 345 888
rect 249 808 265 872
rect 329 808 345 872
rect 249 792 345 808
rect 249 728 265 792
rect 329 728 345 792
rect 249 712 345 728
rect 249 648 265 712
rect 329 648 345 712
rect 249 632 345 648
rect 249 568 265 632
rect 329 568 345 632
rect 249 552 345 568
rect 249 488 265 552
rect 329 488 345 552
rect 249 472 345 488
rect 249 408 265 472
rect 329 408 345 472
rect 249 392 345 408
rect 249 328 265 392
rect 329 328 345 392
rect 249 312 345 328
rect 249 248 265 312
rect 329 248 345 312
rect 249 232 345 248
rect 249 168 265 232
rect 329 168 345 232
rect 249 152 345 168
rect 249 88 265 152
rect 329 88 345 152
rect 249 72 345 88
rect 249 8 265 72
rect 329 8 345 72
rect 249 -8 345 8
rect 249 -72 265 -8
rect 329 -72 345 -8
rect 249 -88 345 -72
rect 249 -152 265 -88
rect 329 -152 345 -88
rect 249 -168 345 -152
rect 249 -232 265 -168
rect 329 -232 345 -168
rect 249 -248 345 -232
rect 249 -312 265 -248
rect 329 -312 345 -248
rect 249 -328 345 -312
rect 249 -392 265 -328
rect 329 -392 345 -328
rect 249 -408 345 -392
rect 249 -472 265 -408
rect 329 -472 345 -408
rect 249 -488 345 -472
rect 249 -552 265 -488
rect 329 -552 345 -488
rect 249 -568 345 -552
rect 249 -632 265 -568
rect 329 -632 345 -568
rect 249 -648 345 -632
rect 249 -712 265 -648
rect 329 -712 345 -648
rect 249 -728 345 -712
rect 249 -792 265 -728
rect 329 -792 345 -728
rect 249 -808 345 -792
rect 249 -872 265 -808
rect 329 -872 345 -808
rect 249 -888 345 -872
rect 249 -952 265 -888
rect 329 -952 345 -888
rect 249 -968 345 -952
rect 249 -1032 265 -968
rect 329 -1032 345 -968
rect 249 -1048 345 -1032
rect 249 -1112 265 -1048
rect 329 -1112 345 -1048
rect 249 -1128 345 -1112
rect 249 -1192 265 -1128
rect 329 -1192 345 -1128
rect 249 -1208 345 -1192
rect 249 -1272 265 -1208
rect 329 -1272 345 -1208
rect 249 -1288 345 -1272
<< properties >>
string FIXED_BBOX -350 -1300 250 1300
<< end >>
