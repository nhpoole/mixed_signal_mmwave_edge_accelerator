magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -3726 3906 40003 18838
rect 6034 -25186 40003 3906
<< metal1 >>
rect 27146 14172 27258 14196
rect 23080 14160 23140 14166
rect 23080 14156 24468 14160
rect 23080 14104 23084 14156
rect 23136 14104 24468 14156
rect 23080 14100 24468 14104
rect 27146 14120 27176 14172
rect 27228 14120 27258 14172
rect 23080 14094 23140 14100
rect 27146 14096 27258 14120
rect 32380 14118 32930 14178
rect 29948 8646 30222 8706
<< via1 >>
rect 23084 14104 23136 14156
rect 27176 14120 27228 14172
<< metal2 >>
rect 27152 14191 27252 14202
rect 27148 14174 27256 14191
rect 23074 14156 23146 14160
rect 23074 14104 23084 14156
rect 23136 14104 23146 14156
rect 23074 14100 23146 14104
rect 27148 14118 27174 14174
rect 27230 14118 27256 14174
rect 27148 14101 27256 14118
rect 23080 9432 23140 14100
rect 27152 14090 27252 14101
rect 34621 13640 34699 13642
rect 34621 13584 34632 13640
rect 34688 13584 34699 13640
rect 34621 13582 34699 13584
rect 30988 12438 32238 12498
rect 34630 8592 34690 13582
<< via2 >>
rect 27174 14172 27230 14174
rect 27174 14120 27176 14172
rect 27176 14120 27228 14172
rect 27228 14120 27230 14172
rect 27174 14118 27230 14120
rect 34632 13584 34688 13640
<< metal3 >>
rect 27152 14174 27252 14196
rect 27152 14118 27174 14174
rect 27230 14118 27252 14174
rect 27152 13664 27252 14118
rect 27152 13640 34698 13664
rect 27152 13584 34632 13640
rect 34688 13584 34698 13640
rect 27152 13564 34698 13584
<< metal4 >>
rect 32818 17455 38736 17578
rect 32818 16899 38059 17455
rect 38615 16899 38736 17455
rect 32818 16778 38736 16899
rect 23256 10806 32856 11076
rect 30394 8472 30514 10240
rect 35772 8584 35892 10308
rect 33074 5166 33194 6154
<< via4 >>
rect 38059 16899 38615 17455
<< metal5 >>
rect 37936 17455 38736 17578
rect 37936 16899 38059 17455
rect 38615 16899 38736 17455
rect 37936 6956 38736 16899
use cs_ring_osc  cs_ring_osc_0
timestamp 1626486988
transform 1 0 -2466 0 1 6424
box 9760 -28686 41209 4472
use freq_div  freq_div_0
timestamp 1626486988
transform 1 0 32794 0 1 8554
box -2674 -2906 3321 454
use pfd_cp_lpf  pfd_cp_lpf_0
timestamp 1626486988
transform -1 0 30256 0 1 14838
box -2600 -3860 7000 2740
<< labels >>
flabel metal1 s 32888 14140 32900 14154 1 FreeSans 600 0 0 0 vsigin
flabel metal2 s 32196 12456 32208 12470 1 FreeSans 600 0 0 0 ibiasn
flabel metal4 s 30452 9650 30462 9664 1 FreeSans 600 0 0 0 VSS
flabel metal4 s 33486 17114 33506 17132 1 FreeSans 600 0 0 0 VDD
flabel metal1 s 23198 14118 23210 14134 1 FreeSans 600 0 0 0 vcp
<< end >>
