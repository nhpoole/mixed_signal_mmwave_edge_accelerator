magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -1454 -1760 1454 1760
<< nwell >>
rect -194 -500 194 500
<< pmoshvt >>
rect -100 -400 100 400
<< pdiff >>
rect -158 357 -100 400
rect -158 323 -146 357
rect -112 323 -100 357
rect -158 289 -100 323
rect -158 255 -146 289
rect -112 255 -100 289
rect -158 221 -100 255
rect -158 187 -146 221
rect -112 187 -100 221
rect -158 153 -100 187
rect -158 119 -146 153
rect -112 119 -100 153
rect -158 85 -100 119
rect -158 51 -146 85
rect -112 51 -100 85
rect -158 17 -100 51
rect -158 -17 -146 17
rect -112 -17 -100 17
rect -158 -51 -100 -17
rect -158 -85 -146 -51
rect -112 -85 -100 -51
rect -158 -119 -100 -85
rect -158 -153 -146 -119
rect -112 -153 -100 -119
rect -158 -187 -100 -153
rect -158 -221 -146 -187
rect -112 -221 -100 -187
rect -158 -255 -100 -221
rect -158 -289 -146 -255
rect -112 -289 -100 -255
rect -158 -323 -100 -289
rect -158 -357 -146 -323
rect -112 -357 -100 -323
rect -158 -400 -100 -357
rect 100 357 158 400
rect 100 323 112 357
rect 146 323 158 357
rect 100 289 158 323
rect 100 255 112 289
rect 146 255 158 289
rect 100 221 158 255
rect 100 187 112 221
rect 146 187 158 221
rect 100 153 158 187
rect 100 119 112 153
rect 146 119 158 153
rect 100 85 158 119
rect 100 51 112 85
rect 146 51 158 85
rect 100 17 158 51
rect 100 -17 112 17
rect 146 -17 158 17
rect 100 -51 158 -17
rect 100 -85 112 -51
rect 146 -85 158 -51
rect 100 -119 158 -85
rect 100 -153 112 -119
rect 146 -153 158 -119
rect 100 -187 158 -153
rect 100 -221 112 -187
rect 146 -221 158 -187
rect 100 -255 158 -221
rect 100 -289 112 -255
rect 146 -289 158 -255
rect 100 -323 158 -289
rect 100 -357 112 -323
rect 146 -357 158 -323
rect 100 -400 158 -357
<< pdiffc >>
rect -146 323 -112 357
rect -146 255 -112 289
rect -146 187 -112 221
rect -146 119 -112 153
rect -146 51 -112 85
rect -146 -17 -112 17
rect -146 -85 -112 -51
rect -146 -153 -112 -119
rect -146 -221 -112 -187
rect -146 -289 -112 -255
rect -146 -357 -112 -323
rect 112 323 146 357
rect 112 255 146 289
rect 112 187 146 221
rect 112 119 146 153
rect 112 51 146 85
rect 112 -17 146 17
rect 112 -85 146 -51
rect 112 -153 146 -119
rect 112 -221 146 -187
rect 112 -289 146 -255
rect 112 -357 146 -323
<< poly >>
rect -66 481 66 497
rect -66 464 -17 481
rect -100 447 -17 464
rect 17 464 66 481
rect 17 447 100 464
rect -100 400 100 447
rect -100 -447 100 -400
rect -100 -464 -17 -447
rect -66 -481 -17 -464
rect 17 -464 100 -447
rect 17 -481 66 -464
rect -66 -497 66 -481
<< polycont >>
rect -17 447 17 481
rect -17 -481 17 -447
<< locali >>
rect -66 447 -17 481
rect 17 447 66 481
rect -146 377 -112 404
rect -146 305 -112 323
rect -146 233 -112 255
rect -146 161 -112 187
rect -146 89 -112 119
rect -146 17 -112 51
rect -146 -51 -112 -17
rect -146 -119 -112 -89
rect -146 -187 -112 -161
rect -146 -255 -112 -233
rect -146 -323 -112 -305
rect -146 -404 -112 -377
rect 112 377 146 404
rect 112 305 146 323
rect 112 233 146 255
rect 112 161 146 187
rect 112 89 146 119
rect 112 17 146 51
rect 112 -51 146 -17
rect 112 -119 146 -89
rect 112 -187 146 -161
rect 112 -255 146 -233
rect 112 -323 146 -305
rect 112 -404 146 -377
rect -66 -481 -17 -447
rect 17 -481 66 -447
<< viali >>
rect -17 447 17 481
rect -146 357 -112 377
rect -146 343 -112 357
rect -146 289 -112 305
rect -146 271 -112 289
rect -146 221 -112 233
rect -146 199 -112 221
rect -146 153 -112 161
rect -146 127 -112 153
rect -146 85 -112 89
rect -146 55 -112 85
rect -146 -17 -112 17
rect -146 -85 -112 -55
rect -146 -89 -112 -85
rect -146 -153 -112 -127
rect -146 -161 -112 -153
rect -146 -221 -112 -199
rect -146 -233 -112 -221
rect -146 -289 -112 -271
rect -146 -305 -112 -289
rect -146 -357 -112 -343
rect -146 -377 -112 -357
rect 112 357 146 377
rect 112 343 146 357
rect 112 289 146 305
rect 112 271 146 289
rect 112 221 146 233
rect 112 199 146 221
rect 112 153 146 161
rect 112 127 146 153
rect 112 85 146 89
rect 112 55 146 85
rect 112 -17 146 17
rect 112 -85 146 -55
rect 112 -89 146 -85
rect 112 -153 146 -127
rect 112 -161 146 -153
rect 112 -221 146 -199
rect 112 -233 146 -221
rect 112 -289 146 -271
rect 112 -305 146 -289
rect 112 -357 146 -343
rect 112 -377 146 -357
rect -17 -481 17 -447
<< metal1 >>
rect -54 481 54 487
rect -54 447 -17 481
rect 17 447 54 481
rect -54 441 54 447
rect -152 377 -106 400
rect -152 343 -146 377
rect -112 343 -106 377
rect -152 305 -106 343
rect -152 271 -146 305
rect -112 271 -106 305
rect -152 233 -106 271
rect -152 199 -146 233
rect -112 199 -106 233
rect -152 161 -106 199
rect -152 127 -146 161
rect -112 127 -106 161
rect -152 89 -106 127
rect -152 55 -146 89
rect -112 55 -106 89
rect -152 17 -106 55
rect -152 -17 -146 17
rect -112 -17 -106 17
rect -152 -55 -106 -17
rect -152 -89 -146 -55
rect -112 -89 -106 -55
rect -152 -127 -106 -89
rect -152 -161 -146 -127
rect -112 -161 -106 -127
rect -152 -199 -106 -161
rect -152 -233 -146 -199
rect -112 -233 -106 -199
rect -152 -271 -106 -233
rect -152 -305 -146 -271
rect -112 -305 -106 -271
rect -152 -343 -106 -305
rect -152 -377 -146 -343
rect -112 -377 -106 -343
rect -152 -400 -106 -377
rect 106 377 152 400
rect 106 343 112 377
rect 146 343 152 377
rect 106 305 152 343
rect 106 271 112 305
rect 146 271 152 305
rect 106 233 152 271
rect 106 199 112 233
rect 146 199 152 233
rect 106 161 152 199
rect 106 127 112 161
rect 146 127 152 161
rect 106 89 152 127
rect 106 55 112 89
rect 146 55 152 89
rect 106 17 152 55
rect 106 -17 112 17
rect 146 -17 152 17
rect 106 -55 152 -17
rect 106 -89 112 -55
rect 146 -89 152 -55
rect 106 -127 152 -89
rect 106 -161 112 -127
rect 146 -161 152 -127
rect 106 -199 152 -161
rect 106 -233 112 -199
rect 146 -233 152 -199
rect 106 -271 152 -233
rect 106 -305 112 -271
rect 146 -305 152 -271
rect 106 -343 152 -305
rect 106 -377 112 -343
rect 146 -377 152 -343
rect 106 -400 152 -377
rect -54 -447 54 -441
rect -54 -481 -17 -447
rect 17 -481 54 -447
rect -54 -487 54 -481
<< end >>
