magic
tech sky130A
magscale 1 2
timestamp 1622100421
<< nwell >>
rect -3497 -200 3497 200
<< pmos >>
rect -3403 -100 -2603 100
rect -2545 -100 -1745 100
rect -1687 -100 -887 100
rect -829 -100 -29 100
rect 29 -100 829 100
rect 887 -100 1687 100
rect 1745 -100 2545 100
rect 2603 -100 3403 100
<< pdiff >>
rect -3461 88 -3403 100
rect -3461 -88 -3449 88
rect -3415 -88 -3403 88
rect -3461 -100 -3403 -88
rect -2603 88 -2545 100
rect -2603 -88 -2591 88
rect -2557 -88 -2545 88
rect -2603 -100 -2545 -88
rect -1745 88 -1687 100
rect -1745 -88 -1733 88
rect -1699 -88 -1687 88
rect -1745 -100 -1687 -88
rect -887 88 -829 100
rect -887 -88 -875 88
rect -841 -88 -829 88
rect -887 -100 -829 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 829 88 887 100
rect 829 -88 841 88
rect 875 -88 887 88
rect 829 -100 887 -88
rect 1687 88 1745 100
rect 1687 -88 1699 88
rect 1733 -88 1745 88
rect 1687 -100 1745 -88
rect 2545 88 2603 100
rect 2545 -88 2557 88
rect 2591 -88 2603 88
rect 2545 -100 2603 -88
rect 3403 88 3461 100
rect 3403 -88 3415 88
rect 3449 -88 3461 88
rect 3403 -100 3461 -88
<< pdiffc >>
rect -3449 -88 -3415 88
rect -2591 -88 -2557 88
rect -1733 -88 -1699 88
rect -875 -88 -841 88
rect -17 -88 17 88
rect 841 -88 875 88
rect 1699 -88 1733 88
rect 2557 -88 2591 88
rect 3415 -88 3449 88
<< poly >>
rect -3211 181 -2795 197
rect -3211 164 -3195 181
rect -3403 147 -3195 164
rect -2811 164 -2795 181
rect -2353 181 -1937 197
rect -2353 164 -2337 181
rect -2811 147 -2603 164
rect -3403 100 -2603 147
rect -2545 147 -2337 164
rect -1953 164 -1937 181
rect -1495 181 -1079 197
rect -1495 164 -1479 181
rect -1953 147 -1745 164
rect -2545 100 -1745 147
rect -1687 147 -1479 164
rect -1095 164 -1079 181
rect -637 181 -221 197
rect -637 164 -621 181
rect -1095 147 -887 164
rect -1687 100 -887 147
rect -829 147 -621 164
rect -237 164 -221 181
rect 221 181 637 197
rect 221 164 237 181
rect -237 147 -29 164
rect -829 100 -29 147
rect 29 147 237 164
rect 621 164 637 181
rect 1079 181 1495 197
rect 1079 164 1095 181
rect 621 147 829 164
rect 29 100 829 147
rect 887 147 1095 164
rect 1479 164 1495 181
rect 1937 181 2353 197
rect 1937 164 1953 181
rect 1479 147 1687 164
rect 887 100 1687 147
rect 1745 147 1953 164
rect 2337 164 2353 181
rect 2795 181 3211 197
rect 2795 164 2811 181
rect 2337 147 2545 164
rect 1745 100 2545 147
rect 2603 147 2811 164
rect 3195 164 3211 181
rect 3195 147 3403 164
rect 2603 100 3403 147
rect -3403 -147 -2603 -100
rect -3403 -164 -3195 -147
rect -3211 -181 -3195 -164
rect -2811 -164 -2603 -147
rect -2545 -147 -1745 -100
rect -2545 -164 -2337 -147
rect -2811 -181 -2795 -164
rect -3211 -197 -2795 -181
rect -2353 -181 -2337 -164
rect -1953 -164 -1745 -147
rect -1687 -147 -887 -100
rect -1687 -164 -1479 -147
rect -1953 -181 -1937 -164
rect -2353 -197 -1937 -181
rect -1495 -181 -1479 -164
rect -1095 -164 -887 -147
rect -829 -147 -29 -100
rect -829 -164 -621 -147
rect -1095 -181 -1079 -164
rect -1495 -197 -1079 -181
rect -637 -181 -621 -164
rect -237 -164 -29 -147
rect 29 -147 829 -100
rect 29 -164 237 -147
rect -237 -181 -221 -164
rect -637 -197 -221 -181
rect 221 -181 237 -164
rect 621 -164 829 -147
rect 887 -147 1687 -100
rect 887 -164 1095 -147
rect 621 -181 637 -164
rect 221 -197 637 -181
rect 1079 -181 1095 -164
rect 1479 -164 1687 -147
rect 1745 -147 2545 -100
rect 1745 -164 1953 -147
rect 1479 -181 1495 -164
rect 1079 -197 1495 -181
rect 1937 -181 1953 -164
rect 2337 -164 2545 -147
rect 2603 -147 3403 -100
rect 2603 -164 2811 -147
rect 2337 -181 2353 -164
rect 1937 -197 2353 -181
rect 2795 -181 2811 -164
rect 3195 -164 3403 -147
rect 3195 -181 3211 -164
rect 2795 -197 3211 -181
<< polycont >>
rect -3195 147 -2811 181
rect -2337 147 -1953 181
rect -1479 147 -1095 181
rect -621 147 -237 181
rect 237 147 621 181
rect 1095 147 1479 181
rect 1953 147 2337 181
rect 2811 147 3195 181
rect -3195 -181 -2811 -147
rect -2337 -181 -1953 -147
rect -1479 -181 -1095 -147
rect -621 -181 -237 -147
rect 237 -181 621 -147
rect 1095 -181 1479 -147
rect 1953 -181 2337 -147
rect 2811 -181 3195 -147
<< locali >>
rect -3211 147 -3195 181
rect -2811 147 -2795 181
rect -2353 147 -2337 181
rect -1953 147 -1937 181
rect -1495 147 -1479 181
rect -1095 147 -1079 181
rect -637 147 -621 181
rect -237 147 -221 181
rect 221 147 237 181
rect 621 147 637 181
rect 1079 147 1095 181
rect 1479 147 1495 181
rect 1937 147 1953 181
rect 2337 147 2353 181
rect 2795 147 2811 181
rect 3195 147 3211 181
rect -3449 88 -3415 104
rect -3449 -104 -3415 -88
rect -2591 88 -2557 104
rect -2591 -104 -2557 -88
rect -1733 88 -1699 104
rect -1733 -104 -1699 -88
rect -875 88 -841 104
rect -875 -104 -841 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 841 88 875 104
rect 841 -104 875 -88
rect 1699 88 1733 104
rect 1699 -104 1733 -88
rect 2557 88 2591 104
rect 2557 -104 2591 -88
rect 3415 88 3449 104
rect 3415 -104 3449 -88
rect -3211 -181 -3195 -147
rect -2811 -181 -2795 -147
rect -2353 -181 -2337 -147
rect -1953 -181 -1937 -147
rect -1495 -181 -1479 -147
rect -1095 -181 -1079 -147
rect -637 -181 -621 -147
rect -237 -181 -221 -147
rect 221 -181 237 -147
rect 621 -181 637 -147
rect 1079 -181 1095 -147
rect 1479 -181 1495 -147
rect 1937 -181 1953 -147
rect 2337 -181 2353 -147
rect 2795 -181 2811 -147
rect 3195 -181 3211 -147
<< viali >>
rect -3195 147 -2811 181
rect -2337 147 -1953 181
rect -1479 147 -1095 181
rect -621 147 -237 181
rect 237 147 621 181
rect 1095 147 1479 181
rect 1953 147 2337 181
rect 2811 147 3195 181
rect -3449 -88 -3415 88
rect -2591 -88 -2557 88
rect -1733 -88 -1699 88
rect -875 -88 -841 88
rect -17 -88 17 88
rect 841 -88 875 88
rect 1699 -88 1733 88
rect 2557 -88 2591 88
rect 3415 -88 3449 88
rect -3195 -181 -2811 -147
rect -2337 -181 -1953 -147
rect -1479 -181 -1095 -147
rect -621 -181 -237 -147
rect 237 -181 621 -147
rect 1095 -181 1479 -147
rect 1953 -181 2337 -147
rect 2811 -181 3195 -147
<< metal1 >>
rect -3207 181 -2799 187
rect -3207 147 -3195 181
rect -2811 147 -2799 181
rect -3207 141 -2799 147
rect -2349 181 -1941 187
rect -2349 147 -2337 181
rect -1953 147 -1941 181
rect -2349 141 -1941 147
rect -1491 181 -1083 187
rect -1491 147 -1479 181
rect -1095 147 -1083 181
rect -1491 141 -1083 147
rect -633 181 -225 187
rect -633 147 -621 181
rect -237 147 -225 181
rect -633 141 -225 147
rect 225 181 633 187
rect 225 147 237 181
rect 621 147 633 181
rect 225 141 633 147
rect 1083 181 1491 187
rect 1083 147 1095 181
rect 1479 147 1491 181
rect 1083 141 1491 147
rect 1941 181 2349 187
rect 1941 147 1953 181
rect 2337 147 2349 181
rect 1941 141 2349 147
rect 2799 181 3207 187
rect 2799 147 2811 181
rect 3195 147 3207 181
rect 2799 141 3207 147
rect -3455 88 -3409 100
rect -3455 -88 -3449 88
rect -3415 -88 -3409 88
rect -3455 -100 -3409 -88
rect -2597 88 -2551 100
rect -2597 -88 -2591 88
rect -2557 -88 -2551 88
rect -2597 -100 -2551 -88
rect -1739 88 -1693 100
rect -1739 -88 -1733 88
rect -1699 -88 -1693 88
rect -1739 -100 -1693 -88
rect -881 88 -835 100
rect -881 -88 -875 88
rect -841 -88 -835 88
rect -881 -100 -835 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 835 88 881 100
rect 835 -88 841 88
rect 875 -88 881 88
rect 835 -100 881 -88
rect 1693 88 1739 100
rect 1693 -88 1699 88
rect 1733 -88 1739 88
rect 1693 -100 1739 -88
rect 2551 88 2597 100
rect 2551 -88 2557 88
rect 2591 -88 2597 88
rect 2551 -100 2597 -88
rect 3409 88 3455 100
rect 3409 -88 3415 88
rect 3449 -88 3455 88
rect 3409 -100 3455 -88
rect -3207 -147 -2799 -141
rect -3207 -181 -3195 -147
rect -2811 -181 -2799 -147
rect -3207 -187 -2799 -181
rect -2349 -147 -1941 -141
rect -2349 -181 -2337 -147
rect -1953 -181 -1941 -147
rect -2349 -187 -1941 -181
rect -1491 -147 -1083 -141
rect -1491 -181 -1479 -147
rect -1095 -181 -1083 -147
rect -1491 -187 -1083 -181
rect -633 -147 -225 -141
rect -633 -181 -621 -147
rect -237 -181 -225 -147
rect -633 -187 -225 -181
rect 225 -147 633 -141
rect 225 -181 237 -147
rect 621 -181 633 -147
rect 225 -187 633 -181
rect 1083 -147 1491 -141
rect 1083 -181 1095 -147
rect 1479 -181 1491 -147
rect 1083 -187 1491 -181
rect 1941 -147 2349 -141
rect 1941 -181 1953 -147
rect 2337 -181 2349 -147
rect 1941 -187 2349 -181
rect 2799 -147 3207 -141
rect 2799 -181 2811 -147
rect 3195 -181 3207 -147
rect 2799 -187 3207 -181
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 1 l 4 m 1 nf 8 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
