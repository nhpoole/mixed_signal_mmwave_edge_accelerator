magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< error_p >>
rect -1609 -500 -1551 500
rect -1451 -500 -1393 500
rect -1293 -500 -1235 500
rect -1135 -500 -1077 500
rect -977 -500 -919 500
rect -819 -500 -761 500
rect -661 -500 -603 500
rect -503 -500 -445 500
rect -345 -500 -287 500
rect -187 -500 -129 500
rect -29 -500 29 500
rect 129 -500 187 500
rect 287 -500 345 500
rect 445 -500 503 500
rect 603 -500 661 500
rect 761 -500 819 500
rect 919 -500 977 500
rect 1077 -500 1135 500
rect 1235 -500 1293 500
rect 1393 -500 1451 500
rect 1551 -500 1609 500
<< mvnmos >>
rect -1551 -500 -1451 500
rect -1393 -500 -1293 500
rect -1235 -500 -1135 500
rect -1077 -500 -977 500
rect -919 -500 -819 500
rect -761 -500 -661 500
rect -603 -500 -503 500
rect -445 -500 -345 500
rect -287 -500 -187 500
rect -129 -500 -29 500
rect 29 -500 129 500
rect 187 -500 287 500
rect 345 -500 445 500
rect 503 -500 603 500
rect 661 -500 761 500
rect 819 -500 919 500
rect 977 -500 1077 500
rect 1135 -500 1235 500
rect 1293 -500 1393 500
rect 1451 -500 1551 500
<< mvndiff >>
rect -1609 488 -1551 500
rect -1609 -488 -1597 488
rect -1563 -488 -1551 488
rect -1609 -500 -1551 -488
rect -1451 488 -1393 500
rect -1451 -488 -1439 488
rect -1405 -488 -1393 488
rect -1451 -500 -1393 -488
rect -1293 488 -1235 500
rect -1293 -488 -1281 488
rect -1247 -488 -1235 488
rect -1293 -500 -1235 -488
rect -1135 488 -1077 500
rect -1135 -488 -1123 488
rect -1089 -488 -1077 488
rect -1135 -500 -1077 -488
rect -977 488 -919 500
rect -977 -488 -965 488
rect -931 -488 -919 488
rect -977 -500 -919 -488
rect -819 488 -761 500
rect -819 -488 -807 488
rect -773 -488 -761 488
rect -819 -500 -761 -488
rect -661 488 -603 500
rect -661 -488 -649 488
rect -615 -488 -603 488
rect -661 -500 -603 -488
rect -503 488 -445 500
rect -503 -488 -491 488
rect -457 -488 -445 488
rect -503 -500 -445 -488
rect -345 488 -287 500
rect -345 -488 -333 488
rect -299 -488 -287 488
rect -345 -500 -287 -488
rect -187 488 -129 500
rect -187 -488 -175 488
rect -141 -488 -129 488
rect -187 -500 -129 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 129 488 187 500
rect 129 -488 141 488
rect 175 -488 187 488
rect 129 -500 187 -488
rect 287 488 345 500
rect 287 -488 299 488
rect 333 -488 345 488
rect 287 -500 345 -488
rect 445 488 503 500
rect 445 -488 457 488
rect 491 -488 503 488
rect 445 -500 503 -488
rect 603 488 661 500
rect 603 -488 615 488
rect 649 -488 661 488
rect 603 -500 661 -488
rect 761 488 819 500
rect 761 -488 773 488
rect 807 -488 819 488
rect 761 -500 819 -488
rect 919 488 977 500
rect 919 -488 931 488
rect 965 -488 977 488
rect 919 -500 977 -488
rect 1077 488 1135 500
rect 1077 -488 1089 488
rect 1123 -488 1135 488
rect 1077 -500 1135 -488
rect 1235 488 1293 500
rect 1235 -488 1247 488
rect 1281 -488 1293 488
rect 1235 -500 1293 -488
rect 1393 488 1451 500
rect 1393 -488 1405 488
rect 1439 -488 1451 488
rect 1393 -500 1451 -488
rect 1551 488 1609 500
rect 1551 -488 1563 488
rect 1597 -488 1609 488
rect 1551 -500 1609 -488
<< mvndiffc >>
rect -1597 -488 -1563 488
rect -1439 -488 -1405 488
rect -1281 -488 -1247 488
rect -1123 -488 -1089 488
rect -965 -488 -931 488
rect -807 -488 -773 488
rect -649 -488 -615 488
rect -491 -488 -457 488
rect -333 -488 -299 488
rect -175 -488 -141 488
rect -17 -488 17 488
rect 141 -488 175 488
rect 299 -488 333 488
rect 457 -488 491 488
rect 615 -488 649 488
rect 773 -488 807 488
rect 931 -488 965 488
rect 1089 -488 1123 488
rect 1247 -488 1281 488
rect 1405 -488 1439 488
rect 1563 -488 1597 488
<< poly >>
rect -1537 572 -1465 588
rect -1537 555 -1521 572
rect -1551 538 -1521 555
rect -1481 555 -1465 572
rect -1379 572 -1307 588
rect -1379 555 -1363 572
rect -1481 538 -1451 555
rect -1551 500 -1451 538
rect -1393 538 -1363 555
rect -1323 555 -1307 572
rect -1221 572 -1149 588
rect -1221 555 -1205 572
rect -1323 538 -1293 555
rect -1393 500 -1293 538
rect -1235 538 -1205 555
rect -1165 555 -1149 572
rect -1063 572 -991 588
rect -1063 555 -1047 572
rect -1165 538 -1135 555
rect -1235 500 -1135 538
rect -1077 538 -1047 555
rect -1007 555 -991 572
rect -905 572 -833 588
rect -905 555 -889 572
rect -1007 538 -977 555
rect -1077 500 -977 538
rect -919 538 -889 555
rect -849 555 -833 572
rect -747 572 -675 588
rect -747 555 -731 572
rect -849 538 -819 555
rect -919 500 -819 538
rect -761 538 -731 555
rect -691 555 -675 572
rect -589 572 -517 588
rect -589 555 -573 572
rect -691 538 -661 555
rect -761 500 -661 538
rect -603 538 -573 555
rect -533 555 -517 572
rect -431 572 -359 588
rect -431 555 -415 572
rect -533 538 -503 555
rect -603 500 -503 538
rect -445 538 -415 555
rect -375 555 -359 572
rect -273 572 -201 588
rect -273 555 -257 572
rect -375 538 -345 555
rect -445 500 -345 538
rect -287 538 -257 555
rect -217 555 -201 572
rect -115 572 -43 588
rect -115 555 -99 572
rect -217 538 -187 555
rect -287 500 -187 538
rect -129 538 -99 555
rect -59 555 -43 572
rect 43 572 115 588
rect 43 555 59 572
rect -59 538 -29 555
rect -129 500 -29 538
rect 29 538 59 555
rect 99 555 115 572
rect 201 572 273 588
rect 201 555 217 572
rect 99 538 129 555
rect 29 500 129 538
rect 187 538 217 555
rect 257 555 273 572
rect 359 572 431 588
rect 359 555 375 572
rect 257 538 287 555
rect 187 500 287 538
rect 345 538 375 555
rect 415 555 431 572
rect 517 572 589 588
rect 517 555 533 572
rect 415 538 445 555
rect 345 500 445 538
rect 503 538 533 555
rect 573 555 589 572
rect 675 572 747 588
rect 675 555 691 572
rect 573 538 603 555
rect 503 500 603 538
rect 661 538 691 555
rect 731 555 747 572
rect 833 572 905 588
rect 833 555 849 572
rect 731 538 761 555
rect 661 500 761 538
rect 819 538 849 555
rect 889 555 905 572
rect 991 572 1063 588
rect 991 555 1007 572
rect 889 538 919 555
rect 819 500 919 538
rect 977 538 1007 555
rect 1047 555 1063 572
rect 1149 572 1221 588
rect 1149 555 1165 572
rect 1047 538 1077 555
rect 977 500 1077 538
rect 1135 538 1165 555
rect 1205 555 1221 572
rect 1307 572 1379 588
rect 1307 555 1323 572
rect 1205 538 1235 555
rect 1135 500 1235 538
rect 1293 538 1323 555
rect 1363 555 1379 572
rect 1465 572 1537 588
rect 1465 555 1481 572
rect 1363 538 1393 555
rect 1293 500 1393 538
rect 1451 538 1481 555
rect 1521 555 1537 572
rect 1521 538 1551 555
rect 1451 500 1551 538
rect -1551 -538 -1451 -500
rect -1551 -555 -1521 -538
rect -1537 -572 -1521 -555
rect -1481 -555 -1451 -538
rect -1393 -538 -1293 -500
rect -1393 -555 -1363 -538
rect -1481 -572 -1465 -555
rect -1537 -588 -1465 -572
rect -1379 -572 -1363 -555
rect -1323 -555 -1293 -538
rect -1235 -538 -1135 -500
rect -1235 -555 -1205 -538
rect -1323 -572 -1307 -555
rect -1379 -588 -1307 -572
rect -1221 -572 -1205 -555
rect -1165 -555 -1135 -538
rect -1077 -538 -977 -500
rect -1077 -555 -1047 -538
rect -1165 -572 -1149 -555
rect -1221 -588 -1149 -572
rect -1063 -572 -1047 -555
rect -1007 -555 -977 -538
rect -919 -538 -819 -500
rect -919 -555 -889 -538
rect -1007 -572 -991 -555
rect -1063 -588 -991 -572
rect -905 -572 -889 -555
rect -849 -555 -819 -538
rect -761 -538 -661 -500
rect -761 -555 -731 -538
rect -849 -572 -833 -555
rect -905 -588 -833 -572
rect -747 -572 -731 -555
rect -691 -555 -661 -538
rect -603 -538 -503 -500
rect -603 -555 -573 -538
rect -691 -572 -675 -555
rect -747 -588 -675 -572
rect -589 -572 -573 -555
rect -533 -555 -503 -538
rect -445 -538 -345 -500
rect -445 -555 -415 -538
rect -533 -572 -517 -555
rect -589 -588 -517 -572
rect -431 -572 -415 -555
rect -375 -555 -345 -538
rect -287 -538 -187 -500
rect -287 -555 -257 -538
rect -375 -572 -359 -555
rect -431 -588 -359 -572
rect -273 -572 -257 -555
rect -217 -555 -187 -538
rect -129 -538 -29 -500
rect -129 -555 -99 -538
rect -217 -572 -201 -555
rect -273 -588 -201 -572
rect -115 -572 -99 -555
rect -59 -555 -29 -538
rect 29 -538 129 -500
rect 29 -555 59 -538
rect -59 -572 -43 -555
rect -115 -588 -43 -572
rect 43 -572 59 -555
rect 99 -555 129 -538
rect 187 -538 287 -500
rect 187 -555 217 -538
rect 99 -572 115 -555
rect 43 -588 115 -572
rect 201 -572 217 -555
rect 257 -555 287 -538
rect 345 -538 445 -500
rect 345 -555 375 -538
rect 257 -572 273 -555
rect 201 -588 273 -572
rect 359 -572 375 -555
rect 415 -555 445 -538
rect 503 -538 603 -500
rect 503 -555 533 -538
rect 415 -572 431 -555
rect 359 -588 431 -572
rect 517 -572 533 -555
rect 573 -555 603 -538
rect 661 -538 761 -500
rect 661 -555 691 -538
rect 573 -572 589 -555
rect 517 -588 589 -572
rect 675 -572 691 -555
rect 731 -555 761 -538
rect 819 -538 919 -500
rect 819 -555 849 -538
rect 731 -572 747 -555
rect 675 -588 747 -572
rect 833 -572 849 -555
rect 889 -555 919 -538
rect 977 -538 1077 -500
rect 977 -555 1007 -538
rect 889 -572 905 -555
rect 833 -588 905 -572
rect 991 -572 1007 -555
rect 1047 -555 1077 -538
rect 1135 -538 1235 -500
rect 1135 -555 1165 -538
rect 1047 -572 1063 -555
rect 991 -588 1063 -572
rect 1149 -572 1165 -555
rect 1205 -555 1235 -538
rect 1293 -538 1393 -500
rect 1293 -555 1323 -538
rect 1205 -572 1221 -555
rect 1149 -588 1221 -572
rect 1307 -572 1323 -555
rect 1363 -555 1393 -538
rect 1451 -538 1551 -500
rect 1451 -555 1481 -538
rect 1363 -572 1379 -555
rect 1307 -588 1379 -572
rect 1465 -572 1481 -555
rect 1521 -555 1551 -538
rect 1521 -572 1537 -555
rect 1465 -588 1537 -572
<< polycont >>
rect -1521 538 -1481 572
rect -1363 538 -1323 572
rect -1205 538 -1165 572
rect -1047 538 -1007 572
rect -889 538 -849 572
rect -731 538 -691 572
rect -573 538 -533 572
rect -415 538 -375 572
rect -257 538 -217 572
rect -99 538 -59 572
rect 59 538 99 572
rect 217 538 257 572
rect 375 538 415 572
rect 533 538 573 572
rect 691 538 731 572
rect 849 538 889 572
rect 1007 538 1047 572
rect 1165 538 1205 572
rect 1323 538 1363 572
rect 1481 538 1521 572
rect -1521 -572 -1481 -538
rect -1363 -572 -1323 -538
rect -1205 -572 -1165 -538
rect -1047 -572 -1007 -538
rect -889 -572 -849 -538
rect -731 -572 -691 -538
rect -573 -572 -533 -538
rect -415 -572 -375 -538
rect -257 -572 -217 -538
rect -99 -572 -59 -538
rect 59 -572 99 -538
rect 217 -572 257 -538
rect 375 -572 415 -538
rect 533 -572 573 -538
rect 691 -572 731 -538
rect 849 -572 889 -538
rect 1007 -572 1047 -538
rect 1165 -572 1205 -538
rect 1323 -572 1363 -538
rect 1481 -572 1521 -538
<< locali >>
rect -1537 538 -1521 572
rect -1481 538 -1465 572
rect -1379 538 -1363 572
rect -1323 538 -1307 572
rect -1221 538 -1205 572
rect -1165 538 -1149 572
rect -1063 538 -1047 572
rect -1007 538 -991 572
rect -905 538 -889 572
rect -849 538 -833 572
rect -747 538 -731 572
rect -691 538 -675 572
rect -589 538 -573 572
rect -533 538 -517 572
rect -431 538 -415 572
rect -375 538 -359 572
rect -273 538 -257 572
rect -217 538 -201 572
rect -115 538 -99 572
rect -59 538 -43 572
rect 43 538 59 572
rect 99 538 115 572
rect 201 538 217 572
rect 257 538 273 572
rect 359 538 375 572
rect 415 538 431 572
rect 517 538 533 572
rect 573 538 589 572
rect 675 538 691 572
rect 731 538 747 572
rect 833 538 849 572
rect 889 538 905 572
rect 991 538 1007 572
rect 1047 538 1063 572
rect 1149 538 1165 572
rect 1205 538 1221 572
rect 1307 538 1323 572
rect 1363 538 1379 572
rect 1465 538 1481 572
rect 1521 538 1537 572
rect -1597 488 -1563 504
rect -1597 -504 -1563 -488
rect -1439 488 -1405 504
rect -1439 -504 -1405 -488
rect -1281 488 -1247 504
rect -1281 -504 -1247 -488
rect -1123 488 -1089 504
rect -1123 -504 -1089 -488
rect -965 488 -931 504
rect -965 -504 -931 -488
rect -807 488 -773 504
rect -807 -504 -773 -488
rect -649 488 -615 504
rect -649 -504 -615 -488
rect -491 488 -457 504
rect -491 -504 -457 -488
rect -333 488 -299 504
rect -333 -504 -299 -488
rect -175 488 -141 504
rect -175 -504 -141 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 141 488 175 504
rect 141 -504 175 -488
rect 299 488 333 504
rect 299 -504 333 -488
rect 457 488 491 504
rect 457 -504 491 -488
rect 615 488 649 504
rect 615 -504 649 -488
rect 773 488 807 504
rect 773 -504 807 -488
rect 931 488 965 504
rect 931 -504 965 -488
rect 1089 488 1123 504
rect 1089 -504 1123 -488
rect 1247 488 1281 504
rect 1247 -504 1281 -488
rect 1405 488 1439 504
rect 1405 -504 1439 -488
rect 1563 488 1597 504
rect 1563 -504 1597 -488
rect -1537 -572 -1521 -538
rect -1481 -572 -1465 -538
rect -1379 -572 -1363 -538
rect -1323 -572 -1307 -538
rect -1221 -572 -1205 -538
rect -1165 -572 -1149 -538
rect -1063 -572 -1047 -538
rect -1007 -572 -991 -538
rect -905 -572 -889 -538
rect -849 -572 -833 -538
rect -747 -572 -731 -538
rect -691 -572 -675 -538
rect -589 -572 -573 -538
rect -533 -572 -517 -538
rect -431 -572 -415 -538
rect -375 -572 -359 -538
rect -273 -572 -257 -538
rect -217 -572 -201 -538
rect -115 -572 -99 -538
rect -59 -572 -43 -538
rect 43 -572 59 -538
rect 99 -572 115 -538
rect 201 -572 217 -538
rect 257 -572 273 -538
rect 359 -572 375 -538
rect 415 -572 431 -538
rect 517 -572 533 -538
rect 573 -572 589 -538
rect 675 -572 691 -538
rect 731 -572 747 -538
rect 833 -572 849 -538
rect 889 -572 905 -538
rect 991 -572 1007 -538
rect 1047 -572 1063 -538
rect 1149 -572 1165 -538
rect 1205 -572 1221 -538
rect 1307 -572 1323 -538
rect 1363 -572 1379 -538
rect 1465 -572 1481 -538
rect 1521 -572 1537 -538
<< viali >>
rect -1597 -488 -1563 488
rect -1439 -488 -1405 488
rect -1281 -488 -1247 488
rect -1123 -488 -1089 488
rect -965 -488 -931 488
rect -807 -488 -773 488
rect -649 -488 -615 488
rect -491 -488 -457 488
rect -333 -488 -299 488
rect -175 -488 -141 488
rect -17 -488 17 488
rect 141 -488 175 488
rect 299 -488 333 488
rect 457 -488 491 488
rect 615 -488 649 488
rect 773 -488 807 488
rect 931 -488 965 488
rect 1089 -488 1123 488
rect 1247 -488 1281 488
rect 1405 -488 1439 488
rect 1563 -488 1597 488
<< metal1 >>
rect -1603 488 -1557 500
rect -1603 -488 -1597 488
rect -1563 -488 -1557 488
rect -1603 -500 -1557 -488
rect -1445 488 -1399 500
rect -1445 -488 -1439 488
rect -1405 -488 -1399 488
rect -1445 -500 -1399 -488
rect -1287 488 -1241 500
rect -1287 -488 -1281 488
rect -1247 -488 -1241 488
rect -1287 -500 -1241 -488
rect -1129 488 -1083 500
rect -1129 -488 -1123 488
rect -1089 -488 -1083 488
rect -1129 -500 -1083 -488
rect -971 488 -925 500
rect -971 -488 -965 488
rect -931 -488 -925 488
rect -971 -500 -925 -488
rect -813 488 -767 500
rect -813 -488 -807 488
rect -773 -488 -767 488
rect -813 -500 -767 -488
rect -655 488 -609 500
rect -655 -488 -649 488
rect -615 -488 -609 488
rect -655 -500 -609 -488
rect -497 488 -451 500
rect -497 -488 -491 488
rect -457 -488 -451 488
rect -497 -500 -451 -488
rect -339 488 -293 500
rect -339 -488 -333 488
rect -299 -488 -293 488
rect -339 -500 -293 -488
rect -181 488 -135 500
rect -181 -488 -175 488
rect -141 -488 -135 488
rect -181 -500 -135 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 135 488 181 500
rect 135 -488 141 488
rect 175 -488 181 488
rect 135 -500 181 -488
rect 293 488 339 500
rect 293 -488 299 488
rect 333 -488 339 488
rect 293 -500 339 -488
rect 451 488 497 500
rect 451 -488 457 488
rect 491 -488 497 488
rect 451 -500 497 -488
rect 609 488 655 500
rect 609 -488 615 488
rect 649 -488 655 488
rect 609 -500 655 -488
rect 767 488 813 500
rect 767 -488 773 488
rect 807 -488 813 488
rect 767 -500 813 -488
rect 925 488 971 500
rect 925 -488 931 488
rect 965 -488 971 488
rect 925 -500 971 -488
rect 1083 488 1129 500
rect 1083 -488 1089 488
rect 1123 -488 1129 488
rect 1083 -500 1129 -488
rect 1241 488 1287 500
rect 1241 -488 1247 488
rect 1281 -488 1287 488
rect 1241 -500 1287 -488
rect 1399 488 1445 500
rect 1399 -488 1405 488
rect 1439 -488 1445 488
rect 1399 -500 1445 -488
rect 1557 488 1603 500
rect 1557 -488 1563 488
rect 1597 -488 1603 488
rect 1557 -500 1603 -488
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string parameters w 5 l 0.5 m 1 nf 20 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
