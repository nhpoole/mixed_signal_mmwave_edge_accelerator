magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect 3116 -7662 92653 2722
<< metal2 >>
rect 13914 1401 13970 1449
rect 16410 1401 16466 1449
rect 18906 1401 18962 1449
rect 21402 1401 21458 1449
rect 23898 1401 23954 1449
rect 26394 1401 26450 1449
rect 28890 1401 28946 1449
rect 31386 1401 31442 1449
rect 33882 1401 33938 1449
rect 36378 1401 36434 1449
rect 38874 1401 38930 1449
rect 41370 1401 41426 1449
rect 43866 1401 43922 1449
rect 46362 1401 46418 1449
rect 48858 1401 48914 1449
rect 51354 1401 51410 1449
rect 53850 1401 53906 1449
rect 56346 1401 56402 1449
rect 58842 1401 58898 1449
rect 61338 1401 61394 1449
rect 63834 1401 63890 1449
rect 66330 1401 66386 1449
rect 68826 1401 68882 1449
rect 71322 1401 71378 1449
rect 73818 1401 73874 1449
rect 76314 1401 76370 1449
rect 78810 1401 78866 1449
rect 81306 1401 81362 1449
rect 83802 1401 83858 1449
rect 86298 1401 86354 1449
rect 88794 1401 88850 1449
rect 91290 1401 91346 1449
<< metal3 >>
rect 13867 1393 14017 1457
rect 16363 1393 16513 1457
rect 18859 1393 19009 1457
rect 21355 1393 21505 1457
rect 23851 1393 24001 1457
rect 26347 1393 26497 1457
rect 28843 1393 28993 1457
rect 31339 1393 31489 1457
rect 33835 1393 33985 1457
rect 36331 1393 36481 1457
rect 38827 1393 38977 1457
rect 41323 1393 41473 1457
rect 43819 1393 43969 1457
rect 46315 1393 46465 1457
rect 48811 1393 48961 1457
rect 51307 1393 51457 1457
rect 53803 1393 53953 1457
rect 56299 1393 56449 1457
rect 58795 1393 58945 1457
rect 61291 1393 61441 1457
rect 63787 1393 63937 1457
rect 66283 1393 66433 1457
rect 68779 1393 68929 1457
rect 71275 1393 71425 1457
rect 73771 1393 73921 1457
rect 76267 1393 76417 1457
rect 78763 1393 78913 1457
rect 81259 1393 81409 1457
rect 83755 1393 83905 1457
rect 86251 1393 86401 1457
rect 88747 1393 88897 1457
rect 91243 1393 91393 1457
rect 13582 273 13732 337
rect 33550 273 33700 337
rect 53518 273 53668 337
rect 73486 273 73636 337
rect 44163 -514 88822 -454
rect 42995 -758 86326 -698
rect 40659 -1002 81334 -942
rect 38323 -1246 76342 -1186
rect 5619 -1490 33625 -1430
rect 35987 -1490 71350 -1430
rect 33651 -1734 66358 -1674
rect 17299 -1978 31414 -1918
rect 32483 -1978 63862 -1918
rect 31315 -2222 61366 -2162
rect 16131 -2466 28918 -2406
rect 30147 -2466 58870 -2406
rect 28979 -2710 56374 -2650
rect 14963 -2954 26422 -2894
rect 27811 -2954 53878 -2894
rect 26643 -3198 51382 -3138
rect 25475 -3442 48886 -3382
rect 9123 -3686 13942 -3626
rect 23139 -3686 43894 -3626
rect 45331 -3686 91318 -3626
rect 4451 -3930 13657 -3870
rect 20803 -3930 38902 -3870
rect 39491 -3930 78838 -3870
rect 13795 -4174 23926 -4114
rect 24307 -4174 46390 -4114
rect 12627 -4418 21430 -4358
rect 21971 -4418 41398 -4358
rect 41827 -4418 83830 -4358
rect 11459 -4662 18934 -4602
rect 19635 -4662 36406 -4602
rect 37155 -4662 73846 -4602
rect 10291 -4906 16438 -4846
rect 18467 -4906 33910 -4846
rect 34819 -4906 68854 -4846
rect 7955 -5150 73561 -5090
rect 6787 -5394 53593 -5334
rect 4376 -6397 4526 -6333
rect 5544 -6397 5694 -6333
rect 6712 -6397 6862 -6333
rect 7880 -6397 8030 -6333
rect 9048 -6397 9198 -6333
rect 10216 -6397 10366 -6333
rect 11384 -6397 11534 -6333
rect 12552 -6397 12702 -6333
rect 13720 -6397 13870 -6333
rect 14888 -6397 15038 -6333
rect 16056 -6397 16206 -6333
rect 17224 -6397 17374 -6333
rect 18392 -6397 18542 -6333
rect 19560 -6397 19710 -6333
rect 20728 -6397 20878 -6333
rect 21896 -6397 22046 -6333
rect 23064 -6397 23214 -6333
rect 24232 -6397 24382 -6333
rect 25400 -6397 25550 -6333
rect 26568 -6397 26718 -6333
rect 27736 -6397 27886 -6333
rect 28904 -6397 29054 -6333
rect 30072 -6397 30222 -6333
rect 31240 -6397 31390 -6333
rect 32408 -6397 32558 -6333
rect 33576 -6397 33726 -6333
rect 34744 -6397 34894 -6333
rect 35912 -6397 36062 -6333
rect 37080 -6397 37230 -6333
rect 38248 -6397 38398 -6333
rect 39416 -6397 39566 -6333
rect 40584 -6397 40734 -6333
rect 41752 -6397 41902 -6333
rect 42920 -6397 43070 -6333
rect 44088 -6397 44238 -6333
rect 45256 -6397 45406 -6333
<< metal4 >>
rect 4421 -6365 4481 -3900
rect 5589 -6365 5649 -1460
rect 6757 -6365 6817 -5364
rect 7925 -6365 7985 -5120
rect 9093 -6365 9153 -3656
rect 13627 -3900 13687 305
rect 13912 -3656 13972 1425
rect 10261 -6365 10321 -4876
rect 11429 -6365 11489 -4632
rect 12597 -6365 12657 -4388
rect 13765 -6365 13825 -4144
rect 14933 -6365 14993 -2924
rect 16101 -6365 16161 -2436
rect 16408 -4876 16468 1425
rect 17269 -6365 17329 -1948
rect 18904 -4632 18964 1425
rect 18437 -6365 18497 -4876
rect 19605 -6365 19665 -4632
rect 20773 -6365 20833 -3900
rect 21400 -4388 21460 1425
rect 21941 -6365 22001 -4388
rect 23109 -6365 23169 -3656
rect 23896 -4144 23956 1425
rect 26392 -2924 26452 1425
rect 28888 -2436 28948 1425
rect 31384 -1948 31444 1425
rect 33595 -1460 33655 305
rect 24277 -6365 24337 -4144
rect 25445 -6365 25505 -3412
rect 26613 -6365 26673 -3168
rect 27781 -6365 27841 -2924
rect 28949 -6365 29009 -2680
rect 30117 -6365 30177 -2436
rect 31285 -6365 31345 -2192
rect 32453 -6365 32513 -1948
rect 33621 -6365 33681 -1704
rect 33880 -4876 33940 1425
rect 34789 -6365 34849 -4876
rect 35957 -6365 36017 -1460
rect 36376 -4632 36436 1425
rect 37125 -6365 37185 -4632
rect 38293 -6365 38353 -1216
rect 38872 -3900 38932 1425
rect 39461 -6365 39521 -3900
rect 40629 -6365 40689 -972
rect 41368 -4388 41428 1425
rect 41797 -6365 41857 -4388
rect 42965 -6365 43025 -728
rect 43864 -3656 43924 1425
rect 44133 -6365 44193 -484
rect 45301 -6365 45361 -3656
rect 46360 -4144 46420 1425
rect 48856 -3412 48916 1425
rect 51352 -3168 51412 1425
rect 53563 -5364 53623 305
rect 53848 -2924 53908 1425
rect 56344 -2680 56404 1425
rect 58840 -2436 58900 1425
rect 61336 -2192 61396 1425
rect 63832 -1948 63892 1425
rect 66328 -1704 66388 1425
rect 68824 -4876 68884 1425
rect 71320 -1460 71380 1425
rect 73531 -5120 73591 305
rect 73816 -4632 73876 1425
rect 76312 -1216 76372 1425
rect 78808 -3900 78868 1425
rect 81304 -972 81364 1425
rect 83800 -4388 83860 1425
rect 86296 -728 86356 1425
rect 88792 -484 88852 1425
rect 91288 -3656 91348 1425
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_71
timestamp 1626486988
transform 1 0 53560 0 1 268
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_70
timestamp 1626486988
transform 1 0 73528 0 1 268
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_69
timestamp 1626486988
transform 1 0 68821 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_68
timestamp 1626486988
transform 1 0 73813 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_67
timestamp 1626486988
transform 1 0 83797 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_66
timestamp 1626486988
transform 1 0 78805 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_65
timestamp 1626486988
transform 1 0 91285 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_64
timestamp 1626486988
transform 1 0 48853 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_63
timestamp 1626486988
transform 1 0 51349 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_62
timestamp 1626486988
transform 1 0 53845 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_61
timestamp 1626486988
transform 1 0 56341 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_60
timestamp 1626486988
transform 1 0 58837 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_59
timestamp 1626486988
transform 1 0 61333 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_58
timestamp 1626486988
transform 1 0 63829 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_57
timestamp 1626486988
transform 1 0 66325 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_56
timestamp 1626486988
transform 1 0 71317 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_55
timestamp 1626486988
transform 1 0 76309 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_54
timestamp 1626486988
transform 1 0 81301 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_53
timestamp 1626486988
transform 1 0 86293 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_52
timestamp 1626486988
transform 1 0 88789 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_51
timestamp 1626486988
transform 1 0 46357 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_50
timestamp 1626486988
transform 1 0 38869 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_49
timestamp 1626486988
transform 1 0 33877 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_48
timestamp 1626486988
transform 1 0 39458 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_47
timestamp 1626486988
transform 1 0 43861 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_46
timestamp 1626486988
transform 1 0 45298 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_45
timestamp 1626486988
transform 1 0 34786 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_44
timestamp 1626486988
transform 1 0 26610 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_43
timestamp 1626486988
transform 1 0 26389 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_42
timestamp 1626486988
transform 1 0 27778 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_41
timestamp 1626486988
transform 1 0 28946 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_40
timestamp 1626486988
transform 1 0 28885 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_39
timestamp 1626486988
transform 1 0 36373 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_38
timestamp 1626486988
transform 1 0 30114 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_37
timestamp 1626486988
transform 1 0 31282 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_36
timestamp 1626486988
transform 1 0 31381 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_35
timestamp 1626486988
transform 1 0 37122 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_34
timestamp 1626486988
transform 1 0 32450 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_33
timestamp 1626486988
transform 1 0 33618 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_32
timestamp 1626486988
transform 1 0 33592 0 1 268
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_31
timestamp 1626486988
transform 1 0 35954 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_30
timestamp 1626486988
transform 1 0 41365 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_29
timestamp 1626486988
transform 1 0 38290 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_28
timestamp 1626486988
transform 1 0 40626 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_27
timestamp 1626486988
transform 1 0 41794 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_26
timestamp 1626486988
transform 1 0 42962 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_25
timestamp 1626486988
transform 1 0 44130 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_24
timestamp 1626486988
transform 1 0 23106 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_23
timestamp 1626486988
transform 1 0 16098 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_22
timestamp 1626486988
transform 1 0 19602 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_21
timestamp 1626486988
transform 1 0 18434 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_20
timestamp 1626486988
transform 1 0 7922 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_19
timestamp 1626486988
transform 1 0 13762 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_18
timestamp 1626486988
transform 1 0 6754 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_17
timestamp 1626486988
transform 1 0 17266 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_16
timestamp 1626486988
transform 1 0 25442 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_15
timestamp 1626486988
transform 1 0 20770 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_14
timestamp 1626486988
transform 1 0 21397 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_13
timestamp 1626486988
transform 1 0 24274 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_12
timestamp 1626486988
transform 1 0 13624 0 1 268
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_11
timestamp 1626486988
transform 1 0 5586 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_10
timestamp 1626486988
transform 1 0 12594 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_9
timestamp 1626486988
transform 1 0 14930 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_8
timestamp 1626486988
transform 1 0 18901 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_7
timestamp 1626486988
transform 1 0 21938 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_6
timestamp 1626486988
transform 1 0 16405 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_5
timestamp 1626486988
transform 1 0 13909 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_4
timestamp 1626486988
transform 1 0 11426 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_3
timestamp 1626486988
transform 1 0 10258 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_2
timestamp 1626486988
transform 1 0 9090 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_1
timestamp 1626486988
transform 1 0 4418 0 1 -6402
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_0
timestamp 1626486988
transform 1 0 23893 0 1 1388
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_31
timestamp 1626486988
transform 1 0 68822 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_30
timestamp 1626486988
transform 1 0 73814 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_29
timestamp 1626486988
transform 1 0 83798 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_28
timestamp 1626486988
transform 1 0 78806 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_27
timestamp 1626486988
transform 1 0 91286 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_26
timestamp 1626486988
transform 1 0 48854 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_25
timestamp 1626486988
transform 1 0 51350 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_24
timestamp 1626486988
transform 1 0 53846 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_23
timestamp 1626486988
transform 1 0 56342 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_22
timestamp 1626486988
transform 1 0 58838 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_21
timestamp 1626486988
transform 1 0 61334 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_20
timestamp 1626486988
transform 1 0 63830 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_19
timestamp 1626486988
transform 1 0 66326 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_18
timestamp 1626486988
transform 1 0 71318 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_17
timestamp 1626486988
transform 1 0 76310 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_16
timestamp 1626486988
transform 1 0 81302 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_15
timestamp 1626486988
transform 1 0 86294 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_14
timestamp 1626486988
transform 1 0 88790 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_13
timestamp 1626486988
transform 1 0 46358 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_12
timestamp 1626486988
transform 1 0 38870 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_11
timestamp 1626486988
transform 1 0 33878 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_10
timestamp 1626486988
transform 1 0 43862 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_9
timestamp 1626486988
transform 1 0 26390 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_8
timestamp 1626486988
transform 1 0 36374 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_7
timestamp 1626486988
transform 1 0 28886 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_6
timestamp 1626486988
transform 1 0 31382 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_5
timestamp 1626486988
transform 1 0 41366 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_4
timestamp 1626486988
transform 1 0 16406 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_3
timestamp 1626486988
transform 1 0 21398 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_2
timestamp 1626486988
transform 1 0 18902 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_1
timestamp 1626486988
transform 1 0 13910 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_0
timestamp 1626486988
transform 1 0 23894 0 1 1393
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_143
timestamp 1626486988
transform 1 0 53555 0 1 -5397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_142
timestamp 1626486988
transform 1 0 53555 0 1 272
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_141
timestamp 1626486988
transform 1 0 73523 0 1 -5153
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_140
timestamp 1626486988
transform 1 0 73523 0 1 272
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_139
timestamp 1626486988
transform 1 0 68816 0 1 -4909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_138
timestamp 1626486988
transform 1 0 68816 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_137
timestamp 1626486988
transform 1 0 73808 0 1 -4665
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_136
timestamp 1626486988
transform 1 0 73808 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_135
timestamp 1626486988
transform 1 0 83792 0 1 -4421
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_134
timestamp 1626486988
transform 1 0 83792 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_133
timestamp 1626486988
transform 1 0 78800 0 1 -3933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_132
timestamp 1626486988
transform 1 0 78800 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_131
timestamp 1626486988
transform 1 0 91280 0 1 -3689
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_130
timestamp 1626486988
transform 1 0 91280 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_129
timestamp 1626486988
transform 1 0 48848 0 1 -3445
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_128
timestamp 1626486988
transform 1 0 48848 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_127
timestamp 1626486988
transform 1 0 51344 0 1 -3201
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_126
timestamp 1626486988
transform 1 0 51344 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_125
timestamp 1626486988
transform 1 0 53840 0 1 -2957
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_124
timestamp 1626486988
transform 1 0 53840 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_123
timestamp 1626486988
transform 1 0 56336 0 1 -2713
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_122
timestamp 1626486988
transform 1 0 56336 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_121
timestamp 1626486988
transform 1 0 58832 0 1 -2469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_120
timestamp 1626486988
transform 1 0 58832 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_119
timestamp 1626486988
transform 1 0 61328 0 1 -2225
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_118
timestamp 1626486988
transform 1 0 61328 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_117
timestamp 1626486988
transform 1 0 63824 0 1 -1981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_116
timestamp 1626486988
transform 1 0 63824 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_115
timestamp 1626486988
transform 1 0 66320 0 1 -1737
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_114
timestamp 1626486988
transform 1 0 66320 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_113
timestamp 1626486988
transform 1 0 71312 0 1 -1493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_112
timestamp 1626486988
transform 1 0 71312 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_111
timestamp 1626486988
transform 1 0 76304 0 1 -1249
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_110
timestamp 1626486988
transform 1 0 76304 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_109
timestamp 1626486988
transform 1 0 81296 0 1 -1005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_108
timestamp 1626486988
transform 1 0 81296 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_107
timestamp 1626486988
transform 1 0 86288 0 1 -761
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_106
timestamp 1626486988
transform 1 0 86288 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_105
timestamp 1626486988
transform 1 0 88784 0 1 -517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_104
timestamp 1626486988
transform 1 0 88784 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_103
timestamp 1626486988
transform 1 0 46352 0 1 -4177
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_102
timestamp 1626486988
transform 1 0 46352 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_101
timestamp 1626486988
transform 1 0 38864 0 1 -3933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_100
timestamp 1626486988
transform 1 0 38864 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_99
timestamp 1626486988
transform 1 0 33872 0 1 -4909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_98
timestamp 1626486988
transform 1 0 39453 0 1 -3933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_97
timestamp 1626486988
transform 1 0 39453 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_96
timestamp 1626486988
transform 1 0 43856 0 1 -3689
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_95
timestamp 1626486988
transform 1 0 43856 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_94
timestamp 1626486988
transform 1 0 33872 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_93
timestamp 1626486988
transform 1 0 45293 0 1 -3689
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_92
timestamp 1626486988
transform 1 0 45293 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_91
timestamp 1626486988
transform 1 0 34781 0 1 -4909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_90
timestamp 1626486988
transform 1 0 34781 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_89
timestamp 1626486988
transform 1 0 26605 0 1 -3201
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_88
timestamp 1626486988
transform 1 0 26605 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_87
timestamp 1626486988
transform 1 0 26384 0 1 -2957
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_86
timestamp 1626486988
transform 1 0 26384 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_85
timestamp 1626486988
transform 1 0 27773 0 1 -2957
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_84
timestamp 1626486988
transform 1 0 27773 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_83
timestamp 1626486988
transform 1 0 36368 0 1 -4665
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_82
timestamp 1626486988
transform 1 0 28941 0 1 -2713
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_81
timestamp 1626486988
transform 1 0 28941 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_80
timestamp 1626486988
transform 1 0 28880 0 1 -2469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_79
timestamp 1626486988
transform 1 0 28880 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_78
timestamp 1626486988
transform 1 0 36368 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_77
timestamp 1626486988
transform 1 0 30109 0 1 -2469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_76
timestamp 1626486988
transform 1 0 30109 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_75
timestamp 1626486988
transform 1 0 31277 0 1 -2225
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_74
timestamp 1626486988
transform 1 0 31277 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_73
timestamp 1626486988
transform 1 0 31376 0 1 -1981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_72
timestamp 1626486988
transform 1 0 31376 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_71
timestamp 1626486988
transform 1 0 37117 0 1 -4665
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_70
timestamp 1626486988
transform 1 0 37117 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_69
timestamp 1626486988
transform 1 0 32445 0 1 -1981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_68
timestamp 1626486988
transform 1 0 32445 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_67
timestamp 1626486988
transform 1 0 33613 0 1 -1737
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_66
timestamp 1626486988
transform 1 0 33613 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_65
timestamp 1626486988
transform 1 0 33587 0 1 -1493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_64
timestamp 1626486988
transform 1 0 33587 0 1 272
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_63
timestamp 1626486988
transform 1 0 41360 0 1 -4421
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_62
timestamp 1626486988
transform 1 0 35949 0 1 -1493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_61
timestamp 1626486988
transform 1 0 35949 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_60
timestamp 1626486988
transform 1 0 41360 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_59
timestamp 1626486988
transform 1 0 38285 0 1 -1249
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_58
timestamp 1626486988
transform 1 0 38285 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_57
timestamp 1626486988
transform 1 0 40621 0 1 -1005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_56
timestamp 1626486988
transform 1 0 40621 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_55
timestamp 1626486988
transform 1 0 41789 0 1 -4421
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_54
timestamp 1626486988
transform 1 0 42957 0 1 -761
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_53
timestamp 1626486988
transform 1 0 42957 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_52
timestamp 1626486988
transform 1 0 41789 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_51
timestamp 1626486988
transform 1 0 44125 0 1 -517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_50
timestamp 1626486988
transform 1 0 44125 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_49
timestamp 1626486988
transform 1 0 16093 0 1 -2469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_48
timestamp 1626486988
transform 1 0 16093 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_47
timestamp 1626486988
transform 1 0 23101 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_46
timestamp 1626486988
transform 1 0 13757 0 1 -4177
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_45
timestamp 1626486988
transform 1 0 19597 0 1 -4665
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_44
timestamp 1626486988
transform 1 0 18429 0 1 -4909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_43
timestamp 1626486988
transform 1 0 18429 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_42
timestamp 1626486988
transform 1 0 19597 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_41
timestamp 1626486988
transform 1 0 7917 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_40
timestamp 1626486988
transform 1 0 16400 0 1 -4909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_39
timestamp 1626486988
transform 1 0 13757 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_38
timestamp 1626486988
transform 1 0 20765 0 1 -3933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_37
timestamp 1626486988
transform 1 0 6749 0 1 -5397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_36
timestamp 1626486988
transform 1 0 6749 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_35
timestamp 1626486988
transform 1 0 7917 0 1 -5153
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_34
timestamp 1626486988
transform 1 0 17261 0 1 -1981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_33
timestamp 1626486988
transform 1 0 17261 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_32
timestamp 1626486988
transform 1 0 25437 0 1 -3445
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_31
timestamp 1626486988
transform 1 0 25437 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_30
timestamp 1626486988
transform 1 0 20765 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_29
timestamp 1626486988
transform 1 0 10253 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_28
timestamp 1626486988
transform 1 0 21392 0 1 -4421
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_27
timestamp 1626486988
transform 1 0 21392 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_26
timestamp 1626486988
transform 1 0 18896 0 1 -4665
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_25
timestamp 1626486988
transform 1 0 24269 0 1 -4177
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_24
timestamp 1626486988
transform 1 0 24269 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_23
timestamp 1626486988
transform 1 0 13619 0 1 -3933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_22
timestamp 1626486988
transform 1 0 5581 0 1 -1493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_21
timestamp 1626486988
transform 1 0 5581 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_20
timestamp 1626486988
transform 1 0 12589 0 1 -4421
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_19
timestamp 1626486988
transform 1 0 12589 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_18
timestamp 1626486988
transform 1 0 13619 0 1 272
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_17
timestamp 1626486988
transform 1 0 13904 0 1 -3689
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_16
timestamp 1626486988
transform 1 0 14925 0 1 -2957
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_15
timestamp 1626486988
transform 1 0 14925 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_14
timestamp 1626486988
transform 1 0 21933 0 1 -4421
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_13
timestamp 1626486988
transform 1 0 18896 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_12
timestamp 1626486988
transform 1 0 11421 0 1 -4665
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_11
timestamp 1626486988
transform 1 0 21933 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_10
timestamp 1626486988
transform 1 0 16400 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_9
timestamp 1626486988
transform 1 0 13904 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_8
timestamp 1626486988
transform 1 0 10253 0 1 -4909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_7
timestamp 1626486988
transform 1 0 11421 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_6
timestamp 1626486988
transform 1 0 9085 0 1 -3689
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_5
timestamp 1626486988
transform 1 0 9085 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_4
timestamp 1626486988
transform 1 0 4413 0 1 -3933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3
timestamp 1626486988
transform 1 0 23888 0 1 -4177
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2
timestamp 1626486988
transform 1 0 4413 0 1 -6398
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1
timestamp 1626486988
transform 1 0 23888 0 1 1392
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_0
timestamp 1626486988
transform 1 0 23101 0 1 -3689
box 0 0 76 66
<< properties >>
string FIXED_BBOX 4376 -6402 91393 1462
<< end >>
