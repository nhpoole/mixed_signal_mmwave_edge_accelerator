magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -1286 -1286 1436 1862
<< pwell >>
rect -26 -26 176 602
<< scnmos >>
rect 60 0 90 576
<< ndiff >>
rect 0 0 60 576
rect 90 0 150 576
<< poly >>
rect 60 576 90 602
rect 60 -26 90 0
<< locali >>
rect 8 255 42 321
rect 108 255 142 321
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_11  sky130_sram_2kbyte_1rw1r_32x512_8_contact_11_0
timestamp 1626065694
transform 1 0 100 0 1 255
box -26 -22 76 88
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_11  sky130_sram_2kbyte_1rw1r_32x512_8_contact_11_1
timestamp 1626065694
transform 1 0 0 0 1 255
box -26 -22 76 88
<< labels >>
rlabel locali s 25 288 25 288 4 S
rlabel locali s 125 288 125 288 4 D
rlabel poly s 75 288 75 288 4 G
<< properties >>
string FIXED_BBOX -25 -26 175 602
<< end >>
