magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< metal1 >>
rect 552 1388 616 1440
rect 1720 1388 1784 1440
rect 2888 1388 2952 1440
rect 4056 1388 4120 1440
rect 552 -26 616 26
rect 1720 -26 1784 26
rect 2888 -26 2952 26
rect 4056 -26 4120 26
<< metal2 >>
rect 137 538 203 590
rect 369 0 397 1414
rect 556 1390 612 1438
rect 1082 609 1148 661
rect 1305 538 1371 590
rect 556 -24 612 24
rect 1537 0 1565 1414
rect 1724 1390 1780 1438
rect 2250 609 2316 661
rect 2473 538 2539 590
rect 1724 -24 1780 24
rect 2705 0 2733 1414
rect 2892 1390 2948 1438
rect 3418 609 3484 661
rect 3641 538 3707 590
rect 2892 -24 2948 24
rect 3873 0 3901 1414
rect 4060 1390 4116 1438
rect 4586 609 4652 661
rect 4060 -24 4116 24
<< metal3 >>
rect 535 1365 633 1463
rect 1703 1365 1801 1463
rect 2871 1365 2969 1463
rect 4039 1365 4137 1463
rect 0 278 4672 338
rect 535 -49 633 49
rect 1703 -49 1801 49
rect 2871 -49 2969 49
rect 4039 -49 4137 49
use contact_9  contact_9_3
timestamp 1624494425
transform 1 0 363 0 1 271
box 0 0 66 74
use contact_9  contact_9_10
timestamp 1624494425
transform 1 0 551 0 1 -37
box 0 0 66 74
use contact_9  contact_9_11
timestamp 1624494425
transform 1 0 551 0 1 1377
box 0 0 66 74
use contact_8  contact_8_6
timestamp 1624494425
transform 1 0 552 0 1 -32
box 0 0 64 64
use contact_8  contact_8_7
timestamp 1624494425
transform 1 0 552 0 1 1382
box 0 0 64 64
use contact_7  contact_7_6
timestamp 1624494425
transform 1 0 555 0 1 -33
box 0 0 58 66
use contact_7  contact_7_7
timestamp 1624494425
transform 1 0 555 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_2
timestamp 1624494425
transform 1 0 1168 0 1 0
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_3
timestamp 1624494425
transform 1 0 0 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_2
timestamp 1624494425
transform 1 0 1531 0 1 271
box 0 0 66 74
use contact_9  contact_9_8
timestamp 1624494425
transform 1 0 1719 0 1 -37
box 0 0 66 74
use contact_9  contact_9_9
timestamp 1624494425
transform 1 0 1719 0 1 1377
box 0 0 66 74
use contact_8  contact_8_4
timestamp 1624494425
transform 1 0 1720 0 1 -32
box 0 0 64 64
use contact_8  contact_8_5
timestamp 1624494425
transform 1 0 1720 0 1 1382
box 0 0 64 64
use contact_7  contact_7_4
timestamp 1624494425
transform 1 0 1723 0 1 -33
box 0 0 58 66
use contact_7  contact_7_5
timestamp 1624494425
transform 1 0 1723 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_1
timestamp 1624494425
transform 1 0 2336 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_1
timestamp 1624494425
transform 1 0 2699 0 1 271
box 0 0 66 74
use contact_9  contact_9_6
timestamp 1624494425
transform 1 0 2887 0 1 -37
box 0 0 66 74
use contact_9  contact_9_7
timestamp 1624494425
transform 1 0 2887 0 1 1377
box 0 0 66 74
use contact_8  contact_8_2
timestamp 1624494425
transform 1 0 2888 0 1 -32
box 0 0 64 64
use contact_8  contact_8_3
timestamp 1624494425
transform 1 0 2888 0 1 1382
box 0 0 64 64
use contact_7  contact_7_2
timestamp 1624494425
transform 1 0 2891 0 1 -33
box 0 0 58 66
use contact_7  contact_7_3
timestamp 1624494425
transform 1 0 2891 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_0
timestamp 1624494425
transform 1 0 3504 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_0
timestamp 1624494425
transform 1 0 3867 0 1 271
box 0 0 66 74
use contact_9  contact_9_4
timestamp 1624494425
transform 1 0 4055 0 1 -37
box 0 0 66 74
use contact_9  contact_9_5
timestamp 1624494425
transform 1 0 4055 0 1 1377
box 0 0 66 74
use contact_8  contact_8_0
timestamp 1624494425
transform 1 0 4056 0 1 -32
box 0 0 64 64
use contact_8  contact_8_1
timestamp 1624494425
transform 1 0 4056 0 1 1382
box 0 0 64 64
use contact_7  contact_7_0
timestamp 1624494425
transform 1 0 4059 0 1 -33
box 0 0 58 66
use contact_7  contact_7_1
timestamp 1624494425
transform 1 0 4059 0 1 1381
box 0 0 58 66
<< labels >>
rlabel metal3 s 4039 1365 4137 1463 4 vdd
rlabel metal3 s 535 1365 633 1463 4 vdd
rlabel metal3 s 1703 1365 1801 1463 4 vdd
rlabel metal3 s 2871 1365 2969 1463 4 vdd
rlabel metal3 s 535 -49 633 49 4 gnd
rlabel metal3 s 1703 -49 1801 49 4 gnd
rlabel metal3 s 2871 -49 2969 49 4 gnd
rlabel metal3 s 4039 -49 4137 49 4 gnd
rlabel metal2 s 137 538 203 590 4 din_0
rlabel metal2 s 1082 609 1148 661 4 dout_0
rlabel metal2 s 1305 538 1371 590 4 din_1
rlabel metal2 s 2250 609 2316 661 4 dout_1
rlabel metal2 s 2473 538 2539 590 4 din_2
rlabel metal2 s 3418 609 3484 661 4 dout_2
rlabel metal2 s 3641 538 3707 590 4 din_3
rlabel metal2 s 4586 609 4652 661 4 dout_3
rlabel metal3 s 0 278 4672 338 4 clk
<< properties >>
string FIXED_BBOX 0 0 4672 1414
<< end >>
